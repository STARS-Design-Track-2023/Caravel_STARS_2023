magic
tech sky130A
magscale 1 2
timestamp 1691529705
<< viali >>
rect 19441 42313 19475 42347
rect 30573 42313 30607 42347
rect 38301 42313 38335 42347
rect 1869 42245 1903 42279
rect 7297 42245 7331 42279
rect 11621 42245 11655 42279
rect 34805 42245 34839 42279
rect 1501 42177 1535 42211
rect 3341 42177 3375 42211
rect 11253 42177 11287 42211
rect 11529 42177 11563 42211
rect 14657 42177 14691 42211
rect 15209 42177 15243 42211
rect 19349 42177 19383 42211
rect 22661 42177 22695 42211
rect 30481 42177 30515 42211
rect 38209 42177 38243 42211
rect 41061 42177 41095 42211
rect 15393 42109 15427 42143
rect 32689 42109 32723 42143
rect 7481 42041 7515 42075
rect 11069 42041 11103 42075
rect 3525 41973 3559 42007
rect 14933 41973 14967 42007
rect 22845 41973 22879 42007
rect 33333 41973 33367 42007
rect 34897 41973 34931 42007
rect 40877 41973 40911 42007
rect 23949 41769 23983 41803
rect 28733 41769 28767 41803
rect 30922 41769 30956 41803
rect 32413 41769 32447 41803
rect 19625 41701 19659 41735
rect 20729 41701 20763 41735
rect 11069 41633 11103 41667
rect 14105 41633 14139 41667
rect 19901 41633 19935 41667
rect 19993 41633 20027 41667
rect 22569 41633 22603 41667
rect 28549 41633 28583 41667
rect 30665 41633 30699 41667
rect 32597 41633 32631 41667
rect 32873 41633 32907 41667
rect 10517 41565 10551 41599
rect 11437 41565 11471 41599
rect 13553 41565 13587 41599
rect 13645 41565 13679 41599
rect 15945 41565 15979 41599
rect 16589 41565 16623 41599
rect 16773 41565 16807 41599
rect 18245 41565 18279 41599
rect 18429 41565 18463 41599
rect 19809 41565 19843 41599
rect 20085 41565 20119 41599
rect 20453 41565 20487 41599
rect 20637 41565 20671 41599
rect 22385 41565 22419 41599
rect 22753 41565 22787 41599
rect 23857 41565 23891 41599
rect 24409 41565 24443 41599
rect 24685 41565 24719 41599
rect 26525 41565 26559 41599
rect 28733 41565 28767 41599
rect 14381 41497 14415 41531
rect 17141 41497 17175 41531
rect 18521 41497 18555 41531
rect 18705 41497 18739 41531
rect 19073 41497 19107 41531
rect 22017 41497 22051 41531
rect 24593 41497 24627 41531
rect 25145 41497 25179 41531
rect 26157 41497 26191 41531
rect 26341 41497 26375 41531
rect 26709 41497 26743 41531
rect 27077 41497 27111 41531
rect 28457 41497 28491 41531
rect 10609 41429 10643 41463
rect 12863 41429 12897 41463
rect 13369 41429 13403 41463
rect 13829 41429 13863 41463
rect 15853 41429 15887 41463
rect 22201 41429 22235 41463
rect 22293 41429 22327 41463
rect 22937 41429 22971 41463
rect 28917 41429 28951 41463
rect 34345 41429 34379 41463
rect 11161 41225 11195 41259
rect 14289 41225 14323 41259
rect 14657 41225 14691 41259
rect 17693 41225 17727 41259
rect 24593 41225 24627 41259
rect 25881 41225 25915 41259
rect 16405 41157 16439 41191
rect 18061 41157 18095 41191
rect 20545 41157 20579 41191
rect 24317 41157 24351 41191
rect 25237 41157 25271 41191
rect 25789 41157 25823 41191
rect 28917 41157 28951 41191
rect 29009 41157 29043 41191
rect 31125 41157 31159 41191
rect 11345 41089 11379 41123
rect 12725 41089 12759 41123
rect 15485 41089 15519 41123
rect 15577 41089 15611 41123
rect 15669 41089 15703 41123
rect 15853 41089 15887 41123
rect 16221 41089 16255 41123
rect 16497 41089 16531 41123
rect 16773 41089 16807 41123
rect 17141 41089 17175 41123
rect 17877 41089 17911 41123
rect 17969 41089 18003 41123
rect 18153 41089 18187 41123
rect 18613 41089 18647 41123
rect 19073 41089 19107 41123
rect 19697 41089 19731 41123
rect 19809 41089 19843 41123
rect 19901 41089 19935 41123
rect 20085 41089 20119 41123
rect 20453 41089 20487 41123
rect 20913 41089 20947 41123
rect 21005 41089 21039 41123
rect 21833 41089 21867 41123
rect 22017 41089 22051 41123
rect 23213 41089 23247 41123
rect 23581 41089 23615 41123
rect 25053 41089 25087 41123
rect 25329 41089 25363 41123
rect 25421 41089 25455 41123
rect 26341 41089 26375 41123
rect 26617 41089 26651 41123
rect 26985 41089 27019 41123
rect 27169 41089 27203 41123
rect 27261 41089 27295 41123
rect 27353 41089 27387 41123
rect 27629 41089 27663 41123
rect 27997 41089 28031 41123
rect 28090 41089 28124 41123
rect 28273 41089 28307 41123
rect 28365 41089 28399 41123
rect 28462 41089 28496 41123
rect 28733 41089 28767 41123
rect 29101 41089 29135 41123
rect 29377 41089 29411 41123
rect 29653 41089 29687 41123
rect 30757 41089 30791 41123
rect 32137 41089 32171 41123
rect 40325 41089 40359 41123
rect 40601 41089 40635 41123
rect 9229 41021 9263 41055
rect 9505 41021 9539 41055
rect 11621 41021 11655 41055
rect 12817 41021 12851 41055
rect 13001 41021 13035 41055
rect 14749 41021 14783 41055
rect 14933 41021 14967 41055
rect 17417 41021 17451 41055
rect 17509 41021 17543 41055
rect 17785 41021 17819 41055
rect 18429 41021 18463 41055
rect 19257 41021 19291 41055
rect 19441 41021 19475 41055
rect 21465 41021 21499 41055
rect 22477 41021 22511 41055
rect 23949 41021 23983 41055
rect 24225 41021 24259 41055
rect 24434 41021 24468 41055
rect 26525 41021 26559 41055
rect 29469 41021 29503 41055
rect 30665 41021 30699 41055
rect 31033 41021 31067 41055
rect 32413 41021 32447 41055
rect 40785 41021 40819 41055
rect 12173 40953 12207 40987
rect 12357 40953 12391 40987
rect 16221 40953 16255 40987
rect 22937 40953 22971 40987
rect 25605 40953 25639 40987
rect 27537 40953 27571 40987
rect 10977 40885 11011 40919
rect 15209 40885 15243 40919
rect 17233 40885 17267 40919
rect 22201 40885 22235 40919
rect 26341 40885 26375 40919
rect 26801 40885 26835 40919
rect 27813 40885 27847 40919
rect 28641 40885 28675 40919
rect 29285 40885 29319 40919
rect 29377 40885 29411 40919
rect 29837 40885 29871 40919
rect 30481 40885 30515 40919
rect 40417 40885 40451 40919
rect 9965 40681 9999 40715
rect 16405 40681 16439 40715
rect 17325 40681 17359 40715
rect 18061 40681 18095 40715
rect 20085 40681 20119 40715
rect 20545 40681 20579 40715
rect 22201 40681 22235 40715
rect 23121 40681 23155 40715
rect 24133 40681 24167 40715
rect 30297 40681 30331 40715
rect 23213 40613 23247 40647
rect 23765 40613 23799 40647
rect 11069 40545 11103 40579
rect 11345 40545 11379 40579
rect 12817 40545 12851 40579
rect 15393 40545 15427 40579
rect 15577 40545 15611 40579
rect 17049 40545 17083 40579
rect 21833 40545 21867 40579
rect 22937 40545 22971 40579
rect 23305 40545 23339 40579
rect 24409 40545 24443 40579
rect 24593 40545 24627 40579
rect 24777 40545 24811 40579
rect 24869 40545 24903 40579
rect 32781 40545 32815 40579
rect 37933 40545 37967 40579
rect 39405 40545 39439 40579
rect 39865 40545 39899 40579
rect 1409 40477 1443 40511
rect 1685 40477 1719 40511
rect 10149 40477 10183 40511
rect 10333 40477 10367 40511
rect 10425 40477 10459 40511
rect 13185 40477 13219 40511
rect 14105 40477 14139 40511
rect 14381 40477 14415 40511
rect 14565 40477 14599 40511
rect 14841 40477 14875 40511
rect 15945 40477 15979 40511
rect 16037 40477 16071 40511
rect 16589 40477 16623 40511
rect 16681 40477 16715 40511
rect 17233 40477 17267 40511
rect 17417 40477 17451 40511
rect 17601 40477 17635 40511
rect 17969 40477 18003 40511
rect 18245 40477 18279 40511
rect 18705 40477 18739 40511
rect 19533 40477 19567 40511
rect 19809 40477 19843 40511
rect 19993 40477 20027 40511
rect 20361 40477 20395 40511
rect 21557 40477 21591 40511
rect 22477 40477 22511 40511
rect 23029 40477 23063 40511
rect 23949 40477 23983 40511
rect 24225 40477 24259 40511
rect 24685 40477 24719 40511
rect 25145 40477 25179 40511
rect 25809 40477 25843 40511
rect 25973 40477 26007 40511
rect 26065 40477 26099 40511
rect 26157 40477 26191 40511
rect 26801 40477 26835 40511
rect 26949 40477 26983 40511
rect 27266 40477 27300 40511
rect 28457 40477 28491 40511
rect 28825 40477 28859 40511
rect 29561 40477 29595 40511
rect 29929 40477 29963 40511
rect 30297 40477 30331 40511
rect 30389 40477 30423 40511
rect 37657 40477 37691 40511
rect 16129 40409 16163 40443
rect 16773 40409 16807 40443
rect 16911 40409 16945 40443
rect 20913 40409 20947 40443
rect 22042 40409 22076 40443
rect 22569 40409 22603 40443
rect 22661 40409 22695 40443
rect 22799 40409 22833 40443
rect 27077 40409 27111 40443
rect 27169 40409 27203 40443
rect 28641 40409 28675 40443
rect 28733 40409 28767 40443
rect 29745 40409 29779 40443
rect 29837 40409 29871 40443
rect 32229 40409 32263 40443
rect 32413 40409 32447 40443
rect 33057 40409 33091 40443
rect 13737 40341 13771 40375
rect 14197 40341 14231 40375
rect 17785 40341 17819 40375
rect 18797 40341 18831 40375
rect 19349 40341 19383 40375
rect 19717 40341 19751 40375
rect 21005 40341 21039 40375
rect 21925 40341 21959 40375
rect 22293 40341 22327 40375
rect 25329 40341 25363 40375
rect 26341 40341 26375 40375
rect 27445 40341 27479 40375
rect 29009 40341 29043 40375
rect 30113 40341 30147 40375
rect 30665 40341 30699 40375
rect 32597 40341 32631 40375
rect 34529 40341 34563 40375
rect 40509 40341 40543 40375
rect 12909 40137 12943 40171
rect 13277 40137 13311 40171
rect 15669 40137 15703 40171
rect 16037 40137 16071 40171
rect 17233 40137 17267 40171
rect 17601 40137 17635 40171
rect 24317 40137 24351 40171
rect 27353 40137 27387 40171
rect 31493 40137 31527 40171
rect 32873 40137 32907 40171
rect 10057 40069 10091 40103
rect 10273 40069 10307 40103
rect 23949 40069 23983 40103
rect 24041 40069 24075 40103
rect 29101 40069 29135 40103
rect 31033 40069 31067 40103
rect 8493 40001 8527 40035
rect 9597 40001 9631 40035
rect 9689 40001 9723 40035
rect 13093 40001 13127 40035
rect 13369 40001 13403 40035
rect 14289 40001 14323 40035
rect 14381 40001 14415 40035
rect 14565 40001 14599 40035
rect 14657 40001 14691 40035
rect 15025 40001 15059 40035
rect 15117 40001 15151 40035
rect 17417 40001 17451 40035
rect 17693 40001 17727 40035
rect 19993 40001 20027 40035
rect 21833 40001 21867 40035
rect 23673 40001 23707 40035
rect 23766 40001 23800 40035
rect 24138 40001 24172 40035
rect 25789 40001 25823 40035
rect 25973 40001 26007 40035
rect 26065 40001 26099 40035
rect 26157 40001 26191 40035
rect 26985 40001 27019 40035
rect 29285 40001 29319 40035
rect 29377 40001 29411 40035
rect 31309 40001 31343 40035
rect 33057 40001 33091 40035
rect 9781 39933 9815 39967
rect 15393 39933 15427 39967
rect 15761 39933 15795 39967
rect 15853 39933 15887 39967
rect 27077 39933 27111 39967
rect 31217 39933 31251 39967
rect 10425 39865 10459 39899
rect 20085 39865 20119 39899
rect 22109 39865 22143 39899
rect 22293 39865 22327 39899
rect 8309 39797 8343 39831
rect 9229 39797 9263 39831
rect 10241 39797 10275 39831
rect 14105 39797 14139 39831
rect 15025 39797 15059 39831
rect 26341 39797 26375 39831
rect 26985 39797 27019 39831
rect 29285 39797 29319 39831
rect 29561 39797 29595 39831
rect 31033 39797 31067 39831
rect 9413 39593 9447 39627
rect 15117 39593 15151 39627
rect 17601 39593 17635 39627
rect 18613 39593 18647 39627
rect 25329 39593 25363 39627
rect 29561 39593 29595 39627
rect 30941 39593 30975 39627
rect 31769 39593 31803 39627
rect 32045 39593 32079 39627
rect 9229 39525 9263 39559
rect 16129 39525 16163 39559
rect 18981 39525 19015 39559
rect 31401 39525 31435 39559
rect 8953 39457 8987 39491
rect 11437 39457 11471 39491
rect 11529 39457 11563 39491
rect 14565 39457 14599 39491
rect 15485 39457 15519 39491
rect 19349 39457 19383 39491
rect 25421 39457 25455 39491
rect 29653 39457 29687 39491
rect 31033 39457 31067 39491
rect 32137 39457 32171 39491
rect 37933 39457 37967 39491
rect 38209 39457 38243 39491
rect 9689 39389 9723 39423
rect 15970 39389 16004 39423
rect 17785 39389 17819 39423
rect 17969 39389 18003 39423
rect 18245 39389 18279 39423
rect 18613 39389 18647 39423
rect 18797 39389 18831 39423
rect 19257 39389 19291 39423
rect 19533 39389 19567 39423
rect 19809 39389 19843 39423
rect 19901 39389 19935 39423
rect 25513 39389 25547 39423
rect 28181 39389 28215 39423
rect 28549 39389 28583 39423
rect 29561 39389 29595 39423
rect 31217 39389 31251 39423
rect 31585 39389 31619 39423
rect 31677 39389 31711 39423
rect 32321 39389 32355 39423
rect 33517 39389 33551 39423
rect 9965 39321 9999 39355
rect 17877 39321 17911 39355
rect 18087 39321 18121 39355
rect 19717 39321 19751 39355
rect 25237 39321 25271 39355
rect 28365 39321 28399 39355
rect 28457 39321 28491 39355
rect 30941 39321 30975 39355
rect 32045 39321 32079 39355
rect 12173 39253 12207 39287
rect 15761 39253 15795 39287
rect 15853 39253 15887 39287
rect 20085 39253 20119 39287
rect 25697 39253 25731 39287
rect 28733 39253 28767 39287
rect 29929 39253 29963 39287
rect 31953 39253 31987 39287
rect 32505 39253 32539 39287
rect 33333 39253 33367 39287
rect 39681 39253 39715 39287
rect 9413 39049 9447 39083
rect 10333 39049 10367 39083
rect 14473 39049 14507 39083
rect 20085 39049 20119 39083
rect 20269 39049 20303 39083
rect 21005 39049 21039 39083
rect 25881 39049 25915 39083
rect 26709 39049 26743 39083
rect 27629 39049 27663 39083
rect 29101 39049 29135 39083
rect 31493 39049 31527 39083
rect 32597 39049 32631 39083
rect 33057 39049 33091 39083
rect 7941 38981 7975 39015
rect 10057 38981 10091 39015
rect 13001 38981 13035 39015
rect 21373 38981 21407 39015
rect 21511 38981 21545 39015
rect 23397 38981 23431 39015
rect 24133 38981 24167 39015
rect 27261 38981 27295 39015
rect 27445 38981 27479 39015
rect 28641 38981 28675 39015
rect 29837 38981 29871 39015
rect 31033 38981 31067 39015
rect 9781 38913 9815 38947
rect 9965 38913 9999 38947
rect 10149 38913 10183 38947
rect 12725 38913 12759 38947
rect 17509 38913 17543 38947
rect 17785 38913 17819 38947
rect 18061 38913 18095 38947
rect 18245 38913 18279 38947
rect 18613 38913 18647 38947
rect 18797 38913 18831 38947
rect 18889 38913 18923 38947
rect 19717 38913 19751 38947
rect 19901 38913 19935 38947
rect 20453 38913 20487 38947
rect 20545 38913 20579 38947
rect 20637 38913 20671 38947
rect 20755 38913 20789 38947
rect 21189 38913 21223 38947
rect 21281 38913 21315 38947
rect 22753 38913 22787 38947
rect 22937 38913 22971 38947
rect 23305 38913 23339 38947
rect 23489 38913 23523 38947
rect 23627 38913 23661 38947
rect 23949 38913 23983 38947
rect 24225 38913 24259 38947
rect 24317 38913 24351 38947
rect 24593 38913 24627 38947
rect 24777 38913 24811 38947
rect 24869 38913 24903 38947
rect 24961 38913 24995 38947
rect 25237 38913 25271 38947
rect 25385 38913 25419 38947
rect 25513 38913 25547 38947
rect 25605 38913 25639 38947
rect 25743 38913 25777 38947
rect 26157 38913 26191 38947
rect 26341 38913 26375 38947
rect 26433 38913 26467 38947
rect 26525 38913 26559 38947
rect 27721 38913 27755 38947
rect 27905 38913 27939 38947
rect 27997 38913 28031 38947
rect 28089 38913 28123 38947
rect 28917 38913 28951 38947
rect 29211 38913 29245 38947
rect 29377 38913 29411 38947
rect 29653 38913 29687 38947
rect 30297 38913 30331 38947
rect 31349 38913 31383 38947
rect 31585 38913 31619 38947
rect 31769 38913 31803 38947
rect 32137 38913 32171 38947
rect 32413 38913 32447 38947
rect 32689 38913 32723 38947
rect 32781 38913 32815 38947
rect 33425 38913 33459 38947
rect 33609 38913 33643 38947
rect 7665 38845 7699 38879
rect 17969 38845 18003 38879
rect 20913 38845 20947 38879
rect 21649 38845 21683 38879
rect 22661 38845 22695 38879
rect 23765 38845 23799 38879
rect 28733 38845 28767 38879
rect 29561 38845 29595 38879
rect 30389 38845 30423 38879
rect 31125 38845 31159 38879
rect 32229 38845 32263 38879
rect 33885 38845 33919 38879
rect 25145 38777 25179 38811
rect 28273 38777 28307 38811
rect 30021 38777 30055 38811
rect 31953 38777 31987 38811
rect 33241 38777 33275 38811
rect 18429 38709 18463 38743
rect 18613 38709 18647 38743
rect 22201 38709 22235 38743
rect 22477 38709 22511 38743
rect 22569 38709 22603 38743
rect 23121 38709 23155 38743
rect 24501 38709 24535 38743
rect 28641 38709 28675 38743
rect 30297 38709 30331 38743
rect 30665 38709 30699 38743
rect 31033 38709 31067 38743
rect 31585 38709 31619 38743
rect 32137 38709 32171 38743
rect 32689 38709 32723 38743
rect 35357 38709 35391 38743
rect 17325 38505 17359 38539
rect 17969 38505 18003 38539
rect 18153 38505 18187 38539
rect 23489 38505 23523 38539
rect 25881 38505 25915 38539
rect 27077 38505 27111 38539
rect 29009 38505 29043 38539
rect 30665 38505 30699 38539
rect 31309 38505 31343 38539
rect 15393 38437 15427 38471
rect 21465 38437 21499 38471
rect 25605 38437 25639 38471
rect 26341 38437 26375 38471
rect 11529 38369 11563 38403
rect 15945 38369 15979 38403
rect 16037 38369 16071 38403
rect 20913 38369 20947 38403
rect 24409 38369 24443 38403
rect 25973 38369 26007 38403
rect 27077 38369 27111 38403
rect 30481 38369 30515 38403
rect 15577 38301 15611 38335
rect 15669 38301 15703 38335
rect 17233 38301 17267 38335
rect 17877 38301 17911 38335
rect 18153 38301 18187 38335
rect 18337 38301 18371 38335
rect 19993 38301 20027 38335
rect 21097 38301 21131 38335
rect 21373 38301 21407 38335
rect 21465 38301 21499 38335
rect 21649 38301 21683 38335
rect 23121 38301 23155 38335
rect 23305 38301 23339 38335
rect 24593 38301 24627 38335
rect 24777 38301 24811 38335
rect 25053 38301 25087 38335
rect 25421 38301 25455 38335
rect 26157 38301 26191 38335
rect 27261 38301 27295 38335
rect 30665 38301 30699 38335
rect 31125 38301 31159 38335
rect 11805 38233 11839 38267
rect 13553 38233 13587 38267
rect 16221 38233 16255 38267
rect 16405 38233 16439 38267
rect 21281 38233 21315 38267
rect 25237 38233 25271 38267
rect 25329 38233 25363 38267
rect 25881 38233 25915 38267
rect 26985 38233 27019 38267
rect 28641 38233 28675 38267
rect 28825 38233 28859 38267
rect 30389 38233 30423 38267
rect 30941 38233 30975 38267
rect 16497 38165 16531 38199
rect 16589 38165 16623 38199
rect 16773 38165 16807 38199
rect 20177 38165 20211 38199
rect 27445 38165 27479 38199
rect 30849 38165 30883 38199
rect 12909 37961 12943 37995
rect 17141 37961 17175 37995
rect 19457 37961 19491 37995
rect 19625 37961 19659 37995
rect 27629 37961 27663 37995
rect 28641 37961 28675 37995
rect 29653 37961 29687 37995
rect 31953 37961 31987 37995
rect 13395 37893 13429 37927
rect 16313 37893 16347 37927
rect 19257 37893 19291 37927
rect 20085 37893 20119 37927
rect 23397 37893 23431 37927
rect 28273 37893 28307 37927
rect 28361 37893 28395 37927
rect 29285 37893 29319 37927
rect 29377 37893 29411 37927
rect 33793 37893 33827 37927
rect 13093 37825 13127 37859
rect 13185 37825 13219 37859
rect 13277 37825 13311 37859
rect 15209 37825 15243 37859
rect 15577 37825 15611 37859
rect 15945 37825 15979 37859
rect 16129 37825 16163 37859
rect 16221 37825 16255 37859
rect 16405 37825 16439 37859
rect 16957 37825 16991 37859
rect 19901 37825 19935 37859
rect 19993 37825 20027 37859
rect 20223 37825 20257 37859
rect 23213 37825 23247 37859
rect 23305 37825 23339 37859
rect 23515 37825 23549 37859
rect 23673 37825 23707 37859
rect 26985 37825 27019 37859
rect 27078 37825 27112 37859
rect 27261 37825 27295 37859
rect 27353 37825 27387 37859
rect 27450 37825 27484 37859
rect 28089 37825 28123 37859
rect 28457 37825 28491 37859
rect 29009 37825 29043 37859
rect 29102 37825 29136 37859
rect 29515 37825 29549 37859
rect 31493 37825 31527 37859
rect 31769 37825 31803 37859
rect 32229 37825 32263 37859
rect 32321 37825 32355 37859
rect 33517 37825 33551 37859
rect 7297 37757 7331 37791
rect 7573 37757 7607 37791
rect 9597 37757 9631 37791
rect 9873 37757 9907 37791
rect 13553 37757 13587 37791
rect 15485 37757 15519 37791
rect 15853 37757 15887 37791
rect 16773 37757 16807 37791
rect 20361 37757 20395 37791
rect 31585 37757 31619 37791
rect 15025 37689 15059 37723
rect 15669 37689 15703 37723
rect 16037 37689 16071 37723
rect 19717 37689 19751 37723
rect 9045 37621 9079 37655
rect 11345 37621 11379 37655
rect 15393 37621 15427 37655
rect 15761 37621 15795 37655
rect 18889 37621 18923 37655
rect 19441 37621 19475 37655
rect 23029 37621 23063 37655
rect 31493 37621 31527 37655
rect 32229 37621 32263 37655
rect 32597 37621 32631 37655
rect 35265 37621 35299 37655
rect 8309 37417 8343 37451
rect 11529 37417 11563 37451
rect 18245 37417 18279 37451
rect 23029 37417 23063 37451
rect 23489 37417 23523 37451
rect 25973 37417 26007 37451
rect 30113 37417 30147 37451
rect 30297 37417 30331 37451
rect 31769 37417 31803 37451
rect 32137 37417 32171 37451
rect 12725 37349 12759 37383
rect 26801 37349 26835 37383
rect 8769 37281 8803 37315
rect 9597 37281 9631 37315
rect 10333 37281 10367 37315
rect 13645 37281 13679 37315
rect 16221 37281 16255 37315
rect 22845 37281 22879 37315
rect 30297 37281 30331 37315
rect 8493 37213 8527 37247
rect 8677 37213 8711 37247
rect 9045 37213 9079 37247
rect 10977 37213 11011 37247
rect 11345 37213 11379 37247
rect 12541 37213 12575 37247
rect 13001 37213 13035 37247
rect 15025 37213 15059 37247
rect 15209 37213 15243 37247
rect 15301 37213 15335 37247
rect 15761 37213 15795 37247
rect 16129 37213 16163 37247
rect 17417 37213 17451 37247
rect 17601 37213 17635 37247
rect 18521 37213 18555 37247
rect 18705 37213 18739 37247
rect 20453 37213 20487 37247
rect 20637 37213 20671 37247
rect 21925 37213 21959 37247
rect 22017 37213 22051 37247
rect 22385 37213 22419 37247
rect 22477 37213 22511 37247
rect 22569 37213 22603 37247
rect 23029 37213 23063 37247
rect 23213 37213 23247 37247
rect 23305 37213 23339 37247
rect 25421 37213 25455 37247
rect 25605 37213 25639 37247
rect 25697 37213 25731 37247
rect 25789 37213 25823 37247
rect 26249 37213 26283 37247
rect 26617 37213 26651 37247
rect 26893 37213 26927 37247
rect 26986 37213 27020 37247
rect 27399 37213 27433 37247
rect 29561 37213 29595 37247
rect 29929 37213 29963 37247
rect 30481 37213 30515 37247
rect 30849 37213 30883 37247
rect 30942 37213 30976 37247
rect 31314 37213 31348 37247
rect 32321 37213 32355 37247
rect 32413 37213 32447 37247
rect 33609 37213 33643 37247
rect 40785 37213 40819 37247
rect 11161 37145 11195 37179
rect 11253 37145 11287 37179
rect 13553 37145 13587 37179
rect 15117 37145 15151 37179
rect 17785 37145 17819 37179
rect 18061 37145 18095 37179
rect 18277 37145 18311 37179
rect 22707 37145 22741 37179
rect 26433 37145 26467 37179
rect 26525 37145 26559 37179
rect 27169 37145 27203 37179
rect 27261 37145 27295 37179
rect 29745 37145 29779 37179
rect 29837 37145 29871 37179
rect 30205 37145 30239 37179
rect 31125 37145 31159 37179
rect 31217 37145 31251 37179
rect 31677 37145 31711 37179
rect 32137 37145 32171 37179
rect 10885 37077 10919 37111
rect 12909 37077 12943 37111
rect 13093 37077 13127 37111
rect 13461 37077 13495 37111
rect 18429 37077 18463 37111
rect 18613 37077 18647 37111
rect 20545 37077 20579 37111
rect 22201 37077 22235 37111
rect 27537 37077 27571 37111
rect 30665 37077 30699 37111
rect 31493 37077 31527 37111
rect 32597 37077 32631 37111
rect 33425 37077 33459 37111
rect 40969 37077 41003 37111
rect 12081 36873 12115 36907
rect 16221 36873 16255 36907
rect 17877 36873 17911 36907
rect 19165 36873 19199 36907
rect 31953 36873 31987 36907
rect 32505 36873 32539 36907
rect 12541 36805 12575 36839
rect 14289 36805 14323 36839
rect 15761 36805 15795 36839
rect 21557 36805 21591 36839
rect 23857 36805 23891 36839
rect 23949 36805 23983 36839
rect 24087 36805 24121 36839
rect 25697 36805 25731 36839
rect 27905 36805 27939 36839
rect 31217 36805 31251 36839
rect 34069 36805 34103 36839
rect 8033 36737 8067 36771
rect 9873 36737 9907 36771
rect 10609 36737 10643 36771
rect 10793 36737 10827 36771
rect 10885 36737 10919 36771
rect 10977 36737 11011 36771
rect 11529 36737 11563 36771
rect 11713 36737 11747 36771
rect 11805 36737 11839 36771
rect 11897 36737 11931 36771
rect 15393 36737 15427 36771
rect 15577 36737 15611 36771
rect 16129 36737 16163 36771
rect 16681 36737 16715 36771
rect 16865 36737 16899 36771
rect 17141 36737 17175 36771
rect 17601 36737 17635 36771
rect 18064 36759 18098 36793
rect 18153 36737 18187 36771
rect 18337 36737 18371 36771
rect 18429 36737 18463 36771
rect 18521 36737 18555 36771
rect 19073 36737 19107 36771
rect 20177 36737 20211 36771
rect 20361 36737 20395 36771
rect 21465 36737 21499 36771
rect 21649 36737 21683 36771
rect 22293 36737 22327 36771
rect 22753 36737 22787 36771
rect 22845 36737 22879 36771
rect 22937 36737 22971 36771
rect 23765 36737 23799 36771
rect 24501 36737 24535 36771
rect 25421 36737 25455 36771
rect 25514 36737 25548 36771
rect 25789 36737 25823 36771
rect 25886 36737 25920 36771
rect 28181 36737 28215 36771
rect 28825 36737 28859 36771
rect 31033 36737 31067 36771
rect 31493 36737 31527 36771
rect 31769 36737 31803 36771
rect 32137 36737 32171 36771
rect 32229 36737 32263 36771
rect 33241 36737 33275 36771
rect 33793 36737 33827 36771
rect 8309 36669 8343 36703
rect 12265 36669 12299 36703
rect 17693 36669 17727 36703
rect 19257 36669 19291 36703
rect 19533 36669 19567 36703
rect 19901 36669 19935 36703
rect 20085 36669 20119 36703
rect 20269 36669 20303 36703
rect 20637 36669 20671 36703
rect 21005 36669 21039 36703
rect 21097 36669 21131 36703
rect 21925 36669 21959 36703
rect 22109 36669 22143 36703
rect 22201 36669 22235 36703
rect 22385 36669 22419 36703
rect 23029 36669 23063 36703
rect 24225 36669 24259 36703
rect 24317 36669 24351 36703
rect 27997 36669 28031 36703
rect 28917 36669 28951 36703
rect 31585 36669 31619 36703
rect 10057 36601 10091 36635
rect 18981 36601 19015 36635
rect 21281 36601 21315 36635
rect 24685 36601 24719 36635
rect 26065 36601 26099 36635
rect 31401 36601 31435 36635
rect 9781 36533 9815 36567
rect 11161 36533 11195 36567
rect 16681 36533 16715 36567
rect 17417 36533 17451 36567
rect 18705 36533 18739 36567
rect 19441 36533 19475 36567
rect 22569 36533 22603 36567
rect 23581 36533 23615 36567
rect 28181 36533 28215 36567
rect 28365 36533 28399 36567
rect 28825 36533 28859 36567
rect 29193 36533 29227 36567
rect 31493 36533 31527 36567
rect 32137 36533 32171 36567
rect 33057 36533 33091 36567
rect 35541 36533 35575 36567
rect 6732 36329 6766 36363
rect 16313 36329 16347 36363
rect 16497 36329 16531 36363
rect 19441 36329 19475 36363
rect 20177 36329 20211 36363
rect 20637 36329 20671 36363
rect 24869 36329 24903 36363
rect 28089 36329 28123 36363
rect 31217 36329 31251 36363
rect 19993 36261 20027 36295
rect 27169 36261 27203 36295
rect 11437 36193 11471 36227
rect 17969 36193 18003 36227
rect 20269 36193 20303 36227
rect 21097 36193 21131 36227
rect 28273 36193 28307 36227
rect 29009 36193 29043 36227
rect 31401 36193 31435 36227
rect 34253 36193 34287 36227
rect 6469 36125 6503 36159
rect 11713 36125 11747 36159
rect 19809 36125 19843 36159
rect 20453 36125 20487 36159
rect 20913 36125 20947 36159
rect 22293 36125 22327 36159
rect 22477 36125 22511 36159
rect 22661 36125 22695 36159
rect 22753 36125 22787 36159
rect 23581 36125 23615 36159
rect 23674 36125 23708 36159
rect 23949 36125 23983 36159
rect 24087 36125 24121 36159
rect 25053 36125 25087 36159
rect 25375 36125 25409 36159
rect 25513 36125 25547 36159
rect 25973 36125 26007 36159
rect 26121 36125 26155 36159
rect 26479 36125 26513 36159
rect 27353 36125 27387 36159
rect 27445 36125 27479 36159
rect 27629 36125 27663 36159
rect 27721 36125 27755 36159
rect 28089 36125 28123 36159
rect 28365 36125 28399 36159
rect 28641 36125 28675 36159
rect 31493 36125 31527 36159
rect 1501 36057 1535 36091
rect 9045 36057 9079 36091
rect 10701 36057 10735 36091
rect 11989 36057 12023 36091
rect 16129 36057 16163 36091
rect 17693 36057 17727 36091
rect 19257 36057 19291 36091
rect 20177 36057 20211 36091
rect 20729 36057 20763 36091
rect 23857 36057 23891 36091
rect 25145 36057 25179 36091
rect 25237 36057 25271 36091
rect 26249 36057 26283 36091
rect 26341 36057 26375 36091
rect 28825 36057 28859 36091
rect 31217 36057 31251 36091
rect 33517 36057 33551 36091
rect 1593 35989 1627 36023
rect 8217 35989 8251 36023
rect 9137 35989 9171 36023
rect 16329 35989 16363 36023
rect 19441 35989 19475 36023
rect 19625 35989 19659 36023
rect 24225 35989 24259 36023
rect 26617 35989 26651 36023
rect 28549 35989 28583 36023
rect 31677 35989 31711 36023
rect 9045 35785 9079 35819
rect 10977 35785 11011 35819
rect 13093 35785 13127 35819
rect 23029 35785 23063 35819
rect 24317 35785 24351 35819
rect 25881 35785 25915 35819
rect 27721 35785 27755 35819
rect 30297 35785 30331 35819
rect 9321 35717 9355 35751
rect 9678 35717 9712 35751
rect 23489 35717 23523 35751
rect 24593 35717 24627 35751
rect 8953 35649 8987 35683
rect 9505 35649 9539 35683
rect 10241 35649 10275 35683
rect 10701 35649 10735 35683
rect 10793 35649 10827 35683
rect 11989 35649 12023 35683
rect 12827 35671 12861 35705
rect 19717 35649 19751 35683
rect 22661 35649 22695 35683
rect 23121 35649 23155 35683
rect 23213 35649 23247 35683
rect 23306 35649 23340 35683
rect 23581 35649 23615 35683
rect 23719 35649 23753 35683
rect 24501 35649 24535 35683
rect 24685 35649 24719 35683
rect 24803 35649 24837 35683
rect 24961 35649 24995 35683
rect 26065 35649 26099 35683
rect 26203 35649 26237 35683
rect 26341 35649 26375 35683
rect 26433 35649 26467 35683
rect 27077 35649 27111 35683
rect 27170 35649 27204 35683
rect 27353 35649 27387 35683
rect 27445 35649 27479 35683
rect 27542 35649 27576 35683
rect 27813 35649 27847 35683
rect 27997 35649 28031 35683
rect 28089 35649 28123 35683
rect 28181 35649 28215 35683
rect 29469 35649 29503 35683
rect 29617 35649 29651 35683
rect 29745 35649 29779 35683
rect 29837 35649 29871 35683
rect 29975 35649 30009 35683
rect 30757 35649 30791 35683
rect 30849 35649 30883 35683
rect 31033 35649 31067 35683
rect 32505 35649 32539 35683
rect 33333 35649 33367 35683
rect 6377 35581 6411 35615
rect 6745 35581 6779 35615
rect 9137 35581 9171 35615
rect 11805 35581 11839 35615
rect 13093 35581 13127 35615
rect 19993 35581 20027 35615
rect 22385 35581 22419 35615
rect 22845 35581 22879 35615
rect 30665 35581 30699 35615
rect 33609 35581 33643 35615
rect 8171 35513 8205 35547
rect 12909 35513 12943 35547
rect 19533 35513 19567 35547
rect 28365 35513 28399 35547
rect 30113 35513 30147 35547
rect 35081 35513 35115 35547
rect 9229 35445 9263 35479
rect 9873 35445 9907 35479
rect 10057 35445 10091 35479
rect 12173 35445 12207 35479
rect 19901 35445 19935 35479
rect 22753 35445 22787 35479
rect 23857 35445 23891 35479
rect 30573 35445 30607 35479
rect 32321 35445 32355 35479
rect 6745 35241 6779 35275
rect 10057 35241 10091 35275
rect 10425 35241 10459 35275
rect 22477 35241 22511 35275
rect 25145 35241 25179 35275
rect 27445 35241 27479 35275
rect 28641 35241 28675 35275
rect 32670 35241 32704 35275
rect 9689 35173 9723 35207
rect 10885 35173 10919 35207
rect 15945 35173 15979 35207
rect 30113 35173 30147 35207
rect 31033 35173 31067 35207
rect 8033 35105 8067 35139
rect 9965 35105 9999 35139
rect 10517 35105 10551 35139
rect 22385 35105 22419 35139
rect 27813 35105 27847 35139
rect 27905 35105 27939 35139
rect 32413 35105 32447 35139
rect 6929 35037 6963 35071
rect 7757 35037 7791 35071
rect 8401 35037 8435 35071
rect 8677 35037 8711 35071
rect 9873 35037 9907 35071
rect 10425 35037 10459 35071
rect 10701 35037 10735 35071
rect 11253 35037 11287 35071
rect 11345 35037 11379 35071
rect 11529 35037 11563 35071
rect 11621 35037 11655 35071
rect 11897 35037 11931 35071
rect 11989 35037 12023 35071
rect 12173 35037 12207 35071
rect 12265 35037 12299 35071
rect 12633 35037 12667 35071
rect 14105 35037 14139 35071
rect 14749 35037 14783 35071
rect 14933 35037 14967 35071
rect 15025 35037 15059 35071
rect 15117 35037 15151 35071
rect 15301 35037 15335 35071
rect 15393 35037 15427 35071
rect 15813 35037 15847 35071
rect 16129 35037 16163 35071
rect 16277 35037 16311 35071
rect 16497 35037 16531 35071
rect 16635 35037 16669 35071
rect 22293 35037 22327 35071
rect 24593 35037 24627 35071
rect 24961 35037 24995 35071
rect 25237 35037 25271 35071
rect 25421 35037 25455 35071
rect 25605 35037 25639 35071
rect 27629 35037 27663 35071
rect 27721 35037 27755 35071
rect 28825 35037 28859 35071
rect 29009 35037 29043 35071
rect 29285 35037 29319 35071
rect 29561 35037 29595 35071
rect 29745 35037 29779 35071
rect 29929 35037 29963 35071
rect 30396 35037 30430 35071
rect 30537 35037 30571 35071
rect 30854 35037 30888 35071
rect 31217 35037 31251 35071
rect 31310 35037 31344 35071
rect 31682 35037 31716 35071
rect 31953 35037 31987 35071
rect 32137 35037 32171 35071
rect 34805 35037 34839 35071
rect 8585 34969 8619 35003
rect 9413 34969 9447 35003
rect 11713 34969 11747 35003
rect 12909 34969 12943 35003
rect 13461 34969 13495 35003
rect 13645 34969 13679 35003
rect 14197 34969 14231 35003
rect 15209 34969 15243 35003
rect 15577 34969 15611 35003
rect 15669 34969 15703 35003
rect 16405 34969 16439 35003
rect 22569 34969 22603 35003
rect 24777 34969 24811 35003
rect 24869 34969 24903 35003
rect 25513 34969 25547 35003
rect 28917 34969 28951 35003
rect 29147 34969 29181 35003
rect 29837 34969 29871 35003
rect 30665 34969 30699 35003
rect 30757 34969 30791 35003
rect 31493 34969 31527 35003
rect 31582 34969 31616 35003
rect 7389 34901 7423 34935
rect 7849 34901 7883 34935
rect 8217 34901 8251 34935
rect 10241 34901 10275 34935
rect 11069 34901 11103 34935
rect 13829 34901 13863 34935
rect 14565 34901 14599 34935
rect 16773 34901 16807 34935
rect 25789 34901 25823 34935
rect 31861 34901 31895 34935
rect 32045 34901 32079 34935
rect 34161 34901 34195 34935
rect 34897 34901 34931 34935
rect 10241 34697 10275 34731
rect 13093 34697 13127 34731
rect 14473 34697 14507 34731
rect 18889 34697 18923 34731
rect 21465 34697 21499 34731
rect 22201 34697 22235 34731
rect 26065 34697 26099 34731
rect 27997 34697 28031 34731
rect 29837 34697 29871 34731
rect 30573 34697 30607 34731
rect 30849 34697 30883 34731
rect 35081 34697 35115 34731
rect 6653 34629 6687 34663
rect 9321 34629 9355 34663
rect 9873 34629 9907 34663
rect 14105 34629 14139 34663
rect 21005 34629 21039 34663
rect 22477 34629 22511 34663
rect 27629 34629 27663 34663
rect 29561 34629 29595 34663
rect 30205 34629 30239 34663
rect 32229 34629 32263 34663
rect 9505 34561 9539 34595
rect 9597 34561 9631 34595
rect 10057 34561 10091 34595
rect 12633 34561 12667 34595
rect 13369 34561 13403 34595
rect 13461 34561 13495 34595
rect 13553 34561 13587 34595
rect 13737 34561 13771 34595
rect 13829 34561 13863 34595
rect 13977 34561 14011 34595
rect 14197 34561 14231 34595
rect 14294 34561 14328 34595
rect 14565 34561 14599 34595
rect 14749 34561 14783 34595
rect 16957 34561 16991 34595
rect 17233 34561 17267 34595
rect 17417 34561 17451 34595
rect 17509 34561 17543 34595
rect 17602 34561 17636 34595
rect 17785 34561 17819 34595
rect 17877 34561 17911 34595
rect 18015 34561 18049 34595
rect 18337 34561 18371 34595
rect 18521 34561 18555 34595
rect 18613 34561 18647 34595
rect 18705 34561 18739 34595
rect 19165 34561 19199 34595
rect 21281 34561 21315 34595
rect 22201 34561 22235 34595
rect 25973 34561 26007 34595
rect 26157 34561 26191 34595
rect 27445 34561 27479 34595
rect 27721 34561 27755 34595
rect 27813 34561 27847 34595
rect 29285 34561 29319 34595
rect 29469 34561 29503 34595
rect 29653 34561 29687 34595
rect 30021 34561 30055 34595
rect 30297 34561 30331 34595
rect 30389 34561 30423 34595
rect 30665 34561 30699 34595
rect 31493 34561 31527 34595
rect 31677 34561 31711 34595
rect 31769 34561 31803 34595
rect 32137 34561 32171 34595
rect 33885 34561 33919 34595
rect 34437 34561 34471 34595
rect 34713 34561 34747 34595
rect 34897 34561 34931 34595
rect 35173 34561 35207 34595
rect 35541 34561 35575 34595
rect 35633 34561 35667 34595
rect 7389 34493 7423 34527
rect 17049 34493 17083 34527
rect 19441 34493 19475 34527
rect 21189 34493 21223 34527
rect 31309 34493 31343 34527
rect 34069 34493 34103 34527
rect 18153 34425 18187 34459
rect 19349 34425 19383 34459
rect 22293 34425 22327 34459
rect 31585 34425 31619 34459
rect 35817 34425 35851 34459
rect 9321 34357 9355 34391
rect 9781 34357 9815 34391
rect 12725 34357 12759 34391
rect 14565 34357 14599 34391
rect 14933 34357 14967 34391
rect 16681 34357 16715 34391
rect 17141 34357 17175 34391
rect 18981 34357 19015 34391
rect 21281 34357 21315 34391
rect 34529 34357 34563 34391
rect 35357 34357 35391 34391
rect 17049 34153 17083 34187
rect 20821 34153 20855 34187
rect 21741 34153 21775 34187
rect 22937 34153 22971 34187
rect 25329 34153 25363 34187
rect 31769 34153 31803 34187
rect 34253 34153 34287 34187
rect 35173 34153 35207 34187
rect 7941 34085 7975 34119
rect 11161 34085 11195 34119
rect 13553 34085 13587 34119
rect 11713 34017 11747 34051
rect 11805 34017 11839 34051
rect 21281 34017 21315 34051
rect 33701 34017 33735 34051
rect 35081 34017 35115 34051
rect 9413 33949 9447 33983
rect 9561 33949 9595 33983
rect 9781 33949 9815 33983
rect 9878 33949 9912 33983
rect 11342 33949 11376 33983
rect 12725 33949 12759 33983
rect 15301 33949 15335 33983
rect 16865 33949 16899 33983
rect 17601 33949 17635 33983
rect 18429 33949 18463 33983
rect 18521 33949 18555 33983
rect 18705 33949 18739 33983
rect 18797 33949 18831 33983
rect 19257 33949 19291 33983
rect 19533 33949 19567 33983
rect 19625 33949 19659 33983
rect 20085 33949 20119 33983
rect 20178 33949 20212 33983
rect 20591 33949 20625 33983
rect 21005 33949 21039 33983
rect 21189 33949 21223 33983
rect 21741 33949 21775 33983
rect 21925 33949 21959 33983
rect 22937 33949 22971 33983
rect 23121 33949 23155 33983
rect 24961 33949 24995 33983
rect 25145 33949 25179 33983
rect 25421 33949 25455 33983
rect 25605 33949 25639 33983
rect 31769 33949 31803 33983
rect 31953 33949 31987 33983
rect 33517 33949 33551 33983
rect 34713 33949 34747 33983
rect 35173 33949 35207 33983
rect 7573 33881 7607 33915
rect 9689 33881 9723 33915
rect 11989 33881 12023 33915
rect 13277 33881 13311 33915
rect 14105 33881 14139 33915
rect 14289 33881 14323 33915
rect 15577 33881 15611 33915
rect 16681 33881 16715 33915
rect 18245 33881 18279 33915
rect 19441 33881 19475 33915
rect 20361 33881 20395 33915
rect 20453 33881 20487 33915
rect 34161 33881 34195 33915
rect 8033 33813 8067 33847
rect 10057 33813 10091 33847
rect 11345 33813 11379 33847
rect 12081 33813 12115 33847
rect 12817 33813 12851 33847
rect 14473 33813 14507 33847
rect 17693 33813 17727 33847
rect 19809 33813 19843 33847
rect 20729 33813 20763 33847
rect 25513 33813 25547 33847
rect 35357 33813 35391 33847
rect 9597 33609 9631 33643
rect 13461 33609 13495 33643
rect 18889 33609 18923 33643
rect 23489 33609 23523 33643
rect 23949 33609 23983 33643
rect 26709 33609 26743 33643
rect 27077 33609 27111 33643
rect 28181 33609 28215 33643
rect 29377 33609 29411 33643
rect 34713 33609 34747 33643
rect 8769 33541 8803 33575
rect 10149 33541 10183 33575
rect 13185 33541 13219 33575
rect 15945 33541 15979 33575
rect 21925 33541 21959 33575
rect 23029 33541 23063 33575
rect 24317 33541 24351 33575
rect 26249 33541 26283 33575
rect 35173 33541 35207 33575
rect 8217 33473 8251 33507
rect 9459 33473 9493 33507
rect 9689 33473 9723 33507
rect 9965 33473 9999 33507
rect 11529 33473 11563 33507
rect 11621 33473 11655 33507
rect 12633 33473 12667 33507
rect 14013 33473 14047 33507
rect 15485 33473 15519 33507
rect 15669 33473 15703 33507
rect 16221 33473 16255 33507
rect 18705 33473 18739 33507
rect 18981 33473 19015 33507
rect 20637 33473 20671 33507
rect 20913 33473 20947 33507
rect 21833 33473 21867 33507
rect 22017 33473 22051 33507
rect 22201 33473 22235 33507
rect 22385 33473 22419 33507
rect 22569 33473 22603 33507
rect 22845 33473 22879 33507
rect 23581 33473 23615 33507
rect 23765 33473 23799 33507
rect 23857 33473 23891 33507
rect 24041 33473 24075 33507
rect 24225 33473 24259 33507
rect 24409 33473 24443 33507
rect 24501 33479 24535 33513
rect 24961 33473 24995 33507
rect 25145 33473 25179 33507
rect 25329 33473 25363 33507
rect 25605 33473 25639 33507
rect 25881 33473 25915 33507
rect 26065 33473 26099 33507
rect 26617 33473 26651 33507
rect 26801 33473 26835 33507
rect 27077 33473 27111 33507
rect 27169 33473 27203 33507
rect 27445 33473 27479 33507
rect 27629 33473 27663 33507
rect 28089 33473 28123 33507
rect 28273 33473 28307 33507
rect 28917 33473 28951 33507
rect 29233 33473 29267 33507
rect 29549 33473 29583 33507
rect 29745 33473 29779 33507
rect 31401 33473 31435 33507
rect 34621 33473 34655 33507
rect 35449 33473 35483 33507
rect 6377 33405 6411 33439
rect 6745 33405 6779 33439
rect 9045 33405 9079 33439
rect 9781 33405 9815 33439
rect 11805 33405 11839 33439
rect 12725 33405 12759 33439
rect 14105 33405 14139 33439
rect 16129 33405 16163 33439
rect 18245 33405 18279 33439
rect 20821 33405 20855 33439
rect 24593 33405 24627 33439
rect 25513 33405 25547 33439
rect 29009 33405 29043 33439
rect 31585 33405 31619 33439
rect 13001 33337 13035 33371
rect 22385 33337 22419 33371
rect 22845 33337 22879 33371
rect 23305 33337 23339 33371
rect 23581 33337 23615 33371
rect 9229 33269 9263 33303
rect 11713 33269 11747 33303
rect 12633 33269 12667 33303
rect 14013 33269 14047 33303
rect 14381 33269 14415 33303
rect 15853 33269 15887 33303
rect 16221 33269 16255 33303
rect 16405 33269 16439 33303
rect 18521 33269 18555 33303
rect 18613 33269 18647 33303
rect 20821 33269 20855 33303
rect 21097 33269 21131 33303
rect 24501 33269 24535 33303
rect 24869 33269 24903 33303
rect 24961 33269 24995 33303
rect 25605 33269 25639 33303
rect 25789 33269 25823 33303
rect 27445 33269 27479 33303
rect 29193 33269 29227 33303
rect 29561 33269 29595 33303
rect 35265 33269 35299 33303
rect 35633 33269 35667 33303
rect 5549 33065 5583 33099
rect 8125 33065 8159 33099
rect 13645 33065 13679 33099
rect 18613 33065 18647 33099
rect 21557 33065 21591 33099
rect 27629 33065 27663 33099
rect 35265 33065 35299 33099
rect 6837 32997 6871 33031
rect 13185 32997 13219 33031
rect 24685 32997 24719 33031
rect 31309 32997 31343 33031
rect 35449 32997 35483 33031
rect 6009 32929 6043 32963
rect 8677 32929 8711 32963
rect 13277 32929 13311 32963
rect 27261 32929 27295 32963
rect 27997 32929 28031 32963
rect 28549 32929 28583 32963
rect 30481 32929 30515 32963
rect 34069 32929 34103 32963
rect 34805 32929 34839 32963
rect 5733 32861 5767 32895
rect 5825 32861 5859 32895
rect 6101 32861 6135 32895
rect 6285 32861 6319 32895
rect 8401 32861 8435 32895
rect 11437 32861 11471 32895
rect 13461 32861 13495 32895
rect 13737 32861 13771 32895
rect 14105 32861 14139 32895
rect 14253 32861 14287 32895
rect 14381 32861 14415 32895
rect 14570 32861 14604 32895
rect 16037 32861 16071 32895
rect 16129 32861 16163 32895
rect 16313 32861 16347 32895
rect 16405 32861 16439 32895
rect 18061 32861 18095 32895
rect 18245 32861 18279 32895
rect 18337 32861 18371 32895
rect 18429 32861 18463 32895
rect 21373 32861 21407 32895
rect 21465 32861 21499 32895
rect 24409 32861 24443 32895
rect 24685 32861 24719 32895
rect 25237 32861 25271 32895
rect 25329 32861 25363 32895
rect 25421 32861 25455 32895
rect 27445 32861 27479 32895
rect 27721 32861 27755 32895
rect 27813 32861 27847 32895
rect 28365 32861 28399 32895
rect 30021 32861 30055 32895
rect 30205 32861 30239 32895
rect 30757 32861 30791 32895
rect 31033 32861 31067 32895
rect 31677 32861 31711 32895
rect 32045 32861 32079 32895
rect 33885 32861 33919 32895
rect 34897 32861 34931 32895
rect 35265 32861 35299 32895
rect 35541 32861 35575 32895
rect 40785 32861 40819 32895
rect 7849 32793 7883 32827
rect 12817 32793 12851 32827
rect 13001 32793 13035 32827
rect 14473 32793 14507 32827
rect 30573 32793 30607 32827
rect 30941 32793 30975 32827
rect 32321 32793 32355 32827
rect 32873 32793 32907 32827
rect 33609 32793 33643 32827
rect 11713 32725 11747 32759
rect 14749 32725 14783 32759
rect 15853 32725 15887 32759
rect 21741 32725 21775 32759
rect 35725 32725 35759 32759
rect 40969 32725 41003 32759
rect 6101 32521 6135 32555
rect 6469 32521 6503 32555
rect 9045 32521 9079 32555
rect 14381 32521 14415 32555
rect 15853 32521 15887 32555
rect 17325 32521 17359 32555
rect 18521 32521 18555 32555
rect 20177 32521 20211 32555
rect 27353 32521 27387 32555
rect 28917 32521 28951 32555
rect 30205 32521 30239 32555
rect 33977 32521 34011 32555
rect 34805 32521 34839 32555
rect 1501 32453 1535 32487
rect 10517 32453 10551 32487
rect 13277 32453 13311 32487
rect 13645 32453 13679 32487
rect 14013 32453 14047 32487
rect 14749 32453 14783 32487
rect 16681 32453 16715 32487
rect 18153 32453 18187 32487
rect 19165 32453 19199 32487
rect 24317 32453 24351 32487
rect 37381 32453 37415 32487
rect 38117 32453 38151 32487
rect 6377 32385 6411 32419
rect 7757 32385 7791 32419
rect 7941 32385 7975 32419
rect 8125 32385 8159 32419
rect 8309 32385 8343 32419
rect 8585 32385 8619 32419
rect 8769 32385 8803 32419
rect 9137 32385 9171 32419
rect 9321 32385 9355 32419
rect 9597 32385 9631 32419
rect 10701 32385 10735 32419
rect 10793 32385 10827 32419
rect 10977 32385 11011 32419
rect 11069 32385 11103 32419
rect 11713 32385 11747 32419
rect 11897 32385 11931 32419
rect 11989 32385 12023 32419
rect 12541 32385 12575 32419
rect 12633 32385 12667 32419
rect 12725 32385 12759 32419
rect 12909 32385 12943 32419
rect 13461 32385 13495 32419
rect 13737 32385 13771 32419
rect 13830 32385 13864 32419
rect 14105 32385 14139 32419
rect 14202 32385 14236 32419
rect 15025 32385 15059 32419
rect 15301 32385 15335 32419
rect 15485 32385 15519 32419
rect 15577 32385 15611 32419
rect 15669 32385 15703 32419
rect 16129 32385 16163 32419
rect 16221 32385 16255 32419
rect 16405 32385 16439 32419
rect 16497 32385 16531 32419
rect 16957 32385 16991 32419
rect 17417 32385 17451 32419
rect 17693 32385 17727 32419
rect 17877 32385 17911 32419
rect 17969 32385 18003 32419
rect 18245 32385 18279 32419
rect 18337 32385 18371 32419
rect 19349 32385 19383 32419
rect 19717 32385 19751 32419
rect 19993 32385 20027 32419
rect 20453 32385 20487 32419
rect 21833 32385 21867 32419
rect 22109 32385 22143 32419
rect 24041 32385 24075 32419
rect 27169 32385 27203 32419
rect 27353 32385 27387 32419
rect 27537 32385 27571 32419
rect 27721 32385 27755 32419
rect 28813 32385 28847 32419
rect 29009 32385 29043 32419
rect 30113 32385 30147 32419
rect 30297 32385 30331 32419
rect 31033 32385 31067 32419
rect 31677 32385 31711 32419
rect 32689 32385 32723 32419
rect 33425 32385 33459 32419
rect 33793 32385 33827 32419
rect 34253 32385 34287 32419
rect 34621 32385 34655 32419
rect 34989 32385 35023 32419
rect 35081 32385 35115 32419
rect 35449 32385 35483 32419
rect 4353 32317 4387 32351
rect 4629 32317 4663 32351
rect 7849 32317 7883 32351
rect 9045 32317 9079 32351
rect 14841 32317 14875 32351
rect 17049 32317 17083 32351
rect 17509 32317 17543 32351
rect 19625 32317 19659 32351
rect 19809 32317 19843 32351
rect 20269 32317 20303 32351
rect 22017 32317 22051 32351
rect 23857 32317 23891 32351
rect 24409 32317 24443 32351
rect 30389 32317 30423 32351
rect 32873 32317 32907 32351
rect 33333 32317 33367 32351
rect 34161 32317 34195 32351
rect 9413 32249 9447 32283
rect 9505 32249 9539 32283
rect 20637 32249 20671 32283
rect 30665 32249 30699 32283
rect 31309 32249 31343 32283
rect 1593 32181 1627 32215
rect 11529 32181 11563 32215
rect 12265 32181 12299 32215
rect 15025 32181 15059 32215
rect 15209 32181 15243 32215
rect 15945 32181 15979 32215
rect 17141 32181 17175 32215
rect 19533 32181 19567 32215
rect 19993 32181 20027 32215
rect 21925 32181 21959 32215
rect 22293 32181 22327 32215
rect 27537 32181 27571 32215
rect 30849 32181 30883 32215
rect 33793 32181 33827 32215
rect 34621 32181 34655 32215
rect 35449 32181 35483 32215
rect 35633 32181 35667 32215
rect 6193 31977 6227 32011
rect 7941 31977 7975 32011
rect 9045 31977 9079 32011
rect 10609 31977 10643 32011
rect 15945 31977 15979 32011
rect 16681 31977 16715 32011
rect 18429 31977 18463 32011
rect 20821 31977 20855 32011
rect 21189 31977 21223 32011
rect 21281 31977 21315 32011
rect 21649 31977 21683 32011
rect 22201 31977 22235 32011
rect 27813 31977 27847 32011
rect 31861 31977 31895 32011
rect 33793 31977 33827 32011
rect 10793 31909 10827 31943
rect 13829 31909 13863 31943
rect 17049 31909 17083 31943
rect 22109 31909 22143 31943
rect 25973 31909 26007 31943
rect 26341 31909 26375 31943
rect 28181 31909 28215 31943
rect 33977 31909 34011 31943
rect 8585 31841 8619 31875
rect 9689 31841 9723 31875
rect 10333 31841 10367 31875
rect 13461 31841 13495 31875
rect 13921 31841 13955 31875
rect 15853 31841 15887 31875
rect 21741 31841 21775 31875
rect 27905 31841 27939 31875
rect 30573 31841 30607 31875
rect 33701 31841 33735 31875
rect 34897 31841 34931 31875
rect 5641 31773 5675 31807
rect 5917 31773 5951 31807
rect 6009 31773 6043 31807
rect 8125 31773 8159 31807
rect 8217 31773 8251 31807
rect 8309 31773 8343 31807
rect 9229 31773 9263 31807
rect 9321 31773 9355 31807
rect 9490 31773 9524 31807
rect 9607 31751 9641 31785
rect 9873 31773 9907 31807
rect 10195 31773 10229 31807
rect 12449 31773 12483 31807
rect 12542 31773 12576 31807
rect 12725 31773 12759 31807
rect 12817 31773 12851 31807
rect 12914 31773 12948 31807
rect 13645 31773 13679 31807
rect 15669 31773 15703 31807
rect 15945 31773 15979 31807
rect 16865 31773 16899 31807
rect 17141 31773 17175 31807
rect 17969 31773 18003 31807
rect 18245 31773 18279 31807
rect 18337 31773 18371 31807
rect 18521 31773 18555 31807
rect 18705 31773 18739 31807
rect 21097 31773 21131 31807
rect 21373 31773 21407 31807
rect 21557 31773 21591 31807
rect 21649 31773 21683 31807
rect 21925 31773 21959 31807
rect 22201 31773 22235 31807
rect 22477 31773 22511 31807
rect 24501 31773 24535 31807
rect 24961 31773 24995 31807
rect 26157 31773 26191 31807
rect 26249 31773 26283 31807
rect 26433 31773 26467 31807
rect 27813 31773 27847 31807
rect 28549 31773 28583 31807
rect 28733 31773 28767 31807
rect 28917 31773 28951 31807
rect 29009 31773 29043 31807
rect 29101 31773 29135 31807
rect 29217 31773 29251 31807
rect 29377 31773 29411 31807
rect 30297 31773 30331 31807
rect 30481 31773 30515 31807
rect 30941 31773 30975 31807
rect 31401 31773 31435 31807
rect 31769 31773 31803 31807
rect 33333 31773 33367 31807
rect 33793 31773 33827 31807
rect 34713 31773 34747 31807
rect 5825 31705 5859 31739
rect 8447 31705 8481 31739
rect 9965 31705 9999 31739
rect 10057 31705 10091 31739
rect 10425 31705 10459 31739
rect 22385 31705 22419 31739
rect 25145 31705 25179 31739
rect 10635 31637 10669 31671
rect 13093 31637 13127 31671
rect 16129 31637 16163 31671
rect 28641 31637 28675 31671
rect 29285 31637 29319 31671
rect 30941 31637 30975 31671
rect 6193 31433 6227 31467
rect 29101 31433 29135 31467
rect 31033 31433 31067 31467
rect 33977 31433 34011 31467
rect 6653 31365 6687 31399
rect 8401 31365 8435 31399
rect 9597 31365 9631 31399
rect 13001 31365 13035 31399
rect 14473 31365 14507 31399
rect 24961 31365 24995 31399
rect 25697 31365 25731 31399
rect 27721 31365 27755 31399
rect 33517 31365 33551 31399
rect 5641 31297 5675 31331
rect 5825 31297 5859 31331
rect 5917 31297 5951 31331
rect 6009 31297 6043 31331
rect 8493 31297 8527 31331
rect 8677 31297 8711 31331
rect 8769 31297 8803 31331
rect 8862 31297 8896 31331
rect 9321 31297 9355 31331
rect 9505 31297 9539 31331
rect 9689 31297 9723 31331
rect 12633 31297 12667 31331
rect 12726 31297 12760 31331
rect 12909 31297 12943 31331
rect 13098 31297 13132 31331
rect 14105 31297 14139 31331
rect 14253 31297 14287 31331
rect 14381 31297 14415 31331
rect 14611 31297 14645 31331
rect 20453 31297 20487 31331
rect 20821 31297 20855 31331
rect 21097 31297 21131 31331
rect 21189 31297 21223 31331
rect 21557 31297 21591 31331
rect 22017 31297 22051 31331
rect 22282 31297 22316 31331
rect 23765 31297 23799 31331
rect 24133 31297 24167 31331
rect 24409 31297 24443 31331
rect 24777 31297 24811 31331
rect 25053 31297 25087 31331
rect 25145 31297 25179 31331
rect 25605 31297 25639 31331
rect 25789 31297 25823 31331
rect 26157 31297 26191 31331
rect 26433 31297 26467 31331
rect 26617 31297 26651 31331
rect 26985 31297 27019 31331
rect 27997 31297 28031 31331
rect 28549 31297 28583 31331
rect 29009 31297 29043 31331
rect 29285 31297 29319 31331
rect 29653 31297 29687 31331
rect 30205 31297 30239 31331
rect 31033 31297 31067 31331
rect 31217 31297 31251 31331
rect 33793 31297 33827 31331
rect 6377 31229 6411 31263
rect 21833 31229 21867 31263
rect 22109 31229 22143 31263
rect 22201 31229 22235 31263
rect 28457 31229 28491 31263
rect 30113 31229 30147 31263
rect 33609 31229 33643 31263
rect 9137 31161 9171 31195
rect 20545 31161 20579 31195
rect 23673 31161 23707 31195
rect 9873 31093 9907 31127
rect 13277 31093 13311 31127
rect 14749 31093 14783 31127
rect 25329 31093 25363 31127
rect 33793 31093 33827 31127
rect 7297 30889 7331 30923
rect 9781 30889 9815 30923
rect 10149 30889 10183 30923
rect 16497 30889 16531 30923
rect 17693 30889 17727 30923
rect 26065 30889 26099 30923
rect 26249 30889 26283 30923
rect 26617 30889 26651 30923
rect 28917 30889 28951 30923
rect 29193 30889 29227 30923
rect 29653 30889 29687 30923
rect 18061 30821 18095 30855
rect 24501 30821 24535 30855
rect 26985 30821 27019 30855
rect 28641 30821 28675 30855
rect 4169 30753 4203 30787
rect 9689 30753 9723 30787
rect 11437 30753 11471 30787
rect 26433 30753 26467 30787
rect 27813 30753 27847 30787
rect 29101 30753 29135 30787
rect 29837 30753 29871 30787
rect 33609 30753 33643 30787
rect 35541 30753 35575 30787
rect 6285 30685 6319 30719
rect 6469 30685 6503 30719
rect 6653 30685 6687 30719
rect 7205 30685 7239 30719
rect 9413 30685 9447 30719
rect 10057 30685 10091 30719
rect 10241 30685 10275 30719
rect 11345 30685 11379 30719
rect 11805 30685 11839 30719
rect 12357 30685 12391 30719
rect 12633 30685 12667 30719
rect 13001 30685 13035 30719
rect 15209 30685 15243 30719
rect 15393 30685 15427 30719
rect 16497 30685 16531 30719
rect 16681 30685 16715 30719
rect 17877 30685 17911 30719
rect 18153 30685 18187 30719
rect 19257 30685 19291 30719
rect 19441 30685 19475 30719
rect 19717 30685 19751 30719
rect 21465 30685 21499 30719
rect 21557 30685 21591 30719
rect 22937 30685 22971 30719
rect 23121 30685 23155 30719
rect 23213 30685 23247 30719
rect 23765 30685 23799 30719
rect 24041 30685 24075 30719
rect 24593 30685 24627 30719
rect 24961 30685 24995 30719
rect 25237 30685 25271 30719
rect 25881 30685 25915 30719
rect 26065 30685 26099 30719
rect 26341 30685 26375 30719
rect 26525 30685 26559 30719
rect 26617 30685 26651 30719
rect 26801 30685 26835 30719
rect 27629 30685 27663 30719
rect 28365 30685 28399 30719
rect 28641 30685 28675 30719
rect 28825 30685 28859 30719
rect 29193 30685 29227 30719
rect 29377 30685 29411 30719
rect 29561 30685 29595 30719
rect 33425 30685 33459 30719
rect 35265 30685 35299 30719
rect 4445 30617 4479 30651
rect 6193 30617 6227 30651
rect 6561 30617 6595 30651
rect 16037 30617 16071 30651
rect 16221 30617 16255 30651
rect 19809 30617 19843 30651
rect 24225 30617 24259 30651
rect 25605 30617 25639 30651
rect 27169 30617 27203 30651
rect 27537 30617 27571 30651
rect 32965 30617 32999 30651
rect 34805 30617 34839 30651
rect 6837 30549 6871 30583
rect 9965 30549 9999 30583
rect 15301 30549 15335 30583
rect 16405 30549 16439 30583
rect 22753 30549 22787 30583
rect 27261 30549 27295 30583
rect 27353 30549 27387 30583
rect 29101 30549 29135 30583
rect 29837 30549 29871 30583
rect 33241 30549 33275 30583
rect 34897 30549 34931 30583
rect 8677 30345 8711 30379
rect 11253 30345 11287 30379
rect 16037 30345 16071 30379
rect 26065 30345 26099 30379
rect 35909 30345 35943 30379
rect 10885 30277 10919 30311
rect 10977 30277 11011 30311
rect 23305 30277 23339 30311
rect 23673 30277 23707 30311
rect 32413 30277 32447 30311
rect 8493 30209 8527 30243
rect 8953 30209 8987 30243
rect 10609 30209 10643 30243
rect 10702 30209 10736 30243
rect 11074 30209 11108 30243
rect 11713 30209 11747 30243
rect 11989 30209 12023 30243
rect 14289 30209 14323 30243
rect 14841 30209 14875 30243
rect 14933 30209 14967 30243
rect 15301 30209 15335 30243
rect 15669 30209 15703 30243
rect 16681 30209 16715 30243
rect 16865 30209 16899 30243
rect 18245 30209 18279 30243
rect 19165 30209 19199 30243
rect 19349 30209 19383 30243
rect 19625 30209 19659 30243
rect 19993 30209 20027 30243
rect 21281 30209 21315 30243
rect 21373 30209 21407 30243
rect 22017 30209 22051 30243
rect 23029 30209 23063 30243
rect 23213 30209 23247 30243
rect 23489 30209 23523 30243
rect 23765 30209 23799 30243
rect 25145 30209 25179 30243
rect 25329 30209 25363 30243
rect 25605 30209 25639 30243
rect 25881 30209 25915 30243
rect 26065 30209 26099 30243
rect 26157 30209 26191 30243
rect 29653 30209 29687 30243
rect 30297 30209 30331 30243
rect 30757 30209 30791 30243
rect 31217 30209 31251 30243
rect 31585 30209 31619 30243
rect 32689 30209 32723 30243
rect 32873 30209 32907 30243
rect 33149 30209 33183 30243
rect 33425 30209 33459 30243
rect 33977 30209 34011 30243
rect 34437 30209 34471 30243
rect 34805 30209 34839 30243
rect 35357 30209 35391 30243
rect 35725 30209 35759 30243
rect 11529 30141 11563 30175
rect 14381 30141 14415 30175
rect 18521 30141 18555 30175
rect 22293 30141 22327 30175
rect 25697 30141 25731 30175
rect 30389 30141 30423 30175
rect 32137 30141 32171 30175
rect 35265 30141 35299 30175
rect 14657 30073 14691 30107
rect 20269 30073 20303 30107
rect 9045 30005 9079 30039
rect 11897 30005 11931 30039
rect 14473 30005 14507 30039
rect 15301 30005 15335 30039
rect 15485 30005 15519 30039
rect 16037 30005 16071 30039
rect 16221 30005 16255 30039
rect 16865 30005 16899 30039
rect 17049 30005 17083 30039
rect 18337 30005 18371 30039
rect 18797 30005 18831 30039
rect 23029 30005 23063 30039
rect 29929 30005 29963 30039
rect 30113 30005 30147 30039
rect 33701 30005 33735 30039
rect 35633 30005 35667 30039
rect 7665 29801 7699 29835
rect 8585 29801 8619 29835
rect 11437 29801 11471 29835
rect 14381 29801 14415 29835
rect 14473 29801 14507 29835
rect 19349 29801 19383 29835
rect 22661 29801 22695 29835
rect 35265 29801 35299 29835
rect 35449 29801 35483 29835
rect 37565 29801 37599 29835
rect 9137 29733 9171 29767
rect 10333 29733 10367 29767
rect 14565 29733 14599 29767
rect 16221 29733 16255 29767
rect 17877 29733 17911 29767
rect 23029 29733 23063 29767
rect 29837 29733 29871 29767
rect 30573 29733 30607 29767
rect 8033 29665 8067 29699
rect 8677 29665 8711 29699
rect 14933 29665 14967 29699
rect 18705 29665 18739 29699
rect 22109 29665 22143 29699
rect 22477 29665 22511 29699
rect 27445 29665 27479 29699
rect 27721 29665 27755 29699
rect 32045 29665 32079 29699
rect 35817 29665 35851 29699
rect 5457 29597 5491 29631
rect 5733 29597 5767 29631
rect 5825 29597 5859 29631
rect 7849 29597 7883 29631
rect 7941 29597 7975 29631
rect 8125 29597 8159 29631
rect 8401 29597 8435 29631
rect 8493 29597 8527 29631
rect 9321 29597 9355 29631
rect 9413 29597 9447 29631
rect 9689 29597 9723 29631
rect 9782 29597 9816 29631
rect 9965 29597 9999 29631
rect 10057 29597 10091 29631
rect 10195 29597 10229 29631
rect 10517 29597 10551 29631
rect 10793 29597 10827 29631
rect 11345 29597 11379 29631
rect 12725 29597 12759 29631
rect 12817 29597 12851 29631
rect 12909 29597 12943 29631
rect 13093 29597 13127 29631
rect 14841 29597 14875 29631
rect 15117 29597 15151 29631
rect 15393 29597 15427 29631
rect 16037 29597 16071 29631
rect 16129 29597 16163 29631
rect 16313 29597 16347 29631
rect 16497 29597 16531 29631
rect 16589 29597 16623 29631
rect 17049 29597 17083 29631
rect 17509 29597 17543 29631
rect 17877 29597 17911 29631
rect 18245 29597 18279 29631
rect 18889 29597 18923 29631
rect 19257 29597 19291 29631
rect 19533 29597 19567 29631
rect 19901 29597 19935 29631
rect 20085 29597 20119 29631
rect 20361 29597 20395 29631
rect 21557 29597 21591 29631
rect 21741 29597 21775 29631
rect 22017 29597 22051 29631
rect 22661 29597 22695 29631
rect 23029 29597 23063 29631
rect 23305 29597 23339 29631
rect 24869 29597 24903 29631
rect 25047 29597 25081 29631
rect 27629 29597 27663 29631
rect 28089 29597 28123 29631
rect 30297 29597 30331 29631
rect 30389 29597 30423 29631
rect 31309 29597 31343 29631
rect 31493 29597 31527 29631
rect 31794 29594 31828 29628
rect 32597 29597 32631 29631
rect 32965 29597 32999 29631
rect 33241 29597 33275 29631
rect 33609 29597 33643 29631
rect 34069 29597 34103 29631
rect 34345 29597 34379 29631
rect 34805 29597 34839 29631
rect 34897 29597 34931 29631
rect 35265 29597 35299 29631
rect 35725 29597 35759 29631
rect 5641 29529 5675 29563
rect 9137 29529 9171 29563
rect 10701 29529 10735 29563
rect 11253 29529 11287 29563
rect 14105 29529 14139 29563
rect 15301 29529 15335 29563
rect 21005 29529 21039 29563
rect 22385 29529 22419 29563
rect 29837 29529 29871 29563
rect 30849 29529 30883 29563
rect 30941 29529 30975 29563
rect 31401 29529 31435 29563
rect 36093 29529 36127 29563
rect 37749 29529 37783 29563
rect 6009 29461 6043 29495
rect 12449 29461 12483 29495
rect 14749 29461 14783 29495
rect 15853 29461 15887 29495
rect 19073 29461 19107 29495
rect 22845 29461 22879 29495
rect 23213 29461 23247 29495
rect 24961 29461 24995 29495
rect 27813 29461 27847 29495
rect 27997 29461 28031 29495
rect 33885 29461 33919 29495
rect 35541 29461 35575 29495
rect 37841 29461 37875 29495
rect 7573 29257 7607 29291
rect 8217 29257 8251 29291
rect 9137 29257 9171 29291
rect 10333 29257 10367 29291
rect 10625 29257 10659 29291
rect 12265 29257 12299 29291
rect 12909 29257 12943 29291
rect 15393 29257 15427 29291
rect 18245 29257 18279 29291
rect 26065 29257 26099 29291
rect 26525 29257 26559 29291
rect 27261 29257 27295 29291
rect 30481 29257 30515 29291
rect 31677 29257 31711 29291
rect 36001 29257 36035 29291
rect 36369 29257 36403 29291
rect 40969 29257 41003 29291
rect 6101 29189 6135 29223
rect 9965 29189 9999 29223
rect 10425 29189 10459 29223
rect 14473 29189 14507 29223
rect 15025 29189 15059 29223
rect 15241 29189 15275 29223
rect 21005 29189 21039 29223
rect 21189 29189 21223 29223
rect 23213 29189 23247 29223
rect 23995 29189 24029 29223
rect 30322 29189 30356 29223
rect 31585 29189 31619 29223
rect 7481 29121 7515 29155
rect 7665 29121 7699 29155
rect 8309 29121 8343 29155
rect 8677 29121 8711 29155
rect 8953 29121 8987 29155
rect 9689 29121 9723 29155
rect 9782 29121 9816 29155
rect 10057 29121 10091 29155
rect 10195 29121 10229 29155
rect 14749 29121 14783 29155
rect 15945 29121 15979 29155
rect 16957 29121 16991 29155
rect 17141 29121 17175 29155
rect 17233 29121 17267 29155
rect 18429 29121 18463 29155
rect 18613 29121 18647 29155
rect 18981 29121 19015 29155
rect 19441 29121 19475 29155
rect 19717 29121 19751 29155
rect 20269 29121 20303 29155
rect 20361 29121 20395 29155
rect 20453 29121 20487 29155
rect 20545 29121 20579 29155
rect 21373 29121 21407 29155
rect 22201 29121 22235 29155
rect 22477 29121 22511 29155
rect 22661 29121 22695 29155
rect 22753 29121 22787 29155
rect 23121 29121 23155 29155
rect 23581 29121 23615 29155
rect 24225 29121 24259 29155
rect 24317 29121 24351 29155
rect 24501 29121 24535 29155
rect 25145 29121 25179 29155
rect 25329 29121 25363 29155
rect 25421 29121 25455 29155
rect 25513 29121 25547 29155
rect 25881 29121 25915 29155
rect 26157 29121 26191 29155
rect 26525 29121 26559 29155
rect 26617 29121 26651 29155
rect 27445 29121 27479 29155
rect 27629 29121 27663 29155
rect 28181 29121 28215 29155
rect 28549 29121 28583 29155
rect 29561 29121 29595 29155
rect 30205 29121 30239 29155
rect 30573 29121 30607 29155
rect 31309 29121 31343 29155
rect 31794 29121 31828 29155
rect 32781 29121 32815 29155
rect 33609 29121 33643 29155
rect 33885 29121 33919 29155
rect 34161 29121 34195 29155
rect 40785 29121 40819 29155
rect 4077 29053 4111 29087
rect 7757 29053 7791 29087
rect 12633 29053 12667 29087
rect 12725 29053 12759 29087
rect 14657 29053 14691 29087
rect 15761 29053 15795 29087
rect 18153 29053 18187 29087
rect 18889 29053 18923 29087
rect 20085 29053 20119 29087
rect 22385 29053 22419 29087
rect 23029 29053 23063 29087
rect 24869 29053 24903 29087
rect 29745 29053 29779 29087
rect 29837 29053 29871 29087
rect 30113 29053 30147 29087
rect 36461 29053 36495 29087
rect 36553 29053 36587 29087
rect 8033 28985 8067 29019
rect 8493 28985 8527 29019
rect 8769 28985 8803 29019
rect 14933 28985 14967 29019
rect 16129 28985 16163 29019
rect 16957 28985 16991 29019
rect 19257 28985 19291 29019
rect 19625 28985 19659 29019
rect 22017 28985 22051 29019
rect 22293 28985 22327 29019
rect 24777 28985 24811 29019
rect 25697 28985 25731 29019
rect 28089 28985 28123 29019
rect 30849 28985 30883 29019
rect 31953 28985 31987 29019
rect 4340 28917 4374 28951
rect 10609 28917 10643 28951
rect 10793 28917 10827 28951
rect 14473 28917 14507 28951
rect 15209 28917 15243 28951
rect 23397 28917 23431 28951
rect 23949 28917 23983 28951
rect 25881 28917 25915 28951
rect 31033 28917 31067 28951
rect 33057 28917 33091 28951
rect 5549 28713 5583 28747
rect 5898 28713 5932 28747
rect 7389 28713 7423 28747
rect 9229 28713 9263 28747
rect 14381 28713 14415 28747
rect 19533 28713 19567 28747
rect 22845 28713 22879 28747
rect 29561 28713 29595 28747
rect 39129 28713 39163 28747
rect 25881 28645 25915 28679
rect 25973 28645 26007 28679
rect 28181 28645 28215 28679
rect 13093 28577 13127 28611
rect 19441 28577 19475 28611
rect 24961 28577 24995 28611
rect 37381 28577 37415 28611
rect 4997 28509 5031 28543
rect 5181 28509 5215 28543
rect 5365 28509 5399 28543
rect 5641 28509 5675 28543
rect 8953 28509 8987 28543
rect 9137 28509 9171 28543
rect 10333 28509 10367 28543
rect 10793 28509 10827 28543
rect 11897 28509 11931 28543
rect 11989 28509 12023 28543
rect 12173 28509 12207 28543
rect 12265 28509 12299 28543
rect 12725 28509 12759 28543
rect 12909 28509 12943 28543
rect 14289 28509 14323 28543
rect 19533 28509 19567 28543
rect 20361 28509 20395 28543
rect 20545 28509 20579 28543
rect 21281 28509 21315 28543
rect 21649 28509 21683 28543
rect 24409 28509 24443 28543
rect 24593 28509 24627 28543
rect 26617 28509 26651 28543
rect 26985 28509 27019 28543
rect 27169 28509 27203 28543
rect 27813 28509 27847 28543
rect 27997 28509 28031 28543
rect 28641 28509 28675 28543
rect 29101 28509 29135 28543
rect 29561 28509 29595 28543
rect 29745 28509 29779 28543
rect 30113 28509 30147 28543
rect 30297 28509 30331 28543
rect 37289 28509 37323 28543
rect 5273 28441 5307 28475
rect 10517 28441 10551 28475
rect 11529 28441 11563 28475
rect 14105 28441 14139 28475
rect 19257 28441 19291 28475
rect 20729 28441 20763 28475
rect 21465 28441 21499 28475
rect 21557 28441 21591 28475
rect 22661 28441 22695 28475
rect 22877 28441 22911 28475
rect 37657 28441 37691 28475
rect 10701 28373 10735 28407
rect 12357 28373 12391 28407
rect 19717 28373 19751 28407
rect 21833 28373 21867 28407
rect 23029 28373 23063 28407
rect 24593 28373 24627 28407
rect 28733 28373 28767 28407
rect 30297 28373 30331 28407
rect 37105 28373 37139 28407
rect 8953 28169 8987 28203
rect 11069 28169 11103 28203
rect 18797 28169 18831 28203
rect 27169 28169 27203 28203
rect 32689 28169 32723 28203
rect 32873 28169 32907 28203
rect 33425 28169 33459 28203
rect 33609 28169 33643 28203
rect 34529 28169 34563 28203
rect 34897 28169 34931 28203
rect 37381 28169 37415 28203
rect 37749 28169 37783 28203
rect 39129 28169 39163 28203
rect 8309 28101 8343 28135
rect 9597 28101 9631 28135
rect 12541 28101 12575 28135
rect 17969 28101 18003 28135
rect 19257 28101 19291 28135
rect 30665 28101 30699 28135
rect 30849 28101 30883 28135
rect 31033 28101 31067 28135
rect 33057 28101 33091 28135
rect 37841 28101 37875 28135
rect 1409 28033 1443 28067
rect 4261 28033 4295 28067
rect 8033 28033 8067 28067
rect 8861 28033 8895 28067
rect 9229 28033 9263 28067
rect 9321 28033 9355 28067
rect 9413 28033 9447 28067
rect 12265 28033 12299 28067
rect 12413 28033 12447 28067
rect 12633 28033 12667 28067
rect 12771 28033 12805 28067
rect 14841 28033 14875 28067
rect 14933 28033 14967 28067
rect 15117 28033 15151 28067
rect 15761 28033 15795 28067
rect 15945 28033 15979 28067
rect 16313 28033 16347 28067
rect 17693 28033 17727 28067
rect 18245 28033 18279 28067
rect 18613 28033 18647 28067
rect 18889 28033 18923 28067
rect 18982 28033 19016 28067
rect 19165 28033 19199 28067
rect 19354 28033 19388 28067
rect 27353 28033 27387 28067
rect 27537 28033 27571 28067
rect 29837 28033 29871 28067
rect 31677 28033 31711 28067
rect 31861 28033 31895 28067
rect 32321 28033 32355 28067
rect 32505 28033 32539 28067
rect 32597 28033 32631 28067
rect 33241 28033 33275 28067
rect 33333 28033 33367 28067
rect 33977 28033 34011 28067
rect 38577 28033 38611 28067
rect 4997 27965 5031 27999
rect 9045 27965 9079 27999
rect 9597 27965 9631 27999
rect 10609 27965 10643 27999
rect 15025 27965 15059 27999
rect 17969 27965 18003 27999
rect 18153 27965 18187 27999
rect 29929 27965 29963 27999
rect 31953 27965 31987 27999
rect 32965 27965 32999 27999
rect 33701 27965 33735 27999
rect 34253 27965 34287 27999
rect 35265 27965 35299 27999
rect 35357 27965 35391 27999
rect 37933 27965 37967 27999
rect 1593 27897 1627 27931
rect 9229 27897 9263 27931
rect 10885 27897 10919 27931
rect 14657 27897 14691 27931
rect 12909 27829 12943 27863
rect 16221 27829 16255 27863
rect 17785 27829 17819 27863
rect 18521 27829 18555 27863
rect 19533 27829 19567 27863
rect 29929 27829 29963 27863
rect 30205 27829 30239 27863
rect 34345 27829 34379 27863
rect 35541 27829 35575 27863
rect 5549 27625 5583 27659
rect 12265 27625 12299 27659
rect 12909 27625 12943 27659
rect 13461 27625 13495 27659
rect 14105 27625 14139 27659
rect 19073 27625 19107 27659
rect 20913 27625 20947 27659
rect 22845 27625 22879 27659
rect 23121 27625 23155 27659
rect 28457 27625 28491 27659
rect 30297 27625 30331 27659
rect 31125 27625 31159 27659
rect 35068 27625 35102 27659
rect 12633 27557 12667 27591
rect 15025 27557 15059 27591
rect 22109 27557 22143 27591
rect 23305 27557 23339 27591
rect 28641 27557 28675 27591
rect 29101 27557 29135 27591
rect 5641 27489 5675 27523
rect 14381 27489 14415 27523
rect 17144 27489 17178 27523
rect 27077 27489 27111 27523
rect 27261 27489 27295 27523
rect 28733 27489 28767 27523
rect 30205 27489 30239 27523
rect 30941 27489 30975 27523
rect 31677 27489 31711 27523
rect 34805 27489 34839 27523
rect 36829 27489 36863 27523
rect 3801 27421 3835 27455
rect 6377 27421 6411 27455
rect 6561 27421 6595 27455
rect 6745 27421 6779 27455
rect 8953 27421 8987 27455
rect 9229 27421 9263 27455
rect 9321 27421 9355 27455
rect 12265 27421 12299 27455
rect 12357 27421 12391 27455
rect 14289 27421 14323 27455
rect 14473 27421 14507 27455
rect 14565 27421 14599 27455
rect 15209 27421 15243 27455
rect 15301 27421 15335 27455
rect 15577 27421 15611 27455
rect 15669 27421 15703 27455
rect 16129 27421 16163 27455
rect 16865 27421 16899 27455
rect 16957 27421 16991 27455
rect 17233 27421 17267 27455
rect 17417 27421 17451 27455
rect 18521 27421 18555 27455
rect 18705 27421 18739 27455
rect 18797 27421 18831 27455
rect 18889 27421 18923 27455
rect 21097 27421 21131 27455
rect 21189 27421 21223 27455
rect 21373 27421 21407 27455
rect 21465 27421 21499 27455
rect 22569 27421 22603 27455
rect 23673 27421 23707 27455
rect 23857 27421 23891 27455
rect 24225 27421 24259 27455
rect 25053 27421 25087 27455
rect 25237 27421 25271 27455
rect 25513 27421 25547 27455
rect 25605 27421 25639 27455
rect 25973 27421 26007 27455
rect 26525 27421 26559 27455
rect 26617 27421 26651 27455
rect 26709 27421 26743 27455
rect 26801 27421 26835 27455
rect 26985 27421 27019 27455
rect 27537 27421 27571 27455
rect 28917 27421 28951 27455
rect 29009 27421 29043 27455
rect 29193 27421 29227 27455
rect 29377 27421 29411 27455
rect 30389 27421 30423 27455
rect 31125 27421 31159 27455
rect 31401 27421 31435 27455
rect 33517 27421 33551 27455
rect 4077 27353 4111 27387
rect 6653 27353 6687 27387
rect 9137 27353 9171 27387
rect 12734 27353 12768 27387
rect 12909 27353 12943 27387
rect 13277 27353 13311 27387
rect 13461 27353 13495 27387
rect 15393 27353 15427 27387
rect 22109 27353 22143 27387
rect 22937 27353 22971 27387
rect 28273 27353 28307 27387
rect 29929 27353 29963 27387
rect 30665 27353 30699 27387
rect 6285 27285 6319 27319
rect 6929 27285 6963 27319
rect 9505 27285 9539 27319
rect 13093 27285 13127 27319
rect 13645 27285 13679 27319
rect 16313 27285 16347 27319
rect 17141 27285 17175 27319
rect 17417 27285 17451 27319
rect 22661 27285 22695 27319
rect 23137 27285 23171 27319
rect 24133 27285 24167 27319
rect 25973 27285 26007 27319
rect 28473 27285 28507 27319
rect 30573 27285 30607 27319
rect 31309 27285 31343 27319
rect 34069 27285 34103 27319
rect 3985 27081 4019 27115
rect 4905 27081 4939 27115
rect 12925 27081 12959 27115
rect 14473 27081 14507 27115
rect 15485 27081 15519 27115
rect 18731 27081 18765 27115
rect 27169 27081 27203 27115
rect 27905 27081 27939 27115
rect 28549 27081 28583 27115
rect 28917 27081 28951 27115
rect 30297 27081 30331 27115
rect 6653 27013 6687 27047
rect 8401 27013 8435 27047
rect 12725 27013 12759 27047
rect 15301 27013 15335 27047
rect 17141 27013 17175 27047
rect 18521 27013 18555 27047
rect 33333 27013 33367 27047
rect 17371 26979 17405 27013
rect 4169 26945 4203 26979
rect 6377 26945 6411 26979
rect 8585 26945 8619 26979
rect 8769 26945 8803 26979
rect 9045 26945 9079 26979
rect 9321 26945 9355 26979
rect 9689 26945 9723 26979
rect 9781 26945 9815 26979
rect 9965 26945 9999 26979
rect 10057 26945 10091 26979
rect 11713 26945 11747 26979
rect 12081 26945 12115 26979
rect 12173 26945 12207 26979
rect 14105 26945 14139 26979
rect 14933 26945 14967 26979
rect 15485 26945 15519 26979
rect 15945 26945 15979 26979
rect 16313 26945 16347 26979
rect 16681 26945 16715 26979
rect 19165 26945 19199 26979
rect 20637 26945 20671 26979
rect 20821 26945 20855 26979
rect 21189 26945 21223 26979
rect 21465 26945 21499 26979
rect 21649 26945 21683 26979
rect 22845 26945 22879 26979
rect 23213 26945 23247 26979
rect 23581 26945 23615 26979
rect 24409 26945 24443 26979
rect 24593 26945 24627 26979
rect 24961 26945 24995 26979
rect 25145 26945 25179 26979
rect 25329 26945 25363 26979
rect 25697 26945 25731 26979
rect 27169 26945 27203 26979
rect 27721 26945 27755 26979
rect 27813 26945 27847 26979
rect 28089 26945 28123 26979
rect 28273 26945 28307 26979
rect 28549 26945 28583 26979
rect 28917 26945 28951 26979
rect 29009 26945 29043 26979
rect 30205 26945 30239 26979
rect 33057 26945 33091 26979
rect 33241 26945 33275 26979
rect 33425 26945 33459 26979
rect 33701 26945 33735 26979
rect 4997 26877 5031 26911
rect 5181 26877 5215 26911
rect 9137 26877 9171 26911
rect 9229 26877 9263 26911
rect 11529 26877 11563 26911
rect 14197 26877 14231 26911
rect 14749 26877 14783 26911
rect 15209 26877 15243 26911
rect 19257 26877 19291 26911
rect 20453 26877 20487 26911
rect 23765 26877 23799 26911
rect 24869 26877 24903 26911
rect 25973 26877 26007 26911
rect 26985 26877 27019 26911
rect 27537 26877 27571 26911
rect 28825 26877 28859 26911
rect 29193 26877 29227 26911
rect 30481 26877 30515 26911
rect 33977 26877 34011 26911
rect 35449 26877 35483 26911
rect 4537 26809 4571 26843
rect 20085 26809 20119 26843
rect 20545 26809 20579 26843
rect 24041 26809 24075 26843
rect 24593 26809 24627 26843
rect 24685 26809 24719 26843
rect 25881 26809 25915 26843
rect 28365 26809 28399 26843
rect 28641 26809 28675 26843
rect 30573 26809 30607 26843
rect 33609 26809 33643 26843
rect 8677 26741 8711 26775
rect 8861 26741 8895 26775
rect 9505 26741 9539 26775
rect 11989 26741 12023 26775
rect 12265 26741 12299 26775
rect 12633 26741 12667 26775
rect 12909 26741 12943 26775
rect 13093 26741 13127 26775
rect 14105 26741 14139 26775
rect 16773 26741 16807 26775
rect 17325 26741 17359 26775
rect 17509 26741 17543 26775
rect 18705 26741 18739 26775
rect 18889 26741 18923 26775
rect 19349 26741 19383 26775
rect 19533 26741 19567 26775
rect 20361 26741 20395 26775
rect 20913 26741 20947 26775
rect 21281 26741 21315 26775
rect 21373 26741 21407 26775
rect 30021 26741 30055 26775
rect 30765 26741 30799 26775
rect 7941 26537 7975 26571
rect 19717 26537 19751 26571
rect 33149 26537 33183 26571
rect 35541 26537 35575 26571
rect 5365 26469 5399 26503
rect 10517 26469 10551 26503
rect 11437 26469 11471 26503
rect 22201 26469 22235 26503
rect 22845 26469 22879 26503
rect 26525 26469 26559 26503
rect 33241 26469 33275 26503
rect 6009 26401 6043 26435
rect 9597 26401 9631 26435
rect 15117 26401 15151 26435
rect 15393 26401 15427 26435
rect 15761 26401 15795 26435
rect 18245 26401 18279 26435
rect 19625 26401 19659 26435
rect 19809 26401 19843 26435
rect 23121 26401 23155 26435
rect 25605 26401 25639 26435
rect 5273 26333 5307 26367
rect 7665 26333 7699 26367
rect 9137 26333 9171 26367
rect 9229 26333 9263 26367
rect 9439 26333 9473 26367
rect 10701 26333 10735 26367
rect 10793 26333 10827 26367
rect 11345 26333 11379 26367
rect 11529 26333 11563 26367
rect 15301 26333 15335 26367
rect 15485 26333 15519 26367
rect 15577 26333 15611 26367
rect 15945 26333 15979 26367
rect 17969 26333 18003 26367
rect 18705 26333 18739 26367
rect 18797 26333 18831 26367
rect 18889 26333 18923 26367
rect 19073 26333 19107 26367
rect 19901 26333 19935 26367
rect 20085 26333 20119 26367
rect 20637 26333 20671 26367
rect 20729 26333 20763 26367
rect 20913 26333 20947 26367
rect 21005 26333 21039 26367
rect 22109 26333 22143 26367
rect 22845 26333 22879 26367
rect 22937 26333 22971 26367
rect 24593 26333 24627 26367
rect 24961 26333 24995 26367
rect 25421 26333 25455 26367
rect 25789 26333 25823 26367
rect 25881 26333 25915 26367
rect 26050 26333 26084 26367
rect 26157 26333 26191 26367
rect 26433 26333 26467 26367
rect 26617 26333 26651 26367
rect 26709 26333 26743 26367
rect 32137 26333 32171 26367
rect 32505 26333 32539 26367
rect 33425 26333 33459 26367
rect 33517 26333 33551 26367
rect 34713 26333 34747 26367
rect 35449 26333 35483 26367
rect 35817 26333 35851 26367
rect 35909 26333 35943 26367
rect 5733 26265 5767 26299
rect 8953 26265 8987 26299
rect 9321 26265 9355 26299
rect 10517 26265 10551 26299
rect 18429 26265 18463 26299
rect 32321 26265 32355 26299
rect 32413 26265 32447 26299
rect 32781 26265 32815 26299
rect 32973 26265 33007 26299
rect 33241 26265 33275 26299
rect 35357 26265 35391 26299
rect 5089 26197 5123 26231
rect 5825 26197 5859 26231
rect 16129 26197 16163 26231
rect 19349 26197 19383 26231
rect 20453 26197 20487 26231
rect 24501 26197 24535 26231
rect 26249 26197 26283 26231
rect 32689 26197 32723 26231
rect 36093 26197 36127 26231
rect 8401 25993 8435 26027
rect 11161 25993 11195 26027
rect 14289 25993 14323 26027
rect 27997 25993 28031 26027
rect 28565 25993 28599 26027
rect 31309 25993 31343 26027
rect 31953 25993 31987 26027
rect 32965 25993 32999 26027
rect 35449 25993 35483 26027
rect 4721 25925 4755 25959
rect 10057 25925 10091 25959
rect 11805 25925 11839 25959
rect 19073 25925 19107 25959
rect 25145 25925 25179 25959
rect 28365 25925 28399 25959
rect 30757 25925 30791 25959
rect 33425 25925 33459 25959
rect 33885 25925 33919 25959
rect 7205 25857 7239 25891
rect 8125 25857 8159 25891
rect 8769 25857 8803 25891
rect 8861 25857 8895 25891
rect 9413 25857 9447 25891
rect 9781 25857 9815 25891
rect 9929 25857 9963 25891
rect 10149 25857 10183 25891
rect 10287 25857 10321 25891
rect 11069 25857 11103 25891
rect 12817 25857 12851 25891
rect 14473 25857 14507 25891
rect 17049 25857 17083 25891
rect 17233 25857 17267 25891
rect 17326 25879 17360 25913
rect 17451 25857 17485 25891
rect 18337 25857 18371 25891
rect 18521 25857 18555 25891
rect 19809 25857 19843 25891
rect 19993 25857 20027 25891
rect 20085 25857 20119 25891
rect 24869 25857 24903 25891
rect 24962 25857 24996 25891
rect 25237 25857 25271 25891
rect 25334 25857 25368 25891
rect 26341 25857 26375 25891
rect 26433 25857 26467 25891
rect 26617 25857 26651 25891
rect 27445 25857 27479 25891
rect 27537 25857 27571 25891
rect 27905 25857 27939 25891
rect 30573 25857 30607 25891
rect 30941 25857 30975 25891
rect 31585 25857 31619 25891
rect 32505 25857 32539 25891
rect 32781 25857 32815 25891
rect 33333 25857 33367 25891
rect 33517 25857 33551 25891
rect 35817 25857 35851 25891
rect 36829 25857 36863 25891
rect 4445 25789 4479 25823
rect 6193 25789 6227 25823
rect 6469 25789 6503 25823
rect 7113 25789 7147 25823
rect 9045 25789 9079 25823
rect 9689 25789 9723 25823
rect 12633 25789 12667 25823
rect 13093 25789 13127 25823
rect 14749 25789 14783 25823
rect 18245 25789 18279 25823
rect 18429 25789 18463 25823
rect 19625 25789 19659 25823
rect 25697 25789 25731 25823
rect 26157 25789 26191 25823
rect 27353 25789 27387 25823
rect 27629 25789 27663 25823
rect 31677 25789 31711 25823
rect 33609 25789 33643 25823
rect 35909 25789 35943 25823
rect 36185 25789 36219 25823
rect 17693 25721 17727 25755
rect 25513 25721 25547 25755
rect 32597 25721 32631 25755
rect 7297 25653 7331 25687
rect 8953 25653 8987 25687
rect 9229 25653 9263 25687
rect 9597 25653 9631 25687
rect 10425 25653 10459 25687
rect 12909 25653 12943 25687
rect 13001 25653 13035 25687
rect 14657 25653 14691 25687
rect 18061 25653 18095 25687
rect 27169 25653 27203 25687
rect 28549 25653 28583 25687
rect 28733 25653 28767 25687
rect 31585 25653 31619 25687
rect 35357 25653 35391 25687
rect 36093 25653 36127 25687
rect 5549 25449 5583 25483
rect 9137 25449 9171 25483
rect 9689 25449 9723 25483
rect 15393 25449 15427 25483
rect 15577 25449 15611 25483
rect 16681 25449 16715 25483
rect 28089 25449 28123 25483
rect 31033 25449 31067 25483
rect 7849 25381 7883 25415
rect 9505 25381 9539 25415
rect 18245 25381 18279 25415
rect 28181 25381 28215 25415
rect 3801 25313 3835 25347
rect 6653 25313 6687 25347
rect 6745 25313 6779 25347
rect 14565 25313 14599 25347
rect 14933 25313 14967 25347
rect 15669 25313 15703 25347
rect 16037 25313 16071 25347
rect 16865 25313 16899 25347
rect 17049 25313 17083 25347
rect 17969 25313 18003 25347
rect 18337 25313 18371 25347
rect 28365 25313 28399 25347
rect 29653 25313 29687 25347
rect 31309 25313 31343 25347
rect 32505 25313 32539 25347
rect 34529 25313 34563 25347
rect 35081 25313 35115 25347
rect 6561 25245 6595 25279
rect 6837 25245 6871 25279
rect 7849 25245 7883 25279
rect 8125 25245 8159 25279
rect 8677 25245 8711 25279
rect 9321 25245 9355 25279
rect 9597 25245 9631 25279
rect 9689 25245 9723 25279
rect 9873 25245 9907 25279
rect 11161 25245 11195 25279
rect 11345 25245 11379 25279
rect 14749 25245 14783 25279
rect 15209 25245 15243 25279
rect 15485 25245 15519 25279
rect 15577 25245 15611 25279
rect 16221 25245 16255 25279
rect 16957 25245 16991 25279
rect 17141 25245 17175 25279
rect 18153 25245 18187 25279
rect 18429 25245 18463 25279
rect 18613 25245 18647 25279
rect 21005 25245 21039 25279
rect 21281 25245 21315 25279
rect 21373 25245 21407 25279
rect 22661 25245 22695 25279
rect 22753 25245 22787 25279
rect 22937 25245 22971 25279
rect 23029 25245 23063 25279
rect 25145 25245 25179 25279
rect 25237 25245 25271 25279
rect 25421 25245 25455 25279
rect 25513 25245 25547 25279
rect 28089 25245 28123 25279
rect 29009 25245 29043 25279
rect 29269 25239 29303 25273
rect 29561 25245 29595 25279
rect 29745 25245 29779 25279
rect 30297 25245 30331 25279
rect 30481 25245 30515 25279
rect 31033 25245 31067 25279
rect 31125 25245 31159 25279
rect 34805 25245 34839 25279
rect 36829 25245 36863 25279
rect 4077 25177 4111 25211
rect 8309 25177 8343 25211
rect 16497 25177 16531 25211
rect 16589 25177 16623 25211
rect 21189 25177 21223 25211
rect 32781 25177 32815 25211
rect 6377 25109 6411 25143
rect 8033 25109 8067 25143
rect 11345 25109 11379 25143
rect 15025 25109 15059 25143
rect 15945 25109 15979 25143
rect 21557 25109 21591 25143
rect 22477 25109 22511 25143
rect 24961 25109 24995 25143
rect 28825 25109 28859 25143
rect 29193 25109 29227 25143
rect 30389 25109 30423 25143
rect 3709 24905 3743 24939
rect 4629 24905 4663 24939
rect 12265 24837 12299 24871
rect 12357 24837 12391 24871
rect 13645 24837 13679 24871
rect 13737 24837 13771 24871
rect 15577 24837 15611 24871
rect 15669 24837 15703 24871
rect 28365 24837 28399 24871
rect 3893 24769 3927 24803
rect 8033 24769 8067 24803
rect 8125 24769 8159 24803
rect 8309 24769 8343 24803
rect 8401 24769 8435 24803
rect 8493 24769 8527 24803
rect 8641 24769 8675 24803
rect 8769 24769 8803 24803
rect 8861 24769 8895 24803
rect 8999 24769 9033 24803
rect 11989 24769 12023 24803
rect 12137 24769 12171 24803
rect 12454 24769 12488 24803
rect 12725 24769 12759 24803
rect 12818 24769 12852 24803
rect 13001 24769 13035 24803
rect 13093 24769 13127 24803
rect 13190 24769 13224 24803
rect 13461 24769 13495 24803
rect 13829 24769 13863 24803
rect 14289 24769 14323 24803
rect 14381 24769 14415 24803
rect 14565 24769 14599 24803
rect 14657 24769 14691 24803
rect 15301 24769 15335 24803
rect 15394 24769 15428 24803
rect 15766 24769 15800 24803
rect 17325 24769 17359 24803
rect 19165 24769 19199 24803
rect 19349 24769 19383 24803
rect 19993 24769 20027 24803
rect 20361 24769 20395 24803
rect 20729 24769 20763 24803
rect 21097 24769 21131 24803
rect 21649 24769 21683 24803
rect 21925 24769 21959 24803
rect 22385 24769 22419 24803
rect 23949 24769 23983 24803
rect 24225 24769 24259 24803
rect 27077 24769 27111 24803
rect 27261 24769 27295 24803
rect 28549 24769 28583 24803
rect 28641 24769 28675 24803
rect 31309 24769 31343 24803
rect 40877 24769 40911 24803
rect 4721 24701 4755 24735
rect 4905 24701 4939 24735
rect 17601 24701 17635 24735
rect 19717 24701 19751 24735
rect 20821 24701 20855 24735
rect 22109 24701 22143 24735
rect 22293 24701 22327 24735
rect 22661 24701 22695 24735
rect 27445 24701 27479 24735
rect 27537 24701 27571 24735
rect 31125 24701 31159 24735
rect 4261 24633 4295 24667
rect 17509 24633 17543 24667
rect 19625 24633 19659 24667
rect 22201 24633 22235 24667
rect 22937 24633 22971 24667
rect 24041 24633 24075 24667
rect 24133 24633 24167 24667
rect 7849 24565 7883 24599
rect 9137 24565 9171 24599
rect 12633 24565 12667 24599
rect 13369 24565 13403 24599
rect 14013 24565 14047 24599
rect 14105 24565 14139 24599
rect 15945 24565 15979 24599
rect 17141 24565 17175 24599
rect 21925 24565 21959 24599
rect 22477 24565 22511 24599
rect 23765 24565 23799 24599
rect 28365 24565 28399 24599
rect 31493 24565 31527 24599
rect 41061 24565 41095 24599
rect 13369 24361 13403 24395
rect 15945 24361 15979 24395
rect 18153 24361 18187 24395
rect 19625 24361 19659 24395
rect 23213 24361 23247 24395
rect 26065 24361 26099 24395
rect 38025 24361 38059 24395
rect 11897 24293 11931 24327
rect 17785 24293 17819 24327
rect 19809 24293 19843 24327
rect 21373 24293 21407 24327
rect 22293 24293 22327 24327
rect 23397 24293 23431 24327
rect 23765 24293 23799 24327
rect 23857 24293 23891 24327
rect 24777 24293 24811 24327
rect 26893 24293 26927 24327
rect 27537 24293 27571 24327
rect 30205 24293 30239 24327
rect 30941 24293 30975 24327
rect 8953 24225 8987 24259
rect 9413 24225 9447 24259
rect 10793 24225 10827 24259
rect 11345 24225 11379 24259
rect 16037 24225 16071 24259
rect 16589 24225 16623 24259
rect 18889 24225 18923 24259
rect 21465 24225 21499 24259
rect 22385 24225 22419 24259
rect 26709 24225 26743 24259
rect 27629 24225 27663 24259
rect 29285 24225 29319 24259
rect 30297 24225 30331 24259
rect 36277 24225 36311 24259
rect 1501 24157 1535 24191
rect 6193 24157 6227 24191
rect 7113 24157 7147 24191
rect 9321 24157 9355 24191
rect 10333 24157 10367 24191
rect 10609 24157 10643 24191
rect 11437 24157 11471 24191
rect 11529 24157 11563 24191
rect 11621 24157 11655 24191
rect 11897 24157 11931 24191
rect 12081 24157 12115 24191
rect 12357 24157 12391 24191
rect 12541 24157 12575 24191
rect 12633 24157 12667 24191
rect 12817 24157 12851 24191
rect 12909 24157 12943 24191
rect 13001 24157 13035 24191
rect 13277 24157 13311 24191
rect 15853 24157 15887 24191
rect 16129 24157 16163 24191
rect 16313 24157 16347 24191
rect 16773 24157 16807 24191
rect 17049 24157 17083 24191
rect 17141 24157 17175 24191
rect 17325 24157 17359 24191
rect 17999 24157 18033 24191
rect 18245 24157 18279 24191
rect 18705 24157 18739 24191
rect 19533 24157 19567 24191
rect 19717 24157 19751 24191
rect 19993 24157 20027 24191
rect 20545 24157 20579 24191
rect 20769 24157 20803 24191
rect 21189 24157 21223 24191
rect 22201 24157 22235 24191
rect 22477 24157 22511 24191
rect 22661 24157 22695 24191
rect 22753 24157 22787 24191
rect 23121 24157 23155 24191
rect 23213 24157 23247 24191
rect 23673 24157 23707 24191
rect 23949 24157 23983 24191
rect 24409 24157 24443 24191
rect 24593 24157 24627 24191
rect 24685 24157 24719 24191
rect 24869 24157 24903 24191
rect 25053 24157 25087 24191
rect 26893 24157 26927 24191
rect 27169 24157 27203 24191
rect 27445 24157 27479 24191
rect 27721 24157 27755 24191
rect 27902 24135 27936 24169
rect 29193 24157 29227 24191
rect 30205 24157 30239 24191
rect 30757 24157 30791 24191
rect 30941 24157 30975 24191
rect 31953 24157 31987 24191
rect 14197 24089 14231 24123
rect 17233 24089 17267 24123
rect 18521 24089 18555 24123
rect 20361 24089 20395 24123
rect 20913 24089 20947 24123
rect 21005 24089 21039 24123
rect 27261 24089 27295 24123
rect 30573 24089 30607 24123
rect 36553 24089 36587 24123
rect 1593 24021 1627 24055
rect 6837 24021 6871 24055
rect 6929 24021 6963 24055
rect 9597 24021 9631 24055
rect 11161 24021 11195 24055
rect 13553 24021 13587 24055
rect 14473 24021 14507 24055
rect 15577 24021 15611 24055
rect 16957 24021 16991 24055
rect 19257 24021 19291 24055
rect 20637 24021 20671 24055
rect 22017 24021 22051 24055
rect 23489 24021 23523 24055
rect 26433 24021 26467 24055
rect 26525 24021 26559 24055
rect 27077 24021 27111 24055
rect 31769 24021 31803 24055
rect 6101 23817 6135 23851
rect 12173 23817 12207 23851
rect 15301 23817 15335 23851
rect 16221 23817 16255 23851
rect 26985 23817 27019 23851
rect 29837 23817 29871 23851
rect 36001 23817 36035 23851
rect 37289 23817 37323 23851
rect 4629 23749 4663 23783
rect 10057 23749 10091 23783
rect 10257 23749 10291 23783
rect 17056 23749 17090 23783
rect 20821 23749 20855 23783
rect 27721 23749 27755 23783
rect 37749 23749 37783 23783
rect 8309 23681 8343 23715
rect 10701 23681 10735 23715
rect 11621 23681 11655 23715
rect 11989 23681 12023 23715
rect 12725 23681 12759 23715
rect 12817 23681 12851 23715
rect 13001 23681 13035 23715
rect 13093 23681 13127 23715
rect 14933 23681 14967 23715
rect 16129 23681 16163 23715
rect 16313 23681 16347 23715
rect 17365 23681 17399 23715
rect 18613 23681 18647 23715
rect 18797 23681 18831 23715
rect 18889 23681 18923 23715
rect 20269 23681 20303 23715
rect 21005 23681 21039 23715
rect 21281 23681 21315 23715
rect 24225 23681 24259 23715
rect 24409 23681 24443 23715
rect 25145 23681 25179 23715
rect 25697 23681 25731 23715
rect 25973 23681 26007 23715
rect 26525 23681 26559 23715
rect 27905 23681 27939 23715
rect 29745 23681 29779 23715
rect 32137 23681 32171 23715
rect 34253 23681 34287 23715
rect 36553 23681 36587 23715
rect 37473 23681 37507 23715
rect 4353 23613 4387 23647
rect 6377 23613 6411 23647
rect 6653 23613 6687 23647
rect 8125 23613 8159 23647
rect 10517 23613 10551 23647
rect 10885 23613 10919 23647
rect 17233 23613 17267 23647
rect 20545 23613 20579 23647
rect 21097 23613 21131 23647
rect 21189 23613 21223 23647
rect 25421 23613 25455 23647
rect 25513 23613 25547 23647
rect 26801 23613 26835 23647
rect 27353 23613 27387 23647
rect 27445 23613 27479 23647
rect 30021 23613 30055 23647
rect 30297 23613 30331 23647
rect 32505 23613 32539 23647
rect 34529 23613 34563 23647
rect 36645 23613 36679 23647
rect 36737 23613 36771 23647
rect 38485 23613 38519 23647
rect 18705 23545 18739 23579
rect 20361 23545 20395 23579
rect 24593 23545 24627 23579
rect 25789 23545 25823 23579
rect 25881 23545 25915 23579
rect 27629 23545 27663 23579
rect 31769 23545 31803 23579
rect 36185 23545 36219 23579
rect 8861 23477 8895 23511
rect 10241 23477 10275 23511
rect 10425 23477 10459 23511
rect 11713 23477 11747 23511
rect 12541 23477 12575 23511
rect 15301 23477 15335 23511
rect 15485 23477 15519 23511
rect 17049 23477 17083 23511
rect 17509 23477 17543 23511
rect 18429 23477 18463 23511
rect 20453 23477 20487 23511
rect 24225 23477 24259 23511
rect 24961 23477 24995 23511
rect 25329 23477 25363 23511
rect 26341 23477 26375 23511
rect 26709 23477 26743 23511
rect 28089 23477 28123 23511
rect 33885 23477 33919 23511
rect 2053 23273 2087 23307
rect 5089 23273 5123 23307
rect 7113 23273 7147 23307
rect 11437 23273 11471 23307
rect 14841 23273 14875 23307
rect 20729 23273 20763 23307
rect 10425 23205 10459 23239
rect 20085 23205 20119 23239
rect 20453 23205 20487 23239
rect 25053 23205 25087 23239
rect 25237 23205 25271 23239
rect 27905 23205 27939 23239
rect 29837 23205 29871 23239
rect 30665 23205 30699 23239
rect 31585 23205 31619 23239
rect 6377 23137 6411 23171
rect 7757 23137 7791 23171
rect 16313 23137 16347 23171
rect 27445 23137 27479 23171
rect 30297 23137 30331 23171
rect 30389 23137 30423 23171
rect 32965 23137 32999 23171
rect 35357 23137 35391 23171
rect 1869 23069 1903 23103
rect 5273 23069 5307 23103
rect 6101 23069 6135 23103
rect 7573 23069 7607 23103
rect 9045 23069 9079 23103
rect 10609 23069 10643 23103
rect 10701 23069 10735 23103
rect 10793 23069 10827 23103
rect 14749 23069 14783 23103
rect 14933 23069 14967 23103
rect 15025 23069 15059 23103
rect 15209 23069 15243 23103
rect 15485 23069 15519 23103
rect 15577 23069 15611 23103
rect 15761 23069 15795 23103
rect 15853 23069 15887 23103
rect 16037 23069 16071 23103
rect 16129 23069 16163 23103
rect 17785 23069 17819 23103
rect 17969 23069 18003 23103
rect 20269 23069 20303 23103
rect 20361 23069 20395 23103
rect 20545 23069 20579 23103
rect 20913 23069 20947 23103
rect 21005 23069 21039 23103
rect 21097 23069 21131 23103
rect 21189 23069 21223 23103
rect 23213 23069 23247 23103
rect 23397 23069 23431 23103
rect 23489 23069 23523 23103
rect 24961 23069 24995 23103
rect 25145 23069 25179 23103
rect 25421 23069 25455 23103
rect 26985 23069 27019 23103
rect 27261 23069 27295 23103
rect 27537 23069 27571 23103
rect 27721 23069 27755 23103
rect 27997 23069 28031 23103
rect 28181 23069 28215 23103
rect 28733 23069 28767 23103
rect 28825 23069 28859 23103
rect 28917 23069 28951 23103
rect 29101 23069 29135 23103
rect 30849 23069 30883 23103
rect 31677 23069 31711 23103
rect 31861 23069 31895 23103
rect 32137 23069 32171 23103
rect 32413 23069 32447 23103
rect 32689 23069 32723 23103
rect 35081 23069 35115 23103
rect 11161 23001 11195 23035
rect 23029 23001 23063 23035
rect 26433 23001 26467 23035
rect 5733 22933 5767 22967
rect 6193 22933 6227 22967
rect 7481 22933 7515 22967
rect 9229 22933 9263 22967
rect 10977 22933 11011 22967
rect 14473 22933 14507 22967
rect 15301 22933 15335 22967
rect 18153 22933 18187 22967
rect 24685 22933 24719 22967
rect 28181 22933 28215 22967
rect 28457 22933 28491 22967
rect 30205 22933 30239 22967
rect 34437 22933 34471 22967
rect 34713 22933 34747 22967
rect 35173 22933 35207 22967
rect 11805 22729 11839 22763
rect 12357 22729 12391 22763
rect 16865 22729 16899 22763
rect 20913 22729 20947 22763
rect 24133 22729 24167 22763
rect 29285 22729 29319 22763
rect 34621 22729 34655 22763
rect 13001 22661 13035 22695
rect 13645 22661 13679 22695
rect 14841 22661 14875 22695
rect 16681 22661 16715 22695
rect 21833 22661 21867 22695
rect 23673 22661 23707 22695
rect 5273 22593 5307 22627
rect 10517 22593 10551 22627
rect 11713 22593 11747 22627
rect 11897 22593 11931 22627
rect 12081 22593 12115 22627
rect 12817 22593 12851 22627
rect 13185 22593 13219 22627
rect 13461 22593 13495 22627
rect 14381 22593 14415 22627
rect 15025 22593 15059 22627
rect 15117 22593 15151 22627
rect 15485 22593 15519 22627
rect 15761 22593 15795 22627
rect 16957 22593 16991 22627
rect 18245 22593 18279 22627
rect 18705 22593 18739 22627
rect 18889 22593 18923 22627
rect 19073 22593 19107 22627
rect 19993 22593 20027 22627
rect 20262 22593 20296 22627
rect 20545 22593 20579 22627
rect 20729 22593 20763 22627
rect 23857 22593 23891 22627
rect 24317 22593 24351 22627
rect 24501 22593 24535 22627
rect 29469 22593 29503 22627
rect 29561 22593 29595 22627
rect 29745 22593 29779 22627
rect 29837 22593 29871 22627
rect 34805 22593 34839 22627
rect 4629 22525 4663 22559
rect 7481 22525 7515 22559
rect 7757 22525 7791 22559
rect 9229 22525 9263 22559
rect 9781 22525 9815 22559
rect 10793 22525 10827 22559
rect 13277 22525 13311 22559
rect 15577 22525 15611 22559
rect 18337 22525 18371 22559
rect 20085 22525 20119 22559
rect 24041 22525 24075 22559
rect 24593 22525 24627 22559
rect 37289 22525 37323 22559
rect 37565 22525 37599 22559
rect 39313 22525 39347 22559
rect 5181 22457 5215 22491
rect 5549 22457 5583 22491
rect 23305 22457 23339 22491
rect 5733 22389 5767 22423
rect 10425 22389 10459 22423
rect 14473 22389 14507 22423
rect 15117 22389 15151 22423
rect 15301 22389 15335 22423
rect 15485 22389 15519 22423
rect 15945 22389 15979 22423
rect 16681 22389 16715 22423
rect 18245 22389 18279 22423
rect 18613 22389 18647 22423
rect 19993 22389 20027 22423
rect 20453 22389 20487 22423
rect 2513 22185 2547 22219
rect 5549 22185 5583 22219
rect 15761 22185 15795 22219
rect 17509 22185 17543 22219
rect 18613 22185 18647 22219
rect 23121 22185 23155 22219
rect 23673 22185 23707 22219
rect 37933 22185 37967 22219
rect 13645 22117 13679 22151
rect 17785 22117 17819 22151
rect 18797 22117 18831 22151
rect 20177 22117 20211 22151
rect 21097 22117 21131 22151
rect 22569 22117 22603 22151
rect 24961 22117 24995 22151
rect 3801 22049 3835 22083
rect 8585 22049 8619 22083
rect 11897 22049 11931 22083
rect 14473 22049 14507 22083
rect 18521 22049 18555 22083
rect 22937 22049 22971 22083
rect 23489 22049 23523 22083
rect 24133 22049 24167 22083
rect 24777 22049 24811 22083
rect 24869 22049 24903 22083
rect 28733 22049 28767 22083
rect 35633 22049 35667 22083
rect 36093 22049 36127 22083
rect 37657 22049 37691 22083
rect 2237 21981 2271 22015
rect 2329 21981 2363 22015
rect 7849 21981 7883 22015
rect 8033 21981 8067 22015
rect 9873 21981 9907 22015
rect 10057 21981 10091 22015
rect 10149 21981 10183 22015
rect 10241 21981 10275 22015
rect 10609 21981 10643 22015
rect 11713 21981 11747 22015
rect 11989 21981 12023 22015
rect 12173 21981 12207 22015
rect 12541 21981 12575 22015
rect 12725 21981 12759 22015
rect 13001 21981 13035 22015
rect 13185 21981 13219 22015
rect 13645 21981 13679 22015
rect 14381 21981 14415 22015
rect 14565 21981 14599 22015
rect 17417 21981 17451 22015
rect 17693 21981 17727 22015
rect 17969 21981 18003 22015
rect 18613 21981 18647 22015
rect 18889 21981 18923 22015
rect 19073 21981 19107 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 20361 21981 20395 22015
rect 20453 21981 20487 22015
rect 20637 21981 20671 22015
rect 20729 21981 20763 22015
rect 20821 21981 20855 22015
rect 21005 21981 21039 22015
rect 22753 21981 22787 22015
rect 23029 21981 23063 22015
rect 23305 21981 23339 22015
rect 23581 21981 23615 22015
rect 23857 21981 23891 22015
rect 24041 21981 24075 22015
rect 24685 21981 24719 22015
rect 25145 21981 25179 22015
rect 28457 21981 28491 22015
rect 29561 21981 29595 22015
rect 35725 21981 35759 22015
rect 37565 21981 37599 22015
rect 38117 21981 38151 22015
rect 4077 21913 4111 21947
rect 8217 21913 8251 21947
rect 8401 21913 8435 21947
rect 11345 21913 11379 21947
rect 11621 21913 11655 21947
rect 15393 21913 15427 21947
rect 15577 21913 15611 21947
rect 18153 21913 18187 21947
rect 18981 21913 19015 21947
rect 21373 21913 21407 21947
rect 27537 21913 27571 21947
rect 30297 21913 30331 21947
rect 7941 21845 7975 21879
rect 10425 21845 10459 21879
rect 11253 21845 11287 21879
rect 11529 21845 11563 21879
rect 12081 21845 12115 21879
rect 12633 21845 12667 21879
rect 19349 21845 19383 21879
rect 24409 21845 24443 21879
rect 27629 21845 27663 21879
rect 28089 21845 28123 21879
rect 28549 21845 28583 21879
rect 37105 21845 37139 21879
rect 37473 21845 37507 21879
rect 10241 21641 10275 21675
rect 17233 21641 17267 21675
rect 21465 21641 21499 21675
rect 31585 21641 31619 21675
rect 37013 21641 37047 21675
rect 5365 21573 5399 21607
rect 10977 21573 11011 21607
rect 14013 21573 14047 21607
rect 23489 21573 23523 21607
rect 25973 21573 26007 21607
rect 29285 21573 29319 21607
rect 30967 21573 31001 21607
rect 31141 21573 31175 21607
rect 31401 21573 31435 21607
rect 31861 21573 31895 21607
rect 36001 21573 36035 21607
rect 36369 21573 36403 21607
rect 36645 21573 36679 21607
rect 4629 21505 4663 21539
rect 5641 21505 5675 21539
rect 5825 21505 5859 21539
rect 6377 21505 6411 21539
rect 8401 21505 8435 21539
rect 10609 21505 10643 21539
rect 10701 21505 10735 21539
rect 11069 21505 11103 21539
rect 11529 21505 11563 21539
rect 13277 21505 13311 21539
rect 13461 21505 13495 21539
rect 13737 21505 13771 21539
rect 17049 21505 17083 21539
rect 17233 21505 17267 21539
rect 17509 21505 17543 21539
rect 17877 21505 17911 21539
rect 18245 21505 18279 21539
rect 18429 21505 18463 21539
rect 18521 21505 18555 21539
rect 18797 21505 18831 21539
rect 19073 21505 19107 21539
rect 21097 21505 21131 21539
rect 21833 21505 21867 21539
rect 22201 21505 22235 21539
rect 22661 21505 22695 21539
rect 23857 21505 23891 21539
rect 25605 21505 25639 21539
rect 25698 21505 25732 21539
rect 25881 21505 25915 21539
rect 26111 21505 26145 21539
rect 26341 21505 26375 21539
rect 30665 21505 30699 21539
rect 30849 21505 30883 21539
rect 31677 21505 31711 21539
rect 31769 21505 31803 21539
rect 32137 21505 32171 21539
rect 35633 21505 35667 21539
rect 35817 21505 35851 21539
rect 35909 21505 35943 21539
rect 36185 21505 36219 21539
rect 36461 21505 36495 21539
rect 36737 21505 36771 21539
rect 36829 21505 36863 21539
rect 2697 21437 2731 21471
rect 2973 21437 3007 21471
rect 4445 21437 4479 21471
rect 6653 21437 6687 21471
rect 8493 21437 8527 21471
rect 8769 21437 8803 21471
rect 17325 21437 17359 21471
rect 18889 21437 18923 21471
rect 18981 21437 19015 21471
rect 21189 21437 21223 21471
rect 23673 21437 23707 21471
rect 26617 21437 26651 21471
rect 26985 21437 27019 21471
rect 27261 21437 27295 21471
rect 29377 21437 29411 21471
rect 29469 21437 29503 21471
rect 32413 21437 32447 21471
rect 34161 21437 34195 21471
rect 10425 21369 10459 21403
rect 14013 21369 14047 21403
rect 17785 21369 17819 21403
rect 22661 21369 22695 21403
rect 23765 21369 23799 21403
rect 26249 21369 26283 21403
rect 35633 21369 35667 21403
rect 5917 21301 5951 21335
rect 11713 21301 11747 21335
rect 18061 21301 18095 21335
rect 18613 21301 18647 21335
rect 21281 21301 21315 21335
rect 23489 21301 23523 21335
rect 28733 21301 28767 21335
rect 28917 21301 28951 21335
rect 30757 21301 30791 21335
rect 31125 21301 31159 21335
rect 31309 21301 31343 21335
rect 31401 21301 31435 21335
rect 4537 21097 4571 21131
rect 6285 21097 6319 21131
rect 7849 21097 7883 21131
rect 10609 21097 10643 21131
rect 10793 21097 10827 21131
rect 13369 21097 13403 21131
rect 28089 21097 28123 21131
rect 28273 21097 28307 21131
rect 29929 21097 29963 21131
rect 7113 21029 7147 21063
rect 27721 21029 27755 21063
rect 6469 20961 6503 20995
rect 6837 20961 6871 20995
rect 7481 20961 7515 20995
rect 9965 20961 9999 20995
rect 12173 20961 12207 20995
rect 12265 20961 12299 20995
rect 12541 20961 12575 20995
rect 12817 20961 12851 20995
rect 16037 20961 16071 20995
rect 17233 20961 17267 20995
rect 24685 20961 24719 20995
rect 29561 20961 29595 20995
rect 31953 20961 31987 20995
rect 34713 20961 34747 20995
rect 35541 20961 35575 20995
rect 4721 20893 4755 20927
rect 5733 20893 5767 20927
rect 6561 20893 6595 20927
rect 6929 20893 6963 20927
rect 7113 20893 7147 20927
rect 7297 20893 7331 20927
rect 7665 20893 7699 20927
rect 9689 20893 9723 20927
rect 10425 20893 10459 20927
rect 10517 20893 10551 20927
rect 12909 20893 12943 20927
rect 16405 20893 16439 20927
rect 16773 20893 16807 20927
rect 16957 20893 16991 20927
rect 19533 20893 19567 20927
rect 19809 20893 19843 20927
rect 19993 20893 20027 20927
rect 24869 20893 24903 20927
rect 27077 20893 27111 20927
rect 27261 20893 27295 20927
rect 28733 20893 28767 20927
rect 29009 20893 29043 20927
rect 29745 20893 29779 20927
rect 30757 20893 30791 20927
rect 30941 20893 30975 20927
rect 31033 20893 31067 20927
rect 31401 20893 31435 20927
rect 31677 20893 31711 20927
rect 32045 20893 32079 20927
rect 35173 20893 35207 20927
rect 35455 20893 35489 20927
rect 35633 20893 35667 20927
rect 35731 20893 35765 20927
rect 35903 20893 35937 20927
rect 36001 20893 36035 20927
rect 36185 20893 36219 20927
rect 40693 20893 40727 20927
rect 5825 20825 5859 20859
rect 13093 20825 13127 20859
rect 15853 20825 15887 20859
rect 28089 20825 28123 20859
rect 31309 20825 31343 20859
rect 38393 20825 38427 20859
rect 38853 20825 38887 20859
rect 39037 20825 39071 20859
rect 6745 20757 6779 20791
rect 19717 20757 19751 20791
rect 19901 20757 19935 20791
rect 25053 20757 25087 20791
rect 27169 20757 27203 20791
rect 28549 20757 28583 20791
rect 28917 20757 28951 20791
rect 30849 20757 30883 20791
rect 32413 20757 32447 20791
rect 34989 20757 35023 20791
rect 35081 20757 35115 20791
rect 35817 20757 35851 20791
rect 36093 20757 36127 20791
rect 38485 20757 38519 20791
rect 39221 20757 39255 20791
rect 40969 20757 41003 20791
rect 15025 20553 15059 20587
rect 19441 20553 19475 20587
rect 22201 20553 22235 20587
rect 22661 20553 22695 20587
rect 25973 20553 26007 20587
rect 26157 20553 26191 20587
rect 32781 20553 32815 20587
rect 36185 20553 36219 20587
rect 5089 20485 5123 20519
rect 13001 20485 13035 20519
rect 14657 20485 14691 20519
rect 17141 20485 17175 20519
rect 17417 20485 17451 20519
rect 21005 20485 21039 20519
rect 21833 20485 21867 20519
rect 22109 20485 22143 20519
rect 22477 20485 22511 20519
rect 25145 20485 25179 20519
rect 28549 20485 28583 20519
rect 30297 20485 30331 20519
rect 40417 20485 40451 20519
rect 4905 20417 4939 20451
rect 5365 20417 5399 20451
rect 5549 20417 5583 20451
rect 12173 20417 12207 20451
rect 12265 20417 12299 20451
rect 12357 20417 12391 20451
rect 12725 20417 12759 20451
rect 13277 20417 13311 20451
rect 13461 20417 13495 20451
rect 14473 20417 14507 20451
rect 14749 20417 14783 20451
rect 14841 20417 14875 20451
rect 15025 20417 15059 20451
rect 16129 20417 16163 20451
rect 16957 20417 16991 20451
rect 17233 20417 17267 20451
rect 17325 20417 17359 20451
rect 17693 20417 17727 20451
rect 19073 20417 19107 20451
rect 19349 20417 19383 20451
rect 19533 20417 19567 20451
rect 19809 20417 19843 20451
rect 20177 20417 20211 20451
rect 20269 20417 20303 20451
rect 20361 20417 20395 20451
rect 20545 20417 20579 20451
rect 21373 20417 21407 20451
rect 22017 20417 22051 20451
rect 22385 20417 22419 20451
rect 23029 20417 23063 20451
rect 26098 20417 26132 20451
rect 26525 20417 26559 20451
rect 28273 20417 28307 20451
rect 32137 20417 32171 20451
rect 32230 20417 32264 20451
rect 32413 20417 32447 20451
rect 32505 20417 32539 20451
rect 32602 20417 32636 20451
rect 33333 20417 33367 20451
rect 36369 20417 36403 20451
rect 36461 20417 36495 20451
rect 36553 20417 36587 20451
rect 36737 20417 36771 20451
rect 36829 20417 36863 20451
rect 37289 20417 37323 20451
rect 37473 20417 37507 20451
rect 37565 20417 37599 20451
rect 37933 20417 37967 20451
rect 12449 20349 12483 20383
rect 15393 20349 15427 20383
rect 16221 20349 16255 20383
rect 16313 20349 16347 20383
rect 16405 20349 16439 20383
rect 17969 20349 18003 20383
rect 19717 20349 19751 20383
rect 26617 20349 26651 20383
rect 33609 20349 33643 20383
rect 35357 20349 35391 20383
rect 35449 20349 35483 20383
rect 37841 20349 37875 20383
rect 38393 20349 38427 20383
rect 38669 20349 38703 20383
rect 5365 20281 5399 20315
rect 11989 20281 12023 20315
rect 37289 20281 37323 20315
rect 5273 20213 5307 20247
rect 13277 20213 13311 20247
rect 14289 20213 14323 20247
rect 15945 20213 15979 20247
rect 16773 20213 16807 20247
rect 19901 20213 19935 20247
rect 22661 20213 22695 20247
rect 22845 20213 22879 20247
rect 23213 20213 23247 20247
rect 25421 20213 25455 20247
rect 36093 20213 36127 20247
rect 38301 20213 38335 20247
rect 6653 20009 6687 20043
rect 11345 20009 11379 20043
rect 12081 20009 12115 20043
rect 16405 20009 16439 20043
rect 16497 20009 16531 20043
rect 21189 20009 21223 20043
rect 23673 20009 23707 20043
rect 25375 20009 25409 20043
rect 27537 20009 27571 20043
rect 31493 20009 31527 20043
rect 34161 20009 34195 20043
rect 35725 20009 35759 20043
rect 36185 20009 36219 20043
rect 36645 20009 36679 20043
rect 38301 20009 38335 20043
rect 13645 19941 13679 19975
rect 23765 19941 23799 19975
rect 39037 19941 39071 19975
rect 7113 19873 7147 19907
rect 7849 19873 7883 19907
rect 14105 19873 14139 19907
rect 14289 19873 14323 19907
rect 14933 19873 14967 19907
rect 19625 19873 19659 19907
rect 19717 19873 19751 19907
rect 21005 19873 21039 19907
rect 21741 19873 21775 19907
rect 25789 19873 25823 19907
rect 34713 19873 34747 19907
rect 35173 19873 35207 19907
rect 36277 19873 36311 19907
rect 38485 19873 38519 19907
rect 38577 19873 38611 19907
rect 4445 19805 4479 19839
rect 4905 19805 4939 19839
rect 6561 19805 6595 19839
rect 6745 19805 6779 19839
rect 7021 19805 7055 19839
rect 7205 19805 7239 19839
rect 7297 19805 7331 19839
rect 7481 19805 7515 19839
rect 10333 19805 10367 19839
rect 10517 19805 10551 19839
rect 12541 19805 12575 19839
rect 12817 19805 12851 19839
rect 13645 19805 13679 19839
rect 13829 19805 13863 19839
rect 13921 19805 13955 19839
rect 14565 19805 14599 19839
rect 16589 19805 16623 19839
rect 16681 19805 16715 19839
rect 17509 19805 17543 19839
rect 17601 19805 17635 19839
rect 17785 19805 17819 19839
rect 17877 19805 17911 19839
rect 18153 19805 18187 19839
rect 19809 19805 19843 19839
rect 19901 19805 19935 19839
rect 20085 19805 20119 19839
rect 21465 19805 21499 19839
rect 22109 19805 22143 19839
rect 22569 19805 22603 19839
rect 23489 19805 23523 19839
rect 24593 19805 24627 19839
rect 24895 19805 24929 19839
rect 25053 19805 25087 19839
rect 25237 19805 25271 19839
rect 25513 19805 25547 19839
rect 25697 19805 25731 19839
rect 31401 19805 31435 19839
rect 33517 19805 33551 19839
rect 33665 19805 33699 19839
rect 33982 19805 34016 19839
rect 34897 19805 34931 19839
rect 35081 19805 35115 19839
rect 35357 19805 35391 19839
rect 35541 19805 35575 19839
rect 36001 19805 36035 19839
rect 36461 19805 36495 19839
rect 38669 19805 38703 19839
rect 38761 19805 38795 19839
rect 38945 19805 38979 19839
rect 39129 19805 39163 19839
rect 1501 19737 1535 19771
rect 1685 19737 1719 19771
rect 7665 19737 7699 19771
rect 11161 19737 11195 19771
rect 11345 19737 11379 19771
rect 11805 19737 11839 19771
rect 12357 19737 12391 19771
rect 12725 19737 12759 19771
rect 16221 19737 16255 19771
rect 16773 19737 16807 19771
rect 23857 19737 23891 19771
rect 24685 19737 24719 19771
rect 24777 19737 24811 19771
rect 25605 19737 25639 19771
rect 26065 19737 26099 19771
rect 33793 19737 33827 19771
rect 33885 19737 33919 19771
rect 35817 19737 35851 19771
rect 4721 19669 4755 19703
rect 4813 19669 4847 19703
rect 6837 19669 6871 19703
rect 10425 19669 10459 19703
rect 11529 19669 11563 19703
rect 14381 19669 14415 19703
rect 17325 19669 17359 19703
rect 17969 19669 18003 19703
rect 19441 19669 19475 19703
rect 20177 19669 20211 19703
rect 21373 19669 21407 19703
rect 22671 19669 22705 19703
rect 23581 19669 23615 19703
rect 24409 19669 24443 19703
rect 4537 19465 4571 19499
rect 5365 19465 5399 19499
rect 7021 19465 7055 19499
rect 11187 19465 11221 19499
rect 17325 19465 17359 19499
rect 17693 19465 17727 19499
rect 26065 19465 26099 19499
rect 9689 19397 9723 19431
rect 10977 19397 11011 19431
rect 11529 19397 11563 19431
rect 11713 19397 11747 19431
rect 14105 19397 14139 19431
rect 14473 19397 14507 19431
rect 14749 19397 14783 19431
rect 14933 19397 14967 19431
rect 17509 19397 17543 19431
rect 25421 19397 25455 19431
rect 27445 19397 27479 19431
rect 33885 19397 33919 19431
rect 3893 19329 3927 19363
rect 4077 19329 4111 19363
rect 4445 19329 4479 19363
rect 4629 19329 4663 19363
rect 4905 19329 4939 19363
rect 4997 19329 5031 19363
rect 6469 19329 6503 19363
rect 6653 19329 6687 19363
rect 6959 19329 6993 19363
rect 8309 19329 8343 19363
rect 8769 19329 8803 19363
rect 8953 19329 8987 19363
rect 9321 19329 9355 19363
rect 9597 19329 9631 19363
rect 9781 19329 9815 19363
rect 10241 19329 10275 19363
rect 10425 19329 10459 19363
rect 10609 19329 10643 19363
rect 10793 19329 10827 19363
rect 12633 19329 12667 19363
rect 12817 19329 12851 19363
rect 13001 19329 13035 19363
rect 14289 19329 14323 19363
rect 14381 19329 14415 19363
rect 16957 19329 16991 19363
rect 17417 19329 17451 19363
rect 17785 19329 17819 19363
rect 19533 19329 19567 19363
rect 20177 19329 20211 19363
rect 20269 19329 20303 19363
rect 20637 19329 20671 19363
rect 21833 19329 21867 19363
rect 22017 19329 22051 19363
rect 22293 19329 22327 19363
rect 23029 19329 23063 19363
rect 23305 19329 23339 19363
rect 25789 19329 25823 19363
rect 25881 19329 25915 19363
rect 27353 19329 27387 19363
rect 29929 19329 29963 19363
rect 32137 19329 32171 19363
rect 4813 19261 4847 19295
rect 7481 19261 7515 19295
rect 8401 19261 8435 19295
rect 8585 19261 8619 19295
rect 9045 19261 9079 19295
rect 9137 19261 9171 19295
rect 17049 19261 17083 19295
rect 17141 19261 17175 19295
rect 20913 19261 20947 19295
rect 27537 19261 27571 19295
rect 30205 19261 30239 19295
rect 5549 19193 5583 19227
rect 6561 19193 6595 19227
rect 7389 19193 7423 19227
rect 9505 19193 9539 19227
rect 22569 19193 22603 19227
rect 3893 19125 3927 19159
rect 4169 19125 4203 19159
rect 5365 19125 5399 19159
rect 6837 19125 6871 19159
rect 7941 19125 7975 19159
rect 10333 19125 10367 19159
rect 10609 19125 10643 19159
rect 11161 19125 11195 19159
rect 11345 19125 11379 19159
rect 11713 19125 11747 19159
rect 11897 19125 11931 19159
rect 14657 19125 14691 19159
rect 15117 19125 15151 19159
rect 16681 19125 16715 19159
rect 17509 19125 17543 19159
rect 22201 19125 22235 19159
rect 25789 19125 25823 19159
rect 26985 19125 27019 19159
rect 31677 19125 31711 19159
rect 32229 19125 32263 19159
rect 34161 19125 34195 19159
rect 10241 18921 10275 18955
rect 17417 18921 17451 18955
rect 18705 18921 18739 18955
rect 19901 18921 19935 18955
rect 23029 18921 23063 18955
rect 29285 18921 29319 18955
rect 33517 18921 33551 18955
rect 35357 18921 35391 18955
rect 36645 18921 36679 18955
rect 6285 18853 6319 18887
rect 9781 18853 9815 18887
rect 38853 18853 38887 18887
rect 4537 18785 4571 18819
rect 4905 18785 4939 18819
rect 5181 18785 5215 18819
rect 5365 18785 5399 18819
rect 7849 18785 7883 18819
rect 16405 18785 16439 18819
rect 16589 18785 16623 18819
rect 16681 18785 16715 18819
rect 16773 18785 16807 18819
rect 18797 18785 18831 18819
rect 25145 18785 25179 18819
rect 27537 18785 27571 18819
rect 30205 18785 30239 18819
rect 33241 18785 33275 18819
rect 33609 18785 33643 18819
rect 37289 18785 37323 18819
rect 39497 18785 39531 18819
rect 4353 18717 4387 18751
rect 4997 18717 5031 18751
rect 5089 18717 5123 18751
rect 5549 18717 5583 18751
rect 5825 18717 5859 18751
rect 7113 18717 7147 18751
rect 7389 18717 7423 18751
rect 7665 18717 7699 18751
rect 7941 18717 7975 18751
rect 8493 18717 8527 18751
rect 8585 18717 8619 18751
rect 8953 18717 8987 18751
rect 9229 18717 9263 18751
rect 9413 18717 9447 18751
rect 9873 18717 9907 18751
rect 10057 18717 10091 18751
rect 12449 18717 12483 18751
rect 12633 18717 12667 18751
rect 14289 18717 14323 18751
rect 14749 18717 14783 18751
rect 14933 18717 14967 18751
rect 16129 18717 16163 18751
rect 16865 18717 16899 18751
rect 17141 18717 17175 18751
rect 17601 18717 17635 18751
rect 18521 18717 18555 18751
rect 19809 18717 19843 18751
rect 22201 18717 22235 18751
rect 22385 18717 22419 18751
rect 22845 18717 22879 18751
rect 23213 18717 23247 18751
rect 23765 18717 23799 18751
rect 23949 18717 23983 18751
rect 24225 18717 24259 18751
rect 24593 18717 24627 18751
rect 24685 18717 24719 18751
rect 25053 18717 25087 18751
rect 25329 18717 25363 18751
rect 27445 18717 27479 18751
rect 29929 18717 29963 18751
rect 31309 18717 31343 18751
rect 32045 18717 32079 18751
rect 32229 18717 32263 18751
rect 33149 18717 33183 18751
rect 33793 18717 33827 18751
rect 33977 18717 34011 18751
rect 35265 18717 35299 18751
rect 35449 18717 35483 18751
rect 36829 18717 36863 18751
rect 40049 18717 40083 18751
rect 4261 18649 4295 18683
rect 6469 18649 6503 18683
rect 6571 18649 6605 18683
rect 6837 18649 6871 18683
rect 6929 18649 6963 18683
rect 7481 18649 7515 18683
rect 9321 18649 9355 18683
rect 9597 18649 9631 18683
rect 12725 18649 12759 18683
rect 23857 18649 23891 18683
rect 24087 18649 24121 18683
rect 24777 18649 24811 18683
rect 24915 18649 24949 18683
rect 27813 18649 27847 18683
rect 36921 18649 36955 18683
rect 37013 18649 37047 18683
rect 37131 18649 37165 18683
rect 39313 18649 39347 18683
rect 3893 18581 3927 18615
rect 4721 18581 4755 18615
rect 5733 18581 5767 18615
rect 6653 18581 6687 18615
rect 7297 18581 7331 18615
rect 15577 18581 15611 18615
rect 16313 18581 16347 18615
rect 17785 18581 17819 18615
rect 18337 18581 18371 18615
rect 22385 18581 22419 18615
rect 23305 18581 23339 18615
rect 23581 18581 23615 18615
rect 24409 18581 24443 18615
rect 25513 18581 25547 18615
rect 27261 18581 27295 18615
rect 29561 18581 29595 18615
rect 30021 18581 30055 18615
rect 31585 18581 31619 18615
rect 32045 18581 32079 18615
rect 39221 18581 39255 18615
rect 39865 18581 39899 18615
rect 3157 18377 3191 18411
rect 5825 18377 5859 18411
rect 7205 18377 7239 18411
rect 11989 18377 12023 18411
rect 12633 18377 12667 18411
rect 22937 18377 22971 18411
rect 24041 18377 24075 18411
rect 29929 18377 29963 18411
rect 31585 18377 31619 18411
rect 33517 18377 33551 18411
rect 34161 18377 34195 18411
rect 35005 18377 35039 18411
rect 35173 18377 35207 18411
rect 36645 18377 36679 18411
rect 37105 18377 37139 18411
rect 37841 18377 37875 18411
rect 38761 18377 38795 18411
rect 40969 18377 41003 18411
rect 5457 18309 5491 18343
rect 5657 18309 5691 18343
rect 14841 18309 14875 18343
rect 27905 18309 27939 18343
rect 32229 18309 32263 18343
rect 33149 18309 33183 18343
rect 33365 18309 33399 18343
rect 33701 18309 33735 18343
rect 34805 18309 34839 18343
rect 36921 18309 36955 18343
rect 39497 18309 39531 18343
rect 1409 18241 1443 18275
rect 4721 18241 4755 18275
rect 4997 18241 5031 18275
rect 5365 18241 5399 18275
rect 7113 18241 7147 18275
rect 7297 18241 7331 18275
rect 10517 18241 10551 18275
rect 10977 18241 11011 18275
rect 11529 18241 11563 18275
rect 12173 18241 12207 18275
rect 12357 18241 12391 18275
rect 12449 18241 12483 18275
rect 12541 18241 12575 18275
rect 12725 18241 12759 18275
rect 15301 18241 15335 18275
rect 15577 18241 15611 18275
rect 15761 18241 15795 18275
rect 16681 18241 16715 18275
rect 17049 18241 17083 18275
rect 17693 18241 17727 18275
rect 17785 18241 17819 18275
rect 18245 18241 18279 18275
rect 18429 18241 18463 18275
rect 18521 18241 18555 18275
rect 18613 18241 18647 18275
rect 19073 18241 19107 18275
rect 19165 18241 19199 18275
rect 19257 18241 19291 18275
rect 19993 18241 20027 18275
rect 20177 18241 20211 18275
rect 20269 18241 20303 18275
rect 20453 18241 20487 18275
rect 20637 18241 20671 18275
rect 23029 18241 23063 18275
rect 23765 18241 23799 18275
rect 24133 18241 24167 18275
rect 24409 18241 24443 18275
rect 26985 18241 27019 18275
rect 27078 18241 27112 18275
rect 27261 18241 27295 18275
rect 27353 18241 27387 18275
rect 27491 18241 27525 18275
rect 27721 18241 27755 18275
rect 27997 18241 28031 18275
rect 28089 18241 28123 18275
rect 29561 18241 29595 18275
rect 31493 18241 31527 18275
rect 31677 18241 31711 18275
rect 33609 18241 33643 18275
rect 33793 18241 33827 18275
rect 33885 18241 33919 18275
rect 36461 18241 36495 18275
rect 36645 18241 36679 18275
rect 36737 18241 36771 18275
rect 37473 18241 37507 18275
rect 39221 18241 39255 18275
rect 1685 18173 1719 18207
rect 5089 18173 5123 18207
rect 10609 18173 10643 18207
rect 20821 18173 20855 18207
rect 23673 18173 23707 18207
rect 24225 18173 24259 18207
rect 29469 18173 29503 18207
rect 34161 18173 34195 18207
rect 37565 18173 37599 18207
rect 38853 18173 38887 18207
rect 39037 18173 39071 18207
rect 15117 18105 15151 18139
rect 15577 18105 15611 18139
rect 18061 18105 18095 18139
rect 18889 18105 18923 18139
rect 22569 18105 22603 18139
rect 22661 18105 22695 18139
rect 23857 18105 23891 18139
rect 24593 18105 24627 18139
rect 28273 18105 28307 18139
rect 38393 18105 38427 18139
rect 5641 18037 5675 18071
rect 11161 18037 11195 18071
rect 11713 18037 11747 18071
rect 15945 18037 15979 18071
rect 18797 18037 18831 18071
rect 19441 18037 19475 18071
rect 20269 18037 20303 18071
rect 22293 18037 22327 18071
rect 22753 18037 22787 18071
rect 23397 18037 23431 18071
rect 27629 18037 27663 18071
rect 32321 18037 32355 18071
rect 33333 18037 33367 18071
rect 33977 18037 34011 18071
rect 34989 18037 35023 18071
rect 2697 17833 2731 17867
rect 9413 17833 9447 17867
rect 10149 17833 10183 17867
rect 12817 17833 12851 17867
rect 22385 17833 22419 17867
rect 30941 17833 30975 17867
rect 35541 17833 35575 17867
rect 39589 17833 39623 17867
rect 4261 17765 4295 17799
rect 36829 17765 36863 17799
rect 1961 17697 1995 17731
rect 13461 17697 13495 17731
rect 20085 17697 20119 17731
rect 30757 17697 30791 17731
rect 35909 17697 35943 17731
rect 36553 17697 36587 17731
rect 2881 17629 2915 17663
rect 3157 17629 3191 17663
rect 4445 17629 4479 17663
rect 4721 17629 4755 17663
rect 5365 17629 5399 17663
rect 5549 17629 5583 17663
rect 5825 17629 5859 17663
rect 9321 17629 9355 17663
rect 9505 17629 9539 17663
rect 10057 17629 10091 17663
rect 10241 17629 10275 17663
rect 11345 17629 11379 17663
rect 11621 17629 11655 17663
rect 11713 17629 11747 17663
rect 11897 17629 11931 17663
rect 13645 17629 13679 17663
rect 14105 17629 14139 17663
rect 14657 17629 14691 17663
rect 15117 17629 15151 17663
rect 15393 17629 15427 17663
rect 18245 17629 18279 17663
rect 18337 17629 18371 17663
rect 18521 17629 18555 17663
rect 20177 17629 20211 17663
rect 22569 17629 22603 17663
rect 22661 17629 22695 17663
rect 22753 17629 22787 17663
rect 22871 17629 22905 17663
rect 23029 17629 23063 17663
rect 26893 17629 26927 17663
rect 26985 17629 27019 17663
rect 27169 17629 27203 17663
rect 27261 17629 27295 17663
rect 30665 17629 30699 17663
rect 31125 17629 31159 17663
rect 31309 17629 31343 17663
rect 31585 17629 31619 17663
rect 35817 17629 35851 17663
rect 36461 17629 36495 17663
rect 36921 17629 36955 17663
rect 37105 17629 37139 17663
rect 2605 17561 2639 17595
rect 3065 17561 3099 17595
rect 11161 17561 11195 17595
rect 11805 17561 11839 17595
rect 13185 17561 13219 17595
rect 13737 17561 13771 17595
rect 15945 17561 15979 17595
rect 34989 17561 35023 17595
rect 35265 17561 35299 17595
rect 35357 17561 35391 17595
rect 39221 17561 39255 17595
rect 39405 17561 39439 17595
rect 40693 17561 40727 17595
rect 11529 17493 11563 17527
rect 13277 17493 13311 17527
rect 14197 17493 14231 17527
rect 18705 17493 18739 17527
rect 20545 17493 20579 17527
rect 26709 17493 26743 17527
rect 31493 17493 31527 17527
rect 35173 17493 35207 17527
rect 36185 17493 36219 17527
rect 37105 17493 37139 17527
rect 40969 17493 41003 17527
rect 5457 17289 5491 17323
rect 6745 17289 6779 17323
rect 12541 17289 12575 17323
rect 12909 17289 12943 17323
rect 15485 17289 15519 17323
rect 15669 17289 15703 17323
rect 30113 17289 30147 17323
rect 30665 17289 30699 17323
rect 30941 17289 30975 17323
rect 33149 17289 33183 17323
rect 39405 17289 39439 17323
rect 8493 17221 8527 17255
rect 8953 17221 8987 17255
rect 9413 17221 9447 17255
rect 11529 17221 11563 17255
rect 13001 17221 13035 17255
rect 20729 17221 20763 17255
rect 20913 17221 20947 17255
rect 26525 17221 26559 17255
rect 29929 17221 29963 17255
rect 38761 17221 38795 17255
rect 39218 17221 39252 17255
rect 38991 17187 39025 17221
rect 4629 17153 4663 17187
rect 4813 17153 4847 17187
rect 5089 17153 5123 17187
rect 5273 17153 5307 17187
rect 6929 17153 6963 17187
rect 7849 17153 7883 17187
rect 8033 17153 8067 17187
rect 8217 17153 8251 17187
rect 8309 17153 8343 17187
rect 8861 17153 8895 17187
rect 9045 17153 9079 17187
rect 9163 17153 9197 17187
rect 9597 17153 9631 17187
rect 11713 17153 11747 17187
rect 14841 17153 14875 17187
rect 14934 17153 14968 17187
rect 15117 17153 15151 17187
rect 15209 17153 15243 17187
rect 15306 17153 15340 17187
rect 16129 17153 16163 17187
rect 18061 17153 18095 17187
rect 18337 17153 18371 17187
rect 18521 17153 18555 17187
rect 18797 17153 18831 17187
rect 20085 17153 20119 17187
rect 20269 17153 20303 17187
rect 20453 17153 20487 17187
rect 23121 17153 23155 17187
rect 23305 17153 23339 17187
rect 24041 17153 24075 17187
rect 24225 17153 24259 17187
rect 24317 17153 24351 17187
rect 24777 17153 24811 17187
rect 24961 17153 24995 17187
rect 25053 17153 25087 17187
rect 25329 17153 25363 17187
rect 26433 17153 26467 17187
rect 30389 17153 30423 17187
rect 30665 17153 30699 17187
rect 30849 17153 30883 17187
rect 31033 17153 31067 17187
rect 33425 17153 33459 17187
rect 38485 17153 38519 17187
rect 38669 17153 38703 17187
rect 39497 17153 39531 17187
rect 4721 17085 4755 17119
rect 4905 17085 4939 17119
rect 7205 17085 7239 17119
rect 9321 17085 9355 17119
rect 13185 17085 13219 17119
rect 15853 17085 15887 17119
rect 18613 17085 18647 17119
rect 18981 17085 19015 17119
rect 25145 17085 25179 17119
rect 33333 17085 33367 17119
rect 33517 17085 33551 17119
rect 33609 17085 33643 17119
rect 40509 17085 40543 17119
rect 16037 17017 16071 17051
rect 18337 17017 18371 17051
rect 24317 17017 24351 17051
rect 29561 17017 29595 17051
rect 38577 17017 38611 17051
rect 39129 17017 39163 17051
rect 4445 16949 4479 16983
rect 7113 16949 7147 16983
rect 7941 16949 7975 16983
rect 8677 16949 8711 16983
rect 9781 16949 9815 16983
rect 11897 16949 11931 16983
rect 20913 16949 20947 16983
rect 21097 16949 21131 16983
rect 23489 16949 23523 16983
rect 25513 16949 25547 16983
rect 29929 16949 29963 16983
rect 38945 16949 38979 16983
rect 39221 16949 39255 16983
rect 41061 16949 41095 16983
rect 9137 16745 9171 16779
rect 9413 16745 9447 16779
rect 15393 16745 15427 16779
rect 17785 16745 17819 16779
rect 23581 16745 23615 16779
rect 30757 16745 30791 16779
rect 30941 16745 30975 16779
rect 33241 16745 33275 16779
rect 39221 16745 39255 16779
rect 5365 16677 5399 16711
rect 7941 16677 7975 16711
rect 8401 16677 8435 16711
rect 29745 16677 29779 16711
rect 30481 16677 30515 16711
rect 33057 16677 33091 16711
rect 4721 16609 4755 16643
rect 8033 16609 8067 16643
rect 11897 16609 11931 16643
rect 13093 16609 13127 16643
rect 16681 16609 16715 16643
rect 17233 16609 17267 16643
rect 20545 16609 20579 16643
rect 21741 16609 21775 16643
rect 25605 16609 25639 16643
rect 25697 16609 25731 16643
rect 26801 16609 26835 16643
rect 27445 16609 27479 16643
rect 28733 16609 28767 16643
rect 29009 16609 29043 16643
rect 29101 16609 29135 16643
rect 30205 16609 30239 16643
rect 31033 16609 31067 16643
rect 31401 16609 31435 16643
rect 33517 16609 33551 16643
rect 40509 16609 40543 16643
rect 40601 16609 40635 16643
rect 29285 16575 29319 16609
rect 4077 16541 4111 16575
rect 4169 16541 4203 16575
rect 4261 16541 4295 16575
rect 4445 16541 4479 16575
rect 4905 16541 4939 16575
rect 5089 16541 5123 16575
rect 5457 16541 5491 16575
rect 5547 16519 5581 16553
rect 7849 16541 7883 16575
rect 8125 16541 8159 16575
rect 8309 16541 8343 16575
rect 8401 16541 8435 16575
rect 8585 16541 8619 16575
rect 8953 16541 8987 16575
rect 9321 16541 9355 16575
rect 9505 16541 9539 16575
rect 11437 16541 11471 16575
rect 11529 16541 11563 16575
rect 11621 16541 11655 16575
rect 11805 16541 11839 16575
rect 12081 16541 12115 16575
rect 12173 16541 12207 16575
rect 12357 16541 12391 16575
rect 12449 16541 12483 16575
rect 12909 16541 12943 16575
rect 15577 16541 15611 16575
rect 15669 16541 15703 16575
rect 15853 16541 15887 16575
rect 15945 16541 15979 16575
rect 16037 16541 16071 16575
rect 16221 16541 16255 16575
rect 16313 16541 16347 16575
rect 16405 16541 16439 16575
rect 16957 16541 16991 16575
rect 17509 16541 17543 16575
rect 19901 16541 19935 16575
rect 20085 16541 20119 16575
rect 20269 16541 20303 16575
rect 20821 16541 20855 16575
rect 21189 16541 21223 16575
rect 21281 16541 21315 16575
rect 21465 16541 21499 16575
rect 21925 16541 21959 16575
rect 22385 16541 22419 16575
rect 22569 16541 22603 16575
rect 23305 16541 23339 16575
rect 23398 16541 23432 16575
rect 23673 16541 23707 16575
rect 26157 16541 26191 16575
rect 26525 16541 26559 16575
rect 27537 16541 27571 16575
rect 27721 16541 27755 16575
rect 28457 16541 28491 16575
rect 28552 16541 28586 16575
rect 29193 16541 29227 16575
rect 31217 16541 31251 16575
rect 31493 16541 31527 16575
rect 32321 16541 32355 16575
rect 32781 16541 32815 16575
rect 32965 16541 32999 16575
rect 33149 16541 33183 16575
rect 33413 16541 33447 16575
rect 33885 16541 33919 16575
rect 34253 16541 34287 16575
rect 34437 16541 34471 16575
rect 35909 16541 35943 16575
rect 37749 16541 37783 16575
rect 38577 16541 38611 16575
rect 38853 16541 38887 16575
rect 38945 16541 38979 16575
rect 39129 16541 39163 16575
rect 39221 16541 39255 16575
rect 39405 16541 39439 16575
rect 39681 16541 39715 16575
rect 40417 16541 40451 16575
rect 30803 16507 30837 16541
rect 5181 16473 5215 16507
rect 5273 16473 5307 16507
rect 16523 16473 16557 16507
rect 17141 16473 17175 16507
rect 20453 16473 20487 16507
rect 20913 16473 20947 16507
rect 22201 16473 22235 16507
rect 28181 16473 28215 16507
rect 29745 16473 29779 16507
rect 30573 16473 30607 16507
rect 32413 16473 32447 16507
rect 38761 16473 38795 16507
rect 3801 16405 3835 16439
rect 7665 16405 7699 16439
rect 11161 16405 11195 16439
rect 12541 16405 12575 16439
rect 13001 16405 13035 16439
rect 17969 16405 18003 16439
rect 21005 16405 21039 16439
rect 23121 16405 23155 16439
rect 25145 16405 25179 16439
rect 25513 16405 25547 16439
rect 26065 16405 26099 16439
rect 28825 16405 28859 16439
rect 30297 16405 30331 16439
rect 31677 16405 31711 16439
rect 33609 16405 33643 16439
rect 33793 16405 33827 16439
rect 34437 16405 34471 16439
rect 36001 16405 36035 16439
rect 37933 16405 37967 16439
rect 38675 16405 38709 16439
rect 39037 16405 39071 16439
rect 39497 16405 39531 16439
rect 40049 16405 40083 16439
rect 5273 16201 5307 16235
rect 7389 16201 7423 16235
rect 9413 16201 9447 16235
rect 11897 16201 11931 16235
rect 15761 16201 15795 16235
rect 17049 16201 17083 16235
rect 18337 16201 18371 16235
rect 20637 16201 20671 16235
rect 26709 16201 26743 16235
rect 41061 16201 41095 16235
rect 5089 16133 5123 16167
rect 6009 16133 6043 16167
rect 15393 16133 15427 16167
rect 20729 16133 20763 16167
rect 21189 16133 21223 16167
rect 23305 16133 23339 16167
rect 23521 16133 23555 16167
rect 24501 16133 24535 16167
rect 24685 16133 24719 16167
rect 26433 16133 26467 16167
rect 27353 16133 27387 16167
rect 28917 16133 28951 16167
rect 29377 16133 29411 16167
rect 36921 16133 36955 16167
rect 39589 16133 39623 16167
rect 1409 16065 1443 16099
rect 3801 16065 3835 16099
rect 3893 16065 3927 16099
rect 4077 16065 4111 16099
rect 4169 16065 4203 16099
rect 4261 16065 4295 16099
rect 5273 16065 5307 16099
rect 5365 16065 5399 16099
rect 5733 16065 5767 16099
rect 5917 16065 5951 16099
rect 6745 16065 6779 16099
rect 7205 16065 7239 16099
rect 7481 16065 7515 16099
rect 7573 16065 7607 16099
rect 9229 16065 9263 16099
rect 9413 16065 9447 16099
rect 11161 16065 11195 16099
rect 11529 16065 11563 16099
rect 11713 16065 11747 16099
rect 11989 16065 12023 16099
rect 12173 16065 12207 16099
rect 12265 16065 12299 16099
rect 12357 16065 12391 16099
rect 15209 16065 15243 16099
rect 15485 16065 15519 16099
rect 15577 16065 15611 16099
rect 16681 16065 16715 16099
rect 18153 16063 18187 16097
rect 20545 16065 20579 16099
rect 20913 16065 20947 16099
rect 21005 16065 21039 16099
rect 22845 16065 22879 16099
rect 23121 16065 23155 16099
rect 25513 16065 25547 16099
rect 25697 16065 25731 16099
rect 25881 16065 25915 16099
rect 26341 16065 26375 16099
rect 26617 16065 26651 16099
rect 26801 16065 26835 16099
rect 26985 16065 27019 16099
rect 27078 16065 27112 16099
rect 27261 16065 27295 16099
rect 27450 16065 27484 16099
rect 28825 16065 28859 16099
rect 29009 16065 29043 16099
rect 29544 16065 29578 16099
rect 29654 16065 29688 16099
rect 29929 16065 29963 16099
rect 32583 16065 32617 16099
rect 33517 16065 33551 16099
rect 33609 16065 33643 16099
rect 33885 16065 33919 16099
rect 33977 16065 34011 16099
rect 34161 16065 34195 16099
rect 34621 16065 34655 16099
rect 36461 16065 36495 16099
rect 36829 16065 36863 16099
rect 37013 16065 37047 16099
rect 37473 16065 37507 16099
rect 37749 16065 37783 16099
rect 37841 16065 37875 16099
rect 38761 16065 38795 16099
rect 3617 15997 3651 16031
rect 4537 15997 4571 16031
rect 5549 15997 5583 16031
rect 6837 15997 6871 16031
rect 7849 15997 7883 16031
rect 17969 15997 18003 16031
rect 21373 15997 21407 16031
rect 22937 15997 22971 16031
rect 23029 15997 23063 16031
rect 25605 15997 25639 16031
rect 32413 15997 32447 16031
rect 34529 15997 34563 16031
rect 37289 15997 37323 16031
rect 38577 15997 38611 16031
rect 39313 15997 39347 16031
rect 7205 15929 7239 15963
rect 7665 15929 7699 15963
rect 7757 15929 7791 15963
rect 11253 15929 11287 15963
rect 25973 15929 26007 15963
rect 29837 15929 29871 15963
rect 32873 15929 32907 15963
rect 36645 15929 36679 15963
rect 38117 15929 38151 15963
rect 1593 15861 1627 15895
rect 4629 15861 4663 15895
rect 4813 15861 4847 15895
rect 6929 15861 6963 15895
rect 7113 15861 7147 15895
rect 11989 15861 12023 15895
rect 17049 15861 17083 15895
rect 17233 15861 17267 15895
rect 20269 15861 20303 15895
rect 22661 15861 22695 15895
rect 23489 15861 23523 15895
rect 23673 15861 23707 15895
rect 24869 15861 24903 15895
rect 27629 15861 27663 15895
rect 33333 15861 33367 15895
rect 33793 15861 33827 15895
rect 33977 15861 34011 15895
rect 34989 15861 35023 15895
rect 37657 15861 37691 15895
rect 37749 15861 37783 15895
rect 38945 15861 38979 15895
rect 1593 15657 1627 15691
rect 2040 15657 2074 15691
rect 17601 15657 17635 15691
rect 17969 15657 18003 15691
rect 33425 15657 33459 15691
rect 5273 15589 5307 15623
rect 10793 15589 10827 15623
rect 18705 15589 18739 15623
rect 1777 15521 1811 15555
rect 3525 15521 3559 15555
rect 10425 15521 10459 15555
rect 20361 15521 20395 15555
rect 21281 15521 21315 15555
rect 29653 15521 29687 15555
rect 30113 15521 30147 15555
rect 1409 15453 1443 15487
rect 3985 15453 4019 15487
rect 4721 15453 4755 15487
rect 4905 15453 4939 15487
rect 5089 15453 5123 15487
rect 10977 15453 11011 15487
rect 11161 15453 11195 15487
rect 13737 15453 13771 15487
rect 14105 15453 14139 15487
rect 17601 15453 17635 15487
rect 17693 15453 17727 15487
rect 18153 15453 18187 15487
rect 18429 15453 18463 15487
rect 18521 15453 18555 15487
rect 19993 15453 20027 15487
rect 21465 15453 21499 15487
rect 21613 15453 21647 15487
rect 21741 15453 21775 15487
rect 21930 15453 21964 15487
rect 22569 15453 22603 15487
rect 22753 15453 22787 15487
rect 23029 15453 23063 15487
rect 23122 15453 23156 15487
rect 23494 15453 23528 15487
rect 24409 15453 24443 15487
rect 24557 15453 24591 15487
rect 24874 15453 24908 15487
rect 29745 15453 29779 15487
rect 33609 15453 33643 15487
rect 33885 15453 33919 15487
rect 35541 15453 35575 15487
rect 35725 15453 35759 15487
rect 4997 15385 5031 15419
rect 13829 15385 13863 15419
rect 14381 15385 14415 15419
rect 18337 15385 18371 15419
rect 20177 15385 20211 15419
rect 20453 15385 20487 15419
rect 21833 15385 21867 15419
rect 23305 15385 23339 15419
rect 23397 15385 23431 15419
rect 24685 15385 24719 15419
rect 24777 15385 24811 15419
rect 4629 15317 4663 15351
rect 10885 15317 10919 15351
rect 11345 15317 11379 15351
rect 15853 15317 15887 15351
rect 22109 15317 22143 15351
rect 22661 15317 22695 15351
rect 23673 15317 23707 15351
rect 25053 15317 25087 15351
rect 33793 15317 33827 15351
rect 35633 15317 35667 15351
rect 5549 15113 5583 15147
rect 6929 15113 6963 15147
rect 9873 15113 9907 15147
rect 11713 15113 11747 15147
rect 14105 15113 14139 15147
rect 17233 15113 17267 15147
rect 19533 15113 19567 15147
rect 22845 15113 22879 15147
rect 24409 15113 24443 15147
rect 29929 15113 29963 15147
rect 8953 15045 8987 15079
rect 9045 15045 9079 15079
rect 14473 15045 14507 15079
rect 15025 15045 15059 15079
rect 16957 15045 16991 15079
rect 27169 15045 27203 15079
rect 27261 15045 27295 15079
rect 31217 15045 31251 15079
rect 5365 14977 5399 15011
rect 6653 14977 6687 15011
rect 6745 14977 6779 15011
rect 7297 14977 7331 15011
rect 7481 14977 7515 15011
rect 8309 14977 8343 15011
rect 8861 14977 8895 15011
rect 9163 14977 9197 15011
rect 9689 14977 9723 15011
rect 9965 14977 9999 15011
rect 10241 14977 10275 15011
rect 10885 14977 10919 15011
rect 10977 14977 11011 15011
rect 11253 14977 11287 15011
rect 11529 14977 11563 15011
rect 14933 14977 14967 15011
rect 16681 14977 16715 15011
rect 16865 14977 16899 15011
rect 17049 14977 17083 15011
rect 18153 14977 18187 15011
rect 19441 14977 19475 15011
rect 19625 14977 19659 15011
rect 19717 14977 19751 15011
rect 20177 14977 20211 15011
rect 20453 14977 20487 15011
rect 20913 14977 20947 15011
rect 21649 14977 21683 15011
rect 22753 14977 22787 15011
rect 23857 14977 23891 15011
rect 24041 14977 24075 15011
rect 24133 14977 24167 15011
rect 24225 14977 24259 15011
rect 26985 14977 27019 15011
rect 27353 14977 27387 15011
rect 27629 14977 27663 15011
rect 27813 14977 27847 15011
rect 27905 14977 27939 15011
rect 27997 14977 28031 15011
rect 29745 14977 29779 15011
rect 30021 14977 30055 15011
rect 30757 14977 30791 15011
rect 31401 14977 31435 15011
rect 31493 14977 31527 15011
rect 31585 14977 31619 15011
rect 31723 14977 31757 15011
rect 35357 14977 35391 15011
rect 35541 14977 35575 15011
rect 38688 14999 38722 15033
rect 5181 14909 5215 14943
rect 8125 14909 8159 14943
rect 9321 14909 9355 14943
rect 10149 14909 10183 14943
rect 12173 14909 12207 14943
rect 12449 14909 12483 14943
rect 14565 14909 14599 14943
rect 14657 14909 14691 14943
rect 17969 14909 18003 14943
rect 30849 14909 30883 14943
rect 31861 14909 31895 14943
rect 38945 14909 38979 14943
rect 18337 14841 18371 14875
rect 19809 14841 19843 14875
rect 7389 14773 7423 14807
rect 8493 14773 8527 14807
rect 8677 14773 8711 14807
rect 9505 14773 9539 14807
rect 10609 14773 10643 14807
rect 10701 14773 10735 14807
rect 11161 14773 11195 14807
rect 13921 14773 13955 14807
rect 27537 14773 27571 14807
rect 28181 14773 28215 14807
rect 29561 14773 29595 14807
rect 31125 14773 31159 14807
rect 35449 14773 35483 14807
rect 38761 14773 38795 14807
rect 38853 14773 38887 14807
rect 3433 14569 3467 14603
rect 5641 14569 5675 14603
rect 5825 14569 5859 14603
rect 6101 14569 6135 14603
rect 9321 14569 9355 14603
rect 11161 14569 11195 14603
rect 11897 14569 11931 14603
rect 17233 14569 17267 14603
rect 27261 14569 27295 14603
rect 27353 14569 27387 14603
rect 32045 14569 32079 14603
rect 32229 14569 32263 14603
rect 35357 14569 35391 14603
rect 6561 14501 6595 14535
rect 17693 14501 17727 14535
rect 20729 14501 20763 14535
rect 27445 14501 27479 14535
rect 36185 14501 36219 14535
rect 39497 14501 39531 14535
rect 3617 14433 3651 14467
rect 3985 14433 4019 14467
rect 5549 14433 5583 14467
rect 6193 14433 6227 14467
rect 7665 14433 7699 14467
rect 12909 14433 12943 14467
rect 20545 14433 20579 14467
rect 22937 14433 22971 14467
rect 29561 14433 29595 14467
rect 29837 14433 29871 14467
rect 35173 14433 35207 14467
rect 36553 14433 36587 14467
rect 39129 14433 39163 14467
rect 39865 14433 39899 14467
rect 3341 14365 3375 14399
rect 4169 14365 4203 14399
rect 4373 14365 4407 14399
rect 4537 14365 4571 14399
rect 5457 14365 5491 14399
rect 5917 14359 5951 14393
rect 6009 14365 6043 14399
rect 6285 14365 6319 14399
rect 6469 14365 6503 14399
rect 6745 14365 6779 14399
rect 6837 14365 6871 14399
rect 7205 14365 7239 14399
rect 7757 14365 7791 14399
rect 7941 14365 7975 14399
rect 8033 14365 8067 14399
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 8585 14365 8619 14399
rect 8769 14365 8803 14399
rect 10517 14365 10551 14399
rect 10610 14365 10644 14399
rect 10982 14365 11016 14399
rect 11253 14365 11287 14399
rect 11346 14365 11380 14399
rect 11759 14365 11793 14399
rect 14841 14365 14875 14399
rect 14934 14365 14968 14399
rect 15117 14365 15151 14399
rect 15209 14365 15243 14399
rect 15306 14365 15340 14399
rect 16129 14365 16163 14399
rect 16267 14365 16301 14399
rect 16405 14365 16439 14399
rect 17055 14365 17089 14399
rect 17233 14365 17267 14399
rect 18061 14365 18095 14399
rect 18337 14365 18371 14399
rect 18429 14365 18463 14399
rect 18705 14365 18739 14399
rect 18889 14365 18923 14399
rect 20269 14365 20303 14399
rect 20913 14365 20947 14399
rect 21189 14365 21223 14399
rect 22109 14365 22143 14399
rect 22661 14365 22695 14399
rect 26341 14365 26375 14399
rect 26525 14365 26559 14399
rect 26709 14365 26743 14399
rect 27724 14365 27758 14399
rect 27813 14365 27847 14399
rect 28181 14365 28215 14399
rect 31677 14365 31711 14399
rect 32137 14365 32171 14399
rect 32321 14365 32355 14399
rect 35081 14365 35115 14399
rect 35541 14365 35575 14399
rect 35689 14365 35723 14399
rect 36047 14365 36081 14399
rect 36277 14365 36311 14399
rect 38393 14365 38427 14399
rect 38541 14365 38575 14399
rect 38669 14365 38703 14399
rect 38761 14365 38795 14399
rect 38858 14365 38892 14399
rect 39313 14365 39347 14399
rect 39405 14365 39439 14399
rect 39589 14365 39623 14399
rect 3985 14297 4019 14331
rect 4261 14297 4295 14331
rect 5181 14297 5215 14331
rect 6929 14297 6963 14331
rect 7047 14297 7081 14331
rect 7297 14297 7331 14331
rect 7481 14297 7515 14331
rect 8953 14297 8987 14331
rect 9137 14297 9171 14331
rect 10793 14297 10827 14331
rect 10885 14297 10919 14331
rect 11529 14297 11563 14331
rect 11621 14297 11655 14331
rect 13461 14297 13495 14331
rect 15577 14297 15611 14331
rect 26617 14297 26651 14331
rect 27997 14297 28031 14331
rect 28089 14297 28123 14331
rect 31585 14297 31619 14331
rect 31861 14297 31895 14331
rect 35817 14297 35851 14331
rect 35909 14297 35943 14331
rect 38301 14297 38335 14331
rect 40509 14297 40543 14331
rect 3617 14229 3651 14263
rect 6469 14229 6503 14263
rect 8677 14229 8711 14263
rect 15485 14229 15519 14263
rect 17417 14229 17451 14263
rect 21097 14229 21131 14263
rect 22017 14229 22051 14263
rect 26893 14229 26927 14263
rect 26985 14229 27019 14263
rect 27629 14229 27663 14263
rect 28365 14229 28399 14263
rect 39037 14229 39071 14263
rect 4445 14025 4479 14059
rect 11529 14025 11563 14059
rect 11989 14025 12023 14059
rect 15117 14025 15151 14059
rect 18797 14025 18831 14059
rect 22201 14025 22235 14059
rect 27721 14025 27755 14059
rect 31309 14025 31343 14059
rect 33057 14025 33091 14059
rect 33333 14025 33367 14059
rect 34713 14025 34747 14059
rect 37013 14025 37047 14059
rect 2973 13957 3007 13991
rect 15945 13957 15979 13991
rect 16957 13957 16991 13991
rect 17693 13957 17727 13991
rect 18521 13957 18555 13991
rect 28089 13957 28123 13991
rect 30849 13957 30883 13991
rect 31677 13957 31711 13991
rect 35173 13957 35207 13991
rect 35265 13957 35299 13991
rect 35633 13957 35667 13991
rect 39313 13957 39347 13991
rect 11897 13889 11931 13923
rect 15577 13889 15611 13923
rect 15669 13889 15703 13923
rect 16865 13889 16899 13923
rect 17049 13889 17083 13923
rect 17233 13889 17267 13923
rect 17509 13889 17543 13923
rect 17785 13889 17819 13923
rect 17877 13889 17911 13923
rect 18153 13889 18187 13923
rect 18246 13889 18280 13923
rect 18429 13889 18463 13923
rect 18618 13889 18652 13923
rect 19809 13889 19843 13923
rect 19993 13889 20027 13923
rect 20361 13889 20395 13923
rect 20913 13889 20947 13923
rect 21101 13891 21135 13925
rect 21281 13889 21315 13923
rect 21465 13889 21499 13923
rect 22199 13889 22233 13923
rect 22753 13889 22787 13923
rect 22846 13889 22880 13923
rect 23029 13889 23063 13923
rect 23121 13889 23155 13923
rect 23259 13889 23293 13923
rect 23489 13889 23523 13923
rect 23673 13889 23707 13923
rect 23949 13889 23983 13923
rect 24133 13889 24167 13923
rect 24317 13889 24351 13923
rect 24501 13889 24535 13923
rect 24777 13889 24811 13923
rect 24961 13889 24995 13923
rect 25053 13889 25087 13923
rect 25145 13889 25179 13923
rect 25329 13889 25363 13923
rect 25605 13889 25639 13923
rect 25793 13895 25827 13929
rect 25881 13889 25915 13923
rect 26157 13889 26191 13923
rect 27445 13889 27479 13923
rect 27816 13889 27850 13923
rect 27905 13889 27939 13923
rect 28181 13889 28215 13923
rect 28273 13889 28307 13923
rect 31033 13889 31067 13923
rect 31217 13889 31251 13923
rect 31493 13889 31527 13923
rect 31585 13889 31619 13923
rect 31861 13889 31895 13923
rect 31953 13889 31987 13923
rect 32137 13889 32171 13923
rect 32321 13889 32355 13923
rect 32781 13889 32815 13923
rect 33330 13889 33364 13923
rect 33793 13889 33827 13923
rect 34069 13889 34103 13923
rect 34161 13889 34195 13923
rect 34345 13889 34379 13923
rect 34437 13889 34471 13923
rect 34621 13889 34655 13923
rect 34805 13889 34839 13923
rect 35081 13889 35115 13923
rect 35449 13889 35483 13923
rect 35541 13889 35575 13923
rect 35817 13889 35851 13923
rect 36001 13889 36035 13923
rect 36093 13889 36127 13923
rect 38577 13889 38611 13923
rect 2697 13821 2731 13855
rect 12173 13821 12207 13855
rect 15301 13821 15335 13855
rect 16681 13821 16715 13855
rect 21189 13821 21223 13855
rect 21649 13821 21683 13855
rect 22661 13821 22695 13855
rect 23581 13821 23615 13855
rect 24225 13821 24259 13855
rect 24685 13821 24719 13855
rect 25973 13821 26007 13855
rect 32505 13821 32539 13855
rect 33057 13821 33091 13855
rect 36369 13821 36403 13855
rect 38485 13821 38519 13855
rect 38945 13821 38979 13855
rect 39037 13821 39071 13855
rect 41061 13821 41095 13855
rect 15485 13753 15519 13787
rect 18061 13753 18095 13787
rect 20269 13753 20303 13787
rect 22569 13753 22603 13787
rect 27353 13753 27387 13787
rect 33149 13753 33183 13787
rect 33885 13753 33919 13787
rect 34897 13753 34931 13787
rect 22017 13685 22051 13719
rect 23397 13685 23431 13719
rect 25513 13685 25547 13719
rect 26341 13685 26375 13719
rect 27077 13685 27111 13719
rect 27537 13685 27571 13719
rect 28457 13685 28491 13719
rect 32873 13685 32907 13719
rect 33701 13685 33735 13719
rect 5733 13481 5767 13515
rect 12081 13481 12115 13515
rect 16865 13481 16899 13515
rect 33425 13481 33459 13515
rect 35081 13481 35115 13515
rect 35541 13481 35575 13515
rect 36001 13481 36035 13515
rect 17601 13413 17635 13447
rect 20729 13413 20763 13447
rect 36185 13413 36219 13447
rect 38669 13413 38703 13447
rect 12725 13345 12759 13379
rect 13369 13345 13403 13379
rect 13553 13345 13587 13379
rect 17233 13345 17267 13379
rect 17417 13345 17451 13379
rect 20545 13345 20579 13379
rect 25329 13345 25363 13379
rect 27353 13345 27387 13379
rect 35633 13345 35667 13379
rect 38945 13345 38979 13379
rect 39589 13345 39623 13379
rect 5917 13277 5951 13311
rect 6193 13277 6227 13311
rect 6285 13277 6319 13311
rect 7941 13277 7975 13311
rect 8125 13277 8159 13311
rect 12449 13277 12483 13311
rect 13277 13277 13311 13311
rect 16221 13277 16255 13311
rect 16314 13277 16348 13311
rect 16727 13277 16761 13311
rect 20821 13277 20855 13311
rect 22293 13277 22327 13311
rect 22385 13277 22419 13311
rect 22569 13277 22603 13311
rect 22661 13277 22695 13311
rect 24593 13277 24627 13311
rect 24685 13277 24719 13311
rect 24869 13277 24903 13311
rect 24961 13277 24995 13311
rect 25053 13277 25087 13311
rect 25237 13277 25271 13311
rect 25421 13277 25455 13311
rect 25605 13277 25639 13311
rect 25973 13277 26007 13311
rect 26066 13277 26100 13311
rect 26438 13277 26472 13311
rect 26893 13277 26927 13311
rect 26985 13277 27019 13311
rect 27169 13277 27203 13311
rect 27261 13277 27295 13311
rect 27537 13277 27571 13311
rect 27813 13277 27847 13311
rect 31493 13277 31527 13311
rect 31585 13277 31619 13311
rect 31953 13277 31987 13311
rect 32045 13277 32079 13311
rect 33425 13277 33459 13311
rect 33609 13277 33643 13311
rect 34345 13277 34379 13311
rect 34437 13277 34471 13311
rect 34529 13277 34563 13311
rect 34713 13277 34747 13311
rect 34897 13277 34931 13311
rect 35173 13277 35207 13311
rect 35817 13277 35851 13311
rect 36185 13277 36219 13311
rect 36369 13277 36403 13311
rect 38485 13277 38519 13311
rect 38669 13277 38703 13311
rect 38853 13277 38887 13311
rect 39497 13277 39531 13311
rect 39957 13277 39991 13311
rect 40509 13277 40543 13311
rect 12541 13209 12575 13243
rect 16497 13209 16531 13243
rect 16589 13209 16623 13243
rect 16957 13209 16991 13243
rect 20361 13209 20395 13243
rect 22845 13209 22879 13243
rect 26249 13209 26283 13243
rect 26341 13209 26375 13243
rect 35357 13209 35391 13243
rect 37657 13209 37691 13243
rect 6101 13141 6135 13175
rect 6377 13141 6411 13175
rect 8033 13141 8067 13175
rect 12909 13141 12943 13175
rect 17325 13141 17359 13175
rect 22109 13141 22143 13175
rect 22937 13141 22971 13175
rect 24409 13141 24443 13175
rect 25789 13141 25823 13175
rect 26617 13141 26651 13175
rect 26709 13141 26743 13175
rect 27721 13141 27755 13175
rect 31769 13141 31803 13175
rect 32229 13141 32263 13175
rect 39497 13141 39531 13175
rect 40049 13141 40083 13175
rect 41061 13141 41095 13175
rect 7941 12937 7975 12971
rect 9229 12937 9263 12971
rect 11897 12937 11931 12971
rect 12357 12937 12391 12971
rect 12725 12937 12759 12971
rect 16497 12937 16531 12971
rect 19717 12937 19751 12971
rect 41061 12937 41095 12971
rect 6101 12869 6135 12903
rect 6377 12869 6411 12903
rect 6561 12869 6595 12903
rect 6837 12869 6871 12903
rect 9965 12869 9999 12903
rect 24133 12869 24167 12903
rect 24225 12869 24259 12903
rect 28825 12869 28859 12903
rect 29561 12869 29595 12903
rect 31493 12869 31527 12903
rect 33333 12869 33367 12903
rect 4905 12801 4939 12835
rect 5089 12801 5123 12835
rect 5181 12801 5215 12835
rect 5273 12801 5307 12835
rect 6653 12801 6687 12835
rect 6745 12801 6779 12835
rect 6929 12801 6963 12835
rect 7389 12801 7423 12835
rect 7849 12801 7883 12835
rect 8125 12801 8159 12835
rect 8217 12801 8251 12835
rect 8493 12801 8527 12835
rect 8585 12801 8619 12835
rect 8733 12801 8767 12835
rect 8861 12801 8895 12835
rect 8953 12801 8987 12835
rect 9091 12801 9125 12835
rect 9689 12801 9723 12835
rect 10149 12801 10183 12835
rect 11713 12801 11747 12835
rect 12817 12801 12851 12835
rect 14749 12801 14783 12835
rect 19073 12801 19107 12835
rect 19441 12801 19475 12835
rect 19533 12801 19567 12835
rect 19993 12801 20027 12835
rect 20085 12801 20119 12835
rect 20177 12801 20211 12835
rect 20361 12801 20395 12835
rect 20729 12801 20763 12835
rect 21005 12801 21039 12835
rect 23765 12801 23799 12835
rect 23857 12801 23891 12835
rect 31217 12801 31251 12835
rect 31309 12801 31343 12835
rect 31585 12801 31619 12835
rect 31769 12801 31803 12835
rect 33057 12801 33091 12835
rect 37473 12801 37507 12835
rect 39313 12801 39347 12835
rect 7757 12733 7791 12767
rect 9505 12733 9539 12767
rect 11529 12733 11563 12767
rect 12909 12733 12943 12767
rect 18981 12733 19015 12767
rect 20821 12733 20855 12767
rect 31493 12733 31527 12767
rect 31677 12733 31711 12767
rect 34805 12733 34839 12767
rect 37381 12733 37415 12767
rect 37841 12733 37875 12767
rect 39589 12733 39623 12767
rect 21189 12665 21223 12699
rect 4905 12597 4939 12631
rect 6377 12597 6411 12631
rect 8401 12597 8435 12631
rect 9873 12597 9907 12631
rect 10333 12597 10367 12631
rect 15012 12597 15046 12631
rect 18521 12597 18555 12631
rect 20729 12597 20763 12631
rect 23581 12597 23615 12631
rect 6377 12393 6411 12427
rect 10793 12393 10827 12427
rect 15117 12393 15151 12427
rect 19717 12393 19751 12427
rect 27445 12393 27479 12427
rect 31861 12393 31895 12427
rect 39497 12393 39531 12427
rect 15485 12325 15519 12359
rect 21741 12325 21775 12359
rect 23857 12325 23891 12359
rect 24685 12325 24719 12359
rect 29377 12325 29411 12359
rect 3801 12257 3835 12291
rect 6285 12257 6319 12291
rect 12449 12257 12483 12291
rect 12633 12257 12667 12291
rect 13277 12257 13311 12291
rect 13461 12257 13495 12291
rect 14565 12257 14599 12291
rect 14749 12257 14783 12291
rect 15945 12257 15979 12291
rect 16129 12257 16163 12291
rect 19809 12257 19843 12291
rect 23949 12257 23983 12291
rect 28917 12257 28951 12291
rect 30205 12257 30239 12291
rect 30297 12257 30331 12291
rect 31585 12257 31619 12291
rect 40509 12257 40543 12291
rect 40601 12257 40635 12291
rect 2605 12189 2639 12223
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 5822 12189 5856 12223
rect 6193 12189 6227 12223
rect 6377 12189 6411 12223
rect 6653 12189 6687 12223
rect 8401 12189 8435 12223
rect 8493 12189 8527 12223
rect 8585 12189 8619 12223
rect 8769 12189 8803 12223
rect 9229 12189 9263 12223
rect 9321 12189 9355 12223
rect 9597 12189 9631 12223
rect 10517 12189 10551 12223
rect 10609 12189 10643 12223
rect 13185 12189 13219 12223
rect 15025 12189 15059 12223
rect 16313 12189 16347 12223
rect 19533 12189 19567 12223
rect 21189 12189 21223 12223
rect 21465 12189 21499 12223
rect 21557 12189 21591 12223
rect 21833 12189 21867 12223
rect 23427 12189 23461 12223
rect 24501 12189 24535 12223
rect 25053 12189 25087 12223
rect 25237 12189 25271 12223
rect 26433 12189 26467 12223
rect 26617 12189 26651 12223
rect 27077 12189 27111 12223
rect 27261 12189 27295 12223
rect 27353 12189 27387 12223
rect 27445 12189 27479 12223
rect 27629 12189 27663 12223
rect 28733 12189 28767 12223
rect 29009 12189 29043 12223
rect 30573 12189 30607 12223
rect 30965 12189 30999 12223
rect 31217 12189 31251 12223
rect 31401 12189 31435 12223
rect 31493 12189 31527 12223
rect 31677 12189 31711 12223
rect 31861 12189 31895 12223
rect 32045 12189 32079 12223
rect 38669 12189 38703 12223
rect 39681 12189 39715 12223
rect 40417 12189 40451 12223
rect 4077 12121 4111 12155
rect 9689 12121 9723 12155
rect 12357 12121 12391 12155
rect 15853 12121 15887 12155
rect 16405 12121 16439 12155
rect 19349 12121 19383 12155
rect 21373 12121 21407 12155
rect 23555 12121 23589 12155
rect 30113 12121 30147 12155
rect 30757 12121 30791 12155
rect 30849 12121 30883 12155
rect 2421 12053 2455 12087
rect 2789 12053 2823 12087
rect 3617 12053 3651 12087
rect 5549 12053 5583 12087
rect 5641 12053 5675 12087
rect 5825 12053 5859 12087
rect 6561 12053 6595 12087
rect 8125 12053 8159 12087
rect 9045 12053 9079 12087
rect 11989 12053 12023 12087
rect 12817 12053 12851 12087
rect 14105 12053 14139 12087
rect 14473 12053 14507 12087
rect 21925 12053 21959 12087
rect 23305 12053 23339 12087
rect 26525 12053 26559 12087
rect 26893 12053 26927 12087
rect 28549 12053 28583 12087
rect 29745 12053 29779 12087
rect 31125 12053 31159 12087
rect 38485 12053 38519 12087
rect 40049 12053 40083 12087
rect 4905 11849 4939 11883
rect 6101 11849 6135 11883
rect 6745 11849 6779 11883
rect 7849 11849 7883 11883
rect 8217 11849 8251 11883
rect 9505 11849 9539 11883
rect 13369 11849 13403 11883
rect 13461 11849 13495 11883
rect 15761 11849 15795 11883
rect 17601 11849 17635 11883
rect 18337 11849 18371 11883
rect 21915 11849 21949 11883
rect 22385 11849 22419 11883
rect 25145 11849 25179 11883
rect 36093 11849 36127 11883
rect 36829 11849 36863 11883
rect 1961 11781 1995 11815
rect 5089 11781 5123 11815
rect 5289 11781 5323 11815
rect 5917 11781 5951 11815
rect 11897 11781 11931 11815
rect 12081 11781 12115 11815
rect 20637 11781 20671 11815
rect 21649 11781 21683 11815
rect 24777 11781 24811 11815
rect 24869 11781 24903 11815
rect 27353 11781 27387 11815
rect 28549 11781 28583 11815
rect 30297 11781 30331 11815
rect 36369 11781 36403 11815
rect 36553 11781 36587 11815
rect 4537 11713 4571 11747
rect 4675 11713 4709 11747
rect 4997 11713 5031 11747
rect 6193 11713 6227 11747
rect 6561 11713 6595 11747
rect 6821 11713 6855 11747
rect 7481 11713 7515 11747
rect 7849 11713 7883 11747
rect 8033 11713 8067 11747
rect 8401 11713 8435 11747
rect 8493 11713 8527 11747
rect 8677 11713 8711 11747
rect 8769 11713 8803 11747
rect 9321 11713 9355 11747
rect 9597 11713 9631 11747
rect 9781 11713 9815 11747
rect 10425 11713 10459 11747
rect 10885 11713 10919 11747
rect 15209 11713 15243 11747
rect 15393 11713 15427 11747
rect 15485 11713 15519 11747
rect 15577 11713 15611 11747
rect 17141 11713 17175 11747
rect 18797 11713 18831 11747
rect 19073 11713 19107 11747
rect 20453 11713 20487 11747
rect 20729 11713 20763 11747
rect 20821 11713 20855 11747
rect 21189 11713 21223 11747
rect 21373 11713 21407 11747
rect 21557 11713 21591 11747
rect 23397 11713 23431 11747
rect 23581 11713 23615 11747
rect 23765 11713 23799 11747
rect 23949 11713 23983 11747
rect 24501 11713 24535 11747
rect 25053 11713 25087 11747
rect 25421 11713 25455 11747
rect 25605 11713 25639 11747
rect 26065 11713 26099 11747
rect 26158 11713 26192 11747
rect 26341 11713 26375 11747
rect 26433 11713 26467 11747
rect 26530 11713 26564 11747
rect 26985 11713 27019 11747
rect 27169 11713 27203 11747
rect 28273 11713 28307 11747
rect 35633 11713 35667 11747
rect 35817 11713 35851 11747
rect 35909 11713 35943 11747
rect 36093 11713 36127 11747
rect 36185 11713 36219 11747
rect 36645 11713 36679 11747
rect 36921 11713 36955 11747
rect 38117 11713 38151 11747
rect 1685 11645 1719 11679
rect 9137 11645 9171 11679
rect 10241 11645 10275 11679
rect 10701 11645 10735 11679
rect 12173 11645 12207 11679
rect 13645 11645 13679 11679
rect 18429 11645 18463 11679
rect 18613 11645 18647 11679
rect 18889 11645 18923 11679
rect 22293 11645 22327 11679
rect 22477 11645 22511 11679
rect 24409 11645 24443 11679
rect 38393 11645 38427 11679
rect 4813 11577 4847 11611
rect 5457 11577 5491 11611
rect 9597 11577 9631 11611
rect 10609 11577 10643 11611
rect 17969 11577 18003 11611
rect 21005 11577 21039 11611
rect 3433 11509 3467 11543
rect 5273 11509 5307 11543
rect 5917 11509 5951 11543
rect 6377 11509 6411 11543
rect 7573 11509 7607 11543
rect 11069 11509 11103 11543
rect 11621 11509 11655 11543
rect 13001 11509 13035 11543
rect 17233 11509 17267 11543
rect 18797 11509 18831 11543
rect 19257 11509 19291 11543
rect 23397 11509 23431 11543
rect 23765 11509 23799 11543
rect 24225 11509 24259 11543
rect 26709 11509 26743 11543
rect 35725 11509 35759 11543
rect 36645 11509 36679 11543
rect 39865 11509 39899 11543
rect 1593 11305 1627 11339
rect 5733 11305 5767 11339
rect 16681 11305 16715 11339
rect 18429 11305 18463 11339
rect 19441 11305 19475 11339
rect 19809 11305 19843 11339
rect 20821 11305 20855 11339
rect 25053 11305 25087 11339
rect 33241 11305 33275 11339
rect 36645 11305 36679 11339
rect 38301 11305 38335 11339
rect 12081 11237 12115 11271
rect 14105 11237 14139 11271
rect 18061 11237 18095 11271
rect 20269 11237 20303 11271
rect 22845 11237 22879 11271
rect 25881 11237 25915 11271
rect 26157 11237 26191 11271
rect 27537 11237 27571 11271
rect 12449 11169 12483 11203
rect 12633 11169 12667 11203
rect 14657 11169 14691 11203
rect 15301 11169 15335 11203
rect 19625 11169 19659 11203
rect 19901 11169 19935 11203
rect 21373 11169 21407 11203
rect 22937 11169 22971 11203
rect 26709 11169 26743 11203
rect 33057 11169 33091 11203
rect 34805 11169 34839 11203
rect 37473 11169 37507 11203
rect 37933 11169 37967 11203
rect 38945 11169 38979 11203
rect 1501 11101 1535 11135
rect 5733 11101 5767 11135
rect 5825 11101 5859 11135
rect 13921 11101 13955 11135
rect 17785 11101 17819 11135
rect 19257 11101 19291 11135
rect 19349 11101 19383 11135
rect 19533 11101 19567 11135
rect 20085 11101 20119 11135
rect 21649 11101 21683 11135
rect 21833 11101 21867 11135
rect 22475 11101 22509 11135
rect 23213 11101 23247 11135
rect 23673 11101 23707 11135
rect 23857 11101 23891 11135
rect 24409 11101 24443 11135
rect 24502 11101 24536 11135
rect 24777 11101 24811 11135
rect 24874 11101 24908 11135
rect 25511 11101 25545 11135
rect 25973 11101 26007 11135
rect 26893 11101 26927 11135
rect 26986 11101 27020 11135
rect 27358 11101 27392 11135
rect 32965 11101 32999 11135
rect 34943 11101 34977 11135
rect 36185 11101 36219 11135
rect 36369 11101 36403 11135
rect 37565 11101 37599 11135
rect 12541 11033 12575 11067
rect 14565 11033 14599 11067
rect 15025 11033 15059 11067
rect 16497 11033 16531 11067
rect 16681 11033 16715 11067
rect 17049 11033 17083 11067
rect 18429 11033 18463 11067
rect 19809 11033 19843 11067
rect 21097 11033 21131 11067
rect 21281 11033 21315 11067
rect 21925 11033 21959 11067
rect 24685 11033 24719 11067
rect 26433 11033 26467 11067
rect 26617 11033 26651 11067
rect 27169 11033 27203 11067
rect 27261 11033 27295 11067
rect 36001 11033 36035 11067
rect 36461 11033 36495 11067
rect 36661 11033 36695 11067
rect 38761 11033 38795 11067
rect 6101 10965 6135 10999
rect 13737 10965 13771 10999
rect 14473 10965 14507 10999
rect 16865 10965 16899 10999
rect 18613 10965 18647 10999
rect 22293 10965 22327 10999
rect 22477 10965 22511 10999
rect 23121 10965 23155 10999
rect 25329 10965 25363 10999
rect 25513 10965 25547 10999
rect 35265 10965 35299 10999
rect 36829 10965 36863 10999
rect 38669 10965 38703 10999
rect 10701 10761 10735 10795
rect 15025 10761 15059 10795
rect 17601 10761 17635 10795
rect 18530 10761 18564 10795
rect 19266 10761 19300 10795
rect 26249 10761 26283 10795
rect 26801 10761 26835 10795
rect 30113 10761 30147 10795
rect 30941 10761 30975 10795
rect 31309 10761 31343 10795
rect 38669 10761 38703 10795
rect 39037 10761 39071 10795
rect 13553 10693 13587 10727
rect 15577 10693 15611 10727
rect 17141 10693 17175 10727
rect 18153 10693 18187 10727
rect 18889 10693 18923 10727
rect 23397 10693 23431 10727
rect 23489 10693 23523 10727
rect 23627 10693 23661 10727
rect 25421 10693 25455 10727
rect 30205 10693 30239 10727
rect 36001 10693 36035 10727
rect 36093 10693 36127 10727
rect 8217 10625 8251 10659
rect 8677 10625 8711 10659
rect 8953 10625 8987 10659
rect 10517 10625 10551 10659
rect 10793 10625 10827 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 15301 10625 15335 10659
rect 15485 10625 15519 10659
rect 15669 10625 15703 10659
rect 18797 10625 18831 10659
rect 19625 10625 19659 10659
rect 19809 10625 19843 10659
rect 23121 10625 23155 10659
rect 23305 10625 23339 10659
rect 23765 10625 23799 10659
rect 25513 10625 25547 10659
rect 25697 10625 25731 10659
rect 25835 10625 25869 10659
rect 25973 10625 26007 10659
rect 26065 10625 26099 10659
rect 26617 10625 26651 10659
rect 32505 10625 32539 10659
rect 33057 10625 33091 10659
rect 33333 10625 33367 10659
rect 33793 10625 33827 10659
rect 35173 10625 35207 10659
rect 35357 10625 35391 10659
rect 35725 10625 35759 10659
rect 35817 10625 35851 10659
rect 36277 10625 36311 10659
rect 36369 10625 36403 10659
rect 8401 10557 8435 10591
rect 8493 10557 8527 10591
rect 9229 10557 9263 10591
rect 13277 10557 13311 10591
rect 19993 10557 20027 10591
rect 25421 10557 25455 10591
rect 26433 10557 26467 10591
rect 30297 10557 30331 10591
rect 31401 10557 31435 10591
rect 31585 10557 31619 10591
rect 32597 10557 32631 10591
rect 33241 10557 33275 10591
rect 33609 10557 33643 10591
rect 36001 10557 36035 10591
rect 39129 10557 39163 10591
rect 39313 10557 39347 10591
rect 8309 10489 8343 10523
rect 8769 10489 8803 10523
rect 10333 10489 10367 10523
rect 17417 10489 17451 10523
rect 24961 10489 24995 10523
rect 33977 10489 34011 10523
rect 8033 10421 8067 10455
rect 9137 10421 9171 10455
rect 11897 10421 11931 10455
rect 15853 10421 15887 10455
rect 18521 10421 18555 10455
rect 19257 10421 19291 10455
rect 19441 10421 19475 10455
rect 29745 10421 29779 10455
rect 32781 10421 32815 10455
rect 33057 10421 33091 10455
rect 33517 10421 33551 10455
rect 35265 10421 35299 10455
rect 36093 10421 36127 10455
rect 4905 10217 4939 10251
rect 8769 10217 8803 10251
rect 12081 10217 12115 10251
rect 18889 10217 18923 10251
rect 22385 10217 22419 10251
rect 23305 10217 23339 10251
rect 26341 10217 26375 10251
rect 30941 10217 30975 10251
rect 32873 10217 32907 10251
rect 40325 10217 40359 10251
rect 6561 10149 6595 10183
rect 32597 10149 32631 10183
rect 33149 10149 33183 10183
rect 35173 10149 35207 10183
rect 5549 10081 5583 10115
rect 11713 10081 11747 10115
rect 16405 10081 16439 10115
rect 30757 10081 30791 10115
rect 32781 10081 32815 10115
rect 34437 10081 34471 10115
rect 39037 10081 39071 10115
rect 40141 10081 40175 10115
rect 4813 10013 4847 10047
rect 4905 10013 4939 10047
rect 5181 10013 5215 10047
rect 5457 10013 5491 10047
rect 5733 10013 5767 10047
rect 5917 10013 5951 10047
rect 6285 10013 6319 10047
rect 6837 10013 6871 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 8033 10013 8067 10047
rect 8125 10013 8159 10047
rect 8218 10013 8252 10047
rect 8493 10013 8527 10047
rect 8631 10013 8665 10047
rect 9597 10013 9631 10047
rect 10333 10013 10367 10047
rect 10977 10013 11011 10047
rect 11125 10013 11159 10047
rect 11345 10013 11379 10047
rect 11442 10013 11476 10047
rect 11897 10013 11931 10047
rect 12173 10013 12207 10047
rect 12265 10013 12299 10047
rect 12449 10013 12483 10047
rect 15669 10013 15703 10047
rect 16589 10013 16623 10047
rect 16865 10013 16899 10047
rect 18613 10013 18647 10047
rect 21741 10013 21775 10047
rect 22293 10013 22327 10047
rect 23213 10013 23247 10047
rect 23397 10013 23431 10047
rect 25789 10013 25823 10047
rect 26065 10013 26099 10047
rect 26157 10013 26191 10047
rect 27997 10013 28031 10047
rect 29377 10013 29411 10047
rect 30665 10013 30699 10047
rect 32505 10013 32539 10047
rect 32873 10013 32907 10047
rect 33057 10013 33091 10047
rect 33149 10013 33183 10047
rect 33333 10013 33367 10047
rect 34345 10013 34379 10047
rect 34529 10013 34563 10047
rect 34713 10013 34747 10047
rect 35357 10013 35391 10047
rect 35449 10013 35483 10047
rect 39221 10013 39255 10047
rect 39497 10013 39531 10047
rect 39681 10013 39715 10047
rect 40049 10013 40083 10047
rect 4629 9945 4663 9979
rect 6101 9945 6135 9979
rect 6469 9945 6503 9979
rect 6561 9945 6595 9979
rect 8401 9945 8435 9979
rect 11253 9945 11287 9979
rect 12633 9945 12667 9979
rect 16773 9945 16807 9979
rect 22017 9945 22051 9979
rect 25973 9945 26007 9979
rect 34897 9945 34931 9979
rect 35173 9945 35207 9979
rect 5089 9877 5123 9911
rect 6745 9877 6779 9911
rect 7941 9877 7975 9911
rect 11621 9877 11655 9911
rect 16313 9877 16347 9911
rect 27813 9877 27847 9911
rect 29193 9877 29227 9911
rect 32781 9877 32815 9911
rect 35081 9877 35115 9911
rect 39405 9877 39439 9911
rect 39589 9877 39623 9911
rect 15393 9673 15427 9707
rect 15853 9673 15887 9707
rect 25053 9673 25087 9707
rect 30389 9673 30423 9707
rect 31125 9673 31159 9707
rect 32413 9673 32447 9707
rect 39865 9673 39899 9707
rect 3985 9605 4019 9639
rect 4905 9605 4939 9639
rect 6745 9605 6779 9639
rect 15945 9605 15979 9639
rect 16865 9605 16899 9639
rect 19349 9605 19383 9639
rect 21005 9605 21039 9639
rect 26085 9605 26119 9639
rect 28917 9605 28951 9639
rect 32229 9605 32263 9639
rect 37289 9605 37323 9639
rect 3893 9537 3927 9571
rect 4077 9537 4111 9571
rect 4169 9537 4203 9571
rect 4353 9537 4387 9571
rect 4813 9537 4847 9571
rect 5457 9537 5491 9571
rect 6837 9537 6871 9571
rect 7665 9537 7699 9571
rect 8125 9537 8159 9571
rect 9873 9537 9907 9571
rect 10333 9537 10367 9571
rect 11989 9537 12023 9571
rect 12173 9537 12207 9571
rect 13645 9537 13679 9571
rect 16681 9537 16715 9571
rect 16957 9537 16991 9571
rect 17049 9537 17083 9571
rect 20913 9537 20947 9571
rect 21373 9537 21407 9571
rect 21925 9537 21959 9571
rect 25237 9537 25271 9571
rect 25697 9537 25731 9571
rect 25790 9537 25824 9571
rect 25927 9537 25961 9571
rect 26162 9537 26196 9571
rect 27353 9537 27387 9571
rect 28641 9537 28675 9571
rect 30757 9537 30791 9571
rect 32505 9537 32539 9571
rect 37473 9537 37507 9571
rect 37749 9537 37783 9571
rect 37933 9537 37967 9571
rect 38945 9537 38979 9571
rect 39497 9537 39531 9571
rect 39589 9537 39623 9571
rect 39773 9537 39807 9571
rect 39957 9537 39991 9571
rect 4997 9469 5031 9503
rect 5365 9469 5399 9503
rect 6929 9469 6963 9503
rect 13921 9469 13955 9503
rect 16129 9469 16163 9503
rect 19441 9469 19475 9503
rect 19625 9469 19659 9503
rect 21189 9469 21223 9503
rect 25421 9469 25455 9503
rect 25513 9469 25547 9503
rect 27445 9469 27479 9503
rect 27629 9469 27663 9503
rect 27905 9469 27939 9503
rect 30665 9469 30699 9503
rect 39129 9469 39163 9503
rect 4445 9401 4479 9435
rect 5825 9401 5859 9435
rect 17233 9401 17267 9435
rect 20545 9401 20579 9435
rect 26985 9401 27019 9435
rect 37657 9401 37691 9435
rect 4169 9333 4203 9367
rect 6377 9333 6411 9367
rect 15485 9333 15519 9367
rect 18981 9333 19015 9367
rect 21465 9333 21499 9367
rect 22017 9333 22051 9367
rect 26341 9333 26375 9367
rect 28457 9333 28491 9367
rect 32229 9333 32263 9367
rect 37841 9333 37875 9367
rect 4905 9129 4939 9163
rect 8585 9129 8619 9163
rect 14289 9129 14323 9163
rect 17509 9129 17543 9163
rect 19533 9129 19567 9163
rect 22293 9129 22327 9163
rect 34253 9129 34287 9163
rect 38761 9129 38795 9163
rect 9597 9061 9631 9095
rect 16865 9061 16899 9095
rect 39221 9061 39255 9095
rect 8217 8993 8251 9027
rect 9229 8993 9263 9027
rect 20545 8993 20579 9027
rect 20821 8993 20855 9027
rect 26893 8993 26927 9027
rect 26985 8993 27019 9027
rect 29009 8993 29043 9027
rect 36461 8993 36495 9027
rect 36553 8993 36587 9027
rect 38577 8993 38611 9027
rect 4629 8925 4663 8959
rect 4721 8925 4755 8959
rect 6561 8925 6595 8959
rect 6653 8925 6687 8959
rect 6745 8925 6779 8959
rect 6929 8925 6963 8959
rect 8401 8925 8435 8959
rect 9413 8925 9447 8959
rect 10701 8925 10735 8959
rect 10866 8925 10900 8959
rect 10977 8925 11011 8959
rect 11069 8925 11103 8959
rect 14473 8925 14507 8959
rect 16313 8925 16347 8959
rect 16497 8925 16531 8959
rect 16589 8925 16623 8959
rect 16681 8925 16715 8959
rect 16957 8925 16991 8959
rect 17325 8925 17359 8959
rect 18613 8925 18647 8959
rect 19441 8925 19475 8959
rect 26801 8925 26835 8959
rect 27261 8925 27295 8959
rect 34161 8925 34195 8959
rect 34345 8925 34379 8959
rect 34713 8925 34747 8959
rect 34897 8925 34931 8959
rect 36277 8925 36311 8959
rect 36645 8925 36679 8959
rect 36738 8925 36772 8959
rect 37110 8925 37144 8959
rect 37381 8925 37415 8959
rect 38485 8925 38519 8959
rect 38853 8925 38887 8959
rect 39037 8925 39071 8959
rect 17141 8857 17175 8891
rect 17233 8857 17267 8891
rect 27537 8857 27571 8891
rect 32965 8857 32999 8891
rect 36921 8857 36955 8891
rect 37013 8857 37047 8891
rect 38025 8857 38059 8891
rect 6285 8789 6319 8823
rect 10517 8789 10551 8823
rect 18705 8789 18739 8823
rect 26433 8789 26467 8823
rect 33057 8789 33091 8823
rect 34805 8789 34839 8823
rect 36093 8789 36127 8823
rect 37289 8789 37323 8823
rect 38117 8789 38151 8823
rect 3801 8585 3835 8619
rect 15117 8585 15151 8619
rect 22109 8585 22143 8619
rect 24133 8585 24167 8619
rect 29101 8585 29135 8619
rect 30573 8585 30607 8619
rect 31677 8585 31711 8619
rect 34069 8585 34103 8619
rect 16957 8517 16991 8551
rect 17049 8517 17083 8551
rect 18245 8517 18279 8551
rect 22661 8517 22695 8551
rect 25237 8517 25271 8551
rect 31125 8517 31159 8551
rect 32505 8517 32539 8551
rect 33517 8517 33551 8551
rect 33701 8517 33735 8551
rect 35173 8517 35207 8551
rect 36185 8517 36219 8551
rect 36921 8517 36955 8551
rect 37565 8517 37599 8551
rect 39313 8517 39347 8551
rect 4169 8449 4203 8483
rect 5549 8449 5583 8483
rect 6745 8449 6779 8483
rect 8861 8449 8895 8483
rect 9045 8449 9079 8483
rect 14565 8449 14599 8483
rect 14749 8449 14783 8483
rect 14841 8449 14875 8483
rect 14933 8449 14967 8483
rect 16681 8449 16715 8483
rect 16774 8449 16808 8483
rect 17146 8449 17180 8483
rect 17969 8449 18003 8483
rect 19809 8449 19843 8483
rect 19957 8449 19991 8483
rect 20085 8449 20119 8483
rect 20177 8449 20211 8483
rect 20315 8449 20349 8483
rect 22293 8449 22327 8483
rect 24961 8449 24995 8483
rect 25145 8449 25179 8483
rect 27169 8449 27203 8483
rect 27353 8449 27387 8483
rect 30297 8449 30331 8483
rect 30481 8449 30515 8483
rect 30757 8449 30791 8483
rect 31309 8449 31343 8483
rect 31585 8449 31619 8483
rect 31781 8449 31815 8483
rect 32137 8449 32171 8483
rect 32285 8449 32319 8483
rect 32413 8449 32447 8483
rect 32643 8449 32677 8483
rect 33885 8449 33919 8483
rect 34345 8449 34379 8483
rect 34805 8449 34839 8483
rect 34953 8449 34987 8483
rect 35081 8449 35115 8483
rect 35311 8449 35345 8483
rect 36829 8449 36863 8483
rect 37013 8449 37047 8483
rect 40693 8449 40727 8483
rect 4261 8381 4295 8415
rect 4997 8381 5031 8415
rect 6653 8381 6687 8415
rect 7113 8381 7147 8415
rect 12081 8381 12115 8415
rect 12357 8381 12391 8415
rect 13829 8381 13863 8415
rect 19717 8381 19751 8415
rect 22385 8381 22419 8415
rect 27629 8381 27663 8415
rect 30389 8381 30423 8415
rect 31033 8381 31067 8415
rect 32873 8381 32907 8415
rect 34253 8381 34287 8415
rect 35541 8381 35575 8415
rect 37289 8381 37323 8415
rect 8953 8313 8987 8347
rect 17325 8313 17359 8347
rect 26985 8313 27019 8347
rect 34713 8313 34747 8347
rect 40969 8313 41003 8347
rect 4445 8245 4479 8279
rect 20453 8245 20487 8279
rect 30941 8245 30975 8279
rect 31493 8245 31527 8279
rect 32781 8245 32815 8279
rect 35449 8245 35483 8279
rect 5549 8041 5583 8075
rect 12541 8041 12575 8075
rect 15209 8041 15243 8075
rect 20913 8041 20947 8075
rect 22293 8041 22327 8075
rect 24869 8041 24903 8075
rect 25053 8041 25087 8075
rect 34253 8041 34287 8075
rect 17877 7973 17911 8007
rect 25421 7973 25455 8007
rect 38117 7973 38151 8007
rect 4077 7905 4111 7939
rect 6285 7905 6319 7939
rect 9597 7905 9631 7939
rect 13553 7905 13587 7939
rect 19257 7905 19291 7939
rect 22937 7905 22971 7939
rect 24777 7905 24811 7939
rect 30573 7905 30607 7939
rect 31125 7905 31159 7939
rect 31677 7905 31711 7939
rect 34713 7905 34747 7939
rect 35081 7905 35115 7939
rect 38669 7905 38703 7939
rect 1409 7837 1443 7871
rect 3801 7837 3835 7871
rect 6101 7837 6135 7871
rect 8217 7837 8251 7871
rect 8309 7837 8343 7871
rect 8493 7837 8527 7871
rect 8585 7837 8619 7871
rect 9045 7837 9079 7871
rect 10057 7837 10091 7871
rect 10241 7837 10275 7871
rect 10425 7837 10459 7871
rect 10977 7837 11011 7871
rect 12725 7837 12759 7871
rect 13277 7837 13311 7871
rect 14657 7837 14691 7871
rect 15025 7837 15059 7871
rect 15577 7837 15611 7871
rect 15853 7837 15887 7871
rect 15945 7837 15979 7871
rect 16681 7837 16715 7871
rect 16957 7837 16991 7871
rect 17049 7837 17083 7871
rect 17325 7837 17359 7871
rect 17601 7837 17635 7871
rect 17693 7837 17727 7871
rect 19441 7837 19475 7871
rect 19533 7837 19567 7871
rect 19717 7837 19751 7871
rect 19809 7837 19843 7871
rect 21097 7837 21131 7871
rect 21281 7837 21315 7871
rect 21373 7837 21407 7871
rect 22661 7837 22695 7871
rect 24593 7837 24627 7871
rect 24961 7837 24995 7871
rect 25237 7837 25271 7871
rect 25329 7837 25363 7871
rect 25513 7837 25547 7871
rect 25697 7837 25731 7871
rect 25845 7837 25879 7871
rect 25973 7837 26007 7871
rect 26162 7837 26196 7871
rect 30757 7837 30791 7871
rect 30941 7837 30975 7871
rect 31217 7837 31251 7871
rect 33701 7837 33735 7871
rect 34437 7837 34471 7871
rect 34529 7837 34563 7871
rect 34897 7837 34931 7871
rect 38577 7837 38611 7871
rect 39129 7837 39163 7871
rect 39957 7837 39991 7871
rect 1685 7769 1719 7803
rect 10333 7769 10367 7803
rect 11529 7769 11563 7803
rect 11713 7769 11747 7803
rect 14841 7769 14875 7803
rect 14933 7769 14967 7803
rect 15761 7769 15795 7803
rect 16865 7769 16899 7803
rect 17509 7769 17543 7803
rect 26065 7769 26099 7803
rect 31953 7769 31987 7803
rect 34253 7769 34287 7803
rect 38485 7769 38519 7803
rect 40509 7769 40543 7803
rect 5733 7701 5767 7735
rect 6193 7701 6227 7735
rect 8033 7701 8067 7735
rect 10609 7701 10643 7735
rect 11805 7701 11839 7735
rect 12909 7701 12943 7735
rect 13369 7701 13403 7735
rect 16129 7701 16163 7735
rect 17233 7701 17267 7735
rect 22753 7701 22787 7735
rect 26341 7701 26375 7735
rect 31585 7701 31619 7735
rect 38945 7701 38979 7735
rect 17601 7497 17635 7531
rect 21649 7497 21683 7531
rect 24869 7497 24903 7531
rect 24961 7497 24995 7531
rect 26433 7497 26467 7531
rect 27445 7497 27479 7531
rect 40601 7497 40635 7531
rect 8033 7429 8067 7463
rect 9873 7429 9907 7463
rect 15209 7429 15243 7463
rect 17969 7429 18003 7463
rect 21925 7429 21959 7463
rect 24501 7429 24535 7463
rect 5733 7361 5767 7395
rect 7757 7361 7791 7395
rect 9597 7361 9631 7395
rect 14933 7361 14967 7395
rect 15117 7361 15151 7395
rect 15301 7361 15335 7395
rect 15577 7361 15611 7395
rect 15761 7361 15795 7395
rect 15853 7361 15887 7395
rect 15945 7361 15979 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 17141 7361 17175 7395
rect 17785 7361 17819 7395
rect 18061 7361 18095 7395
rect 18613 7361 18647 7395
rect 21005 7361 21039 7395
rect 21098 7361 21132 7395
rect 21281 7361 21315 7395
rect 21373 7361 21407 7395
rect 21511 7361 21545 7395
rect 21833 7361 21867 7395
rect 22109 7361 22143 7395
rect 22385 7361 22419 7395
rect 22569 7361 22603 7395
rect 22937 7361 22971 7395
rect 24225 7361 24259 7395
rect 24318 7361 24352 7395
rect 24593 7361 24627 7395
rect 24690 7361 24724 7395
rect 25145 7361 25179 7395
rect 25237 7361 25271 7395
rect 25421 7361 25455 7395
rect 25513 7361 25547 7395
rect 25789 7361 25823 7395
rect 25882 7361 25916 7395
rect 26065 7361 26099 7395
rect 26157 7361 26191 7395
rect 26254 7361 26288 7395
rect 27353 7361 27387 7395
rect 28457 7361 28491 7395
rect 28733 7361 28767 7395
rect 34713 7361 34747 7395
rect 27537 7293 27571 7327
rect 27905 7293 27939 7327
rect 34989 7293 35023 7327
rect 36461 7293 36495 7327
rect 38853 7293 38887 7327
rect 39129 7293 39163 7327
rect 16129 7225 16163 7259
rect 26985 7225 27019 7259
rect 5549 7157 5583 7191
rect 9505 7157 9539 7191
rect 11345 7157 11379 7191
rect 15485 7157 15519 7191
rect 16681 7157 16715 7191
rect 19165 7157 19199 7191
rect 28549 7157 28583 7191
rect 5536 6953 5570 6987
rect 7021 6953 7055 6987
rect 22017 6953 22051 6987
rect 29745 6885 29779 6919
rect 5273 6817 5307 6851
rect 13921 6817 13955 6851
rect 14657 6817 14691 6851
rect 16313 6817 16347 6851
rect 18521 6817 18555 6851
rect 19901 6817 19935 6851
rect 20085 6817 20119 6851
rect 20269 6817 20303 6851
rect 25329 6817 25363 6851
rect 26709 6817 26743 6851
rect 26893 6817 26927 6851
rect 28825 6817 28859 6851
rect 30205 6817 30239 6851
rect 30297 6817 30331 6851
rect 9137 6749 9171 6783
rect 9873 6749 9907 6783
rect 11161 6749 11195 6783
rect 11437 6749 11471 6783
rect 12173 6749 12207 6783
rect 14565 6749 14599 6783
rect 18429 6749 18463 6783
rect 19073 6749 19107 6783
rect 21005 6749 21039 6783
rect 21189 6749 21223 6783
rect 21465 6749 21499 6783
rect 21833 6749 21867 6783
rect 24501 6749 24535 6783
rect 24961 6749 24995 6783
rect 25145 6749 25179 6783
rect 26617 6749 26651 6783
rect 27077 6749 27111 6783
rect 29377 6749 29411 6783
rect 30757 6749 30791 6783
rect 36645 6749 36679 6783
rect 9965 6681 9999 6715
rect 12449 6681 12483 6715
rect 18337 6681 18371 6715
rect 19809 6681 19843 6715
rect 20913 6681 20947 6715
rect 21649 6681 21683 6715
rect 21741 6681 21775 6715
rect 27353 6681 27387 6715
rect 30113 6681 30147 6715
rect 31309 6681 31343 6715
rect 37381 6681 37415 6715
rect 9781 6613 9815 6647
rect 10977 6613 11011 6647
rect 11345 6613 11379 6647
rect 14105 6613 14139 6647
rect 14473 6613 14507 6647
rect 16865 6613 16899 6647
rect 17969 6613 18003 6647
rect 18889 6613 18923 6647
rect 19441 6613 19475 6647
rect 21373 6613 21407 6647
rect 24777 6613 24811 6647
rect 26249 6613 26283 6647
rect 29193 6613 29227 6647
rect 4445 6409 4479 6443
rect 4905 6409 4939 6443
rect 9321 6409 9355 6443
rect 12357 6409 12391 6443
rect 12909 6409 12943 6443
rect 13829 6409 13863 6443
rect 15485 6409 15519 6443
rect 15853 6409 15887 6443
rect 15945 6409 15979 6443
rect 20361 6409 20395 6443
rect 26985 6409 27019 6443
rect 29101 6409 29135 6443
rect 36921 6409 36955 6443
rect 9413 6341 9447 6375
rect 27629 6341 27663 6375
rect 29561 6341 29595 6375
rect 37565 6341 37599 6375
rect 4077 6273 4111 6307
rect 4813 6273 4847 6307
rect 5917 6273 5951 6307
rect 13093 6273 13127 6307
rect 13737 6273 13771 6307
rect 15301 6273 15335 6307
rect 16773 6273 16807 6307
rect 18613 6273 18647 6307
rect 24225 6273 24259 6307
rect 27169 6273 27203 6307
rect 29285 6273 29319 6307
rect 37105 6273 37139 6307
rect 4997 6205 5031 6239
rect 5273 6205 5307 6239
rect 7113 6205 7147 6239
rect 7389 6205 7423 6239
rect 9505 6205 9539 6239
rect 11713 6205 11747 6239
rect 16037 6205 16071 6239
rect 17049 6205 17083 6239
rect 18889 6205 18923 6239
rect 22293 6205 22327 6239
rect 22569 6205 22603 6239
rect 24041 6205 24075 6239
rect 24869 6205 24903 6239
rect 27353 6205 27387 6239
rect 37289 6205 37323 6239
rect 39037 6205 39071 6239
rect 39221 6205 39255 6239
rect 18521 6137 18555 6171
rect 3893 6069 3927 6103
rect 8861 6069 8895 6103
rect 8953 6069 8987 6103
rect 15117 6069 15151 6103
rect 24777 6069 24811 6103
rect 25513 6069 25547 6103
rect 31033 6069 31067 6103
rect 39773 6069 39807 6103
rect 8033 5865 8067 5899
rect 10504 5865 10538 5899
rect 16405 5865 16439 5899
rect 17601 5865 17635 5899
rect 21557 5865 21591 5899
rect 22753 5865 22787 5899
rect 37197 5865 37231 5899
rect 23029 5797 23063 5831
rect 7757 5729 7791 5763
rect 10241 5729 10275 5763
rect 13645 5729 13679 5763
rect 14933 5729 14967 5763
rect 19809 5729 19843 5763
rect 21649 5729 21683 5763
rect 23581 5729 23615 5763
rect 25053 5729 25087 5763
rect 26525 5729 26559 5763
rect 31217 5729 31251 5763
rect 31309 5729 31343 5763
rect 31585 5729 31619 5763
rect 33333 5729 33367 5763
rect 35173 5729 35207 5763
rect 35357 5729 35391 5763
rect 37749 5729 37783 5763
rect 5089 5661 5123 5695
rect 7021 5661 7055 5695
rect 8217 5661 8251 5695
rect 14657 5661 14691 5695
rect 17785 5661 17819 5695
rect 22937 5661 22971 5695
rect 24041 5661 24075 5695
rect 24777 5661 24811 5695
rect 25697 5661 25731 5695
rect 35817 5661 35851 5695
rect 37565 5661 37599 5695
rect 5365 5593 5399 5627
rect 13553 5593 13587 5627
rect 20085 5593 20119 5627
rect 23489 5593 23523 5627
rect 24869 5593 24903 5627
rect 31861 5593 31895 5627
rect 35081 5593 35115 5627
rect 36369 5593 36403 5627
rect 6837 5525 6871 5559
rect 11989 5525 12023 5559
rect 13093 5525 13127 5559
rect 13461 5525 13495 5559
rect 22293 5525 22327 5559
rect 23397 5525 23431 5559
rect 23857 5525 23891 5559
rect 24409 5525 24443 5559
rect 30757 5525 30791 5559
rect 31125 5525 31159 5559
rect 34713 5525 34747 5559
rect 37657 5525 37691 5559
rect 5641 5321 5675 5355
rect 6377 5321 6411 5355
rect 6837 5321 6871 5355
rect 11069 5321 11103 5355
rect 13921 5321 13955 5355
rect 20269 5321 20303 5355
rect 20913 5321 20947 5355
rect 24777 5321 24811 5355
rect 26801 5321 26835 5355
rect 31677 5321 31711 5355
rect 3525 5253 3559 5287
rect 23213 5253 23247 5287
rect 25329 5253 25363 5287
rect 5825 5185 5859 5219
rect 6745 5185 6779 5219
rect 7849 5185 7883 5219
rect 10517 5185 10551 5219
rect 10977 5185 11011 5219
rect 11713 5185 11747 5219
rect 12173 5185 12207 5219
rect 20453 5185 20487 5219
rect 22937 5185 22971 5219
rect 24961 5185 24995 5219
rect 31861 5185 31895 5219
rect 34437 5185 34471 5219
rect 34529 5185 34563 5219
rect 3249 5117 3283 5151
rect 6929 5117 6963 5151
rect 7205 5117 7239 5151
rect 9965 5117 9999 5151
rect 11161 5117 11195 5151
rect 12449 5117 12483 5151
rect 21005 5117 21039 5151
rect 21097 5117 21131 5151
rect 24685 5117 24719 5151
rect 25053 5117 25087 5151
rect 34805 5117 34839 5151
rect 10609 5049 10643 5083
rect 20545 5049 20579 5083
rect 34253 5049 34287 5083
rect 4997 4981 5031 5015
rect 11529 4981 11563 5015
rect 36277 4981 36311 5015
rect 10320 4777 10354 4811
rect 12633 4777 12667 4811
rect 18337 4777 18371 4811
rect 24777 4777 24811 4811
rect 28181 4777 28215 4811
rect 11805 4709 11839 4743
rect 25605 4709 25639 4743
rect 36737 4709 36771 4743
rect 10057 4641 10091 4675
rect 18429 4641 18463 4675
rect 20913 4641 20947 4675
rect 21281 4641 21315 4675
rect 25237 4641 25271 4675
rect 25421 4641 25455 4675
rect 26065 4641 26099 4675
rect 26157 4641 26191 4675
rect 26433 4641 26467 4675
rect 37657 4641 37691 4675
rect 12817 4573 12851 4607
rect 16589 4573 16623 4607
rect 20821 4573 20855 4607
rect 25145 4573 25179 4607
rect 36921 4573 36955 4607
rect 37473 4573 37507 4607
rect 38393 4573 38427 4607
rect 40693 4573 40727 4607
rect 16865 4505 16899 4539
rect 20729 4505 20763 4539
rect 21833 4505 21867 4539
rect 25973 4505 26007 4539
rect 26709 4505 26743 4539
rect 37381 4505 37415 4539
rect 38945 4505 38979 4539
rect 19073 4437 19107 4471
rect 20361 4437 20395 4471
rect 37013 4437 37047 4471
rect 40969 4437 41003 4471
rect 15577 4233 15611 4267
rect 16037 4233 16071 4267
rect 17049 4233 17083 4267
rect 17325 4233 17359 4267
rect 17693 4233 17727 4267
rect 21281 4233 21315 4267
rect 21373 4233 21407 4267
rect 22201 4233 22235 4267
rect 26433 4233 26467 4267
rect 18613 4165 18647 4199
rect 37565 4165 37599 4199
rect 13829 4097 13863 4131
rect 16129 4097 16163 4131
rect 16957 4097 16991 4131
rect 17233 4097 17267 4131
rect 18337 4097 18371 4131
rect 20269 4097 20303 4131
rect 24133 4097 24167 4131
rect 25145 4097 25179 4131
rect 25973 4097 26007 4131
rect 26617 4097 26651 4131
rect 37289 4097 37323 4131
rect 14105 4029 14139 4063
rect 16221 4029 16255 4063
rect 17785 4029 17819 4063
rect 17877 4029 17911 4063
rect 21557 4029 21591 4063
rect 22293 4029 22327 4063
rect 22477 4029 22511 4063
rect 25789 3961 25823 3995
rect 15669 3893 15703 3927
rect 16773 3893 16807 3927
rect 20085 3893 20119 3927
rect 20821 3893 20855 3927
rect 20913 3893 20947 3927
rect 21833 3893 21867 3927
rect 23949 3893 23983 3927
rect 25697 3893 25731 3927
rect 39037 3893 39071 3927
rect 14197 3689 14231 3723
rect 17325 3689 17359 3723
rect 18889 3689 18923 3723
rect 22201 3689 22235 3723
rect 24041 3689 24075 3723
rect 24409 3689 24443 3723
rect 26985 3689 27019 3723
rect 17049 3621 17083 3655
rect 19257 3621 19291 3655
rect 13737 3553 13771 3587
rect 15025 3553 15059 3587
rect 17785 3553 17819 3587
rect 17877 3553 17911 3587
rect 19809 3553 19843 3587
rect 20453 3553 20487 3587
rect 22293 3553 22327 3587
rect 24961 3553 24995 3587
rect 25237 3553 25271 3587
rect 25513 3553 25547 3587
rect 1501 3485 1535 3519
rect 13093 3485 13127 3519
rect 13553 3485 13587 3519
rect 14381 3485 14415 3519
rect 14933 3485 14967 3519
rect 15485 3485 15519 3519
rect 15761 3485 15795 3519
rect 18153 3485 18187 3519
rect 19073 3485 19107 3519
rect 19625 3485 19659 3519
rect 20361 3485 20395 3519
rect 24777 3485 24811 3519
rect 16589 3417 16623 3451
rect 17693 3417 17727 3451
rect 18797 3417 18831 3451
rect 20729 3417 20763 3451
rect 22569 3417 22603 3451
rect 1593 3349 1627 3383
rect 12909 3349 12943 3383
rect 13185 3349 13219 3383
rect 13645 3349 13679 3383
rect 14473 3349 14507 3383
rect 14841 3349 14875 3383
rect 15301 3349 15335 3383
rect 19717 3349 19751 3383
rect 20177 3349 20211 3383
rect 24869 3349 24903 3383
rect 21281 3145 21315 3179
rect 22201 3145 22235 3179
rect 25237 3145 25271 3179
rect 25697 3145 25731 3179
rect 26065 3145 26099 3179
rect 13001 3077 13035 3111
rect 15025 3077 15059 3111
rect 16957 3077 16991 3111
rect 23765 3077 23799 3111
rect 26157 3077 26191 3111
rect 14749 3009 14783 3043
rect 16681 3009 16715 3043
rect 19533 3009 19567 3043
rect 22385 3009 22419 3043
rect 23489 3009 23523 3043
rect 12725 2941 12759 2975
rect 19809 2941 19843 2975
rect 26341 2941 26375 2975
rect 16497 2873 16531 2907
rect 14473 2805 14507 2839
rect 18429 2805 18463 2839
rect 20177 2601 20211 2635
rect 1685 2397 1719 2431
rect 7941 2397 7975 2431
rect 11805 2397 11839 2431
rect 15669 2397 15703 2431
rect 19533 2397 19567 2431
rect 20361 2397 20395 2431
rect 23397 2397 23431 2431
rect 31125 2397 31159 2431
rect 34989 2397 35023 2431
rect 38853 2397 38887 2431
rect 40693 2397 40727 2431
rect 1501 2329 1535 2363
rect 4077 2329 4111 2363
rect 27261 2329 27295 2363
rect 4169 2261 4203 2295
rect 8033 2261 8067 2295
rect 11897 2261 11931 2295
rect 15761 2261 15795 2295
rect 19625 2261 19659 2295
rect 23489 2261 23523 2295
rect 27353 2261 27387 2295
rect 31217 2261 31251 2295
rect 35081 2261 35115 2295
rect 38945 2261 38979 2295
rect 40785 2261 40819 2295
<< metal1 >>
rect 10870 42508 10876 42560
rect 10928 42548 10934 42560
rect 14550 42548 14556 42560
rect 10928 42520 14556 42548
rect 10928 42508 10934 42520
rect 14550 42508 14556 42520
rect 14608 42508 14614 42560
rect 1104 42458 41400 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 41400 42458
rect 1104 42384 41400 42406
rect 11054 42304 11060 42356
rect 11112 42304 11118 42356
rect 11624 42316 12434 42344
rect 1857 42279 1915 42285
rect 1857 42245 1869 42279
rect 1903 42276 1915 42279
rect 2774 42276 2780 42288
rect 1903 42248 2780 42276
rect 1903 42245 1915 42248
rect 1857 42239 1915 42245
rect 2774 42236 2780 42248
rect 2832 42236 2838 42288
rect 7098 42236 7104 42288
rect 7156 42276 7162 42288
rect 7285 42279 7343 42285
rect 7285 42276 7297 42279
rect 7156 42248 7297 42276
rect 7156 42236 7162 42248
rect 7285 42245 7297 42248
rect 7331 42245 7343 42279
rect 7285 42239 7343 42245
rect 1486 42168 1492 42220
rect 1544 42168 1550 42220
rect 3234 42168 3240 42220
rect 3292 42208 3298 42220
rect 3329 42211 3387 42217
rect 3329 42208 3341 42211
rect 3292 42180 3341 42208
rect 3292 42168 3298 42180
rect 3329 42177 3341 42180
rect 3375 42177 3387 42211
rect 11072 42208 11100 42304
rect 11624 42285 11652 42316
rect 11609 42279 11667 42285
rect 11609 42245 11621 42279
rect 11655 42245 11667 42279
rect 12406 42276 12434 42316
rect 18690 42304 18696 42356
rect 18748 42344 18754 42356
rect 19429 42347 19487 42353
rect 19429 42344 19441 42347
rect 18748 42316 19441 42344
rect 18748 42304 18754 42316
rect 19429 42313 19441 42316
rect 19475 42313 19487 42347
rect 29086 42344 29092 42356
rect 19429 42307 19487 42313
rect 22066 42316 29092 42344
rect 22066 42276 22094 42316
rect 29086 42304 29092 42316
rect 29144 42304 29150 42356
rect 30374 42304 30380 42356
rect 30432 42344 30438 42356
rect 30561 42347 30619 42353
rect 30561 42344 30573 42347
rect 30432 42316 30573 42344
rect 30432 42304 30438 42316
rect 30561 42313 30573 42316
rect 30607 42313 30619 42347
rect 30561 42307 30619 42313
rect 32950 42304 32956 42356
rect 33008 42304 33014 42356
rect 38286 42304 38292 42356
rect 38344 42304 38350 42356
rect 41874 42304 41880 42356
rect 41932 42304 41938 42356
rect 32968 42276 32996 42304
rect 12406 42248 22094 42276
rect 22480 42248 32996 42276
rect 11609 42239 11667 42245
rect 11241 42211 11299 42217
rect 11241 42208 11253 42211
rect 11072 42180 11253 42208
rect 3329 42171 3387 42177
rect 11241 42177 11253 42180
rect 11287 42177 11299 42211
rect 11241 42171 11299 42177
rect 11517 42211 11575 42217
rect 11517 42177 11529 42211
rect 11563 42177 11575 42211
rect 11517 42171 11575 42177
rect 11532 42140 11560 42171
rect 14642 42168 14648 42220
rect 14700 42168 14706 42220
rect 14826 42168 14832 42220
rect 14884 42208 14890 42220
rect 15197 42211 15255 42217
rect 15197 42208 15209 42211
rect 14884 42180 15209 42208
rect 14884 42168 14890 42180
rect 15197 42177 15209 42180
rect 15243 42177 15255 42211
rect 16022 42208 16028 42220
rect 15197 42171 15255 42177
rect 15488 42180 16028 42208
rect 6886 42112 10916 42140
rect 3513 42007 3571 42013
rect 3513 41973 3525 42007
rect 3559 42004 3571 42007
rect 6886 42004 6914 42112
rect 10888 42084 10916 42112
rect 11072 42112 11560 42140
rect 14660 42140 14688 42168
rect 15381 42143 15439 42149
rect 15381 42140 15393 42143
rect 14660 42112 15393 42140
rect 7469 42075 7527 42081
rect 7469 42041 7481 42075
rect 7515 42041 7527 42075
rect 7469 42035 7527 42041
rect 3559 41976 6914 42004
rect 7484 42004 7512 42035
rect 10870 42032 10876 42084
rect 10928 42032 10934 42084
rect 11072 42081 11100 42112
rect 15381 42109 15393 42112
rect 15427 42109 15439 42143
rect 15381 42103 15439 42109
rect 11057 42075 11115 42081
rect 11057 42041 11069 42075
rect 11103 42041 11115 42075
rect 15488 42072 15516 42180
rect 16022 42168 16028 42180
rect 16080 42168 16086 42220
rect 19337 42211 19395 42217
rect 19337 42177 19349 42211
rect 19383 42208 19395 42211
rect 22480 42208 22508 42248
rect 34514 42236 34520 42288
rect 34572 42276 34578 42288
rect 34793 42279 34851 42285
rect 34793 42276 34805 42279
rect 34572 42248 34805 42276
rect 34572 42236 34578 42248
rect 34793 42245 34805 42248
rect 34839 42245 34851 42279
rect 34793 42239 34851 42245
rect 19383 42180 22508 42208
rect 19383 42177 19395 42180
rect 19337 42171 19395 42177
rect 22554 42168 22560 42220
rect 22612 42208 22618 42220
rect 22649 42211 22707 42217
rect 22649 42208 22661 42211
rect 22612 42180 22661 42208
rect 22612 42168 22618 42180
rect 22649 42177 22661 42180
rect 22695 42177 22707 42211
rect 22649 42171 22707 42177
rect 30466 42168 30472 42220
rect 30524 42168 30530 42220
rect 38194 42168 38200 42220
rect 38252 42168 38258 42220
rect 41049 42211 41107 42217
rect 41049 42177 41061 42211
rect 41095 42208 41107 42211
rect 41892 42208 41920 42304
rect 41095 42180 41920 42208
rect 41095 42177 41107 42180
rect 41049 42171 41107 42177
rect 31662 42140 31668 42152
rect 11057 42035 11115 42041
rect 13924 42044 15516 42072
rect 15580 42112 31668 42140
rect 13924 42004 13952 42044
rect 7484 41976 13952 42004
rect 3559 41973 3571 41976
rect 3513 41967 3571 41973
rect 13998 41964 14004 42016
rect 14056 42004 14062 42016
rect 14921 42007 14979 42013
rect 14921 42004 14933 42007
rect 14056 41976 14933 42004
rect 14056 41964 14062 41976
rect 14921 41973 14933 41976
rect 14967 42004 14979 42007
rect 15580 42004 15608 42112
rect 31662 42100 31668 42112
rect 31720 42100 31726 42152
rect 32674 42100 32680 42152
rect 32732 42100 32738 42152
rect 16022 42032 16028 42084
rect 16080 42072 16086 42084
rect 23474 42072 23480 42084
rect 16080 42044 23480 42072
rect 16080 42032 16086 42044
rect 23474 42032 23480 42044
rect 23532 42032 23538 42084
rect 24394 42032 24400 42084
rect 24452 42072 24458 42084
rect 24452 42044 34928 42072
rect 24452 42032 24458 42044
rect 14967 41976 15608 42004
rect 14967 41973 14979 41976
rect 14921 41967 14979 41973
rect 20714 41964 20720 42016
rect 20772 42004 20778 42016
rect 22833 42007 22891 42013
rect 22833 42004 22845 42007
rect 20772 41976 22845 42004
rect 20772 41964 20778 41976
rect 22833 41973 22845 41976
rect 22879 41973 22891 42007
rect 22833 41967 22891 41973
rect 33318 41964 33324 42016
rect 33376 41964 33382 42016
rect 34900 42013 34928 42044
rect 34885 42007 34943 42013
rect 34885 41973 34897 42007
rect 34931 41973 34943 42007
rect 34885 41967 34943 41973
rect 40862 41964 40868 42016
rect 40920 41964 40926 42016
rect 1104 41914 41400 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 41400 41914
rect 1104 41840 41400 41862
rect 10980 41772 14044 41800
rect 10505 41599 10563 41605
rect 10505 41596 10517 41599
rect 9646 41568 10517 41596
rect 7190 41488 7196 41540
rect 7248 41528 7254 41540
rect 9646 41528 9674 41568
rect 10505 41565 10517 41568
rect 10551 41596 10563 41599
rect 10980 41596 11008 41772
rect 14016 41744 14044 41772
rect 14550 41760 14556 41812
rect 14608 41800 14614 41812
rect 14608 41772 16804 41800
rect 14608 41760 14614 41772
rect 13998 41692 14004 41744
rect 14056 41692 14062 41744
rect 11054 41624 11060 41676
rect 11112 41664 11118 41676
rect 12710 41664 12716 41676
rect 11112 41636 12716 41664
rect 11112 41624 11118 41636
rect 12710 41624 12716 41636
rect 12768 41664 12774 41676
rect 14093 41667 14151 41673
rect 14093 41664 14105 41667
rect 12768 41636 14105 41664
rect 12768 41624 12774 41636
rect 14093 41633 14105 41636
rect 14139 41633 14151 41667
rect 14093 41627 14151 41633
rect 15010 41624 15016 41676
rect 15068 41664 15074 41676
rect 15068 41636 16620 41664
rect 15068 41624 15074 41636
rect 10551 41568 11008 41596
rect 10551 41565 10563 41568
rect 10505 41559 10563 41565
rect 11422 41556 11428 41608
rect 11480 41556 11486 41608
rect 13446 41596 13452 41608
rect 12452 41568 13452 41596
rect 12452 41540 12480 41568
rect 13446 41556 13452 41568
rect 13504 41556 13510 41608
rect 13538 41556 13544 41608
rect 13596 41556 13602 41608
rect 13633 41599 13691 41605
rect 13633 41565 13645 41599
rect 13679 41596 13691 41599
rect 13998 41596 14004 41608
rect 13679 41568 14004 41596
rect 13679 41565 13691 41568
rect 13633 41559 13691 41565
rect 13998 41556 14004 41568
rect 14056 41556 14062 41608
rect 16592 41605 16620 41636
rect 16776 41605 16804 41772
rect 17770 41760 17776 41812
rect 17828 41800 17834 41812
rect 23937 41803 23995 41809
rect 23937 41800 23949 41803
rect 17828 41772 23949 41800
rect 17828 41760 17834 41772
rect 23937 41769 23949 41772
rect 23983 41769 23995 41803
rect 23937 41763 23995 41769
rect 28721 41803 28779 41809
rect 28721 41769 28733 41803
rect 28767 41800 28779 41803
rect 28994 41800 29000 41812
rect 28767 41772 29000 41800
rect 28767 41769 28779 41772
rect 28721 41763 28779 41769
rect 28994 41760 29000 41772
rect 29052 41760 29058 41812
rect 29086 41760 29092 41812
rect 29144 41800 29150 41812
rect 30910 41803 30968 41809
rect 30910 41800 30922 41803
rect 29144 41772 30922 41800
rect 29144 41760 29150 41772
rect 30910 41769 30922 41772
rect 30956 41769 30968 41803
rect 30910 41763 30968 41769
rect 32401 41803 32459 41809
rect 32401 41769 32413 41803
rect 32447 41800 32459 41803
rect 32674 41800 32680 41812
rect 32447 41772 32680 41800
rect 32447 41769 32459 41772
rect 32401 41763 32459 41769
rect 32674 41760 32680 41772
rect 32732 41760 32738 41812
rect 19426 41692 19432 41744
rect 19484 41732 19490 41744
rect 19613 41735 19671 41741
rect 19613 41732 19625 41735
rect 19484 41704 19625 41732
rect 19484 41692 19490 41704
rect 19613 41701 19625 41704
rect 19659 41701 19671 41735
rect 20254 41732 20260 41744
rect 19613 41695 19671 41701
rect 19996 41704 20260 41732
rect 18690 41664 18696 41676
rect 18248 41636 18696 41664
rect 18248 41605 18276 41636
rect 18690 41624 18696 41636
rect 18748 41624 18754 41676
rect 19058 41624 19064 41676
rect 19116 41624 19122 41676
rect 19886 41624 19892 41676
rect 19944 41624 19950 41676
rect 19996 41673 20024 41704
rect 20254 41692 20260 41704
rect 20312 41692 20318 41744
rect 20717 41735 20775 41741
rect 20717 41701 20729 41735
rect 20763 41732 20775 41735
rect 24486 41732 24492 41744
rect 20763 41704 24492 41732
rect 20763 41701 20775 41704
rect 20717 41695 20775 41701
rect 24486 41692 24492 41704
rect 24544 41692 24550 41744
rect 19981 41667 20039 41673
rect 19981 41633 19993 41667
rect 20027 41633 20039 41667
rect 19981 41627 20039 41633
rect 20162 41624 20168 41676
rect 20220 41664 20226 41676
rect 22557 41667 22615 41673
rect 20220 41636 20576 41664
rect 20220 41624 20226 41636
rect 15933 41599 15991 41605
rect 15933 41596 15945 41599
rect 15856 41568 15945 41596
rect 7248 41500 9674 41528
rect 7248 41488 7254 41500
rect 12434 41488 12440 41540
rect 12492 41488 12498 41540
rect 14369 41531 14427 41537
rect 14369 41528 14381 41531
rect 13372 41500 14381 41528
rect 10594 41420 10600 41472
rect 10652 41420 10658 41472
rect 12851 41463 12909 41469
rect 12851 41429 12863 41463
rect 12897 41460 12909 41463
rect 13262 41460 13268 41472
rect 12897 41432 13268 41460
rect 12897 41429 12909 41432
rect 12851 41423 12909 41429
rect 13262 41420 13268 41432
rect 13320 41420 13326 41472
rect 13372 41469 13400 41500
rect 14369 41497 14381 41500
rect 14415 41497 14427 41531
rect 14369 41491 14427 41497
rect 14476 41500 14858 41528
rect 13357 41463 13415 41469
rect 13357 41429 13369 41463
rect 13403 41429 13415 41463
rect 13357 41423 13415 41429
rect 13446 41420 13452 41472
rect 13504 41460 13510 41472
rect 13817 41463 13875 41469
rect 13817 41460 13829 41463
rect 13504 41432 13829 41460
rect 13504 41420 13510 41432
rect 13817 41429 13829 41432
rect 13863 41460 13875 41463
rect 14476 41460 14504 41500
rect 13863 41432 14504 41460
rect 13863 41429 13875 41432
rect 13817 41423 13875 41429
rect 15102 41420 15108 41472
rect 15160 41460 15166 41472
rect 15856 41469 15884 41568
rect 15933 41565 15945 41568
rect 15979 41565 15991 41599
rect 15933 41559 15991 41565
rect 16577 41599 16635 41605
rect 16577 41565 16589 41599
rect 16623 41565 16635 41599
rect 16577 41559 16635 41565
rect 16761 41599 16819 41605
rect 16761 41565 16773 41599
rect 16807 41565 16819 41599
rect 16761 41559 16819 41565
rect 18233 41599 18291 41605
rect 18233 41565 18245 41599
rect 18279 41565 18291 41599
rect 18233 41559 18291 41565
rect 18417 41599 18475 41605
rect 18417 41565 18429 41599
rect 18463 41596 18475 41599
rect 19076 41596 19104 41624
rect 20548 41608 20576 41636
rect 22557 41633 22569 41667
rect 22603 41664 22615 41667
rect 23290 41664 23296 41676
rect 22603 41636 23296 41664
rect 22603 41633 22615 41636
rect 22557 41627 22615 41633
rect 23290 41624 23296 41636
rect 23348 41624 23354 41676
rect 24302 41624 24308 41676
rect 24360 41664 24366 41676
rect 24360 41636 24716 41664
rect 24360 41624 24366 41636
rect 18463 41568 19104 41596
rect 19797 41599 19855 41605
rect 18463 41565 18475 41568
rect 18417 41559 18475 41565
rect 19797 41565 19809 41599
rect 19843 41565 19855 41599
rect 19797 41559 19855 41565
rect 17129 41531 17187 41537
rect 17129 41497 17141 41531
rect 17175 41528 17187 41531
rect 17494 41528 17500 41540
rect 17175 41500 17500 41528
rect 17175 41497 17187 41500
rect 17129 41491 17187 41497
rect 17494 41488 17500 41500
rect 17552 41528 17558 41540
rect 18432 41528 18460 41559
rect 17552 41500 18460 41528
rect 18509 41531 18567 41537
rect 17552 41488 17558 41500
rect 18509 41497 18521 41531
rect 18555 41497 18567 41531
rect 18509 41491 18567 41497
rect 18693 41531 18751 41537
rect 18693 41497 18705 41531
rect 18739 41528 18751 41531
rect 18966 41528 18972 41540
rect 18739 41500 18972 41528
rect 18739 41497 18751 41500
rect 18693 41491 18751 41497
rect 15841 41463 15899 41469
rect 15841 41460 15853 41463
rect 15160 41432 15853 41460
rect 15160 41420 15166 41432
rect 15841 41429 15853 41432
rect 15887 41429 15899 41463
rect 15841 41423 15899 41429
rect 17954 41420 17960 41472
rect 18012 41460 18018 41472
rect 18524 41460 18552 41491
rect 18966 41488 18972 41500
rect 19024 41488 19030 41540
rect 19061 41531 19119 41537
rect 19061 41497 19073 41531
rect 19107 41528 19119 41531
rect 19812 41528 19840 41559
rect 20070 41556 20076 41608
rect 20128 41556 20134 41608
rect 20441 41599 20499 41605
rect 20441 41565 20453 41599
rect 20487 41565 20499 41599
rect 20441 41559 20499 41565
rect 20162 41528 20168 41540
rect 19107 41500 19334 41528
rect 19812 41500 20168 41528
rect 19107 41497 19119 41500
rect 19061 41491 19119 41497
rect 18012 41432 18552 41460
rect 19306 41460 19334 41500
rect 20162 41488 20168 41500
rect 20220 41488 20226 41540
rect 20456 41528 20484 41559
rect 20530 41556 20536 41608
rect 20588 41596 20594 41608
rect 20625 41599 20683 41605
rect 20625 41596 20637 41599
rect 20588 41568 20637 41596
rect 20588 41556 20594 41568
rect 20625 41565 20637 41568
rect 20671 41565 20683 41599
rect 20625 41559 20683 41565
rect 22373 41599 22431 41605
rect 22373 41565 22385 41599
rect 22419 41596 22431 41599
rect 22646 41596 22652 41608
rect 22419 41568 22652 41596
rect 22419 41565 22431 41568
rect 22373 41559 22431 41565
rect 22646 41556 22652 41568
rect 22704 41556 22710 41608
rect 22741 41599 22799 41605
rect 22741 41565 22753 41599
rect 22787 41565 22799 41599
rect 22741 41559 22799 41565
rect 20456 41500 20852 41528
rect 20456 41460 20484 41500
rect 20824 41472 20852 41500
rect 21450 41488 21456 41540
rect 21508 41528 21514 41540
rect 22005 41531 22063 41537
rect 22005 41528 22017 41531
rect 21508 41500 22017 41528
rect 21508 41488 21514 41500
rect 22005 41497 22017 41500
rect 22051 41497 22063 41531
rect 22005 41491 22063 41497
rect 22094 41488 22100 41540
rect 22152 41528 22158 41540
rect 22152 41500 22324 41528
rect 22152 41488 22158 41500
rect 19306 41432 20484 41460
rect 18012 41420 18018 41432
rect 20806 41420 20812 41472
rect 20864 41460 20870 41472
rect 22296 41469 22324 41500
rect 22462 41488 22468 41540
rect 22520 41528 22526 41540
rect 22756 41528 22784 41559
rect 23474 41556 23480 41608
rect 23532 41596 23538 41608
rect 23845 41599 23903 41605
rect 23845 41596 23857 41599
rect 23532 41568 23857 41596
rect 23532 41556 23538 41568
rect 23845 41565 23857 41568
rect 23891 41565 23903 41599
rect 23845 41559 23903 41565
rect 24118 41556 24124 41608
rect 24176 41596 24182 41608
rect 24688 41605 24716 41636
rect 28534 41624 28540 41676
rect 28592 41624 28598 41676
rect 30653 41667 30711 41673
rect 30653 41633 30665 41667
rect 30699 41664 30711 41667
rect 32582 41664 32588 41676
rect 30699 41636 32588 41664
rect 30699 41633 30711 41636
rect 30653 41627 30711 41633
rect 32582 41624 32588 41636
rect 32640 41624 32646 41676
rect 32861 41667 32919 41673
rect 32861 41633 32873 41667
rect 32907 41664 32919 41667
rect 33318 41664 33324 41676
rect 32907 41636 33324 41664
rect 32907 41633 32919 41636
rect 32861 41627 32919 41633
rect 33318 41624 33324 41636
rect 33376 41624 33382 41676
rect 24397 41599 24455 41605
rect 24397 41596 24409 41599
rect 24176 41568 24409 41596
rect 24176 41556 24182 41568
rect 24397 41565 24409 41568
rect 24443 41565 24455 41599
rect 24397 41559 24455 41565
rect 24673 41599 24731 41605
rect 24673 41565 24685 41599
rect 24719 41565 24731 41599
rect 24673 41559 24731 41565
rect 26513 41599 26571 41605
rect 26513 41565 26525 41599
rect 26559 41596 26571 41599
rect 28721 41599 28779 41605
rect 28721 41596 28733 41599
rect 26559 41568 28733 41596
rect 26559 41565 26571 41568
rect 26513 41559 26571 41565
rect 28721 41565 28733 41568
rect 28767 41596 28779 41599
rect 29270 41596 29276 41608
rect 28767 41568 29276 41596
rect 28767 41565 28779 41568
rect 28721 41559 28779 41565
rect 29270 41556 29276 41568
rect 29328 41556 29334 41608
rect 22520 41500 22784 41528
rect 22520 41488 22526 41500
rect 24026 41488 24032 41540
rect 24084 41528 24090 41540
rect 24581 41531 24639 41537
rect 24581 41528 24593 41531
rect 24084 41500 24593 41528
rect 24084 41488 24090 41500
rect 24581 41497 24593 41500
rect 24627 41497 24639 41531
rect 24581 41491 24639 41497
rect 25133 41531 25191 41537
rect 25133 41497 25145 41531
rect 25179 41528 25191 41531
rect 25590 41528 25596 41540
rect 25179 41500 25596 41528
rect 25179 41497 25191 41500
rect 25133 41491 25191 41497
rect 25590 41488 25596 41500
rect 25648 41488 25654 41540
rect 25866 41488 25872 41540
rect 25924 41528 25930 41540
rect 26145 41531 26203 41537
rect 26145 41528 26157 41531
rect 25924 41500 26157 41528
rect 25924 41488 25930 41500
rect 26145 41497 26157 41500
rect 26191 41497 26203 41531
rect 26145 41491 26203 41497
rect 26234 41488 26240 41540
rect 26292 41528 26298 41540
rect 26329 41531 26387 41537
rect 26329 41528 26341 41531
rect 26292 41500 26341 41528
rect 26292 41488 26298 41500
rect 26329 41497 26341 41500
rect 26375 41497 26387 41531
rect 26329 41491 26387 41497
rect 26602 41488 26608 41540
rect 26660 41528 26666 41540
rect 26697 41531 26755 41537
rect 26697 41528 26709 41531
rect 26660 41500 26709 41528
rect 26660 41488 26666 41500
rect 26697 41497 26709 41500
rect 26743 41497 26755 41531
rect 26697 41491 26755 41497
rect 27065 41531 27123 41537
rect 27065 41497 27077 41531
rect 27111 41528 27123 41531
rect 27111 41500 27384 41528
rect 27111 41497 27123 41500
rect 27065 41491 27123 41497
rect 22189 41463 22247 41469
rect 22189 41460 22201 41463
rect 20864 41432 22201 41460
rect 20864 41420 20870 41432
rect 22189 41429 22201 41432
rect 22235 41429 22247 41463
rect 22189 41423 22247 41429
rect 22281 41463 22339 41469
rect 22281 41429 22293 41463
rect 22327 41429 22339 41463
rect 22281 41423 22339 41429
rect 22830 41420 22836 41472
rect 22888 41460 22894 41472
rect 22925 41463 22983 41469
rect 22925 41460 22937 41463
rect 22888 41432 22937 41460
rect 22888 41420 22894 41432
rect 22925 41429 22937 41432
rect 22971 41429 22983 41463
rect 22925 41423 22983 41429
rect 23198 41420 23204 41472
rect 23256 41460 23262 41472
rect 24394 41460 24400 41472
rect 23256 41432 24400 41460
rect 23256 41420 23262 41432
rect 24394 41420 24400 41432
rect 24452 41420 24458 41472
rect 25608 41460 25636 41488
rect 27246 41460 27252 41472
rect 25608 41432 27252 41460
rect 27246 41420 27252 41432
rect 27304 41420 27310 41472
rect 27356 41460 27384 41500
rect 27430 41488 27436 41540
rect 27488 41528 27494 41540
rect 28445 41531 28503 41537
rect 28445 41528 28457 41531
rect 27488 41500 28457 41528
rect 27488 41488 27494 41500
rect 28445 41497 28457 41500
rect 28491 41497 28503 41531
rect 32398 41528 32404 41540
rect 32154 41500 32404 41528
rect 28445 41491 28503 41497
rect 32398 41488 32404 41500
rect 32456 41488 32462 41540
rect 34422 41528 34428 41540
rect 34086 41500 34428 41528
rect 34422 41488 34428 41500
rect 34480 41488 34486 41540
rect 27706 41460 27712 41472
rect 27356 41432 27712 41460
rect 27706 41420 27712 41432
rect 27764 41420 27770 41472
rect 28905 41463 28963 41469
rect 28905 41429 28917 41463
rect 28951 41460 28963 41463
rect 31570 41460 31576 41472
rect 28951 41432 31576 41460
rect 28951 41429 28963 41432
rect 28905 41423 28963 41429
rect 31570 41420 31576 41432
rect 31628 41420 31634 41472
rect 33870 41420 33876 41472
rect 33928 41460 33934 41472
rect 34333 41463 34391 41469
rect 34333 41460 34345 41463
rect 33928 41432 34345 41460
rect 33928 41420 33934 41432
rect 34333 41429 34345 41432
rect 34379 41429 34391 41463
rect 34333 41423 34391 41429
rect 1104 41370 41400 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 41400 41370
rect 1104 41296 41400 41318
rect 11054 41256 11060 41268
rect 9232 41228 11060 41256
rect 9232 41061 9260 41228
rect 11054 41216 11060 41228
rect 11112 41216 11118 41268
rect 11149 41259 11207 41265
rect 11149 41225 11161 41259
rect 11195 41256 11207 41259
rect 11422 41256 11428 41268
rect 11195 41228 11428 41256
rect 11195 41225 11207 41228
rect 11149 41219 11207 41225
rect 11422 41216 11428 41228
rect 11480 41216 11486 41268
rect 13814 41216 13820 41268
rect 13872 41256 13878 41268
rect 14277 41259 14335 41265
rect 14277 41256 14289 41259
rect 13872 41228 14289 41256
rect 13872 41216 13878 41228
rect 14277 41225 14289 41228
rect 14323 41225 14335 41259
rect 14277 41219 14335 41225
rect 14645 41259 14703 41265
rect 14645 41225 14657 41259
rect 14691 41256 14703 41259
rect 15010 41256 15016 41268
rect 14691 41228 15016 41256
rect 14691 41225 14703 41228
rect 14645 41219 14703 41225
rect 15010 41216 15016 41228
rect 15068 41216 15074 41268
rect 15654 41216 15660 41268
rect 15712 41256 15718 41268
rect 17681 41259 17739 41265
rect 15712 41228 17540 41256
rect 15712 41216 15718 41228
rect 16393 41191 16451 41197
rect 10888 41160 16344 41188
rect 10888 41132 10916 41160
rect 10594 41080 10600 41132
rect 10652 41080 10658 41132
rect 10870 41080 10876 41132
rect 10928 41080 10934 41132
rect 11333 41123 11391 41129
rect 11333 41089 11345 41123
rect 11379 41120 11391 41123
rect 12713 41123 12771 41129
rect 11379 41092 12388 41120
rect 11379 41089 11391 41092
rect 11333 41083 11391 41089
rect 9217 41055 9275 41061
rect 9217 41021 9229 41055
rect 9263 41021 9275 41055
rect 9217 41015 9275 41021
rect 9490 41012 9496 41064
rect 9548 41012 9554 41064
rect 11609 41055 11667 41061
rect 11609 41021 11621 41055
rect 11655 41052 11667 41055
rect 11698 41052 11704 41064
rect 11655 41024 11704 41052
rect 11655 41021 11667 41024
rect 11609 41015 11667 41021
rect 11698 41012 11704 41024
rect 11756 41012 11762 41064
rect 12360 40993 12388 41092
rect 12713 41089 12725 41123
rect 12759 41120 12771 41123
rect 13446 41120 13452 41132
rect 12759 41092 13452 41120
rect 12759 41089 12771 41092
rect 12713 41083 12771 41089
rect 13446 41080 13452 41092
rect 13504 41080 13510 41132
rect 13556 41092 14964 41120
rect 12802 41012 12808 41064
rect 12860 41012 12866 41064
rect 12986 41012 12992 41064
rect 13044 41052 13050 41064
rect 13556 41052 13584 41092
rect 13044 41024 13584 41052
rect 13044 41012 13050 41024
rect 14734 41012 14740 41064
rect 14792 41012 14798 41064
rect 14936 41061 14964 41092
rect 15378 41080 15384 41132
rect 15436 41120 15442 41132
rect 15580 41129 15608 41160
rect 15473 41123 15531 41129
rect 15473 41120 15485 41123
rect 15436 41092 15485 41120
rect 15436 41080 15442 41092
rect 15473 41089 15485 41092
rect 15519 41089 15531 41123
rect 15473 41083 15531 41089
rect 15565 41123 15623 41129
rect 15565 41089 15577 41123
rect 15611 41089 15623 41123
rect 15565 41083 15623 41089
rect 14921 41055 14979 41061
rect 14921 41021 14933 41055
rect 14967 41052 14979 41055
rect 15488 41052 15516 41083
rect 15654 41080 15660 41132
rect 15712 41080 15718 41132
rect 15746 41080 15752 41132
rect 15804 41120 15810 41132
rect 15841 41123 15899 41129
rect 15841 41120 15853 41123
rect 15804 41092 15853 41120
rect 15804 41080 15810 41092
rect 15841 41089 15853 41092
rect 15887 41089 15899 41123
rect 15841 41083 15899 41089
rect 16209 41123 16267 41129
rect 16209 41089 16221 41123
rect 16255 41089 16267 41123
rect 16209 41083 16267 41089
rect 16224 41052 16252 41083
rect 14967 41024 15332 41052
rect 15488 41024 16252 41052
rect 14967 41021 14979 41024
rect 14921 41015 14979 41021
rect 12161 40987 12219 40993
rect 12161 40984 12173 40987
rect 10520 40956 12173 40984
rect 10226 40876 10232 40928
rect 10284 40916 10290 40928
rect 10520 40916 10548 40956
rect 12161 40953 12173 40956
rect 12207 40953 12219 40987
rect 12161 40947 12219 40953
rect 12345 40987 12403 40993
rect 12345 40953 12357 40987
rect 12391 40953 12403 40987
rect 12345 40947 12403 40953
rect 10284 40888 10548 40916
rect 10965 40919 11023 40925
rect 10284 40876 10290 40888
rect 10965 40885 10977 40919
rect 11011 40916 11023 40919
rect 11698 40916 11704 40928
rect 11011 40888 11704 40916
rect 11011 40885 11023 40888
rect 10965 40879 11023 40885
rect 11698 40876 11704 40888
rect 11756 40876 11762 40928
rect 15194 40876 15200 40928
rect 15252 40876 15258 40928
rect 15304 40916 15332 41024
rect 16206 40944 16212 40996
rect 16264 40944 16270 40996
rect 16316 40984 16344 41160
rect 16393 41157 16405 41191
rect 16439 41188 16451 41191
rect 17310 41188 17316 41200
rect 16439 41160 17316 41188
rect 16439 41157 16451 41160
rect 16393 41151 16451 41157
rect 17310 41148 17316 41160
rect 17368 41148 17374 41200
rect 17512 41188 17540 41228
rect 17681 41225 17693 41259
rect 17727 41256 17739 41259
rect 21726 41256 21732 41268
rect 17727 41228 18184 41256
rect 17727 41225 17739 41228
rect 17681 41219 17739 41225
rect 17512 41160 17908 41188
rect 17880 41132 17908 41160
rect 18046 41148 18052 41200
rect 18104 41148 18110 41200
rect 16485 41123 16543 41129
rect 16485 41089 16497 41123
rect 16531 41089 16543 41123
rect 16485 41083 16543 41089
rect 16500 41052 16528 41083
rect 16758 41080 16764 41132
rect 16816 41080 16822 41132
rect 17126 41080 17132 41132
rect 17184 41080 17190 41132
rect 17586 41123 17592 41132
rect 17428 41120 17592 41123
rect 17420 41095 17592 41120
rect 17420 41092 17456 41095
rect 17310 41052 17316 41064
rect 16500 41024 17316 41052
rect 17310 41012 17316 41024
rect 17368 41012 17374 41064
rect 17420 41061 17448 41092
rect 17586 41080 17592 41095
rect 17644 41080 17650 41132
rect 17862 41080 17868 41132
rect 17920 41080 17926 41132
rect 17954 41080 17960 41132
rect 18012 41080 18018 41132
rect 18156 41129 18184 41228
rect 20548 41228 21732 41256
rect 18322 41148 18328 41200
rect 18380 41188 18386 41200
rect 18380 41160 20024 41188
rect 18380 41148 18386 41160
rect 18141 41123 18199 41129
rect 18141 41089 18153 41123
rect 18187 41120 18199 41123
rect 18506 41120 18512 41132
rect 18187 41092 18512 41120
rect 18187 41089 18199 41092
rect 18141 41083 18199 41089
rect 18506 41080 18512 41092
rect 18564 41080 18570 41132
rect 18598 41080 18604 41132
rect 18656 41080 18662 41132
rect 19076 41129 19104 41160
rect 19061 41123 19119 41129
rect 19061 41089 19073 41123
rect 19107 41089 19119 41123
rect 19061 41083 19119 41089
rect 19150 41080 19156 41132
rect 19208 41120 19214 41132
rect 19685 41123 19743 41129
rect 19685 41120 19697 41123
rect 19208 41092 19697 41120
rect 19208 41080 19214 41092
rect 19685 41089 19697 41092
rect 19731 41089 19743 41123
rect 19685 41083 19743 41089
rect 19794 41080 19800 41132
rect 19852 41080 19858 41132
rect 19889 41123 19947 41129
rect 19889 41089 19901 41123
rect 19935 41118 19947 41123
rect 19996 41118 20024 41160
rect 20346 41148 20352 41200
rect 20404 41188 20410 41200
rect 20548 41197 20576 41228
rect 21726 41216 21732 41228
rect 21784 41216 21790 41268
rect 22002 41216 22008 41268
rect 22060 41256 22066 41268
rect 22646 41256 22652 41268
rect 22060 41228 22652 41256
rect 22060 41216 22066 41228
rect 22646 41216 22652 41228
rect 22704 41216 22710 41268
rect 24581 41259 24639 41265
rect 24581 41225 24593 41259
rect 24627 41256 24639 41259
rect 24627 41228 25268 41256
rect 24627 41225 24639 41228
rect 24581 41219 24639 41225
rect 25240 41197 25268 41228
rect 25314 41216 25320 41268
rect 25372 41256 25378 41268
rect 25869 41259 25927 41265
rect 25869 41256 25881 41259
rect 25372 41228 25881 41256
rect 25372 41216 25378 41228
rect 25869 41225 25881 41228
rect 25915 41225 25927 41259
rect 25869 41219 25927 41225
rect 26326 41216 26332 41268
rect 26384 41256 26390 41268
rect 26602 41256 26608 41268
rect 26384 41228 26608 41256
rect 26384 41216 26390 41228
rect 26602 41216 26608 41228
rect 26660 41256 26666 41268
rect 26786 41256 26792 41268
rect 26660 41228 26792 41256
rect 26660 41216 26666 41228
rect 26786 41216 26792 41228
rect 26844 41216 26850 41268
rect 27246 41216 27252 41268
rect 27304 41256 27310 41268
rect 29454 41256 29460 41268
rect 27304 41228 28948 41256
rect 27304 41216 27310 41228
rect 20533 41191 20591 41197
rect 20533 41188 20545 41191
rect 20404 41160 20545 41188
rect 20404 41148 20410 41160
rect 20533 41157 20545 41160
rect 20579 41157 20591 41191
rect 24305 41191 24363 41197
rect 24305 41188 24317 41191
rect 20533 41151 20591 41157
rect 20916 41160 23244 41188
rect 19935 41090 20024 41118
rect 19935 41089 19947 41090
rect 19889 41083 19947 41089
rect 20070 41080 20076 41132
rect 20128 41080 20134 41132
rect 20162 41080 20168 41132
rect 20220 41080 20226 41132
rect 20438 41080 20444 41132
rect 20496 41080 20502 41132
rect 20806 41080 20812 41132
rect 20864 41120 20870 41132
rect 20916 41129 20944 41160
rect 20901 41123 20959 41129
rect 20901 41120 20913 41123
rect 20864 41092 20913 41120
rect 20864 41080 20870 41092
rect 20901 41089 20913 41092
rect 20947 41089 20959 41123
rect 20901 41083 20959 41089
rect 20993 41123 21051 41129
rect 20993 41089 21005 41123
rect 21039 41120 21051 41123
rect 21082 41120 21088 41132
rect 21039 41092 21088 41120
rect 21039 41089 21051 41092
rect 20993 41083 21051 41089
rect 21082 41080 21088 41092
rect 21140 41080 21146 41132
rect 21836 41129 21864 41160
rect 23216 41129 23244 41160
rect 23584 41160 24317 41188
rect 21821 41123 21879 41129
rect 21821 41089 21833 41123
rect 21867 41089 21879 41123
rect 21821 41083 21879 41089
rect 22005 41123 22063 41129
rect 22005 41089 22017 41123
rect 22051 41120 22063 41123
rect 23201 41123 23259 41129
rect 22051 41092 22140 41120
rect 22051 41089 22063 41092
rect 22005 41083 22063 41089
rect 17405 41055 17463 41061
rect 17405 41021 17417 41055
rect 17451 41021 17463 41055
rect 17405 41015 17463 41021
rect 17494 41012 17500 41064
rect 17552 41012 17558 41064
rect 17773 41055 17831 41061
rect 17773 41021 17785 41055
rect 17819 41052 17831 41055
rect 18046 41052 18052 41064
rect 17819 41024 18052 41052
rect 17819 41021 17831 41024
rect 17773 41015 17831 41021
rect 18046 41012 18052 41024
rect 18104 41012 18110 41064
rect 18414 41012 18420 41064
rect 18472 41012 18478 41064
rect 19242 41012 19248 41064
rect 19300 41012 19306 41064
rect 19334 41012 19340 41064
rect 19392 41052 19398 41064
rect 19429 41055 19487 41061
rect 19429 41052 19441 41055
rect 19392 41024 19441 41052
rect 19392 41012 19398 41024
rect 19429 41021 19441 41024
rect 19475 41021 19487 41055
rect 20180 41052 20208 41080
rect 21450 41052 21456 41064
rect 20180 41024 21456 41052
rect 19429 41015 19487 41021
rect 21450 41012 21456 41024
rect 21508 41012 21514 41064
rect 18138 40984 18144 40996
rect 16316 40956 17356 40984
rect 15746 40916 15752 40928
rect 15304 40888 15752 40916
rect 15746 40876 15752 40888
rect 15804 40876 15810 40928
rect 16666 40876 16672 40928
rect 16724 40916 16730 40928
rect 17221 40919 17279 40925
rect 17221 40916 17233 40919
rect 16724 40888 17233 40916
rect 16724 40876 16730 40888
rect 17221 40885 17233 40888
rect 17267 40885 17279 40919
rect 17328 40916 17356 40956
rect 17972 40956 18144 40984
rect 17972 40916 18000 40956
rect 18138 40944 18144 40956
rect 18196 40984 18202 40996
rect 19702 40984 19708 40996
rect 18196 40956 19708 40984
rect 18196 40944 18202 40956
rect 19702 40944 19708 40956
rect 19760 40944 19766 40996
rect 19886 40944 19892 40996
rect 19944 40984 19950 40996
rect 22112 40984 22140 41092
rect 23201 41089 23213 41123
rect 23247 41089 23259 41123
rect 23201 41083 23259 41089
rect 23382 41080 23388 41132
rect 23440 41120 23446 41132
rect 23584 41129 23612 41160
rect 24305 41157 24317 41160
rect 24351 41157 24363 41191
rect 24305 41151 24363 41157
rect 25225 41191 25283 41197
rect 25225 41157 25237 41191
rect 25271 41188 25283 41191
rect 25682 41188 25688 41200
rect 25271 41160 25688 41188
rect 25271 41157 25283 41160
rect 25225 41151 25283 41157
rect 25682 41148 25688 41160
rect 25740 41188 25746 41200
rect 25777 41191 25835 41197
rect 25777 41188 25789 41191
rect 25740 41160 25789 41188
rect 25740 41148 25746 41160
rect 25777 41157 25789 41160
rect 25823 41157 25835 41191
rect 26234 41188 26240 41200
rect 25777 41151 25835 41157
rect 26068 41160 26240 41188
rect 23569 41123 23627 41129
rect 23569 41120 23581 41123
rect 23440 41092 23581 41120
rect 23440 41080 23446 41092
rect 23569 41089 23581 41092
rect 23615 41089 23627 41123
rect 23569 41083 23627 41089
rect 25038 41080 25044 41132
rect 25096 41080 25102 41132
rect 25314 41080 25320 41132
rect 25372 41080 25378 41132
rect 25406 41080 25412 41132
rect 25464 41080 25470 41132
rect 22370 41012 22376 41064
rect 22428 41052 22434 41064
rect 22465 41055 22523 41061
rect 22465 41052 22477 41055
rect 22428 41024 22477 41052
rect 22428 41012 22434 41024
rect 22465 41021 22477 41024
rect 22511 41021 22523 41055
rect 22465 41015 22523 41021
rect 22646 41012 22652 41064
rect 22704 41052 22710 41064
rect 23400 41052 23428 41080
rect 22704 41024 23428 41052
rect 22704 41012 22710 41024
rect 23934 41012 23940 41064
rect 23992 41012 23998 41064
rect 24118 41012 24124 41064
rect 24176 41052 24182 41064
rect 24213 41055 24271 41061
rect 24213 41052 24225 41055
rect 24176 41024 24225 41052
rect 24176 41012 24182 41024
rect 24213 41021 24225 41024
rect 24259 41021 24271 41055
rect 24213 41015 24271 41021
rect 24394 41012 24400 41064
rect 24452 41061 24458 41064
rect 24452 41055 24480 41061
rect 24468 41021 24480 41055
rect 24452 41015 24480 41021
rect 24452 41012 24458 41015
rect 19944 40956 22140 40984
rect 19944 40944 19950 40956
rect 22112 40928 22140 40956
rect 22925 40987 22983 40993
rect 22925 40953 22937 40987
rect 22971 40984 22983 40987
rect 23014 40984 23020 40996
rect 22971 40956 23020 40984
rect 22971 40953 22983 40956
rect 22925 40947 22983 40953
rect 23014 40944 23020 40956
rect 23072 40984 23078 40996
rect 25056 40984 25084 41080
rect 23072 40956 25084 40984
rect 25593 40987 25651 40993
rect 23072 40944 23078 40956
rect 25593 40953 25605 40987
rect 25639 40984 25651 40987
rect 26068 40984 26096 41160
rect 26234 41148 26240 41160
rect 26292 41148 26298 41200
rect 28920 41197 28948 41228
rect 29012 41228 29460 41256
rect 29012 41197 29040 41228
rect 29454 41216 29460 41228
rect 29512 41216 29518 41268
rect 28905 41191 28963 41197
rect 28465 41160 28856 41188
rect 28465 41132 28493 41160
rect 26329 41123 26387 41129
rect 26329 41120 26341 41123
rect 25639 40956 26096 40984
rect 26160 41092 26341 41120
rect 26160 40984 26188 41092
rect 26329 41089 26341 41092
rect 26375 41089 26387 41123
rect 26329 41083 26387 41089
rect 26602 41080 26608 41132
rect 26660 41080 26666 41132
rect 26878 41080 26884 41132
rect 26936 41120 26942 41132
rect 26973 41123 27031 41129
rect 26973 41120 26985 41123
rect 26936 41092 26985 41120
rect 26936 41080 26942 41092
rect 26973 41089 26985 41092
rect 27019 41089 27031 41123
rect 26973 41083 27031 41089
rect 27154 41080 27160 41132
rect 27212 41080 27218 41132
rect 27246 41080 27252 41132
rect 27304 41080 27310 41132
rect 27341 41123 27399 41129
rect 27341 41089 27353 41123
rect 27387 41120 27399 41123
rect 27617 41123 27675 41129
rect 27617 41120 27629 41123
rect 27387 41092 27629 41120
rect 27387 41089 27399 41092
rect 27341 41083 27399 41089
rect 27617 41089 27629 41092
rect 27663 41089 27675 41123
rect 27617 41083 27675 41089
rect 27985 41123 28043 41129
rect 27985 41089 27997 41123
rect 28031 41089 28043 41123
rect 27985 41083 28043 41089
rect 26510 41012 26516 41064
rect 26568 41012 26574 41064
rect 26786 41012 26792 41064
rect 26844 41052 26850 41064
rect 27356 41052 27384 41083
rect 28000 41052 28028 41083
rect 28074 41080 28080 41132
rect 28132 41080 28138 41132
rect 28166 41080 28172 41132
rect 28224 41120 28230 41132
rect 28261 41123 28319 41129
rect 28261 41120 28273 41123
rect 28224 41092 28273 41120
rect 28224 41080 28230 41092
rect 28261 41089 28273 41092
rect 28307 41089 28319 41123
rect 28261 41083 28319 41089
rect 28350 41080 28356 41132
rect 28408 41080 28414 41132
rect 28442 41080 28448 41132
rect 28500 41129 28506 41132
rect 28500 41120 28508 41129
rect 28500 41092 28545 41120
rect 28500 41083 28508 41092
rect 28500 41080 28506 41083
rect 28718 41080 28724 41132
rect 28776 41080 28782 41132
rect 28828 41120 28856 41160
rect 28905 41157 28917 41191
rect 28951 41157 28963 41191
rect 28905 41151 28963 41157
rect 28997 41191 29055 41197
rect 28997 41157 29009 41191
rect 29043 41157 29055 41191
rect 28997 41151 29055 41157
rect 29270 41148 29276 41200
rect 29328 41188 29334 41200
rect 31113 41191 31171 41197
rect 31113 41188 31125 41191
rect 29328 41160 29684 41188
rect 29328 41148 29334 41160
rect 29656 41129 29684 41160
rect 29748 41160 31125 41188
rect 29748 41132 29776 41160
rect 31113 41157 31125 41160
rect 31159 41157 31171 41191
rect 40862 41188 40868 41200
rect 31113 41151 31171 41157
rect 40328 41160 40868 41188
rect 29089 41123 29147 41129
rect 29089 41120 29101 41123
rect 28828 41092 29101 41120
rect 29089 41089 29101 41092
rect 29135 41089 29147 41123
rect 29089 41083 29147 41089
rect 29365 41123 29423 41129
rect 29365 41089 29377 41123
rect 29411 41120 29423 41123
rect 29641 41123 29699 41129
rect 29411 41092 29592 41120
rect 29411 41089 29423 41092
rect 29365 41083 29423 41089
rect 28534 41052 28540 41064
rect 26844 41024 27384 41052
rect 27540 41024 28540 41052
rect 26844 41012 26850 41024
rect 27540 40993 27568 41024
rect 28534 41012 28540 41024
rect 28592 41012 28598 41064
rect 29457 41055 29515 41061
rect 29457 41052 29469 41055
rect 28644 41024 29469 41052
rect 27525 40987 27583 40993
rect 26160 40956 27476 40984
rect 25639 40953 25651 40956
rect 25593 40947 25651 40953
rect 17328 40888 18000 40916
rect 17221 40879 17279 40885
rect 18690 40876 18696 40928
rect 18748 40916 18754 40928
rect 21082 40916 21088 40928
rect 18748 40888 21088 40916
rect 18748 40876 18754 40888
rect 21082 40876 21088 40888
rect 21140 40876 21146 40928
rect 22094 40876 22100 40928
rect 22152 40876 22158 40928
rect 22189 40919 22247 40925
rect 22189 40885 22201 40919
rect 22235 40916 22247 40919
rect 22738 40916 22744 40928
rect 22235 40888 22744 40916
rect 22235 40885 22247 40888
rect 22189 40879 22247 40885
rect 22738 40876 22744 40888
rect 22796 40876 22802 40928
rect 24762 40876 24768 40928
rect 24820 40916 24826 40928
rect 26160 40916 26188 40956
rect 24820 40888 26188 40916
rect 24820 40876 24826 40888
rect 26234 40876 26240 40928
rect 26292 40916 26298 40928
rect 26329 40919 26387 40925
rect 26329 40916 26341 40919
rect 26292 40888 26341 40916
rect 26292 40876 26298 40888
rect 26329 40885 26341 40888
rect 26375 40885 26387 40919
rect 26329 40879 26387 40885
rect 26786 40876 26792 40928
rect 26844 40876 26850 40928
rect 26878 40876 26884 40928
rect 26936 40916 26942 40928
rect 27154 40916 27160 40928
rect 26936 40888 27160 40916
rect 26936 40876 26942 40888
rect 27154 40876 27160 40888
rect 27212 40876 27218 40928
rect 27448 40916 27476 40956
rect 27525 40953 27537 40987
rect 27571 40953 27583 40987
rect 28644 40984 28672 41024
rect 29457 41021 29469 41024
rect 29503 41021 29515 41055
rect 29564 41052 29592 41092
rect 29641 41089 29653 41123
rect 29687 41089 29699 41123
rect 29641 41083 29699 41089
rect 29730 41080 29736 41132
rect 29788 41080 29794 41132
rect 30558 41080 30564 41132
rect 30616 41080 30622 41132
rect 30745 41123 30803 41129
rect 30745 41089 30757 41123
rect 30791 41089 30803 41123
rect 30745 41083 30803 41089
rect 30576 41052 30604 41080
rect 29564 41024 30604 41052
rect 29457 41015 29515 41021
rect 30650 41012 30656 41064
rect 30708 41012 30714 41064
rect 30760 41052 30788 41083
rect 31662 41080 31668 41132
rect 31720 41120 31726 41132
rect 32125 41123 32183 41129
rect 32125 41120 32137 41123
rect 31720 41092 32137 41120
rect 31720 41080 31726 41092
rect 32125 41089 32137 41092
rect 32171 41120 32183 41123
rect 34606 41120 34612 41132
rect 32171 41092 34612 41120
rect 32171 41089 32183 41092
rect 32125 41083 32183 41089
rect 34606 41080 34612 41092
rect 34664 41080 34670 41132
rect 40328 41129 40356 41160
rect 40862 41148 40868 41160
rect 40920 41148 40926 41200
rect 40313 41123 40371 41129
rect 40313 41089 40325 41123
rect 40359 41089 40371 41123
rect 40313 41083 40371 41089
rect 40589 41123 40647 41129
rect 40589 41089 40601 41123
rect 40635 41120 40647 41123
rect 41230 41120 41236 41132
rect 40635 41092 41236 41120
rect 40635 41089 40647 41092
rect 40589 41083 40647 41089
rect 41230 41080 41236 41092
rect 41288 41080 41294 41132
rect 30834 41052 30840 41064
rect 30760 41024 30840 41052
rect 30834 41012 30840 41024
rect 30892 41012 30898 41064
rect 31021 41055 31079 41061
rect 31021 41021 31033 41055
rect 31067 41021 31079 41055
rect 31021 41015 31079 41021
rect 27525 40947 27583 40953
rect 27724 40956 28672 40984
rect 29196 40956 29408 40984
rect 27724 40916 27752 40956
rect 27448 40888 27752 40916
rect 27801 40919 27859 40925
rect 27801 40885 27813 40919
rect 27847 40916 27859 40919
rect 28534 40916 28540 40928
rect 27847 40888 28540 40916
rect 27847 40885 27859 40888
rect 27801 40879 27859 40885
rect 28534 40876 28540 40888
rect 28592 40876 28598 40928
rect 28629 40919 28687 40925
rect 28629 40885 28641 40919
rect 28675 40916 28687 40919
rect 29196 40916 29224 40956
rect 28675 40888 29224 40916
rect 28675 40885 28687 40888
rect 28629 40879 28687 40885
rect 29270 40876 29276 40928
rect 29328 40876 29334 40928
rect 29380 40925 29408 40956
rect 30006 40944 30012 40996
rect 30064 40984 30070 40996
rect 31036 40984 31064 41015
rect 32398 41012 32404 41064
rect 32456 41052 32462 41064
rect 34422 41052 34428 41064
rect 32456 41024 34428 41052
rect 32456 41012 32462 41024
rect 34422 41012 34428 41024
rect 34480 41012 34486 41064
rect 40770 41012 40776 41064
rect 40828 41012 40834 41064
rect 30064 40956 31064 40984
rect 30064 40944 30070 40956
rect 29365 40919 29423 40925
rect 29365 40885 29377 40919
rect 29411 40885 29423 40919
rect 29365 40879 29423 40885
rect 29825 40919 29883 40925
rect 29825 40885 29837 40919
rect 29871 40916 29883 40919
rect 30374 40916 30380 40928
rect 29871 40888 30380 40916
rect 29871 40885 29883 40888
rect 29825 40879 29883 40885
rect 30374 40876 30380 40888
rect 30432 40876 30438 40928
rect 30466 40876 30472 40928
rect 30524 40876 30530 40928
rect 40402 40876 40408 40928
rect 40460 40876 40466 40928
rect 1104 40826 41400 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 41400 40826
rect 1104 40752 41400 40774
rect 9490 40672 9496 40724
rect 9548 40712 9554 40724
rect 9953 40715 10011 40721
rect 9953 40712 9965 40715
rect 9548 40684 9965 40712
rect 9548 40672 9554 40684
rect 9953 40681 9965 40684
rect 9999 40681 10011 40715
rect 9953 40675 10011 40681
rect 14734 40672 14740 40724
rect 14792 40712 14798 40724
rect 16393 40715 16451 40721
rect 16393 40712 16405 40715
rect 14792 40684 16405 40712
rect 14792 40672 14798 40684
rect 16393 40681 16405 40684
rect 16439 40681 16451 40715
rect 16393 40675 16451 40681
rect 17310 40672 17316 40724
rect 17368 40672 17374 40724
rect 18046 40672 18052 40724
rect 18104 40672 18110 40724
rect 19058 40672 19064 40724
rect 19116 40712 19122 40724
rect 20073 40715 20131 40721
rect 20073 40712 20085 40715
rect 19116 40684 20085 40712
rect 19116 40672 19122 40684
rect 20073 40681 20085 40684
rect 20119 40712 20131 40715
rect 20162 40712 20168 40724
rect 20119 40684 20168 40712
rect 20119 40681 20131 40684
rect 20073 40675 20131 40681
rect 20162 40672 20168 40684
rect 20220 40672 20226 40724
rect 20530 40672 20536 40724
rect 20588 40672 20594 40724
rect 21910 40672 21916 40724
rect 21968 40712 21974 40724
rect 21968 40684 22140 40712
rect 21968 40672 21974 40684
rect 15194 40604 15200 40656
rect 15252 40604 15258 40656
rect 15654 40644 15660 40656
rect 15580 40616 15660 40644
rect 11054 40536 11060 40588
rect 11112 40536 11118 40588
rect 11333 40579 11391 40585
rect 11333 40545 11345 40579
rect 11379 40576 11391 40579
rect 12618 40576 12624 40588
rect 11379 40548 12624 40576
rect 11379 40545 11391 40548
rect 11333 40539 11391 40545
rect 12618 40536 12624 40548
rect 12676 40536 12682 40588
rect 12805 40579 12863 40585
rect 12805 40545 12817 40579
rect 12851 40576 12863 40579
rect 12851 40548 13216 40576
rect 12851 40545 12863 40548
rect 12805 40539 12863 40545
rect 934 40468 940 40520
rect 992 40508 998 40520
rect 1397 40511 1455 40517
rect 1397 40508 1409 40511
rect 992 40480 1409 40508
rect 992 40468 998 40480
rect 1397 40477 1409 40480
rect 1443 40477 1455 40511
rect 1397 40471 1455 40477
rect 1670 40468 1676 40520
rect 1728 40468 1734 40520
rect 10137 40511 10195 40517
rect 10137 40477 10149 40511
rect 10183 40477 10195 40511
rect 10137 40471 10195 40477
rect 10152 40440 10180 40471
rect 10226 40468 10232 40520
rect 10284 40508 10290 40520
rect 10321 40511 10379 40517
rect 10321 40508 10333 40511
rect 10284 40480 10333 40508
rect 10284 40468 10290 40480
rect 10321 40477 10333 40480
rect 10367 40477 10379 40511
rect 10321 40471 10379 40477
rect 10410 40468 10416 40520
rect 10468 40508 10474 40520
rect 10468 40480 11008 40508
rect 10468 40468 10474 40480
rect 10980 40452 11008 40480
rect 12434 40468 12440 40520
rect 12492 40468 12498 40520
rect 13188 40517 13216 40548
rect 13446 40536 13452 40588
rect 13504 40576 13510 40588
rect 13504 40548 14412 40576
rect 13504 40536 13510 40548
rect 14384 40517 14412 40548
rect 13173 40511 13231 40517
rect 13173 40477 13185 40511
rect 13219 40508 13231 40511
rect 14093 40511 14151 40517
rect 14093 40508 14105 40511
rect 13219 40480 14105 40508
rect 13219 40477 13231 40480
rect 13173 40471 13231 40477
rect 14093 40477 14105 40480
rect 14139 40477 14151 40511
rect 14093 40471 14151 40477
rect 14369 40511 14427 40517
rect 14369 40477 14381 40511
rect 14415 40477 14427 40511
rect 14369 40471 14427 40477
rect 14550 40468 14556 40520
rect 14608 40468 14614 40520
rect 14829 40511 14887 40517
rect 14829 40477 14841 40511
rect 14875 40508 14887 40511
rect 15102 40508 15108 40520
rect 14875 40480 15108 40508
rect 14875 40477 14887 40480
rect 14829 40471 14887 40477
rect 15102 40468 15108 40480
rect 15160 40468 15166 40520
rect 10152 40412 10456 40440
rect 10428 40372 10456 40412
rect 10962 40400 10968 40452
rect 11020 40400 11026 40452
rect 15212 40440 15240 40604
rect 15381 40579 15439 40585
rect 15381 40545 15393 40579
rect 15427 40576 15439 40579
rect 15470 40576 15476 40588
rect 15427 40548 15476 40576
rect 15427 40545 15439 40548
rect 15381 40539 15439 40545
rect 15470 40536 15476 40548
rect 15528 40536 15534 40588
rect 15580 40585 15608 40616
rect 15654 40604 15660 40616
rect 15712 40604 15718 40656
rect 16574 40644 16580 40656
rect 15764 40616 16580 40644
rect 15565 40579 15623 40585
rect 15565 40545 15577 40579
rect 15611 40545 15623 40579
rect 15565 40539 15623 40545
rect 15764 40508 15792 40616
rect 16574 40604 16580 40616
rect 16632 40604 16638 40656
rect 16758 40604 16764 40656
rect 16816 40644 16822 40656
rect 18322 40644 18328 40656
rect 16816 40616 18328 40644
rect 16816 40604 16822 40616
rect 18322 40604 18328 40616
rect 18380 40604 18386 40656
rect 18506 40604 18512 40656
rect 18564 40644 18570 40656
rect 19610 40644 19616 40656
rect 18564 40616 19616 40644
rect 18564 40604 18570 40616
rect 19610 40604 19616 40616
rect 19668 40644 19674 40656
rect 20438 40644 20444 40656
rect 19668 40616 20444 40644
rect 19668 40604 19674 40616
rect 16776 40576 16804 40604
rect 15948 40548 16804 40576
rect 15948 40520 15976 40548
rect 16942 40536 16948 40588
rect 17000 40536 17006 40588
rect 17037 40579 17095 40585
rect 17037 40545 17049 40579
rect 17083 40576 17095 40579
rect 17126 40576 17132 40588
rect 17083 40548 17132 40576
rect 17083 40545 17095 40548
rect 17037 40539 17095 40545
rect 17126 40536 17132 40548
rect 17184 40536 17190 40588
rect 17862 40576 17868 40588
rect 17236 40548 17868 40576
rect 13648 40412 15240 40440
rect 15304 40480 15792 40508
rect 13648 40372 13676 40412
rect 10428 40344 13676 40372
rect 13722 40332 13728 40384
rect 13780 40332 13786 40384
rect 14182 40332 14188 40384
rect 14240 40332 14246 40384
rect 14458 40332 14464 40384
rect 14516 40372 14522 40384
rect 15304 40372 15332 40480
rect 15930 40468 15936 40520
rect 15988 40468 15994 40520
rect 16022 40468 16028 40520
rect 16080 40468 16086 40520
rect 16574 40468 16580 40520
rect 16632 40468 16638 40520
rect 16669 40511 16727 40517
rect 16669 40477 16681 40511
rect 16715 40508 16727 40511
rect 16960 40508 16988 40536
rect 17236 40517 17264 40548
rect 17862 40536 17868 40548
rect 17920 40576 17926 40588
rect 17920 40548 19564 40576
rect 17920 40536 17926 40548
rect 16715 40480 16988 40508
rect 17221 40511 17279 40517
rect 16715 40477 16727 40480
rect 16669 40471 16727 40477
rect 17221 40477 17233 40511
rect 17267 40477 17279 40511
rect 17405 40511 17463 40517
rect 17405 40508 17417 40511
rect 17221 40471 17279 40477
rect 17328 40480 17417 40508
rect 15562 40400 15568 40452
rect 15620 40440 15626 40452
rect 16117 40443 16175 40449
rect 16117 40440 16129 40443
rect 15620 40412 16129 40440
rect 15620 40400 15626 40412
rect 16117 40409 16129 40412
rect 16163 40409 16175 40443
rect 16117 40403 16175 40409
rect 16482 40400 16488 40452
rect 16540 40440 16546 40452
rect 16761 40443 16819 40449
rect 16761 40440 16773 40443
rect 16540 40412 16773 40440
rect 16540 40400 16546 40412
rect 16761 40409 16773 40412
rect 16807 40409 16819 40443
rect 16761 40403 16819 40409
rect 16899 40443 16957 40449
rect 16899 40409 16911 40443
rect 16945 40440 16957 40443
rect 17126 40440 17132 40452
rect 16945 40412 17132 40440
rect 16945 40409 16957 40412
rect 16899 40403 16957 40409
rect 17126 40400 17132 40412
rect 17184 40400 17190 40452
rect 17328 40384 17356 40480
rect 17405 40477 17417 40480
rect 17451 40477 17463 40511
rect 17405 40471 17463 40477
rect 17589 40511 17647 40517
rect 17589 40477 17601 40511
rect 17635 40508 17647 40511
rect 17770 40508 17776 40520
rect 17635 40480 17776 40508
rect 17635 40477 17647 40480
rect 17589 40471 17647 40477
rect 17770 40468 17776 40480
rect 17828 40468 17834 40520
rect 17957 40511 18015 40517
rect 17957 40477 17969 40511
rect 18003 40508 18015 40511
rect 18138 40508 18144 40520
rect 18003 40480 18144 40508
rect 18003 40477 18015 40480
rect 17957 40471 18015 40477
rect 18138 40468 18144 40480
rect 18196 40468 18202 40520
rect 18233 40511 18291 40517
rect 18233 40477 18245 40511
rect 18279 40477 18291 40511
rect 18233 40471 18291 40477
rect 18248 40440 18276 40471
rect 18690 40468 18696 40520
rect 18748 40468 18754 40520
rect 19242 40508 19248 40520
rect 18800 40480 19248 40508
rect 18800 40440 18828 40480
rect 19242 40468 19248 40480
rect 19300 40468 19306 40520
rect 19536 40517 19564 40548
rect 19521 40511 19579 40517
rect 19521 40477 19533 40511
rect 19567 40508 19579 40511
rect 19702 40508 19708 40520
rect 19567 40480 19708 40508
rect 19567 40477 19579 40480
rect 19521 40471 19579 40477
rect 19702 40468 19708 40480
rect 19760 40468 19766 40520
rect 19797 40511 19855 40517
rect 19797 40477 19809 40511
rect 19843 40477 19855 40511
rect 19904 40508 19932 40616
rect 20438 40604 20444 40616
rect 20496 40604 20502 40656
rect 21450 40604 21456 40656
rect 21508 40644 21514 40656
rect 22112 40644 22140 40684
rect 22186 40672 22192 40724
rect 22244 40672 22250 40724
rect 23109 40715 23167 40721
rect 23109 40712 23121 40715
rect 22296 40684 23121 40712
rect 22296 40644 22324 40684
rect 23109 40681 23121 40684
rect 23155 40681 23167 40715
rect 23109 40675 23167 40681
rect 23382 40672 23388 40724
rect 23440 40672 23446 40724
rect 24118 40712 24124 40724
rect 23492 40684 24124 40712
rect 21508 40616 22048 40644
rect 22112 40616 22324 40644
rect 21508 40604 21514 40616
rect 20456 40576 20484 40604
rect 22020 40588 22048 40616
rect 22370 40604 22376 40656
rect 22428 40644 22434 40656
rect 23201 40647 23259 40653
rect 23201 40644 23213 40647
rect 22428 40616 23213 40644
rect 22428 40604 22434 40616
rect 23201 40613 23213 40616
rect 23247 40613 23259 40647
rect 23201 40607 23259 40613
rect 21821 40579 21879 40585
rect 21821 40576 21833 40579
rect 20456 40548 21833 40576
rect 21821 40545 21833 40548
rect 21867 40576 21879 40579
rect 21910 40576 21916 40588
rect 21867 40548 21916 40576
rect 21867 40545 21879 40548
rect 21821 40539 21879 40545
rect 21910 40536 21916 40548
rect 21968 40536 21974 40588
rect 22002 40536 22008 40588
rect 22060 40536 22066 40588
rect 22925 40579 22983 40585
rect 22925 40545 22937 40579
rect 22971 40576 22983 40579
rect 23293 40579 23351 40585
rect 22971 40548 23244 40576
rect 22971 40545 22983 40548
rect 22925 40539 22983 40545
rect 19981 40511 20039 40517
rect 19981 40508 19993 40511
rect 19904 40480 19993 40508
rect 19797 40471 19855 40477
rect 19981 40477 19993 40480
rect 20027 40477 20039 40511
rect 19981 40471 20039 40477
rect 18248 40412 18828 40440
rect 19812 40440 19840 40471
rect 20070 40468 20076 40520
rect 20128 40508 20134 40520
rect 20349 40511 20407 40517
rect 20349 40510 20361 40511
rect 20272 40508 20361 40510
rect 20128 40482 20361 40508
rect 20128 40480 20300 40482
rect 20128 40468 20134 40480
rect 20349 40477 20361 40482
rect 20395 40477 20407 40511
rect 20349 40471 20407 40477
rect 20806 40468 20812 40520
rect 20864 40508 20870 40520
rect 21545 40511 21603 40517
rect 21545 40508 21557 40511
rect 20864 40480 21557 40508
rect 20864 40468 20870 40480
rect 21545 40477 21557 40480
rect 21591 40477 21603 40511
rect 21545 40471 21603 40477
rect 20254 40440 20260 40452
rect 19812 40412 20260 40440
rect 20254 40400 20260 40412
rect 20312 40400 20318 40452
rect 20824 40440 20852 40468
rect 20640 40412 20852 40440
rect 20901 40443 20959 40449
rect 14516 40344 15332 40372
rect 14516 40332 14522 40344
rect 15470 40332 15476 40384
rect 15528 40372 15534 40384
rect 15838 40372 15844 40384
rect 15528 40344 15844 40372
rect 15528 40332 15534 40344
rect 15838 40332 15844 40344
rect 15896 40332 15902 40384
rect 17310 40332 17316 40384
rect 17368 40332 17374 40384
rect 17402 40332 17408 40384
rect 17460 40372 17466 40384
rect 17770 40372 17776 40384
rect 17460 40344 17776 40372
rect 17460 40332 17466 40344
rect 17770 40332 17776 40344
rect 17828 40332 17834 40384
rect 18322 40332 18328 40384
rect 18380 40372 18386 40384
rect 18785 40375 18843 40381
rect 18785 40372 18797 40375
rect 18380 40344 18797 40372
rect 18380 40332 18386 40344
rect 18785 40341 18797 40344
rect 18831 40341 18843 40375
rect 18785 40335 18843 40341
rect 19337 40375 19395 40381
rect 19337 40341 19349 40375
rect 19383 40372 19395 40375
rect 19610 40372 19616 40384
rect 19383 40344 19616 40372
rect 19383 40341 19395 40344
rect 19337 40335 19395 40341
rect 19610 40332 19616 40344
rect 19668 40332 19674 40384
rect 19705 40375 19763 40381
rect 19705 40341 19717 40375
rect 19751 40372 19763 40375
rect 20640 40372 20668 40412
rect 20901 40409 20913 40443
rect 20947 40440 20959 40443
rect 21450 40440 21456 40452
rect 20947 40412 21456 40440
rect 20947 40409 20959 40412
rect 20901 40403 20959 40409
rect 21450 40400 21456 40412
rect 21508 40400 21514 40452
rect 22020 40449 22048 40536
rect 23216 40520 23244 40548
rect 23293 40545 23305 40579
rect 23339 40576 23351 40579
rect 23400 40576 23428 40672
rect 23492 40588 23520 40684
rect 24118 40672 24124 40684
rect 24176 40672 24182 40724
rect 25314 40712 25320 40724
rect 24437 40684 24808 40712
rect 23750 40604 23756 40656
rect 23808 40604 23814 40656
rect 24026 40604 24032 40656
rect 24084 40644 24090 40656
rect 24437 40644 24465 40684
rect 24084 40616 24465 40644
rect 24084 40604 24090 40616
rect 23339 40548 23428 40576
rect 23339 40545 23351 40548
rect 23293 40539 23351 40545
rect 23474 40536 23480 40588
rect 23532 40536 23538 40588
rect 24397 40579 24455 40585
rect 24397 40576 24409 40579
rect 23952 40548 24409 40576
rect 22462 40468 22468 40520
rect 22520 40468 22526 40520
rect 23017 40511 23075 40517
rect 23017 40477 23029 40511
rect 23063 40508 23075 40511
rect 23106 40508 23112 40520
rect 23063 40480 23112 40508
rect 23063 40477 23075 40480
rect 23017 40471 23075 40477
rect 23106 40468 23112 40480
rect 23164 40468 23170 40520
rect 23198 40468 23204 40520
rect 23256 40468 23262 40520
rect 23952 40517 23980 40548
rect 24397 40545 24409 40548
rect 24443 40545 24455 40579
rect 24397 40539 24455 40545
rect 24578 40536 24584 40588
rect 24636 40536 24642 40588
rect 24780 40585 24808 40684
rect 24872 40684 25320 40712
rect 24872 40585 24900 40684
rect 25314 40672 25320 40684
rect 25372 40672 25378 40724
rect 26970 40672 26976 40724
rect 27028 40712 27034 40724
rect 30006 40712 30012 40724
rect 27028 40684 30012 40712
rect 27028 40672 27034 40684
rect 30006 40672 30012 40684
rect 30064 40672 30070 40724
rect 30282 40672 30288 40724
rect 30340 40672 30346 40724
rect 30466 40672 30472 40724
rect 30524 40672 30530 40724
rect 40402 40712 40408 40724
rect 38948 40684 40408 40712
rect 25056 40616 27384 40644
rect 24765 40579 24823 40585
rect 24765 40545 24777 40579
rect 24811 40545 24823 40579
rect 24765 40539 24823 40545
rect 24857 40579 24915 40585
rect 24857 40545 24869 40579
rect 24903 40545 24915 40579
rect 24857 40539 24915 40545
rect 23937 40511 23995 40517
rect 23937 40477 23949 40511
rect 23983 40477 23995 40511
rect 23937 40471 23995 40477
rect 24210 40468 24216 40520
rect 24268 40468 24274 40520
rect 24670 40468 24676 40520
rect 24728 40468 24734 40520
rect 25056 40508 25084 40616
rect 25682 40536 25688 40588
rect 25740 40576 25746 40588
rect 25740 40548 26004 40576
rect 25740 40536 25746 40548
rect 24780 40480 25084 40508
rect 25133 40511 25191 40517
rect 22020 40443 22088 40449
rect 22020 40412 22042 40443
rect 22030 40409 22042 40412
rect 22076 40409 22088 40443
rect 22030 40403 22088 40409
rect 22370 40400 22376 40452
rect 22428 40400 22434 40452
rect 22557 40443 22615 40449
rect 22557 40409 22569 40443
rect 22603 40409 22615 40443
rect 22557 40403 22615 40409
rect 19751 40344 20668 40372
rect 19751 40341 19763 40344
rect 19705 40335 19763 40341
rect 20714 40332 20720 40384
rect 20772 40372 20778 40384
rect 20993 40375 21051 40381
rect 20993 40372 21005 40375
rect 20772 40344 21005 40372
rect 20772 40332 20778 40344
rect 20993 40341 21005 40344
rect 21039 40341 21051 40375
rect 20993 40335 21051 40341
rect 21082 40332 21088 40384
rect 21140 40372 21146 40384
rect 21910 40372 21916 40384
rect 21140 40344 21916 40372
rect 21140 40332 21146 40344
rect 21910 40332 21916 40344
rect 21968 40332 21974 40384
rect 22278 40332 22284 40384
rect 22336 40332 22342 40384
rect 22388 40372 22416 40400
rect 22572 40372 22600 40403
rect 22646 40400 22652 40452
rect 22704 40400 22710 40452
rect 22787 40443 22845 40449
rect 22787 40409 22799 40443
rect 22833 40440 22845 40443
rect 22922 40440 22928 40452
rect 22833 40412 22928 40440
rect 22833 40409 22845 40412
rect 22787 40403 22845 40409
rect 22922 40400 22928 40412
rect 22980 40400 22986 40452
rect 23290 40400 23296 40452
rect 23348 40440 23354 40452
rect 24780 40440 24808 40480
rect 25133 40477 25145 40511
rect 25179 40508 25191 40511
rect 25406 40508 25412 40520
rect 25179 40480 25412 40508
rect 25179 40477 25191 40480
rect 25133 40471 25191 40477
rect 23348 40412 24808 40440
rect 23348 40400 23354 40412
rect 24854 40400 24860 40452
rect 24912 40440 24918 40452
rect 25148 40440 25176 40471
rect 25406 40468 25412 40480
rect 25464 40468 25470 40520
rect 25774 40468 25780 40520
rect 25832 40517 25838 40520
rect 25976 40517 26004 40548
rect 25832 40511 25855 40517
rect 25843 40477 25855 40511
rect 25832 40471 25855 40477
rect 25961 40511 26019 40517
rect 25961 40477 25973 40511
rect 26007 40477 26019 40511
rect 25961 40471 26019 40477
rect 25832 40468 25838 40471
rect 26050 40468 26056 40520
rect 26108 40468 26114 40520
rect 26145 40511 26203 40517
rect 26145 40477 26157 40511
rect 26191 40477 26203 40511
rect 26145 40471 26203 40477
rect 24912 40412 25176 40440
rect 24912 40400 24918 40412
rect 22388 40344 22600 40372
rect 25317 40375 25375 40381
rect 25317 40341 25329 40375
rect 25363 40372 25375 40375
rect 25406 40372 25412 40384
rect 25363 40344 25412 40372
rect 25363 40341 25375 40344
rect 25317 40335 25375 40341
rect 25406 40332 25412 40344
rect 25464 40372 25470 40384
rect 26160 40372 26188 40471
rect 26510 40468 26516 40520
rect 26568 40508 26574 40520
rect 26970 40517 26976 40520
rect 26789 40511 26847 40517
rect 26789 40508 26801 40511
rect 26568 40480 26801 40508
rect 26568 40468 26574 40480
rect 26789 40477 26801 40480
rect 26835 40477 26847 40511
rect 26789 40471 26847 40477
rect 26937 40511 26976 40517
rect 26937 40477 26949 40511
rect 26937 40471 26976 40477
rect 26970 40468 26976 40471
rect 27028 40468 27034 40520
rect 27254 40511 27312 40517
rect 27254 40477 27266 40511
rect 27300 40477 27312 40511
rect 27356 40508 27384 40616
rect 27706 40604 27712 40656
rect 27764 40644 27770 40656
rect 27764 40616 29960 40644
rect 27764 40604 27770 40616
rect 28460 40548 28994 40576
rect 28460 40517 28488 40548
rect 28445 40511 28503 40517
rect 28445 40508 28457 40511
rect 27356 40480 28457 40508
rect 27254 40471 27312 40477
rect 28445 40477 28457 40480
rect 28491 40477 28503 40511
rect 28445 40471 28503 40477
rect 26694 40400 26700 40452
rect 26752 40440 26758 40452
rect 27065 40443 27123 40449
rect 27065 40440 27077 40443
rect 26752 40412 27077 40440
rect 26752 40400 26758 40412
rect 27065 40409 27077 40412
rect 27111 40409 27123 40443
rect 27065 40403 27123 40409
rect 27154 40400 27160 40452
rect 27212 40400 27218 40452
rect 27269 40440 27297 40471
rect 28534 40468 28540 40520
rect 28592 40508 28598 40520
rect 28813 40511 28871 40517
rect 28813 40508 28825 40511
rect 28592 40480 28825 40508
rect 28592 40468 28598 40480
rect 28813 40477 28825 40480
rect 28859 40477 28871 40511
rect 28966 40508 28994 40548
rect 29362 40508 29368 40520
rect 28966 40480 29368 40508
rect 28813 40471 28871 40477
rect 29362 40468 29368 40480
rect 29420 40508 29426 40520
rect 29932 40517 29960 40616
rect 30484 40576 30512 40672
rect 30300 40548 30512 40576
rect 30300 40517 30328 40548
rect 32582 40536 32588 40588
rect 32640 40576 32646 40588
rect 32769 40579 32827 40585
rect 32769 40576 32781 40579
rect 32640 40548 32781 40576
rect 32640 40536 32646 40548
rect 32769 40545 32781 40548
rect 32815 40576 32827 40579
rect 33594 40576 33600 40588
rect 32815 40548 33600 40576
rect 32815 40545 32827 40548
rect 32769 40539 32827 40545
rect 33594 40536 33600 40548
rect 33652 40536 33658 40588
rect 37921 40579 37979 40585
rect 37921 40545 37933 40579
rect 37967 40576 37979 40579
rect 38948 40576 38976 40684
rect 40402 40672 40408 40684
rect 40460 40672 40466 40724
rect 37967 40548 38976 40576
rect 39393 40579 39451 40585
rect 37967 40545 37979 40548
rect 37921 40539 37979 40545
rect 39393 40545 39405 40579
rect 39439 40576 39451 40579
rect 39853 40579 39911 40585
rect 39853 40576 39865 40579
rect 39439 40548 39865 40576
rect 39439 40545 39451 40548
rect 39393 40539 39451 40545
rect 39853 40545 39865 40548
rect 39899 40545 39911 40579
rect 39853 40539 39911 40545
rect 29549 40511 29607 40517
rect 29549 40508 29561 40511
rect 29420 40480 29561 40508
rect 29420 40468 29426 40480
rect 29549 40477 29561 40480
rect 29595 40477 29607 40511
rect 29549 40471 29607 40477
rect 29917 40511 29975 40517
rect 29917 40477 29929 40511
rect 29963 40477 29975 40511
rect 29917 40471 29975 40477
rect 30285 40511 30343 40517
rect 30285 40477 30297 40511
rect 30331 40477 30343 40511
rect 30285 40471 30343 40477
rect 30377 40511 30435 40517
rect 30377 40477 30389 40511
rect 30423 40477 30435 40511
rect 30377 40471 30435 40477
rect 27706 40440 27712 40452
rect 27269 40412 27712 40440
rect 27706 40400 27712 40412
rect 27764 40400 27770 40452
rect 28074 40400 28080 40452
rect 28132 40440 28138 40452
rect 28629 40443 28687 40449
rect 28629 40440 28641 40443
rect 28132 40412 28641 40440
rect 28132 40400 28138 40412
rect 28629 40409 28641 40412
rect 28675 40409 28687 40443
rect 28629 40403 28687 40409
rect 28718 40400 28724 40452
rect 28776 40400 28782 40452
rect 29730 40400 29736 40452
rect 29788 40400 29794 40452
rect 29822 40400 29828 40452
rect 29880 40400 29886 40452
rect 30392 40440 30420 40471
rect 37642 40468 37648 40520
rect 37700 40468 37706 40520
rect 29932 40412 30420 40440
rect 25464 40344 26188 40372
rect 26329 40375 26387 40381
rect 25464 40332 25470 40344
rect 26329 40341 26341 40375
rect 26375 40372 26387 40375
rect 26970 40372 26976 40384
rect 26375 40344 26976 40372
rect 26375 40341 26387 40344
rect 26329 40335 26387 40341
rect 26970 40332 26976 40344
rect 27028 40332 27034 40384
rect 27433 40375 27491 40381
rect 27433 40341 27445 40375
rect 27479 40372 27491 40375
rect 27522 40372 27528 40384
rect 27479 40344 27528 40372
rect 27479 40341 27491 40344
rect 27433 40335 27491 40341
rect 27522 40332 27528 40344
rect 27580 40332 27586 40384
rect 28997 40375 29055 40381
rect 28997 40341 29009 40375
rect 29043 40372 29055 40375
rect 29178 40372 29184 40384
rect 29043 40344 29184 40372
rect 29043 40341 29055 40344
rect 28997 40335 29055 40341
rect 29178 40332 29184 40344
rect 29236 40372 29242 40384
rect 29932 40372 29960 40412
rect 32214 40400 32220 40452
rect 32272 40400 32278 40452
rect 32401 40443 32459 40449
rect 32401 40409 32413 40443
rect 32447 40440 32459 40443
rect 32766 40440 32772 40452
rect 32447 40412 32772 40440
rect 32447 40409 32459 40412
rect 32401 40403 32459 40409
rect 29236 40344 29960 40372
rect 30101 40375 30159 40381
rect 29236 40332 29242 40344
rect 30101 40341 30113 40375
rect 30147 40372 30159 40375
rect 30466 40372 30472 40384
rect 30147 40344 30472 40372
rect 30147 40341 30159 40344
rect 30101 40335 30159 40341
rect 30466 40332 30472 40344
rect 30524 40332 30530 40384
rect 30653 40375 30711 40381
rect 30653 40341 30665 40375
rect 30699 40372 30711 40375
rect 31202 40372 31208 40384
rect 30699 40344 31208 40372
rect 30699 40341 30711 40344
rect 30653 40335 30711 40341
rect 31202 40332 31208 40344
rect 31260 40332 31266 40384
rect 31478 40332 31484 40384
rect 31536 40372 31542 40384
rect 32416 40372 32444 40403
rect 32766 40400 32772 40412
rect 32824 40400 32830 40452
rect 33042 40400 33048 40452
rect 33100 40400 33106 40452
rect 34422 40440 34428 40452
rect 34270 40412 34428 40440
rect 34422 40400 34428 40412
rect 34480 40400 34486 40452
rect 38654 40400 38660 40452
rect 38712 40400 38718 40452
rect 31536 40344 32444 40372
rect 31536 40332 31542 40344
rect 32582 40332 32588 40384
rect 32640 40332 32646 40384
rect 34514 40332 34520 40384
rect 34572 40332 34578 40384
rect 39298 40332 39304 40384
rect 39356 40372 39362 40384
rect 40497 40375 40555 40381
rect 40497 40372 40509 40375
rect 39356 40344 40509 40372
rect 39356 40332 39362 40344
rect 40497 40341 40509 40344
rect 40543 40341 40555 40375
rect 40497 40335 40555 40341
rect 1104 40282 41400 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 41400 40282
rect 1104 40208 41400 40230
rect 10060 40140 11008 40168
rect 10060 40109 10088 40140
rect 10980 40112 11008 40140
rect 12618 40128 12624 40180
rect 12676 40168 12682 40180
rect 12897 40171 12955 40177
rect 12897 40168 12909 40171
rect 12676 40140 12909 40168
rect 12676 40128 12682 40140
rect 12897 40137 12909 40140
rect 12943 40137 12955 40171
rect 12897 40131 12955 40137
rect 13265 40171 13323 40177
rect 13265 40137 13277 40171
rect 13311 40168 13323 40171
rect 13722 40168 13728 40180
rect 13311 40140 13728 40168
rect 13311 40137 13323 40140
rect 13265 40131 13323 40137
rect 13722 40128 13728 40140
rect 13780 40128 13786 40180
rect 14458 40128 14464 40180
rect 14516 40128 14522 40180
rect 15102 40168 15108 40180
rect 14568 40140 15108 40168
rect 10045 40103 10103 40109
rect 10045 40069 10057 40103
rect 10091 40069 10103 40103
rect 10045 40063 10103 40069
rect 10261 40103 10319 40109
rect 10261 40069 10273 40103
rect 10307 40100 10319 40103
rect 10870 40100 10876 40112
rect 10307 40072 10876 40100
rect 10307 40069 10319 40072
rect 10261 40063 10319 40069
rect 10870 40060 10876 40072
rect 10928 40060 10934 40112
rect 10962 40060 10968 40112
rect 11020 40060 11026 40112
rect 11054 40060 11060 40112
rect 11112 40100 11118 40112
rect 12434 40100 12440 40112
rect 11112 40072 12440 40100
rect 11112 40060 11118 40072
rect 12434 40060 12440 40072
rect 12492 40100 12498 40112
rect 14476 40100 14504 40128
rect 12492 40072 14504 40100
rect 12492 40060 12498 40072
rect 8478 39992 8484 40044
rect 8536 39992 8542 40044
rect 9582 39992 9588 40044
rect 9640 39992 9646 40044
rect 13372 40041 13400 40072
rect 14292 40041 14320 40072
rect 9677 40035 9735 40041
rect 9677 40001 9689 40035
rect 9723 40032 9735 40035
rect 13081 40035 13139 40041
rect 9723 40004 11008 40032
rect 9723 40001 9735 40004
rect 9677 39995 9735 40001
rect 10980 39976 11008 40004
rect 13081 40001 13093 40035
rect 13127 40001 13139 40035
rect 13081 39995 13139 40001
rect 13357 40035 13415 40041
rect 13357 40001 13369 40035
rect 13403 40001 13415 40035
rect 13357 39995 13415 40001
rect 14277 40035 14335 40041
rect 14277 40001 14289 40035
rect 14323 40001 14335 40035
rect 14277 39995 14335 40001
rect 9769 39967 9827 39973
rect 9769 39933 9781 39967
rect 9815 39933 9827 39967
rect 9769 39927 9827 39933
rect 8294 39788 8300 39840
rect 8352 39788 8358 39840
rect 9214 39788 9220 39840
rect 9272 39788 9278 39840
rect 9306 39788 9312 39840
rect 9364 39828 9370 39840
rect 9784 39828 9812 39927
rect 10962 39924 10968 39976
rect 11020 39924 11026 39976
rect 9858 39856 9864 39908
rect 9916 39896 9922 39908
rect 10413 39899 10471 39905
rect 10413 39896 10425 39899
rect 9916 39868 10425 39896
rect 9916 39856 9922 39868
rect 10413 39865 10425 39868
rect 10459 39865 10471 39899
rect 13096 39896 13124 39995
rect 14366 39992 14372 40044
rect 14424 39992 14430 40044
rect 14568 40041 14596 40140
rect 15102 40128 15108 40140
rect 15160 40128 15166 40180
rect 15657 40171 15715 40177
rect 15657 40137 15669 40171
rect 15703 40168 15715 40171
rect 15930 40168 15936 40180
rect 15703 40140 15936 40168
rect 15703 40137 15715 40140
rect 15657 40131 15715 40137
rect 15930 40128 15936 40140
rect 15988 40128 15994 40180
rect 16025 40171 16083 40177
rect 16025 40137 16037 40171
rect 16071 40168 16083 40171
rect 16114 40168 16120 40180
rect 16071 40140 16120 40168
rect 16071 40137 16083 40140
rect 16025 40131 16083 40137
rect 16114 40128 16120 40140
rect 16172 40168 16178 40180
rect 16172 40140 17080 40168
rect 16172 40128 16178 40140
rect 16574 40100 16580 40112
rect 14660 40072 16580 40100
rect 14660 40041 14688 40072
rect 16574 40060 16580 40072
rect 16632 40060 16638 40112
rect 16942 40060 16948 40112
rect 17000 40060 17006 40112
rect 17052 40100 17080 40140
rect 17126 40128 17132 40180
rect 17184 40168 17190 40180
rect 17221 40171 17279 40177
rect 17221 40168 17233 40171
rect 17184 40140 17233 40168
rect 17184 40128 17190 40140
rect 17221 40137 17233 40140
rect 17267 40137 17279 40171
rect 17221 40131 17279 40137
rect 17310 40128 17316 40180
rect 17368 40168 17374 40180
rect 17589 40171 17647 40177
rect 17589 40168 17601 40171
rect 17368 40140 17601 40168
rect 17368 40128 17374 40140
rect 17589 40137 17601 40140
rect 17635 40168 17647 40171
rect 17954 40168 17960 40180
rect 17635 40140 17960 40168
rect 17635 40137 17647 40140
rect 17589 40131 17647 40137
rect 17954 40128 17960 40140
rect 18012 40168 18018 40180
rect 18012 40140 18644 40168
rect 18012 40128 18018 40140
rect 18138 40100 18144 40112
rect 17052 40072 17356 40100
rect 14553 40035 14611 40041
rect 14553 40001 14565 40035
rect 14599 40001 14611 40035
rect 14553 39995 14611 40001
rect 14645 40035 14703 40041
rect 14645 40001 14657 40035
rect 14691 40001 14703 40035
rect 14645 39995 14703 40001
rect 15013 40035 15071 40041
rect 15013 40001 15025 40035
rect 15059 40001 15071 40035
rect 15013 39995 15071 40001
rect 15028 39964 15056 39995
rect 15102 39992 15108 40044
rect 15160 39992 15166 40044
rect 15930 40032 15936 40044
rect 15212 40004 15936 40032
rect 15212 39964 15240 40004
rect 15930 39992 15936 40004
rect 15988 39992 15994 40044
rect 16960 40032 16988 40060
rect 16316 40004 16988 40032
rect 15028 39936 15240 39964
rect 15381 39967 15439 39973
rect 15381 39933 15393 39967
rect 15427 39964 15439 39967
rect 15562 39964 15568 39976
rect 15427 39936 15568 39964
rect 15427 39933 15439 39936
rect 15381 39927 15439 39933
rect 15562 39924 15568 39936
rect 15620 39924 15626 39976
rect 15749 39967 15807 39973
rect 15749 39933 15761 39967
rect 15795 39933 15807 39967
rect 15749 39927 15807 39933
rect 15194 39896 15200 39908
rect 13096 39868 15200 39896
rect 10413 39859 10471 39865
rect 15194 39856 15200 39868
rect 15252 39856 15258 39908
rect 15764 39896 15792 39927
rect 15838 39924 15844 39976
rect 15896 39964 15902 39976
rect 16316 39964 16344 40004
rect 15896 39936 16344 39964
rect 17328 39964 17356 40072
rect 17420 40072 18144 40100
rect 17420 40041 17448 40072
rect 18138 40060 18144 40072
rect 18196 40060 18202 40112
rect 18616 40044 18644 40140
rect 19242 40128 19248 40180
rect 19300 40168 19306 40180
rect 20070 40168 20076 40180
rect 19300 40140 20076 40168
rect 19300 40128 19306 40140
rect 20070 40128 20076 40140
rect 20128 40128 20134 40180
rect 20254 40128 20260 40180
rect 20312 40168 20318 40180
rect 20438 40168 20444 40180
rect 20312 40140 20444 40168
rect 20312 40128 20318 40140
rect 20438 40128 20444 40140
rect 20496 40128 20502 40180
rect 22646 40128 22652 40180
rect 22704 40168 22710 40180
rect 24305 40171 24363 40177
rect 22704 40140 23980 40168
rect 22704 40128 22710 40140
rect 19996 40072 20208 40100
rect 17405 40035 17463 40041
rect 17405 40001 17417 40035
rect 17451 40001 17463 40035
rect 17405 39995 17463 40001
rect 17586 39992 17592 40044
rect 17644 40032 17650 40044
rect 17681 40035 17739 40041
rect 17681 40032 17693 40035
rect 17644 40004 17693 40032
rect 17644 39992 17650 40004
rect 17681 40001 17693 40004
rect 17727 40001 17739 40035
rect 17681 39995 17739 40001
rect 18598 39992 18604 40044
rect 18656 39992 18662 40044
rect 19996 40041 20024 40072
rect 19981 40035 20039 40041
rect 19981 40001 19993 40035
rect 20027 40001 20039 40035
rect 20180 40032 20208 40072
rect 20346 40060 20352 40112
rect 20404 40060 20410 40112
rect 20364 40032 20392 40060
rect 20180 40004 20392 40032
rect 19981 39995 20039 40001
rect 20456 39964 20484 40128
rect 20898 40060 20904 40112
rect 20956 40100 20962 40112
rect 23952 40109 23980 40140
rect 24305 40137 24317 40171
rect 24351 40137 24363 40171
rect 24305 40131 24363 40137
rect 23937 40103 23995 40109
rect 20956 40072 23796 40100
rect 20956 40060 20962 40072
rect 20806 39992 20812 40044
rect 20864 40032 20870 40044
rect 21821 40035 21879 40041
rect 21821 40032 21833 40035
rect 20864 40004 21833 40032
rect 20864 39992 20870 40004
rect 21821 40001 21833 40004
rect 21867 40001 21879 40035
rect 21821 39995 21879 40001
rect 23658 39992 23664 40044
rect 23716 39992 23722 40044
rect 23768 40041 23796 40072
rect 23937 40069 23949 40103
rect 23983 40069 23995 40103
rect 23937 40063 23995 40069
rect 24026 40060 24032 40112
rect 24084 40060 24090 40112
rect 24320 40100 24348 40131
rect 27338 40128 27344 40180
rect 27396 40128 27402 40180
rect 31481 40171 31539 40177
rect 28460 40140 29408 40168
rect 28460 40112 28488 40140
rect 24320 40072 27016 40100
rect 23754 40035 23812 40041
rect 23754 40001 23766 40035
rect 23800 40001 23812 40035
rect 23754 39995 23812 40001
rect 24118 39992 24124 40044
rect 24176 40041 24182 40044
rect 24176 40032 24184 40041
rect 24176 40004 24221 40032
rect 24176 39995 24184 40004
rect 24176 39992 24182 39995
rect 24578 39992 24584 40044
rect 24636 40032 24642 40044
rect 25777 40035 25835 40041
rect 25777 40032 25789 40035
rect 24636 40004 25789 40032
rect 24636 39992 24642 40004
rect 25777 40001 25789 40004
rect 25823 40001 25835 40035
rect 25777 39995 25835 40001
rect 25961 40035 26019 40041
rect 25961 40001 25973 40035
rect 26007 40001 26019 40035
rect 25961 39995 26019 40001
rect 17328 39936 20484 39964
rect 15896 39924 15902 39936
rect 25498 39924 25504 39976
rect 25556 39964 25562 39976
rect 25976 39964 26004 39995
rect 26050 39992 26056 40044
rect 26108 39992 26114 40044
rect 26145 40035 26203 40041
rect 26145 40001 26157 40035
rect 26191 40032 26203 40035
rect 26326 40032 26332 40044
rect 26191 40004 26332 40032
rect 26191 40001 26203 40004
rect 26145 39995 26203 40001
rect 26326 39992 26332 40004
rect 26384 39992 26390 40044
rect 26878 39992 26884 40044
rect 26936 39992 26942 40044
rect 26988 40041 27016 40072
rect 28442 40060 28448 40112
rect 28500 40060 28506 40112
rect 29086 40060 29092 40112
rect 29144 40060 29150 40112
rect 26973 40035 27031 40041
rect 26973 40001 26985 40035
rect 27019 40001 27031 40035
rect 26973 39995 27031 40001
rect 29178 39992 29184 40044
rect 29236 40032 29242 40044
rect 29380 40041 29408 40140
rect 31481 40137 31493 40171
rect 31527 40168 31539 40171
rect 32214 40168 32220 40180
rect 31527 40140 32220 40168
rect 31527 40137 31539 40140
rect 31481 40131 31539 40137
rect 32214 40128 32220 40140
rect 32272 40128 32278 40180
rect 32582 40128 32588 40180
rect 32640 40128 32646 40180
rect 32861 40171 32919 40177
rect 32861 40137 32873 40171
rect 32907 40168 32919 40171
rect 33042 40168 33048 40180
rect 32907 40140 33048 40168
rect 32907 40137 32919 40140
rect 32861 40131 32919 40137
rect 33042 40128 33048 40140
rect 33100 40128 33106 40180
rect 30742 40060 30748 40112
rect 30800 40100 30806 40112
rect 31021 40103 31079 40109
rect 31021 40100 31033 40103
rect 30800 40072 31033 40100
rect 30800 40060 30806 40072
rect 31021 40069 31033 40072
rect 31067 40069 31079 40103
rect 32600 40100 32628 40128
rect 32600 40072 33088 40100
rect 31021 40063 31079 40069
rect 29273 40035 29331 40041
rect 29273 40032 29285 40035
rect 29236 40004 29285 40032
rect 29236 39992 29242 40004
rect 29273 40001 29285 40004
rect 29319 40001 29331 40035
rect 29273 39995 29331 40001
rect 29365 40035 29423 40041
rect 29365 40001 29377 40035
rect 29411 40001 29423 40035
rect 29365 39995 29423 40001
rect 30190 39992 30196 40044
rect 30248 40032 30254 40044
rect 33060 40041 33088 40072
rect 31297 40035 31355 40041
rect 31297 40032 31309 40035
rect 30248 40004 31309 40032
rect 30248 39992 30254 40004
rect 31297 40001 31309 40004
rect 31343 40032 31355 40035
rect 33045 40035 33103 40041
rect 31343 40004 32076 40032
rect 31343 40001 31355 40004
rect 31297 39995 31355 40001
rect 26896 39964 26924 39992
rect 25556 39936 26924 39964
rect 25556 39924 25562 39936
rect 27062 39924 27068 39976
rect 27120 39924 27126 39976
rect 27890 39924 27896 39976
rect 27948 39964 27954 39976
rect 28626 39964 28632 39976
rect 27948 39936 28632 39964
rect 27948 39924 27954 39936
rect 28626 39924 28632 39936
rect 28684 39924 28690 39976
rect 31202 39924 31208 39976
rect 31260 39964 31266 39976
rect 31662 39964 31668 39976
rect 31260 39936 31668 39964
rect 31260 39924 31266 39936
rect 31662 39924 31668 39936
rect 31720 39924 31726 39976
rect 16022 39896 16028 39908
rect 15764 39868 16028 39896
rect 16022 39856 16028 39868
rect 16080 39896 16086 39908
rect 16206 39896 16212 39908
rect 16080 39868 16212 39896
rect 16080 39856 16086 39868
rect 16206 39856 16212 39868
rect 16264 39856 16270 39908
rect 17494 39856 17500 39908
rect 17552 39896 17558 39908
rect 19794 39896 19800 39908
rect 17552 39868 19800 39896
rect 17552 39856 17558 39868
rect 19794 39856 19800 39868
rect 19852 39856 19858 39908
rect 20073 39899 20131 39905
rect 20073 39865 20085 39899
rect 20119 39896 20131 39899
rect 20162 39896 20168 39908
rect 20119 39868 20168 39896
rect 20119 39865 20131 39868
rect 20073 39859 20131 39865
rect 20162 39856 20168 39868
rect 20220 39856 20226 39908
rect 22094 39856 22100 39908
rect 22152 39856 22158 39908
rect 22281 39899 22339 39905
rect 22281 39865 22293 39899
rect 22327 39896 22339 39899
rect 23382 39896 23388 39908
rect 22327 39868 23388 39896
rect 22327 39865 22339 39868
rect 22281 39859 22339 39865
rect 23382 39856 23388 39868
rect 23440 39896 23446 39908
rect 23440 39868 27936 39896
rect 23440 39856 23446 39868
rect 27908 39840 27936 39868
rect 32048 39840 32076 40004
rect 33045 40001 33057 40035
rect 33091 40001 33103 40035
rect 33045 39995 33103 40001
rect 10229 39831 10287 39837
rect 10229 39828 10241 39831
rect 9364 39800 10241 39828
rect 9364 39788 9370 39800
rect 10229 39797 10241 39800
rect 10275 39828 10287 39831
rect 12986 39828 12992 39840
rect 10275 39800 12992 39828
rect 10275 39797 10287 39800
rect 10229 39791 10287 39797
rect 12986 39788 12992 39800
rect 13044 39788 13050 39840
rect 13630 39788 13636 39840
rect 13688 39828 13694 39840
rect 14093 39831 14151 39837
rect 14093 39828 14105 39831
rect 13688 39800 14105 39828
rect 13688 39788 13694 39800
rect 14093 39797 14105 39800
rect 14139 39797 14151 39831
rect 14093 39791 14151 39797
rect 15013 39831 15071 39837
rect 15013 39797 15025 39831
rect 15059 39828 15071 39831
rect 15378 39828 15384 39840
rect 15059 39800 15384 39828
rect 15059 39797 15071 39800
rect 15013 39791 15071 39797
rect 15378 39788 15384 39800
rect 15436 39788 15442 39840
rect 17586 39788 17592 39840
rect 17644 39828 17650 39840
rect 19886 39828 19892 39840
rect 17644 39800 19892 39828
rect 17644 39788 17650 39800
rect 19886 39788 19892 39800
rect 19944 39788 19950 39840
rect 20530 39788 20536 39840
rect 20588 39828 20594 39840
rect 20806 39828 20812 39840
rect 20588 39800 20812 39828
rect 20588 39788 20594 39800
rect 20806 39788 20812 39800
rect 20864 39788 20870 39840
rect 22738 39788 22744 39840
rect 22796 39828 22802 39840
rect 25774 39828 25780 39840
rect 22796 39800 25780 39828
rect 22796 39788 22802 39800
rect 25774 39788 25780 39800
rect 25832 39828 25838 39840
rect 25958 39828 25964 39840
rect 25832 39800 25964 39828
rect 25832 39788 25838 39800
rect 25958 39788 25964 39800
rect 26016 39788 26022 39840
rect 26329 39831 26387 39837
rect 26329 39797 26341 39831
rect 26375 39828 26387 39831
rect 26510 39828 26516 39840
rect 26375 39800 26516 39828
rect 26375 39797 26387 39800
rect 26329 39791 26387 39797
rect 26510 39788 26516 39800
rect 26568 39788 26574 39840
rect 26786 39788 26792 39840
rect 26844 39828 26850 39840
rect 26973 39831 27031 39837
rect 26973 39828 26985 39831
rect 26844 39800 26985 39828
rect 26844 39788 26850 39800
rect 26973 39797 26985 39800
rect 27019 39797 27031 39831
rect 26973 39791 27031 39797
rect 27890 39788 27896 39840
rect 27948 39788 27954 39840
rect 29270 39788 29276 39840
rect 29328 39788 29334 39840
rect 29549 39831 29607 39837
rect 29549 39797 29561 39831
rect 29595 39828 29607 39831
rect 29638 39828 29644 39840
rect 29595 39800 29644 39828
rect 29595 39797 29607 39800
rect 29549 39791 29607 39797
rect 29638 39788 29644 39800
rect 29696 39788 29702 39840
rect 30374 39788 30380 39840
rect 30432 39828 30438 39840
rect 31021 39831 31079 39837
rect 31021 39828 31033 39831
rect 30432 39800 31033 39828
rect 30432 39788 30438 39800
rect 31021 39797 31033 39800
rect 31067 39797 31079 39831
rect 31021 39791 31079 39797
rect 32030 39788 32036 39840
rect 32088 39788 32094 39840
rect 1104 39738 41400 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 41400 39738
rect 1104 39664 41400 39686
rect 8478 39584 8484 39636
rect 8536 39624 8542 39636
rect 9401 39627 9459 39633
rect 9401 39624 9413 39627
rect 8536 39596 9413 39624
rect 8536 39584 8542 39596
rect 9401 39593 9413 39596
rect 9447 39593 9459 39627
rect 9401 39587 9459 39593
rect 9766 39584 9772 39636
rect 9824 39584 9830 39636
rect 14366 39584 14372 39636
rect 14424 39624 14430 39636
rect 15105 39627 15163 39633
rect 15105 39624 15117 39627
rect 14424 39596 15117 39624
rect 14424 39584 14430 39596
rect 15105 39593 15117 39596
rect 15151 39593 15163 39627
rect 15105 39587 15163 39593
rect 15286 39584 15292 39636
rect 15344 39624 15350 39636
rect 15654 39624 15660 39636
rect 15344 39596 15660 39624
rect 15344 39584 15350 39596
rect 15654 39584 15660 39596
rect 15712 39624 15718 39636
rect 16482 39624 16488 39636
rect 15712 39596 16488 39624
rect 15712 39584 15718 39596
rect 16482 39584 16488 39596
rect 16540 39584 16546 39636
rect 16574 39584 16580 39636
rect 16632 39624 16638 39636
rect 17589 39627 17647 39633
rect 17589 39624 17601 39627
rect 16632 39596 17601 39624
rect 16632 39584 16638 39596
rect 17589 39593 17601 39596
rect 17635 39593 17647 39627
rect 17589 39587 17647 39593
rect 18506 39584 18512 39636
rect 18564 39624 18570 39636
rect 18601 39627 18659 39633
rect 18601 39624 18613 39627
rect 18564 39596 18613 39624
rect 18564 39584 18570 39596
rect 18601 39593 18613 39596
rect 18647 39593 18659 39627
rect 18601 39587 18659 39593
rect 18690 39584 18696 39636
rect 18748 39624 18754 39636
rect 25222 39624 25228 39636
rect 18748 39596 25228 39624
rect 18748 39584 18754 39596
rect 25222 39584 25228 39596
rect 25280 39584 25286 39636
rect 25314 39584 25320 39636
rect 25372 39584 25378 39636
rect 25590 39624 25596 39636
rect 25424 39596 25596 39624
rect 9214 39516 9220 39568
rect 9272 39516 9278 39568
rect 8941 39491 8999 39497
rect 8941 39457 8953 39491
rect 8987 39488 8999 39491
rect 9784 39488 9812 39584
rect 10962 39516 10968 39568
rect 11020 39556 11026 39568
rect 15930 39556 15936 39568
rect 11020 39528 15936 39556
rect 11020 39516 11026 39528
rect 15930 39516 15936 39528
rect 15988 39556 15994 39568
rect 16117 39559 16175 39565
rect 16117 39556 16129 39559
rect 15988 39528 16129 39556
rect 15988 39516 15994 39528
rect 16117 39525 16129 39528
rect 16163 39525 16175 39559
rect 16117 39519 16175 39525
rect 17678 39516 17684 39568
rect 17736 39556 17742 39568
rect 18969 39559 19027 39565
rect 18969 39556 18981 39559
rect 17736 39528 18981 39556
rect 17736 39516 17742 39528
rect 18969 39525 18981 39528
rect 19015 39556 19027 39559
rect 19015 39528 20116 39556
rect 19015 39525 19027 39528
rect 18969 39519 19027 39525
rect 8987 39460 9812 39488
rect 11425 39491 11483 39497
rect 8987 39457 8999 39460
rect 8941 39451 8999 39457
rect 11425 39457 11437 39491
rect 11471 39488 11483 39491
rect 11517 39491 11575 39497
rect 11517 39488 11529 39491
rect 11471 39460 11529 39488
rect 11471 39457 11483 39460
rect 11425 39451 11483 39457
rect 11517 39457 11529 39460
rect 11563 39488 11575 39491
rect 11606 39488 11612 39500
rect 11563 39460 11612 39488
rect 11563 39457 11575 39460
rect 11517 39451 11575 39457
rect 11606 39448 11612 39460
rect 11664 39448 11670 39500
rect 14550 39448 14556 39500
rect 14608 39448 14614 39500
rect 15473 39491 15531 39497
rect 15473 39457 15485 39491
rect 15519 39488 15531 39491
rect 15838 39488 15844 39500
rect 15519 39460 15844 39488
rect 15519 39457 15531 39460
rect 15473 39451 15531 39457
rect 15838 39448 15844 39460
rect 15896 39488 15902 39500
rect 16298 39488 16304 39500
rect 15896 39460 16304 39488
rect 15896 39448 15902 39460
rect 16298 39448 16304 39460
rect 16356 39448 16362 39500
rect 16574 39448 16580 39500
rect 16632 39488 16638 39500
rect 17586 39488 17592 39500
rect 16632 39460 17592 39488
rect 16632 39448 16638 39460
rect 17586 39448 17592 39460
rect 17644 39488 17650 39500
rect 19337 39491 19395 39497
rect 19337 39488 19349 39491
rect 17644 39460 17816 39488
rect 17644 39448 17650 39460
rect 9674 39380 9680 39432
rect 9732 39380 9738 39432
rect 15958 39423 16016 39429
rect 15958 39389 15970 39423
rect 16004 39420 16016 39423
rect 16206 39420 16212 39432
rect 16004 39392 16212 39420
rect 16004 39389 16016 39392
rect 15958 39383 16016 39389
rect 16206 39380 16212 39392
rect 16264 39420 16270 39432
rect 16390 39420 16396 39432
rect 16264 39392 16396 39420
rect 16264 39380 16270 39392
rect 16390 39380 16396 39392
rect 16448 39380 16454 39432
rect 17788 39429 17816 39460
rect 19076 39460 19349 39488
rect 17773 39423 17831 39429
rect 17773 39389 17785 39423
rect 17819 39389 17831 39423
rect 17773 39383 17831 39389
rect 17954 39380 17960 39432
rect 18012 39380 18018 39432
rect 18230 39380 18236 39432
rect 18288 39380 18294 39432
rect 18598 39380 18604 39432
rect 18656 39380 18662 39432
rect 18782 39380 18788 39432
rect 18840 39380 18846 39432
rect 18966 39380 18972 39432
rect 19024 39422 19030 39432
rect 19076 39422 19104 39460
rect 19337 39457 19349 39460
rect 19383 39488 19395 39491
rect 19383 39460 19840 39488
rect 19383 39457 19395 39460
rect 19337 39451 19395 39457
rect 19024 39394 19104 39422
rect 19024 39380 19030 39394
rect 19150 39380 19156 39432
rect 19208 39420 19214 39432
rect 19812 39429 19840 39460
rect 19245 39423 19303 39429
rect 19245 39420 19257 39423
rect 19208 39392 19257 39420
rect 19208 39380 19214 39392
rect 19245 39389 19257 39392
rect 19291 39389 19303 39423
rect 19245 39383 19303 39389
rect 19521 39423 19579 39429
rect 19521 39389 19533 39423
rect 19567 39389 19579 39423
rect 19521 39383 19579 39389
rect 19797 39423 19855 39429
rect 19797 39389 19809 39423
rect 19843 39389 19855 39423
rect 19797 39383 19855 39389
rect 9950 39312 9956 39364
rect 10008 39312 10014 39364
rect 10594 39312 10600 39364
rect 10652 39312 10658 39364
rect 17865 39355 17923 39361
rect 17865 39321 17877 39355
rect 17911 39321 17923 39355
rect 17865 39315 17923 39321
rect 18075 39355 18133 39361
rect 18075 39321 18087 39355
rect 18121 39352 18133 39355
rect 18322 39352 18328 39364
rect 18121 39324 18328 39352
rect 18121 39321 18133 39324
rect 18075 39315 18133 39321
rect 12158 39244 12164 39296
rect 12216 39244 12222 39296
rect 15286 39244 15292 39296
rect 15344 39284 15350 39296
rect 15562 39284 15568 39296
rect 15344 39256 15568 39284
rect 15344 39244 15350 39256
rect 15562 39244 15568 39256
rect 15620 39284 15626 39296
rect 15749 39287 15807 39293
rect 15749 39284 15761 39287
rect 15620 39256 15761 39284
rect 15620 39244 15626 39256
rect 15749 39253 15761 39256
rect 15795 39253 15807 39287
rect 15749 39247 15807 39253
rect 15841 39287 15899 39293
rect 15841 39253 15853 39287
rect 15887 39284 15899 39287
rect 16482 39284 16488 39296
rect 15887 39256 16488 39284
rect 15887 39253 15899 39256
rect 15841 39247 15899 39253
rect 16482 39244 16488 39256
rect 16540 39244 16546 39296
rect 17880 39284 17908 39315
rect 18322 39312 18328 39324
rect 18380 39312 18386 39364
rect 19426 39352 19432 39364
rect 19168 39324 19432 39352
rect 17954 39284 17960 39296
rect 17880 39256 17960 39284
rect 17954 39244 17960 39256
rect 18012 39244 18018 39296
rect 18340 39284 18368 39312
rect 18690 39284 18696 39296
rect 18340 39256 18696 39284
rect 18690 39244 18696 39256
rect 18748 39244 18754 39296
rect 18782 39244 18788 39296
rect 18840 39284 18846 39296
rect 19168 39284 19196 39324
rect 19426 39312 19432 39324
rect 19484 39312 19490 39364
rect 18840 39256 19196 39284
rect 18840 39244 18846 39256
rect 19334 39244 19340 39296
rect 19392 39284 19398 39296
rect 19536 39284 19564 39383
rect 19886 39380 19892 39432
rect 19944 39380 19950 39432
rect 19705 39355 19763 39361
rect 19705 39321 19717 39355
rect 19751 39352 19763 39355
rect 20088 39352 20116 39528
rect 20806 39516 20812 39568
rect 20864 39556 20870 39568
rect 23198 39556 23204 39568
rect 20864 39528 23204 39556
rect 20864 39516 20870 39528
rect 23198 39516 23204 39528
rect 23256 39516 23262 39568
rect 23750 39516 23756 39568
rect 23808 39556 23814 39568
rect 24762 39556 24768 39568
rect 23808 39528 24768 39556
rect 23808 39516 23814 39528
rect 24762 39516 24768 39528
rect 24820 39516 24826 39568
rect 23014 39448 23020 39500
rect 23072 39488 23078 39500
rect 24302 39488 24308 39500
rect 23072 39460 24308 39488
rect 23072 39448 23078 39460
rect 24302 39448 24308 39460
rect 24360 39448 24366 39500
rect 25424 39497 25452 39596
rect 25590 39584 25596 39596
rect 25648 39584 25654 39636
rect 25682 39584 25688 39636
rect 25740 39624 25746 39636
rect 26510 39624 26516 39636
rect 25740 39596 26516 39624
rect 25740 39584 25746 39596
rect 26510 39584 26516 39596
rect 26568 39584 26574 39636
rect 28350 39584 28356 39636
rect 28408 39624 28414 39636
rect 29270 39624 29276 39636
rect 28408 39596 29276 39624
rect 28408 39584 28414 39596
rect 29270 39584 29276 39596
rect 29328 39584 29334 39636
rect 29546 39584 29552 39636
rect 29604 39584 29610 39636
rect 30466 39584 30472 39636
rect 30524 39624 30530 39636
rect 30929 39627 30987 39633
rect 30929 39624 30941 39627
rect 30524 39596 30941 39624
rect 30524 39584 30530 39596
rect 30929 39593 30941 39596
rect 30975 39593 30987 39627
rect 30929 39587 30987 39593
rect 31757 39627 31815 39633
rect 31757 39593 31769 39627
rect 31803 39624 31815 39627
rect 31846 39624 31852 39636
rect 31803 39596 31852 39624
rect 31803 39593 31815 39596
rect 31757 39587 31815 39593
rect 31846 39584 31852 39596
rect 31904 39584 31910 39636
rect 32030 39584 32036 39636
rect 32088 39584 32094 39636
rect 39298 39584 39304 39636
rect 39356 39584 39362 39636
rect 26234 39556 26240 39568
rect 25516 39528 26240 39556
rect 25409 39491 25467 39497
rect 25409 39457 25421 39491
rect 25455 39457 25467 39491
rect 25409 39451 25467 39457
rect 20254 39380 20260 39432
rect 20312 39420 20318 39432
rect 25516 39429 25544 39528
rect 26234 39516 26240 39528
rect 26292 39556 26298 39568
rect 26602 39556 26608 39568
rect 26292 39528 26608 39556
rect 26292 39516 26298 39528
rect 26602 39516 26608 39528
rect 26660 39556 26666 39568
rect 31202 39556 31208 39568
rect 26660 39528 31208 39556
rect 26660 39516 26666 39528
rect 31202 39516 31208 39528
rect 31260 39516 31266 39568
rect 31389 39559 31447 39565
rect 31389 39525 31401 39559
rect 31435 39556 31447 39559
rect 31435 39528 32168 39556
rect 31435 39525 31447 39528
rect 31389 39519 31447 39525
rect 29178 39488 29184 39500
rect 26160 39460 29184 39488
rect 26160 39432 26188 39460
rect 29178 39448 29184 39460
rect 29236 39448 29242 39500
rect 29638 39448 29644 39500
rect 29696 39448 29702 39500
rect 29730 39448 29736 39500
rect 29788 39488 29794 39500
rect 32140 39497 32168 39528
rect 31021 39491 31079 39497
rect 31021 39488 31033 39491
rect 29788 39460 31033 39488
rect 29788 39448 29794 39460
rect 31021 39457 31033 39460
rect 31067 39457 31079 39491
rect 32125 39491 32183 39497
rect 31021 39451 31079 39457
rect 31128 39460 32076 39488
rect 25501 39423 25559 39429
rect 20312 39392 25360 39420
rect 20312 39380 20318 39392
rect 20162 39352 20168 39364
rect 19751 39324 20168 39352
rect 19751 39321 19763 39324
rect 19705 39315 19763 39321
rect 20162 39312 20168 39324
rect 20220 39312 20226 39364
rect 24946 39312 24952 39364
rect 25004 39352 25010 39364
rect 25225 39355 25283 39361
rect 25225 39352 25237 39355
rect 25004 39324 25237 39352
rect 25004 39312 25010 39324
rect 25225 39321 25237 39324
rect 25271 39321 25283 39355
rect 25332 39352 25360 39392
rect 25501 39389 25513 39423
rect 25547 39389 25559 39423
rect 25501 39383 25559 39389
rect 25866 39380 25872 39432
rect 25924 39380 25930 39432
rect 26142 39380 26148 39432
rect 26200 39380 26206 39432
rect 27706 39380 27712 39432
rect 27764 39420 27770 39432
rect 28074 39420 28080 39432
rect 27764 39392 28080 39420
rect 27764 39380 27770 39392
rect 28074 39380 28080 39392
rect 28132 39420 28138 39432
rect 28169 39423 28227 39429
rect 28169 39420 28181 39423
rect 28132 39392 28181 39420
rect 28132 39380 28138 39392
rect 28169 39389 28181 39392
rect 28215 39389 28227 39423
rect 28169 39383 28227 39389
rect 28258 39380 28264 39432
rect 28316 39420 28322 39432
rect 28316 39392 28488 39420
rect 28316 39380 28322 39392
rect 25884 39352 25912 39380
rect 28350 39352 28356 39364
rect 25332 39324 25912 39352
rect 27540 39324 28356 39352
rect 25225 39315 25283 39321
rect 19392 39256 19564 39284
rect 19392 39244 19398 39256
rect 20070 39244 20076 39296
rect 20128 39244 20134 39296
rect 23566 39244 23572 39296
rect 23624 39284 23630 39296
rect 24026 39284 24032 39296
rect 23624 39256 24032 39284
rect 23624 39244 23630 39256
rect 24026 39244 24032 39256
rect 24084 39244 24090 39296
rect 24302 39244 24308 39296
rect 24360 39284 24366 39296
rect 24854 39284 24860 39296
rect 24360 39256 24860 39284
rect 24360 39244 24366 39256
rect 24854 39244 24860 39256
rect 24912 39244 24918 39296
rect 25682 39244 25688 39296
rect 25740 39244 25746 39296
rect 25774 39244 25780 39296
rect 25832 39284 25838 39296
rect 27540 39284 27568 39324
rect 28350 39312 28356 39324
rect 28408 39312 28414 39364
rect 28460 39361 28488 39392
rect 28534 39380 28540 39432
rect 28592 39380 28598 39432
rect 28994 39380 29000 39432
rect 29052 39420 29058 39432
rect 29549 39423 29607 39429
rect 29549 39420 29561 39423
rect 29052 39392 29561 39420
rect 29052 39380 29058 39392
rect 29549 39389 29561 39392
rect 29595 39389 29607 39423
rect 29549 39383 29607 39389
rect 30650 39380 30656 39432
rect 30708 39420 30714 39432
rect 31128 39420 31156 39460
rect 30708 39392 31156 39420
rect 31205 39423 31263 39429
rect 30708 39380 30714 39392
rect 31205 39389 31217 39423
rect 31251 39389 31263 39423
rect 31205 39383 31263 39389
rect 28445 39355 28503 39361
rect 28445 39321 28457 39355
rect 28491 39321 28503 39355
rect 30558 39352 30564 39364
rect 28445 39315 28503 39321
rect 28644 39324 30564 39352
rect 25832 39256 27568 39284
rect 25832 39244 25838 39256
rect 27614 39244 27620 39296
rect 27672 39284 27678 39296
rect 28644 39284 28672 39324
rect 30558 39312 30564 39324
rect 30616 39312 30622 39364
rect 30926 39312 30932 39364
rect 30984 39312 30990 39364
rect 27672 39256 28672 39284
rect 28721 39287 28779 39293
rect 27672 39244 27678 39256
rect 28721 39253 28733 39287
rect 28767 39284 28779 39287
rect 28810 39284 28816 39296
rect 28767 39256 28816 39284
rect 28767 39253 28779 39256
rect 28721 39247 28779 39253
rect 28810 39244 28816 39256
rect 28868 39244 28874 39296
rect 28902 39244 28908 39296
rect 28960 39284 28966 39296
rect 29638 39284 29644 39296
rect 28960 39256 29644 39284
rect 28960 39244 28966 39256
rect 29638 39244 29644 39256
rect 29696 39244 29702 39296
rect 29914 39244 29920 39296
rect 29972 39244 29978 39296
rect 31220 39284 31248 39383
rect 31570 39380 31576 39432
rect 31628 39380 31634 39432
rect 31665 39423 31723 39429
rect 31665 39389 31677 39423
rect 31711 39389 31723 39423
rect 32048 39420 32076 39460
rect 32125 39457 32137 39491
rect 32171 39457 32183 39491
rect 32125 39451 32183 39457
rect 37642 39448 37648 39500
rect 37700 39488 37706 39500
rect 37921 39491 37979 39497
rect 37921 39488 37933 39491
rect 37700 39460 37933 39488
rect 37700 39448 37706 39460
rect 37921 39457 37933 39460
rect 37967 39457 37979 39491
rect 37921 39451 37979 39457
rect 38197 39491 38255 39497
rect 38197 39457 38209 39491
rect 38243 39488 38255 39491
rect 39316 39488 39344 39584
rect 38243 39460 39344 39488
rect 38243 39457 38255 39460
rect 38197 39451 38255 39457
rect 32309 39423 32367 39429
rect 32309 39420 32321 39423
rect 32048 39392 32321 39420
rect 31665 39383 31723 39389
rect 32309 39389 32321 39392
rect 32355 39420 32367 39423
rect 32355 39392 32720 39420
rect 32355 39389 32367 39392
rect 32309 39383 32367 39389
rect 31386 39312 31392 39364
rect 31444 39352 31450 39364
rect 31680 39352 31708 39383
rect 31444 39324 31708 39352
rect 32033 39355 32091 39361
rect 31444 39312 31450 39324
rect 32033 39321 32045 39355
rect 32079 39352 32091 39355
rect 32582 39352 32588 39364
rect 32079 39324 32588 39352
rect 32079 39321 32091 39324
rect 32033 39315 32091 39321
rect 32582 39312 32588 39324
rect 32640 39312 32646 39364
rect 32692 39296 32720 39392
rect 33502 39380 33508 39432
rect 33560 39380 33566 39432
rect 38654 39312 38660 39364
rect 38712 39312 38718 39364
rect 31570 39284 31576 39296
rect 31220 39256 31576 39284
rect 31570 39244 31576 39256
rect 31628 39244 31634 39296
rect 31938 39244 31944 39296
rect 31996 39244 32002 39296
rect 32490 39244 32496 39296
rect 32548 39244 32554 39296
rect 32674 39244 32680 39296
rect 32732 39244 32738 39296
rect 33321 39287 33379 39293
rect 33321 39253 33333 39287
rect 33367 39284 33379 39287
rect 33686 39284 33692 39296
rect 33367 39256 33692 39284
rect 33367 39253 33379 39256
rect 33321 39247 33379 39253
rect 33686 39244 33692 39256
rect 33744 39244 33750 39296
rect 39666 39244 39672 39296
rect 39724 39244 39730 39296
rect 1104 39194 41400 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 41400 39194
rect 1104 39120 41400 39142
rect 8294 39040 8300 39092
rect 8352 39040 8358 39092
rect 9401 39083 9459 39089
rect 9401 39049 9413 39083
rect 9447 39080 9459 39083
rect 9582 39080 9588 39092
rect 9447 39052 9588 39080
rect 9447 39049 9459 39052
rect 9401 39043 9459 39049
rect 9582 39040 9588 39052
rect 9640 39040 9646 39092
rect 9858 39040 9864 39092
rect 9916 39040 9922 39092
rect 9950 39040 9956 39092
rect 10008 39080 10014 39092
rect 10321 39083 10379 39089
rect 10321 39080 10333 39083
rect 10008 39052 10333 39080
rect 10008 39040 10014 39052
rect 10321 39049 10333 39052
rect 10367 39049 10379 39083
rect 10321 39043 10379 39049
rect 12158 39040 12164 39092
rect 12216 39040 12222 39092
rect 13630 39080 13636 39092
rect 13004 39052 13636 39080
rect 7929 39015 7987 39021
rect 7929 38981 7941 39015
rect 7975 39012 7987 39015
rect 8312 39012 8340 39040
rect 7975 38984 8340 39012
rect 7975 38981 7987 38984
rect 7929 38975 7987 38981
rect 9769 38947 9827 38953
rect 6914 38836 6920 38888
rect 6972 38876 6978 38888
rect 7653 38879 7711 38885
rect 7653 38876 7665 38879
rect 6972 38848 7665 38876
rect 6972 38836 6978 38848
rect 7653 38845 7665 38848
rect 7699 38845 7711 38879
rect 7653 38839 7711 38845
rect 9048 38820 9076 38930
rect 9769 38913 9781 38947
rect 9815 38944 9827 38947
rect 9876 38944 9904 39040
rect 10045 39015 10103 39021
rect 10045 38981 10057 39015
rect 10091 39012 10103 39015
rect 12176 39012 12204 39040
rect 13004 39021 13032 39052
rect 13630 39040 13636 39052
rect 13688 39040 13694 39092
rect 14461 39083 14519 39089
rect 14461 39049 14473 39083
rect 14507 39080 14519 39083
rect 14550 39080 14556 39092
rect 14507 39052 14556 39080
rect 14507 39049 14519 39052
rect 14461 39043 14519 39049
rect 14550 39040 14556 39052
rect 14608 39040 14614 39092
rect 16482 39040 16488 39092
rect 16540 39080 16546 39092
rect 18874 39080 18880 39092
rect 16540 39052 18880 39080
rect 16540 39040 16546 39052
rect 18874 39040 18880 39052
rect 18932 39040 18938 39092
rect 19794 39040 19800 39092
rect 19852 39080 19858 39092
rect 20073 39083 20131 39089
rect 20073 39080 20085 39083
rect 19852 39052 20085 39080
rect 19852 39040 19858 39052
rect 20073 39049 20085 39052
rect 20119 39049 20131 39083
rect 20073 39043 20131 39049
rect 20254 39040 20260 39092
rect 20312 39040 20318 39092
rect 20530 39040 20536 39092
rect 20588 39040 20594 39092
rect 20993 39083 21051 39089
rect 20993 39049 21005 39083
rect 21039 39080 21051 39083
rect 22370 39080 22376 39092
rect 21039 39052 22376 39080
rect 21039 39049 21051 39052
rect 20993 39043 21051 39049
rect 22370 39040 22376 39052
rect 22428 39040 22434 39092
rect 25498 39080 25504 39092
rect 24872 39052 25504 39080
rect 10091 38984 12204 39012
rect 12989 39015 13047 39021
rect 10091 38981 10103 38984
rect 10045 38975 10103 38981
rect 12989 38981 13001 39015
rect 13035 38981 13047 39015
rect 12989 38975 13047 38981
rect 13538 38972 13544 39024
rect 13596 38972 13602 39024
rect 17954 39012 17960 39024
rect 17512 38984 17960 39012
rect 9815 38916 9904 38944
rect 9953 38947 10011 38953
rect 9815 38913 9827 38916
rect 9769 38907 9827 38913
rect 9953 38913 9965 38947
rect 9999 38913 10011 38947
rect 9953 38907 10011 38913
rect 10137 38947 10195 38953
rect 10137 38913 10149 38947
rect 10183 38944 10195 38947
rect 10410 38944 10416 38956
rect 10183 38916 10416 38944
rect 10183 38913 10195 38916
rect 10137 38907 10195 38913
rect 9968 38876 9996 38907
rect 10410 38904 10416 38916
rect 10468 38904 10474 38956
rect 10962 38904 10968 38956
rect 11020 38904 11026 38956
rect 11422 38904 11428 38956
rect 11480 38944 11486 38956
rect 12710 38944 12716 38956
rect 11480 38916 12716 38944
rect 11480 38904 11486 38916
rect 12710 38904 12716 38916
rect 12768 38904 12774 38956
rect 17512 38953 17540 38984
rect 17954 38972 17960 38984
rect 18012 38972 18018 39024
rect 18138 38972 18144 39024
rect 18196 38972 18202 39024
rect 17497 38947 17555 38953
rect 17497 38913 17509 38947
rect 17543 38913 17555 38947
rect 17497 38907 17555 38913
rect 17770 38904 17776 38956
rect 17828 38904 17834 38956
rect 18046 38944 18052 38956
rect 17880 38916 18052 38944
rect 10980 38876 11008 38904
rect 9968 38848 11008 38876
rect 15286 38836 15292 38888
rect 15344 38876 15350 38888
rect 17880 38876 17908 38916
rect 18046 38904 18052 38916
rect 18104 38904 18110 38956
rect 18156 38944 18184 38972
rect 18892 38953 18920 39040
rect 20548 39012 20576 39040
rect 21361 39015 21419 39021
rect 21361 39012 21373 39015
rect 19720 38984 20576 39012
rect 20640 38984 21373 39012
rect 18233 38947 18291 38953
rect 18233 38944 18245 38947
rect 18156 38916 18245 38944
rect 18233 38913 18245 38916
rect 18279 38944 18291 38947
rect 18601 38947 18659 38953
rect 18601 38944 18613 38947
rect 18279 38916 18613 38944
rect 18279 38913 18291 38916
rect 18233 38907 18291 38913
rect 18601 38913 18613 38916
rect 18647 38913 18659 38947
rect 18601 38907 18659 38913
rect 18785 38947 18843 38953
rect 18785 38913 18797 38947
rect 18831 38913 18843 38947
rect 18785 38907 18843 38913
rect 18877 38947 18935 38953
rect 18877 38913 18889 38947
rect 18923 38913 18935 38947
rect 18877 38907 18935 38913
rect 15344 38848 17908 38876
rect 17957 38879 18015 38885
rect 15344 38836 15350 38848
rect 17957 38845 17969 38879
rect 18003 38845 18015 38879
rect 18064 38876 18092 38904
rect 18800 38876 18828 38907
rect 19426 38904 19432 38956
rect 19484 38944 19490 38956
rect 19720 38953 19748 38984
rect 19705 38947 19763 38953
rect 19705 38944 19717 38947
rect 19484 38916 19717 38944
rect 19484 38904 19490 38916
rect 19705 38913 19717 38916
rect 19751 38913 19763 38947
rect 19705 38907 19763 38913
rect 19889 38947 19947 38953
rect 19889 38913 19901 38947
rect 19935 38944 19947 38947
rect 19978 38944 19984 38956
rect 19935 38916 19984 38944
rect 19935 38913 19947 38916
rect 19889 38907 19947 38913
rect 19978 38904 19984 38916
rect 20036 38904 20042 38956
rect 20070 38904 20076 38956
rect 20128 38944 20134 38956
rect 20441 38947 20499 38953
rect 20441 38944 20453 38947
rect 20128 38916 20453 38944
rect 20128 38904 20134 38916
rect 20441 38913 20453 38916
rect 20487 38913 20499 38947
rect 20441 38907 20499 38913
rect 20530 38904 20536 38956
rect 20588 38904 20594 38956
rect 20640 38953 20668 38984
rect 21361 38981 21373 38984
rect 21407 38981 21419 39015
rect 21361 38975 21419 38981
rect 20625 38947 20683 38953
rect 20625 38913 20637 38947
rect 20671 38913 20683 38947
rect 20625 38907 20683 38913
rect 18064 38848 18828 38876
rect 17957 38839 18015 38845
rect 9030 38768 9036 38820
rect 9088 38808 9094 38820
rect 10594 38808 10600 38820
rect 9088 38780 10600 38808
rect 9088 38768 9094 38780
rect 10594 38768 10600 38780
rect 10652 38768 10658 38820
rect 17972 38808 18000 38839
rect 20162 38836 20168 38888
rect 20220 38876 20226 38888
rect 20640 38876 20668 38907
rect 20714 38904 20720 38956
rect 20772 38953 20778 38956
rect 20772 38947 20801 38953
rect 20789 38913 20801 38947
rect 20772 38907 20801 38913
rect 21177 38947 21235 38953
rect 21177 38913 21189 38947
rect 21223 38913 21235 38947
rect 21177 38907 21235 38913
rect 21269 38947 21327 38953
rect 21269 38913 21281 38947
rect 21315 38913 21327 38947
rect 21376 38944 21404 38975
rect 21450 38972 21456 39024
rect 21508 39021 21514 39024
rect 21508 39015 21557 39021
rect 21508 38981 21511 39015
rect 21545 39012 21557 39015
rect 23014 39012 23020 39024
rect 21545 38984 23020 39012
rect 21545 38981 21557 38984
rect 21508 38975 21557 38981
rect 21508 38972 21514 38975
rect 23014 38972 23020 38984
rect 23072 38972 23078 39024
rect 23385 39015 23443 39021
rect 23385 39012 23397 39015
rect 23216 38984 23397 39012
rect 23216 38956 23244 38984
rect 23385 38981 23397 38984
rect 23431 38981 23443 39015
rect 24121 39015 24179 39021
rect 24121 39012 24133 39015
rect 23385 38975 23443 38981
rect 23492 38984 24133 39012
rect 23492 38956 23520 38984
rect 24121 38981 24133 38984
rect 24167 38981 24179 39015
rect 24872 39012 24900 39052
rect 25498 39040 25504 39052
rect 25556 39040 25562 39092
rect 25869 39083 25927 39089
rect 25869 39049 25881 39083
rect 25915 39049 25927 39083
rect 25869 39043 25927 39049
rect 26697 39083 26755 39089
rect 26697 39049 26709 39083
rect 26743 39080 26755 39083
rect 27062 39080 27068 39092
rect 26743 39052 27068 39080
rect 26743 39049 26755 39052
rect 26697 39043 26755 39049
rect 24121 38975 24179 38981
rect 24780 38984 24900 39012
rect 21726 38944 21732 38956
rect 21376 38916 21732 38944
rect 21269 38907 21327 38913
rect 20772 38904 20778 38907
rect 20220 38848 20668 38876
rect 20901 38879 20959 38885
rect 20220 38836 20226 38848
rect 20901 38845 20913 38879
rect 20947 38876 20959 38879
rect 21082 38876 21088 38888
rect 20947 38848 21088 38876
rect 20947 38845 20959 38848
rect 20901 38839 20959 38845
rect 21082 38836 21088 38848
rect 21140 38836 21146 38888
rect 20622 38808 20628 38820
rect 17972 38780 20628 38808
rect 20622 38768 20628 38780
rect 20680 38768 20686 38820
rect 21192 38752 21220 38907
rect 21284 38876 21312 38907
rect 21726 38904 21732 38916
rect 21784 38904 21790 38956
rect 22186 38904 22192 38956
rect 22244 38944 22250 38956
rect 22741 38947 22799 38953
rect 22741 38944 22753 38947
rect 22244 38916 22753 38944
rect 22244 38904 22250 38916
rect 22741 38913 22753 38916
rect 22787 38913 22799 38947
rect 22741 38907 22799 38913
rect 22925 38947 22983 38953
rect 22925 38913 22937 38947
rect 22971 38944 22983 38947
rect 22971 38916 23152 38944
rect 22971 38913 22983 38916
rect 22925 38907 22983 38913
rect 21542 38876 21548 38888
rect 21284 38848 21548 38876
rect 21542 38836 21548 38848
rect 21600 38836 21606 38888
rect 21634 38836 21640 38888
rect 21692 38836 21698 38888
rect 22278 38836 22284 38888
rect 22336 38876 22342 38888
rect 22649 38879 22707 38885
rect 22649 38876 22661 38879
rect 22336 38848 22661 38876
rect 22336 38836 22342 38848
rect 22649 38845 22661 38848
rect 22695 38876 22707 38879
rect 23014 38876 23020 38888
rect 22695 38848 23020 38876
rect 22695 38845 22707 38848
rect 22649 38839 22707 38845
rect 23014 38836 23020 38848
rect 23072 38836 23078 38888
rect 23124 38876 23152 38916
rect 23198 38904 23204 38956
rect 23256 38904 23262 38956
rect 23290 38904 23296 38956
rect 23348 38904 23354 38956
rect 23474 38904 23480 38956
rect 23532 38904 23538 38956
rect 23615 38947 23673 38953
rect 23615 38913 23627 38947
rect 23661 38944 23673 38947
rect 23842 38944 23848 38956
rect 23661 38916 23848 38944
rect 23661 38913 23673 38916
rect 23615 38907 23673 38913
rect 23842 38904 23848 38916
rect 23900 38904 23906 38956
rect 23934 38904 23940 38956
rect 23992 38904 23998 38956
rect 24213 38947 24271 38953
rect 24213 38913 24225 38947
rect 24259 38913 24271 38947
rect 24213 38907 24271 38913
rect 23382 38876 23388 38888
rect 23124 38848 23388 38876
rect 23382 38836 23388 38848
rect 23440 38836 23446 38888
rect 23753 38879 23811 38885
rect 23753 38845 23765 38879
rect 23799 38876 23811 38879
rect 24026 38876 24032 38888
rect 23799 38848 24032 38876
rect 23799 38845 23811 38848
rect 23753 38839 23811 38845
rect 24026 38836 24032 38848
rect 24084 38836 24090 38888
rect 22002 38768 22008 38820
rect 22060 38808 22066 38820
rect 24228 38808 24256 38907
rect 24302 38904 24308 38956
rect 24360 38904 24366 38956
rect 24780 38953 24808 38984
rect 25038 38972 25044 39024
rect 25096 39012 25102 39024
rect 25884 39012 25912 39043
rect 27062 39040 27068 39052
rect 27120 39080 27126 39092
rect 27120 39052 27476 39080
rect 27120 39040 27126 39052
rect 27448 39021 27476 39052
rect 27614 39040 27620 39092
rect 27672 39040 27678 39092
rect 28534 39080 28540 39092
rect 28092 39052 28540 39080
rect 27249 39015 27307 39021
rect 27249 39012 27261 39015
rect 25096 38984 25636 39012
rect 25884 38984 27261 39012
rect 25096 38972 25102 38984
rect 24581 38947 24639 38953
rect 24581 38913 24593 38947
rect 24627 38913 24639 38947
rect 24581 38907 24639 38913
rect 24765 38947 24823 38953
rect 24765 38913 24777 38947
rect 24811 38913 24823 38947
rect 24765 38907 24823 38913
rect 24857 38947 24915 38953
rect 24857 38913 24869 38947
rect 24903 38913 24915 38947
rect 24857 38907 24915 38913
rect 24596 38876 24624 38907
rect 24596 38848 24808 38876
rect 24780 38820 24808 38848
rect 22060 38780 24256 38808
rect 22060 38768 22066 38780
rect 24762 38768 24768 38820
rect 24820 38768 24826 38820
rect 24872 38808 24900 38907
rect 24946 38904 24952 38956
rect 25004 38904 25010 38956
rect 25222 38904 25228 38956
rect 25280 38904 25286 38956
rect 25373 38950 25431 38953
rect 25373 38947 25452 38950
rect 25373 38913 25385 38947
rect 25419 38913 25452 38947
rect 25373 38907 25452 38913
rect 25424 38876 25452 38907
rect 25498 38904 25504 38956
rect 25556 38904 25562 38956
rect 25608 38953 25636 38984
rect 27249 38981 27261 38984
rect 27295 38981 27307 39015
rect 27249 38975 27307 38981
rect 27433 39015 27491 39021
rect 27433 38981 27445 39015
rect 27479 38981 27491 39015
rect 27433 38975 27491 38981
rect 25593 38947 25651 38953
rect 25593 38913 25605 38947
rect 25639 38913 25651 38947
rect 25593 38907 25651 38913
rect 25731 38947 25789 38953
rect 25731 38913 25743 38947
rect 25777 38944 25789 38947
rect 26050 38944 26056 38956
rect 25777 38916 26056 38944
rect 25777 38913 25789 38916
rect 25731 38907 25789 38913
rect 26050 38904 26056 38916
rect 26108 38904 26114 38956
rect 26142 38904 26148 38956
rect 26200 38904 26206 38956
rect 26329 38947 26387 38953
rect 26329 38913 26341 38947
rect 26375 38913 26387 38947
rect 26329 38907 26387 38913
rect 26421 38947 26479 38953
rect 26421 38913 26433 38947
rect 26467 38913 26479 38947
rect 26421 38907 26479 38913
rect 25958 38876 25964 38888
rect 25424 38848 25964 38876
rect 25958 38836 25964 38848
rect 26016 38836 26022 38888
rect 26068 38876 26096 38904
rect 26344 38876 26372 38907
rect 26068 38848 26372 38876
rect 26436 38876 26464 38907
rect 26510 38904 26516 38956
rect 26568 38904 26574 38956
rect 26694 38876 26700 38888
rect 26436 38848 26700 38876
rect 26528 38820 26556 38848
rect 26694 38836 26700 38848
rect 26752 38836 26758 38888
rect 25038 38808 25044 38820
rect 24872 38780 25044 38808
rect 25038 38768 25044 38780
rect 25096 38768 25102 38820
rect 25133 38811 25191 38817
rect 25133 38777 25145 38811
rect 25179 38808 25191 38811
rect 26142 38808 26148 38820
rect 25179 38780 26148 38808
rect 25179 38777 25191 38780
rect 25133 38771 25191 38777
rect 26142 38768 26148 38780
rect 26200 38808 26206 38820
rect 26200 38780 26372 38808
rect 26200 38768 26206 38780
rect 17586 38700 17592 38752
rect 17644 38740 17650 38752
rect 18417 38743 18475 38749
rect 18417 38740 18429 38743
rect 17644 38712 18429 38740
rect 17644 38700 17650 38712
rect 18417 38709 18429 38712
rect 18463 38709 18475 38743
rect 18417 38703 18475 38709
rect 18601 38743 18659 38749
rect 18601 38709 18613 38743
rect 18647 38740 18659 38743
rect 21174 38740 21180 38752
rect 18647 38712 21180 38740
rect 18647 38709 18659 38712
rect 18601 38703 18659 38709
rect 21174 38700 21180 38712
rect 21232 38700 21238 38752
rect 22094 38700 22100 38752
rect 22152 38740 22158 38752
rect 22189 38743 22247 38749
rect 22189 38740 22201 38743
rect 22152 38712 22201 38740
rect 22152 38700 22158 38712
rect 22189 38709 22201 38712
rect 22235 38709 22247 38743
rect 22189 38703 22247 38709
rect 22370 38700 22376 38752
rect 22428 38740 22434 38752
rect 22465 38743 22523 38749
rect 22465 38740 22477 38743
rect 22428 38712 22477 38740
rect 22428 38700 22434 38712
rect 22465 38709 22477 38712
rect 22511 38709 22523 38743
rect 22465 38703 22523 38709
rect 22554 38700 22560 38752
rect 22612 38700 22618 38752
rect 23109 38743 23167 38749
rect 23109 38709 23121 38743
rect 23155 38740 23167 38743
rect 23750 38740 23756 38752
rect 23155 38712 23756 38740
rect 23155 38709 23167 38712
rect 23109 38703 23167 38709
rect 23750 38700 23756 38712
rect 23808 38700 23814 38752
rect 24489 38743 24547 38749
rect 24489 38709 24501 38743
rect 24535 38740 24547 38743
rect 26234 38740 26240 38752
rect 24535 38712 26240 38740
rect 24535 38709 24547 38712
rect 24489 38703 24547 38709
rect 26234 38700 26240 38712
rect 26292 38700 26298 38752
rect 26344 38740 26372 38780
rect 26510 38768 26516 38820
rect 26568 38768 26574 38820
rect 27264 38808 27292 38975
rect 27706 38904 27712 38956
rect 27764 38904 27770 38956
rect 27890 38904 27896 38956
rect 27948 38904 27954 38956
rect 27982 38904 27988 38956
rect 28040 38904 28046 38956
rect 28092 38953 28120 39052
rect 28534 39040 28540 39052
rect 28592 39040 28598 39092
rect 29089 39083 29147 39089
rect 29089 39049 29101 39083
rect 29135 39080 29147 39083
rect 29546 39080 29552 39092
rect 29135 39052 29552 39080
rect 29135 39049 29147 39052
rect 29089 39043 29147 39049
rect 29546 39040 29552 39052
rect 29604 39040 29610 39092
rect 31478 39040 31484 39092
rect 31536 39040 31542 39092
rect 31570 39040 31576 39092
rect 31628 39080 31634 39092
rect 31628 39052 31708 39080
rect 31628 39040 31634 39052
rect 28626 38972 28632 39024
rect 28684 38972 28690 39024
rect 28810 38972 28816 39024
rect 28868 39012 28874 39024
rect 29825 39015 29883 39021
rect 29825 39012 29837 39015
rect 28868 38984 29837 39012
rect 28868 38972 28874 38984
rect 29825 38981 29837 38984
rect 29871 38981 29883 39015
rect 31018 39012 31024 39024
rect 29825 38975 29883 38981
rect 30024 38984 31024 39012
rect 28077 38947 28135 38953
rect 28077 38913 28089 38947
rect 28123 38913 28135 38947
rect 28905 38947 28963 38953
rect 29199 38950 29257 38953
rect 28905 38944 28917 38947
rect 28077 38907 28135 38913
rect 28184 38942 28580 38944
rect 28644 38942 28917 38944
rect 28184 38916 28917 38942
rect 27614 38836 27620 38888
rect 27672 38876 27678 38888
rect 28092 38876 28120 38907
rect 27672 38848 28120 38876
rect 27672 38836 27678 38848
rect 28184 38808 28212 38916
rect 28552 38914 28672 38916
rect 28905 38913 28917 38916
rect 28951 38913 28963 38947
rect 29105 38947 29257 38950
rect 29105 38944 29211 38947
rect 28905 38907 28963 38913
rect 29012 38922 29211 38944
rect 29012 38916 29133 38922
rect 29196 38916 29211 38922
rect 28721 38879 28779 38885
rect 28721 38876 28733 38879
rect 28276 38848 28733 38876
rect 28276 38817 28304 38848
rect 28721 38845 28733 38848
rect 28767 38876 28779 38879
rect 29012 38876 29040 38916
rect 29199 38913 29211 38916
rect 29245 38913 29257 38947
rect 29365 38947 29423 38953
rect 29365 38944 29377 38947
rect 29199 38907 29257 38913
rect 29288 38916 29377 38944
rect 28767 38848 29040 38876
rect 28767 38845 28779 38848
rect 28721 38839 28779 38845
rect 27264 38780 28212 38808
rect 28261 38811 28319 38817
rect 28261 38777 28273 38811
rect 28307 38777 28319 38811
rect 28261 38771 28319 38777
rect 28465 38780 28764 38808
rect 28465 38740 28493 38780
rect 28736 38752 28764 38780
rect 26344 38712 28493 38740
rect 28534 38700 28540 38752
rect 28592 38740 28598 38752
rect 28629 38743 28687 38749
rect 28629 38740 28641 38743
rect 28592 38712 28641 38740
rect 28592 38700 28598 38712
rect 28629 38709 28641 38712
rect 28675 38709 28687 38743
rect 28629 38703 28687 38709
rect 28718 38700 28724 38752
rect 28776 38700 28782 38752
rect 28810 38700 28816 38752
rect 28868 38740 28874 38752
rect 29288 38740 29316 38916
rect 29365 38913 29377 38916
rect 29411 38913 29423 38947
rect 29365 38907 29423 38913
rect 29638 38904 29644 38956
rect 29696 38904 29702 38956
rect 29549 38879 29607 38885
rect 29549 38845 29561 38879
rect 29595 38876 29607 38879
rect 30024 38876 30052 38984
rect 31018 38972 31024 38984
rect 31076 38972 31082 39024
rect 31680 39012 31708 39052
rect 32490 39040 32496 39092
rect 32548 39040 32554 39092
rect 32582 39040 32588 39092
rect 32640 39040 32646 39092
rect 33045 39083 33103 39089
rect 33045 39049 33057 39083
rect 33091 39080 33103 39083
rect 33502 39080 33508 39092
rect 33091 39052 33508 39080
rect 33091 39049 33103 39052
rect 33045 39043 33103 39049
rect 33502 39040 33508 39052
rect 33560 39040 33566 39092
rect 31496 38984 31708 39012
rect 30098 38904 30104 38956
rect 30156 38944 30162 38956
rect 30285 38947 30343 38953
rect 30285 38944 30297 38947
rect 30156 38916 30297 38944
rect 30156 38904 30162 38916
rect 30285 38913 30297 38916
rect 30331 38913 30343 38947
rect 30285 38907 30343 38913
rect 31337 38947 31395 38953
rect 31337 38913 31349 38947
rect 31383 38944 31395 38947
rect 31496 38944 31524 38984
rect 31383 38916 31524 38944
rect 31383 38913 31395 38916
rect 31337 38907 31395 38913
rect 31570 38904 31576 38956
rect 31628 38904 31634 38956
rect 29595 38848 30052 38876
rect 30377 38879 30435 38885
rect 29595 38845 29607 38848
rect 29549 38839 29607 38845
rect 30377 38845 30389 38879
rect 30423 38876 30435 38879
rect 30466 38876 30472 38888
rect 30423 38848 30472 38876
rect 30423 38845 30435 38848
rect 30377 38839 30435 38845
rect 30466 38836 30472 38848
rect 30524 38836 30530 38888
rect 31110 38836 31116 38888
rect 31168 38836 31174 38888
rect 30009 38811 30067 38817
rect 30009 38777 30021 38811
rect 30055 38808 30067 38811
rect 31680 38808 31708 38984
rect 31938 38972 31944 39024
rect 31996 39012 32002 39024
rect 32508 39012 32536 39040
rect 31996 38984 32352 39012
rect 32508 38984 33456 39012
rect 31996 38972 32002 38984
rect 31754 38904 31760 38956
rect 31812 38904 31818 38956
rect 32122 38904 32128 38956
rect 32180 38904 32186 38956
rect 32214 38836 32220 38888
rect 32272 38836 32278 38888
rect 32324 38876 32352 38984
rect 32398 38904 32404 38956
rect 32456 38904 32462 38956
rect 32677 38947 32735 38953
rect 32677 38913 32689 38947
rect 32723 38913 32735 38947
rect 32677 38907 32735 38913
rect 32692 38876 32720 38907
rect 32766 38904 32772 38956
rect 32824 38904 32830 38956
rect 33428 38953 33456 38984
rect 34606 38972 34612 39024
rect 34664 38972 34670 39024
rect 33413 38947 33471 38953
rect 33413 38913 33425 38947
rect 33459 38913 33471 38947
rect 33413 38907 33471 38913
rect 33594 38904 33600 38956
rect 33652 38904 33658 38956
rect 33873 38879 33931 38885
rect 33873 38876 33885 38879
rect 32324 38848 32720 38876
rect 33244 38848 33885 38876
rect 33244 38817 33272 38848
rect 33873 38845 33885 38848
rect 33919 38845 33931 38879
rect 33873 38839 33931 38845
rect 31941 38811 31999 38817
rect 31941 38808 31953 38811
rect 30055 38780 31064 38808
rect 31680 38780 31953 38808
rect 30055 38777 30067 38780
rect 30009 38771 30067 38777
rect 31036 38752 31064 38780
rect 31941 38777 31953 38780
rect 31987 38777 31999 38811
rect 31941 38771 31999 38777
rect 33229 38811 33287 38817
rect 33229 38777 33241 38811
rect 33275 38777 33287 38811
rect 33229 38771 33287 38777
rect 28868 38712 29316 38740
rect 28868 38700 28874 38712
rect 30282 38700 30288 38752
rect 30340 38700 30346 38752
rect 30650 38700 30656 38752
rect 30708 38700 30714 38752
rect 31018 38700 31024 38752
rect 31076 38700 31082 38752
rect 31202 38700 31208 38752
rect 31260 38740 31266 38752
rect 31573 38743 31631 38749
rect 31573 38740 31585 38743
rect 31260 38712 31585 38740
rect 31260 38700 31266 38712
rect 31573 38709 31585 38712
rect 31619 38709 31631 38743
rect 31573 38703 31631 38709
rect 31846 38700 31852 38752
rect 31904 38740 31910 38752
rect 32125 38743 32183 38749
rect 32125 38740 32137 38743
rect 31904 38712 32137 38740
rect 31904 38700 31910 38712
rect 32125 38709 32137 38712
rect 32171 38709 32183 38743
rect 32125 38703 32183 38709
rect 32674 38700 32680 38752
rect 32732 38700 32738 38752
rect 35342 38700 35348 38752
rect 35400 38700 35406 38752
rect 1104 38650 41400 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 41400 38650
rect 1104 38576 41400 38598
rect 17313 38539 17371 38545
rect 17313 38536 17325 38539
rect 13004 38508 17325 38536
rect 13004 38480 13032 38508
rect 17313 38505 17325 38508
rect 17359 38536 17371 38539
rect 17862 38536 17868 38548
rect 17359 38508 17868 38536
rect 17359 38505 17371 38508
rect 17313 38499 17371 38505
rect 17862 38496 17868 38508
rect 17920 38496 17926 38548
rect 17954 38496 17960 38548
rect 18012 38496 18018 38548
rect 18141 38539 18199 38545
rect 18141 38505 18153 38539
rect 18187 38536 18199 38539
rect 18230 38536 18236 38548
rect 18187 38508 18236 38536
rect 18187 38505 18199 38508
rect 18141 38499 18199 38505
rect 18230 38496 18236 38508
rect 18288 38536 18294 38548
rect 23477 38539 23535 38545
rect 18288 38508 21588 38536
rect 18288 38496 18294 38508
rect 12986 38428 12992 38480
rect 13044 38428 13050 38480
rect 15381 38471 15439 38477
rect 15381 38437 15393 38471
rect 15427 38468 15439 38471
rect 15427 38440 20208 38468
rect 15427 38437 15439 38440
rect 15381 38431 15439 38437
rect 9582 38360 9588 38412
rect 9640 38400 9646 38412
rect 11422 38400 11428 38412
rect 9640 38372 11428 38400
rect 9640 38360 9646 38372
rect 11422 38360 11428 38372
rect 11480 38400 11486 38412
rect 11517 38403 11575 38409
rect 11517 38400 11529 38403
rect 11480 38372 11529 38400
rect 11480 38360 11486 38372
rect 11517 38369 11529 38372
rect 11563 38369 11575 38403
rect 11517 38363 11575 38369
rect 12250 38360 12256 38412
rect 12308 38400 12314 38412
rect 12308 38372 15884 38400
rect 12308 38360 12314 38372
rect 13446 38332 13452 38344
rect 12926 38304 13452 38332
rect 13446 38292 13452 38304
rect 13504 38292 13510 38344
rect 15565 38335 15623 38341
rect 15565 38301 15577 38335
rect 15611 38301 15623 38335
rect 15565 38295 15623 38301
rect 15657 38335 15715 38341
rect 15657 38301 15669 38335
rect 15703 38301 15715 38335
rect 15856 38332 15884 38372
rect 15930 38360 15936 38412
rect 15988 38360 15994 38412
rect 16025 38403 16083 38409
rect 16025 38369 16037 38403
rect 16071 38400 16083 38403
rect 17678 38400 17684 38412
rect 16071 38372 17684 38400
rect 16071 38369 16083 38372
rect 16025 38363 16083 38369
rect 17678 38360 17684 38372
rect 17736 38360 17742 38412
rect 17770 38360 17776 38412
rect 17828 38400 17834 38412
rect 17828 38372 18184 38400
rect 17828 38360 17834 38372
rect 15856 38304 16804 38332
rect 15657 38295 15715 38301
rect 11790 38224 11796 38276
rect 11848 38224 11854 38276
rect 13538 38224 13544 38276
rect 13596 38224 13602 38276
rect 15580 38208 15608 38295
rect 15672 38208 15700 38295
rect 16209 38267 16267 38273
rect 16209 38233 16221 38267
rect 16255 38233 16267 38267
rect 16209 38227 16267 38233
rect 16393 38267 16451 38273
rect 16393 38233 16405 38267
rect 16439 38264 16451 38267
rect 16776 38264 16804 38304
rect 17218 38292 17224 38344
rect 17276 38332 17282 38344
rect 18156 38341 18184 38372
rect 18414 38360 18420 38412
rect 18472 38400 18478 38412
rect 19426 38400 19432 38412
rect 18472 38372 19432 38400
rect 18472 38360 18478 38372
rect 19426 38360 19432 38372
rect 19484 38360 19490 38412
rect 17865 38335 17923 38341
rect 17865 38332 17877 38335
rect 17276 38304 17877 38332
rect 17276 38292 17282 38304
rect 17865 38301 17877 38304
rect 17911 38301 17923 38335
rect 17865 38295 17923 38301
rect 18141 38335 18199 38341
rect 18141 38301 18153 38335
rect 18187 38301 18199 38335
rect 18141 38295 18199 38301
rect 18230 38292 18236 38344
rect 18288 38332 18294 38344
rect 18325 38335 18383 38341
rect 18325 38332 18337 38335
rect 18288 38304 18337 38332
rect 18288 38292 18294 38304
rect 18325 38301 18337 38304
rect 18371 38301 18383 38335
rect 18325 38295 18383 38301
rect 19794 38292 19800 38344
rect 19852 38332 19858 38344
rect 19981 38335 20039 38341
rect 19981 38332 19993 38335
rect 19852 38304 19993 38332
rect 19852 38292 19858 38304
rect 19981 38301 19993 38304
rect 20027 38301 20039 38335
rect 20180 38332 20208 38440
rect 20530 38428 20536 38480
rect 20588 38468 20594 38480
rect 21453 38471 21511 38477
rect 21453 38468 21465 38471
rect 20588 38440 21465 38468
rect 20588 38428 20594 38440
rect 21453 38437 21465 38440
rect 21499 38437 21511 38471
rect 21453 38431 21511 38437
rect 20898 38360 20904 38412
rect 20956 38360 20962 38412
rect 21174 38360 21180 38412
rect 21232 38400 21238 38412
rect 21560 38400 21588 38508
rect 23477 38505 23489 38539
rect 23523 38536 23535 38539
rect 23934 38536 23940 38548
rect 23523 38508 23940 38536
rect 23523 38505 23535 38508
rect 23477 38499 23535 38505
rect 23934 38496 23940 38508
rect 23992 38496 23998 38548
rect 25130 38496 25136 38548
rect 25188 38536 25194 38548
rect 25774 38536 25780 38548
rect 25188 38508 25780 38536
rect 25188 38496 25194 38508
rect 25774 38496 25780 38508
rect 25832 38496 25838 38548
rect 25866 38496 25872 38548
rect 25924 38496 25930 38548
rect 25958 38496 25964 38548
rect 26016 38536 26022 38548
rect 26016 38508 27023 38536
rect 26016 38496 26022 38508
rect 22830 38428 22836 38480
rect 22888 38468 22894 38480
rect 22888 38440 24716 38468
rect 22888 38428 22894 38440
rect 24688 38412 24716 38440
rect 25590 38428 25596 38480
rect 25648 38468 25654 38480
rect 26329 38471 26387 38477
rect 25648 38440 26152 38468
rect 25648 38428 25654 38440
rect 23474 38400 23480 38412
rect 21232 38372 21404 38400
rect 21560 38372 23480 38400
rect 21232 38360 21238 38372
rect 21376 38341 21404 38372
rect 23474 38360 23480 38372
rect 23532 38400 23538 38412
rect 24397 38403 24455 38409
rect 24397 38400 24409 38403
rect 23532 38372 24409 38400
rect 23532 38360 23538 38372
rect 24397 38369 24409 38372
rect 24443 38369 24455 38403
rect 24397 38363 24455 38369
rect 24670 38360 24676 38412
rect 24728 38360 24734 38412
rect 24854 38360 24860 38412
rect 24912 38400 24918 38412
rect 24912 38372 25452 38400
rect 24912 38360 24918 38372
rect 21085 38335 21143 38341
rect 21085 38332 21097 38335
rect 20180 38304 21097 38332
rect 19981 38295 20039 38301
rect 21085 38301 21097 38304
rect 21131 38301 21143 38335
rect 21085 38295 21143 38301
rect 21361 38335 21419 38341
rect 21361 38301 21373 38335
rect 21407 38301 21419 38335
rect 21361 38295 21419 38301
rect 21453 38335 21511 38341
rect 21453 38301 21465 38335
rect 21499 38332 21511 38335
rect 21542 38332 21548 38344
rect 21499 38304 21548 38332
rect 21499 38301 21511 38304
rect 21453 38295 21511 38301
rect 21542 38292 21548 38304
rect 21600 38292 21606 38344
rect 21637 38335 21695 38341
rect 21637 38301 21649 38335
rect 21683 38332 21695 38335
rect 22738 38332 22744 38344
rect 21683 38304 22744 38332
rect 21683 38301 21695 38304
rect 21637 38295 21695 38301
rect 21174 38264 21180 38276
rect 16439 38236 16712 38264
rect 16776 38236 21180 38264
rect 16439 38233 16451 38236
rect 16393 38227 16451 38233
rect 15562 38156 15568 38208
rect 15620 38156 15626 38208
rect 15654 38156 15660 38208
rect 15712 38156 15718 38208
rect 15746 38156 15752 38208
rect 15804 38196 15810 38208
rect 16224 38196 16252 38227
rect 16684 38208 16712 38236
rect 21174 38224 21180 38236
rect 21232 38224 21238 38276
rect 21269 38267 21327 38273
rect 21269 38233 21281 38267
rect 21315 38264 21327 38267
rect 21652 38264 21680 38295
rect 22738 38292 22744 38304
rect 22796 38292 22802 38344
rect 23109 38335 23167 38341
rect 23109 38301 23121 38335
rect 23155 38332 23167 38335
rect 23198 38332 23204 38344
rect 23155 38304 23204 38332
rect 23155 38301 23167 38304
rect 23109 38295 23167 38301
rect 21315 38236 21680 38264
rect 21315 38233 21327 38236
rect 21269 38227 21327 38233
rect 22554 38224 22560 38276
rect 22612 38264 22618 38276
rect 23124 38264 23152 38295
rect 23198 38292 23204 38304
rect 23256 38292 23262 38344
rect 23290 38292 23296 38344
rect 23348 38292 23354 38344
rect 24581 38335 24639 38341
rect 24581 38301 24593 38335
rect 24627 38301 24639 38335
rect 24581 38295 24639 38301
rect 24765 38335 24823 38341
rect 24765 38301 24777 38335
rect 24811 38332 24823 38335
rect 25038 38332 25044 38344
rect 24811 38304 25044 38332
rect 24811 38301 24823 38304
rect 24765 38295 24823 38301
rect 24596 38264 24624 38295
rect 25038 38292 25044 38304
rect 25096 38292 25102 38344
rect 25424 38341 25452 38372
rect 25682 38360 25688 38412
rect 25740 38400 25746 38412
rect 25961 38403 26019 38409
rect 25961 38400 25973 38403
rect 25740 38372 25973 38400
rect 25740 38360 25746 38372
rect 25961 38369 25973 38372
rect 26007 38369 26019 38403
rect 26124 38400 26152 38440
rect 26329 38437 26341 38471
rect 26375 38468 26387 38471
rect 26878 38468 26884 38480
rect 26375 38440 26884 38468
rect 26375 38437 26387 38440
rect 26329 38431 26387 38437
rect 26878 38428 26884 38440
rect 26936 38428 26942 38480
rect 26995 38468 27023 38508
rect 27062 38496 27068 38548
rect 27120 38496 27126 38548
rect 27798 38536 27804 38548
rect 27545 38508 27804 38536
rect 27545 38468 27573 38508
rect 27798 38496 27804 38508
rect 27856 38496 27862 38548
rect 28997 38539 29055 38545
rect 28997 38505 29009 38539
rect 29043 38536 29055 38539
rect 29086 38536 29092 38548
rect 29043 38508 29092 38536
rect 29043 38505 29055 38508
rect 28997 38499 29055 38505
rect 29086 38496 29092 38508
rect 29144 38536 29150 38548
rect 29144 38508 29224 38536
rect 29144 38496 29150 38508
rect 26995 38440 27573 38468
rect 27614 38428 27620 38480
rect 27672 38468 27678 38480
rect 27672 38440 27936 38468
rect 27672 38428 27678 38440
rect 27065 38403 27123 38409
rect 27065 38400 27077 38403
rect 26124 38372 27077 38400
rect 25961 38363 26019 38369
rect 27065 38369 27077 38372
rect 27111 38369 27123 38403
rect 27908 38400 27936 38440
rect 28074 38428 28080 38480
rect 28132 38468 28138 38480
rect 28534 38468 28540 38480
rect 28132 38440 28540 38468
rect 28132 38428 28138 38440
rect 28534 38428 28540 38440
rect 28592 38468 28598 38480
rect 29196 38468 29224 38508
rect 29270 38496 29276 38548
rect 29328 38536 29334 38548
rect 29638 38536 29644 38548
rect 29328 38508 29644 38536
rect 29328 38496 29334 38508
rect 29638 38496 29644 38508
rect 29696 38496 29702 38548
rect 30653 38539 30711 38545
rect 30653 38505 30665 38539
rect 30699 38536 30711 38539
rect 31018 38536 31024 38548
rect 30699 38508 31024 38536
rect 30699 38505 30711 38508
rect 30653 38499 30711 38505
rect 31018 38496 31024 38508
rect 31076 38496 31082 38548
rect 31297 38539 31355 38545
rect 31297 38505 31309 38539
rect 31343 38536 31355 38539
rect 31478 38536 31484 38548
rect 31343 38508 31484 38536
rect 31343 38505 31355 38508
rect 31297 38499 31355 38505
rect 31478 38496 31484 38508
rect 31536 38536 31542 38548
rect 32122 38536 32128 38548
rect 31536 38508 32128 38536
rect 31536 38496 31542 38508
rect 32122 38496 32128 38508
rect 32180 38496 32186 38548
rect 28592 38440 29158 38468
rect 29196 38440 31248 38468
rect 28592 38428 28598 38440
rect 28994 38400 29000 38412
rect 27908 38372 29000 38400
rect 27065 38363 27123 38369
rect 28994 38360 29000 38372
rect 29052 38360 29058 38412
rect 29130 38400 29158 38440
rect 29270 38400 29276 38412
rect 29130 38372 29276 38400
rect 29270 38360 29276 38372
rect 29328 38360 29334 38412
rect 30466 38360 30472 38412
rect 30524 38360 30530 38412
rect 25409 38335 25467 38341
rect 25409 38301 25421 38335
rect 25455 38332 25467 38335
rect 25774 38332 25780 38344
rect 25455 38304 25780 38332
rect 25455 38301 25467 38304
rect 25409 38295 25467 38301
rect 25774 38292 25780 38304
rect 25832 38292 25838 38344
rect 26142 38292 26148 38344
rect 26200 38292 26206 38344
rect 27246 38292 27252 38344
rect 27304 38292 27310 38344
rect 27614 38332 27620 38344
rect 27356 38304 27620 38332
rect 22612 38236 24624 38264
rect 22612 38224 22618 38236
rect 25130 38224 25136 38276
rect 25188 38264 25194 38276
rect 25225 38267 25283 38273
rect 25225 38264 25237 38267
rect 25188 38236 25237 38264
rect 25188 38224 25194 38236
rect 25225 38233 25237 38236
rect 25271 38233 25283 38267
rect 25225 38227 25283 38233
rect 25314 38224 25320 38276
rect 25372 38224 25378 38276
rect 25866 38224 25872 38276
rect 25924 38224 25930 38276
rect 26973 38267 27031 38273
rect 26973 38233 26985 38267
rect 27019 38264 27031 38267
rect 27356 38264 27384 38304
rect 27614 38292 27620 38304
rect 27672 38292 27678 38344
rect 27890 38292 27896 38344
rect 27948 38332 27954 38344
rect 30484 38332 30512 38360
rect 27948 38304 30512 38332
rect 27948 38292 27954 38304
rect 30558 38292 30564 38344
rect 30616 38332 30622 38344
rect 30653 38335 30711 38341
rect 30653 38332 30665 38335
rect 30616 38304 30665 38332
rect 30616 38292 30622 38304
rect 30653 38301 30665 38304
rect 30699 38301 30711 38335
rect 31113 38335 31171 38341
rect 31113 38332 31125 38335
rect 30653 38295 30711 38301
rect 30760 38304 31125 38332
rect 27019 38236 27384 38264
rect 27019 38233 27031 38236
rect 26973 38227 27031 38233
rect 27706 38224 27712 38276
rect 27764 38264 27770 38276
rect 28629 38267 28687 38273
rect 28629 38264 28641 38267
rect 27764 38236 28641 38264
rect 27764 38224 27770 38236
rect 28629 38233 28641 38236
rect 28675 38233 28687 38267
rect 28629 38227 28687 38233
rect 28718 38224 28724 38276
rect 28776 38264 28782 38276
rect 28813 38267 28871 38273
rect 28813 38264 28825 38267
rect 28776 38236 28825 38264
rect 28776 38224 28782 38236
rect 28813 38233 28825 38236
rect 28859 38233 28871 38267
rect 28813 38227 28871 38233
rect 29822 38224 29828 38276
rect 29880 38264 29886 38276
rect 30006 38264 30012 38276
rect 29880 38236 30012 38264
rect 29880 38224 29886 38236
rect 30006 38224 30012 38236
rect 30064 38224 30070 38276
rect 30374 38224 30380 38276
rect 30432 38224 30438 38276
rect 15804 38168 16252 38196
rect 15804 38156 15810 38168
rect 16482 38156 16488 38208
rect 16540 38156 16546 38208
rect 16574 38156 16580 38208
rect 16632 38156 16638 38208
rect 16666 38156 16672 38208
rect 16724 38156 16730 38208
rect 16758 38156 16764 38208
rect 16816 38156 16822 38208
rect 19334 38156 19340 38208
rect 19392 38196 19398 38208
rect 20165 38199 20223 38205
rect 20165 38196 20177 38199
rect 19392 38168 20177 38196
rect 19392 38156 19398 38168
rect 20165 38165 20177 38168
rect 20211 38196 20223 38199
rect 21542 38196 21548 38208
rect 20211 38168 21548 38196
rect 20211 38165 20223 38168
rect 20165 38159 20223 38165
rect 21542 38156 21548 38168
rect 21600 38156 21606 38208
rect 22278 38156 22284 38208
rect 22336 38196 22342 38208
rect 23290 38196 23296 38208
rect 22336 38168 23296 38196
rect 22336 38156 22342 38168
rect 23290 38156 23296 38168
rect 23348 38156 23354 38208
rect 24946 38156 24952 38208
rect 25004 38196 25010 38208
rect 26878 38196 26884 38208
rect 25004 38168 26884 38196
rect 25004 38156 25010 38168
rect 26878 38156 26884 38168
rect 26936 38156 26942 38208
rect 27433 38199 27491 38205
rect 27433 38165 27445 38199
rect 27479 38196 27491 38199
rect 30190 38196 30196 38208
rect 27479 38168 30196 38196
rect 27479 38165 27491 38168
rect 27433 38159 27491 38165
rect 30190 38156 30196 38168
rect 30248 38156 30254 38208
rect 30282 38156 30288 38208
rect 30340 38196 30346 38208
rect 30760 38196 30788 38304
rect 31113 38301 31125 38304
rect 31159 38301 31171 38335
rect 31113 38295 31171 38301
rect 30929 38267 30987 38273
rect 30929 38233 30941 38267
rect 30975 38264 30987 38267
rect 31220 38264 31248 38440
rect 30975 38236 31248 38264
rect 30975 38233 30987 38236
rect 30929 38227 30987 38233
rect 30340 38168 30788 38196
rect 30340 38156 30346 38168
rect 30834 38156 30840 38208
rect 30892 38156 30898 38208
rect 1104 38106 41400 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 41400 38106
rect 1104 38032 41400 38054
rect 11790 37952 11796 38004
rect 11848 37992 11854 38004
rect 12897 37995 12955 38001
rect 12897 37992 12909 37995
rect 11848 37964 12909 37992
rect 11848 37952 11854 37964
rect 12897 37961 12909 37964
rect 12943 37961 12955 37995
rect 12897 37955 12955 37961
rect 13078 37952 13084 38004
rect 13136 37992 13142 38004
rect 17129 37995 17187 38001
rect 13136 37964 16896 37992
rect 13136 37952 13142 37964
rect 9030 37924 9036 37936
rect 8786 37896 9036 37924
rect 9030 37884 9036 37896
rect 9088 37884 9094 37936
rect 10594 37884 10600 37936
rect 10652 37884 10658 37936
rect 11974 37884 11980 37936
rect 12032 37924 12038 37936
rect 12434 37924 12440 37936
rect 12032 37896 12440 37924
rect 12032 37884 12038 37896
rect 12434 37884 12440 37896
rect 12492 37924 12498 37936
rect 13383 37927 13441 37933
rect 13383 37924 13395 37927
rect 12492 37896 13395 37924
rect 12492 37884 12498 37896
rect 13383 37893 13395 37896
rect 13429 37893 13441 37927
rect 13383 37887 13441 37893
rect 14274 37884 14280 37936
rect 14332 37884 14338 37936
rect 15654 37924 15660 37936
rect 15212 37896 15660 37924
rect 12986 37816 12992 37868
rect 13044 37816 13050 37868
rect 13078 37816 13084 37868
rect 13136 37816 13142 37868
rect 13173 37859 13231 37865
rect 13173 37825 13185 37859
rect 13219 37825 13231 37859
rect 13173 37819 13231 37825
rect 13265 37859 13323 37865
rect 13265 37825 13277 37859
rect 13311 37856 13323 37859
rect 13630 37856 13636 37868
rect 13311 37828 13636 37856
rect 13311 37825 13323 37828
rect 13265 37819 13323 37825
rect 6914 37748 6920 37800
rect 6972 37788 6978 37800
rect 7285 37791 7343 37797
rect 7285 37788 7297 37791
rect 6972 37760 7297 37788
rect 6972 37748 6978 37760
rect 7285 37757 7297 37760
rect 7331 37757 7343 37791
rect 7285 37751 7343 37757
rect 7558 37748 7564 37800
rect 7616 37748 7622 37800
rect 8570 37748 8576 37800
rect 8628 37788 8634 37800
rect 9582 37788 9588 37800
rect 8628 37760 9588 37788
rect 8628 37748 8634 37760
rect 9582 37748 9588 37760
rect 9640 37748 9646 37800
rect 9861 37791 9919 37797
rect 9861 37757 9873 37791
rect 9907 37788 9919 37791
rect 11514 37788 11520 37800
rect 9907 37760 11520 37788
rect 9907 37757 9919 37760
rect 9861 37751 9919 37757
rect 11514 37748 11520 37760
rect 11572 37748 11578 37800
rect 12434 37748 12440 37800
rect 12492 37748 12498 37800
rect 13004 37788 13032 37816
rect 13188 37788 13216 37819
rect 13630 37816 13636 37828
rect 13688 37856 13694 37868
rect 14292 37856 14320 37884
rect 13688 37828 14320 37856
rect 13688 37816 13694 37828
rect 15010 37816 15016 37868
rect 15068 37816 15074 37868
rect 15212 37865 15240 37896
rect 15654 37884 15660 37896
rect 15712 37924 15718 37936
rect 16301 37927 16359 37933
rect 16301 37924 16313 37927
rect 15712 37896 16313 37924
rect 15712 37884 15718 37896
rect 16301 37893 16313 37896
rect 16347 37893 16359 37927
rect 16301 37887 16359 37893
rect 15197 37859 15255 37865
rect 15197 37825 15209 37859
rect 15243 37825 15255 37859
rect 15562 37856 15568 37868
rect 15197 37819 15255 37825
rect 15304 37828 15568 37856
rect 13004 37760 13216 37788
rect 13538 37748 13544 37800
rect 13596 37748 13602 37800
rect 15028 37788 15056 37816
rect 15304 37788 15332 37828
rect 15562 37816 15568 37828
rect 15620 37816 15626 37868
rect 15933 37859 15991 37865
rect 15933 37825 15945 37859
rect 15979 37856 15991 37859
rect 16022 37856 16028 37868
rect 15979 37828 16028 37856
rect 15979 37825 15991 37828
rect 15933 37819 15991 37825
rect 16022 37816 16028 37828
rect 16080 37816 16086 37868
rect 16114 37816 16120 37868
rect 16172 37816 16178 37868
rect 16209 37859 16267 37865
rect 16209 37825 16221 37859
rect 16255 37856 16267 37859
rect 16255 37828 16344 37856
rect 16255 37825 16267 37828
rect 16209 37819 16267 37825
rect 15028 37760 15332 37788
rect 15378 37748 15384 37800
rect 15436 37788 15442 37800
rect 15473 37791 15531 37797
rect 15473 37788 15485 37791
rect 15436 37760 15485 37788
rect 15436 37748 15442 37760
rect 15473 37757 15485 37760
rect 15519 37757 15531 37791
rect 15580 37788 15608 37816
rect 16316 37800 16344 37828
rect 16390 37816 16396 37868
rect 16448 37816 16454 37868
rect 15580 37760 15792 37788
rect 15473 37751 15531 37757
rect 12452 37720 12480 37748
rect 13556 37720 13584 37748
rect 12452 37692 13584 37720
rect 15013 37723 15071 37729
rect 15013 37689 15025 37723
rect 15059 37720 15071 37723
rect 15657 37723 15715 37729
rect 15657 37720 15669 37723
rect 15059 37692 15669 37720
rect 15059 37689 15071 37692
rect 15013 37683 15071 37689
rect 15657 37689 15669 37692
rect 15703 37689 15715 37723
rect 15764 37720 15792 37760
rect 15838 37748 15844 37800
rect 15896 37788 15902 37800
rect 15896 37760 16160 37788
rect 15896 37748 15902 37760
rect 16025 37723 16083 37729
rect 16025 37720 16037 37723
rect 15764 37692 16037 37720
rect 15657 37683 15715 37689
rect 16025 37689 16037 37692
rect 16071 37689 16083 37723
rect 16132 37720 16160 37760
rect 16298 37748 16304 37800
rect 16356 37748 16362 37800
rect 16666 37748 16672 37800
rect 16724 37788 16730 37800
rect 16761 37791 16819 37797
rect 16761 37788 16773 37791
rect 16724 37760 16773 37788
rect 16724 37748 16730 37760
rect 16761 37757 16773 37760
rect 16807 37757 16819 37791
rect 16868 37788 16896 37964
rect 17129 37961 17141 37995
rect 17175 37992 17187 37995
rect 17218 37992 17224 38004
rect 17175 37964 17224 37992
rect 17175 37961 17187 37964
rect 17129 37955 17187 37961
rect 17218 37952 17224 37964
rect 17276 37952 17282 38004
rect 17862 37952 17868 38004
rect 17920 37992 17926 38004
rect 17920 37964 19380 37992
rect 17920 37952 17926 37964
rect 19245 37927 19303 37933
rect 19245 37893 19257 37927
rect 19291 37893 19303 37927
rect 19245 37887 19303 37893
rect 16942 37816 16948 37868
rect 17000 37816 17006 37868
rect 18874 37816 18880 37868
rect 18932 37856 18938 37868
rect 19260 37856 19288 37887
rect 18932 37828 19288 37856
rect 19352 37856 19380 37964
rect 19426 37952 19432 38004
rect 19484 38001 19490 38004
rect 19484 37995 19503 38001
rect 19491 37961 19503 37995
rect 19484 37955 19503 37961
rect 19613 37995 19671 38001
rect 19613 37961 19625 37995
rect 19659 37992 19671 37995
rect 19978 37992 19984 38004
rect 19659 37964 19984 37992
rect 19659 37961 19671 37964
rect 19613 37955 19671 37961
rect 19484 37952 19490 37955
rect 19978 37952 19984 37964
rect 20036 37952 20042 38004
rect 23290 37992 23296 38004
rect 21560 37964 23296 37992
rect 19996 37924 20024 37952
rect 21560 37936 21588 37964
rect 23290 37952 23296 37964
rect 23348 37992 23354 38004
rect 25590 37992 25596 38004
rect 23348 37964 25596 37992
rect 23348 37952 23354 37964
rect 25590 37952 25596 37964
rect 25648 37992 25654 38004
rect 26510 37992 26516 38004
rect 25648 37964 26516 37992
rect 25648 37952 25654 37964
rect 26510 37952 26516 37964
rect 26568 37952 26574 38004
rect 26878 37952 26884 38004
rect 26936 37992 26942 38004
rect 27522 37992 27528 38004
rect 26936 37964 27528 37992
rect 26936 37952 26942 37964
rect 19904 37896 20024 37924
rect 20073 37927 20131 37933
rect 19904 37865 19932 37896
rect 20073 37893 20085 37927
rect 20119 37924 20131 37927
rect 20438 37924 20444 37936
rect 20119 37896 20444 37924
rect 20119 37893 20131 37896
rect 20073 37887 20131 37893
rect 20438 37884 20444 37896
rect 20496 37884 20502 37936
rect 21542 37884 21548 37936
rect 21600 37884 21606 37936
rect 21726 37884 21732 37936
rect 21784 37924 21790 37936
rect 22646 37924 22652 37936
rect 21784 37896 22652 37924
rect 21784 37884 21790 37896
rect 22646 37884 22652 37896
rect 22704 37924 22710 37936
rect 23106 37924 23112 37936
rect 22704 37896 23112 37924
rect 22704 37884 22710 37896
rect 23106 37884 23112 37896
rect 23164 37924 23170 37936
rect 23385 37927 23443 37933
rect 23385 37924 23397 37927
rect 23164 37896 23397 37924
rect 23164 37884 23170 37896
rect 23385 37893 23397 37896
rect 23431 37893 23443 37927
rect 27453 37924 27481 37964
rect 27522 37952 27528 37964
rect 27580 37952 27586 38004
rect 27614 37952 27620 38004
rect 27672 37952 27678 38004
rect 27822 37964 28580 37992
rect 27822 37924 27850 37964
rect 28350 37933 28356 37936
rect 28261 37927 28319 37933
rect 28261 37924 28273 37927
rect 23385 37887 23443 37893
rect 26896 37896 27109 37924
rect 19889 37859 19947 37865
rect 19352 37828 19840 37856
rect 18932 37816 18938 37828
rect 19334 37788 19340 37800
rect 16868 37760 19340 37788
rect 16761 37751 16819 37757
rect 19334 37748 19340 37760
rect 19392 37748 19398 37800
rect 19812 37788 19840 37828
rect 19889 37825 19901 37859
rect 19935 37825 19947 37859
rect 19889 37819 19947 37825
rect 19978 37816 19984 37868
rect 20036 37816 20042 37868
rect 20211 37859 20269 37865
rect 20211 37825 20223 37859
rect 20257 37856 20269 37859
rect 20714 37856 20720 37868
rect 20257 37828 20720 37856
rect 20257 37825 20269 37828
rect 20211 37819 20269 37825
rect 20714 37816 20720 37828
rect 20772 37816 20778 37868
rect 22370 37816 22376 37868
rect 22428 37856 22434 37868
rect 22830 37856 22836 37868
rect 22428 37828 22836 37856
rect 22428 37816 22434 37828
rect 22830 37816 22836 37828
rect 22888 37856 22894 37868
rect 23201 37859 23259 37865
rect 23201 37856 23213 37859
rect 22888 37828 23213 37856
rect 22888 37816 22894 37828
rect 23201 37825 23213 37828
rect 23247 37825 23259 37859
rect 23201 37819 23259 37825
rect 23290 37816 23296 37868
rect 23348 37816 23354 37868
rect 23503 37859 23561 37865
rect 23503 37825 23515 37859
rect 23549 37825 23561 37859
rect 23503 37819 23561 37825
rect 23661 37859 23719 37865
rect 23661 37825 23673 37859
rect 23707 37856 23719 37859
rect 24118 37856 24124 37868
rect 23707 37828 24124 37856
rect 23707 37825 23719 37828
rect 23661 37819 23719 37825
rect 19996 37788 20024 37816
rect 19812 37760 20024 37788
rect 20070 37748 20076 37800
rect 20128 37788 20134 37800
rect 20349 37791 20407 37797
rect 20349 37788 20361 37791
rect 20128 37760 20361 37788
rect 20128 37748 20134 37760
rect 20349 37757 20361 37760
rect 20395 37757 20407 37791
rect 20349 37751 20407 37757
rect 21726 37748 21732 37800
rect 21784 37788 21790 37800
rect 22186 37788 22192 37800
rect 21784 37760 22192 37788
rect 21784 37748 21790 37760
rect 22186 37748 22192 37760
rect 22244 37748 22250 37800
rect 22738 37748 22744 37800
rect 22796 37788 22802 37800
rect 23518 37788 23546 37819
rect 24118 37816 24124 37828
rect 24176 37816 24182 37868
rect 24486 37816 24492 37868
rect 24544 37856 24550 37868
rect 24670 37856 24676 37868
rect 24544 37828 24676 37856
rect 24544 37816 24550 37828
rect 24670 37816 24676 37828
rect 24728 37816 24734 37868
rect 26694 37816 26700 37868
rect 26752 37856 26758 37868
rect 26896 37856 26924 37896
rect 26752 37828 26924 37856
rect 26752 37816 26758 37828
rect 26970 37816 26976 37868
rect 27028 37816 27034 37868
rect 27081 37865 27109 37896
rect 27453 37896 27850 37924
rect 27908 37896 28273 37924
rect 27453 37865 27481 37896
rect 27066 37859 27124 37865
rect 27066 37825 27078 37859
rect 27112 37825 27124 37859
rect 27066 37819 27124 37825
rect 27249 37859 27307 37865
rect 27249 37825 27261 37859
rect 27295 37825 27307 37859
rect 27249 37819 27307 37825
rect 27341 37859 27399 37865
rect 27341 37825 27353 37859
rect 27387 37825 27399 37859
rect 27341 37819 27399 37825
rect 27438 37859 27496 37865
rect 27438 37825 27450 37859
rect 27484 37825 27496 37859
rect 27438 37819 27496 37825
rect 24946 37788 24952 37800
rect 22796 37760 24952 37788
rect 22796 37748 22802 37760
rect 24946 37748 24952 37760
rect 25004 37748 25010 37800
rect 25130 37748 25136 37800
rect 25188 37788 25194 37800
rect 25958 37788 25964 37800
rect 25188 37760 25964 37788
rect 25188 37748 25194 37760
rect 25958 37748 25964 37760
rect 26016 37748 26022 37800
rect 26418 37748 26424 37800
rect 26476 37788 26482 37800
rect 27264 37788 27292 37819
rect 26476 37760 27292 37788
rect 27356 37788 27384 37819
rect 27706 37816 27712 37868
rect 27764 37816 27770 37868
rect 27798 37816 27804 37868
rect 27856 37856 27862 37868
rect 27908 37856 27936 37896
rect 28261 37893 28273 37896
rect 28307 37893 28319 37927
rect 28261 37887 28319 37893
rect 28349 37887 28356 37933
rect 28350 37884 28356 37887
rect 28408 37884 28414 37936
rect 27856 37828 27936 37856
rect 28077 37859 28135 37865
rect 27856 37816 27862 37828
rect 28077 37825 28089 37859
rect 28123 37856 28135 37859
rect 28445 37859 28503 37865
rect 28123 37828 28304 37856
rect 28123 37825 28135 37828
rect 28077 37819 28135 37825
rect 27522 37788 27528 37800
rect 27356 37760 27528 37788
rect 26476 37748 26482 37760
rect 27522 37748 27528 37760
rect 27580 37748 27586 37800
rect 18414 37720 18420 37732
rect 16132 37692 18420 37720
rect 16025 37683 16083 37689
rect 18414 37680 18420 37692
rect 18472 37680 18478 37732
rect 18506 37680 18512 37732
rect 18564 37720 18570 37732
rect 19705 37723 19763 37729
rect 18564 37692 19472 37720
rect 18564 37680 18570 37692
rect 18800 37664 18828 37692
rect 9030 37612 9036 37664
rect 9088 37612 9094 37664
rect 10318 37612 10324 37664
rect 10376 37652 10382 37664
rect 11333 37655 11391 37661
rect 11333 37652 11345 37655
rect 10376 37624 11345 37652
rect 10376 37612 10382 37624
rect 11333 37621 11345 37624
rect 11379 37652 11391 37655
rect 12158 37652 12164 37664
rect 11379 37624 12164 37652
rect 11379 37621 11391 37624
rect 11333 37615 11391 37621
rect 12158 37612 12164 37624
rect 12216 37612 12222 37664
rect 15381 37655 15439 37661
rect 15381 37621 15393 37655
rect 15427 37652 15439 37655
rect 15470 37652 15476 37664
rect 15427 37624 15476 37652
rect 15427 37621 15439 37624
rect 15381 37615 15439 37621
rect 15470 37612 15476 37624
rect 15528 37612 15534 37664
rect 15746 37612 15752 37664
rect 15804 37612 15810 37664
rect 18782 37612 18788 37664
rect 18840 37612 18846 37664
rect 18874 37612 18880 37664
rect 18932 37612 18938 37664
rect 19444 37661 19472 37692
rect 19705 37689 19717 37723
rect 19751 37720 19763 37723
rect 27724 37720 27752 37816
rect 28276 37800 28304 37828
rect 28445 37825 28457 37859
rect 28491 37846 28503 37859
rect 28552 37846 28580 37964
rect 28626 37952 28632 38004
rect 28684 37952 28690 38004
rect 28994 37952 29000 38004
rect 29052 37992 29058 38004
rect 29641 37995 29699 38001
rect 29052 37964 29408 37992
rect 29052 37952 29058 37964
rect 28491 37825 28580 37846
rect 28644 37856 28672 37952
rect 29270 37884 29276 37936
rect 29328 37884 29334 37936
rect 29380 37933 29408 37964
rect 29641 37961 29653 37995
rect 29687 37992 29699 37995
rect 30098 37992 30104 38004
rect 29687 37964 30104 37992
rect 29687 37961 29699 37964
rect 29641 37955 29699 37961
rect 30098 37952 30104 37964
rect 30156 37952 30162 38004
rect 30834 37952 30840 38004
rect 30892 37952 30898 38004
rect 31941 37995 31999 38001
rect 31941 37961 31953 37995
rect 31987 37961 31999 37995
rect 31941 37955 31999 37961
rect 29365 37927 29423 37933
rect 29365 37893 29377 37927
rect 29411 37893 29423 37927
rect 29365 37887 29423 37893
rect 28997 37859 29055 37865
rect 28997 37856 29009 37859
rect 28644 37828 29009 37856
rect 28445 37819 28580 37825
rect 28997 37825 29009 37828
rect 29043 37825 29055 37859
rect 28997 37819 29055 37825
rect 28460 37818 28580 37819
rect 29086 37816 29092 37868
rect 29144 37856 29150 37868
rect 29503 37859 29561 37865
rect 29144 37828 29189 37856
rect 29144 37816 29150 37828
rect 29503 37825 29515 37859
rect 29549 37856 29561 37859
rect 30006 37856 30012 37868
rect 29549 37828 30012 37856
rect 29549 37825 29561 37828
rect 29503 37819 29561 37825
rect 30006 37816 30012 37828
rect 30064 37816 30070 37868
rect 28258 37748 28264 37800
rect 28316 37748 28322 37800
rect 28626 37748 28632 37800
rect 28684 37788 28690 37800
rect 30558 37788 30564 37800
rect 28684 37760 30564 37788
rect 28684 37748 28690 37760
rect 30558 37748 30564 37760
rect 30616 37748 30622 37800
rect 19751 37692 27752 37720
rect 19751 37689 19763 37692
rect 19705 37683 19763 37689
rect 27798 37680 27804 37732
rect 27856 37720 27862 37732
rect 30466 37720 30472 37732
rect 27856 37692 30472 37720
rect 27856 37680 27862 37692
rect 30466 37680 30472 37692
rect 30524 37680 30530 37732
rect 30852 37720 30880 37952
rect 31956 37924 31984 37955
rect 33594 37952 33600 38004
rect 33652 37952 33658 38004
rect 34422 37952 34428 38004
rect 34480 37992 34486 38004
rect 34480 37964 35112 37992
rect 34480 37952 34486 37964
rect 33612 37924 33640 37952
rect 31956 37896 32352 37924
rect 31294 37816 31300 37868
rect 31352 37856 31358 37868
rect 31481 37859 31539 37865
rect 31481 37856 31493 37859
rect 31352 37828 31493 37856
rect 31352 37816 31358 37828
rect 31481 37825 31493 37828
rect 31527 37825 31539 37859
rect 31481 37819 31539 37825
rect 31662 37816 31668 37868
rect 31720 37856 31726 37868
rect 31757 37859 31815 37865
rect 31757 37856 31769 37859
rect 31720 37828 31769 37856
rect 31720 37816 31726 37828
rect 31757 37825 31769 37828
rect 31803 37825 31815 37859
rect 31757 37819 31815 37825
rect 32214 37816 32220 37868
rect 32272 37816 32278 37868
rect 32324 37865 32352 37896
rect 33520 37896 33640 37924
rect 33520 37865 33548 37896
rect 33686 37884 33692 37936
rect 33744 37924 33750 37936
rect 33781 37927 33839 37933
rect 33781 37924 33793 37927
rect 33744 37896 33793 37924
rect 33744 37884 33750 37896
rect 33781 37893 33793 37896
rect 33827 37893 33839 37927
rect 35084 37924 35112 37964
rect 38562 37924 38568 37936
rect 35006 37896 38568 37924
rect 33781 37887 33839 37893
rect 38562 37884 38568 37896
rect 38620 37884 38626 37936
rect 32309 37859 32367 37865
rect 32309 37825 32321 37859
rect 32355 37825 32367 37859
rect 32309 37819 32367 37825
rect 33505 37859 33563 37865
rect 33505 37825 33517 37859
rect 33551 37825 33563 37859
rect 33505 37819 33563 37825
rect 31202 37748 31208 37800
rect 31260 37788 31266 37800
rect 31573 37791 31631 37797
rect 31573 37788 31585 37791
rect 31260 37760 31585 37788
rect 31260 37748 31266 37760
rect 31573 37757 31585 37760
rect 31619 37788 31631 37791
rect 31938 37788 31944 37800
rect 31619 37760 31944 37788
rect 31619 37757 31631 37760
rect 31573 37751 31631 37757
rect 31938 37748 31944 37760
rect 31996 37748 32002 37800
rect 30852 37692 32260 37720
rect 19429 37655 19487 37661
rect 19429 37621 19441 37655
rect 19475 37621 19487 37655
rect 19429 37615 19487 37621
rect 23017 37655 23075 37661
rect 23017 37621 23029 37655
rect 23063 37652 23075 37655
rect 23382 37652 23388 37664
rect 23063 37624 23388 37652
rect 23063 37621 23075 37624
rect 23017 37615 23075 37621
rect 23382 37612 23388 37624
rect 23440 37612 23446 37664
rect 23474 37612 23480 37664
rect 23532 37652 23538 37664
rect 31110 37652 31116 37664
rect 23532 37624 31116 37652
rect 23532 37612 23538 37624
rect 31110 37612 31116 37624
rect 31168 37612 31174 37664
rect 31478 37612 31484 37664
rect 31536 37612 31542 37664
rect 32232 37661 32260 37692
rect 32217 37655 32275 37661
rect 32217 37621 32229 37655
rect 32263 37621 32275 37655
rect 32217 37615 32275 37621
rect 32585 37655 32643 37661
rect 32585 37621 32597 37655
rect 32631 37652 32643 37655
rect 33134 37652 33140 37664
rect 32631 37624 33140 37652
rect 32631 37621 32643 37624
rect 32585 37615 32643 37621
rect 33134 37612 33140 37624
rect 33192 37612 33198 37664
rect 34790 37612 34796 37664
rect 34848 37652 34854 37664
rect 35253 37655 35311 37661
rect 35253 37652 35265 37655
rect 34848 37624 35265 37652
rect 34848 37612 34854 37624
rect 35253 37621 35265 37624
rect 35299 37621 35311 37655
rect 35253 37615 35311 37621
rect 1104 37562 41400 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 41400 37562
rect 1104 37488 41400 37510
rect 7558 37408 7564 37460
rect 7616 37448 7622 37460
rect 8297 37451 8355 37457
rect 8297 37448 8309 37451
rect 7616 37420 8309 37448
rect 7616 37408 7622 37420
rect 8297 37417 8309 37420
rect 8343 37417 8355 37451
rect 8297 37411 8355 37417
rect 11514 37408 11520 37460
rect 11572 37408 11578 37460
rect 15746 37448 15752 37460
rect 12406 37420 15752 37448
rect 12406 37380 12434 37420
rect 15746 37408 15752 37420
rect 15804 37408 15810 37460
rect 16298 37408 16304 37460
rect 16356 37448 16362 37460
rect 18233 37451 18291 37457
rect 18233 37448 18245 37451
rect 16356 37420 18245 37448
rect 16356 37408 16362 37420
rect 18233 37417 18245 37420
rect 18279 37448 18291 37451
rect 18322 37448 18328 37460
rect 18279 37420 18328 37448
rect 18279 37417 18291 37420
rect 18233 37411 18291 37417
rect 18322 37408 18328 37420
rect 18380 37408 18386 37460
rect 20714 37408 20720 37460
rect 20772 37448 20778 37460
rect 21358 37448 21364 37460
rect 20772 37420 21364 37448
rect 20772 37408 20778 37420
rect 21358 37408 21364 37420
rect 21416 37408 21422 37460
rect 22278 37408 22284 37460
rect 22336 37448 22342 37460
rect 23017 37451 23075 37457
rect 23017 37448 23029 37451
rect 22336 37420 23029 37448
rect 22336 37408 22342 37420
rect 23017 37417 23029 37420
rect 23063 37417 23075 37451
rect 23017 37411 23075 37417
rect 23382 37408 23388 37460
rect 23440 37408 23446 37460
rect 23474 37408 23480 37460
rect 23532 37408 23538 37460
rect 25958 37408 25964 37460
rect 26016 37408 26022 37460
rect 26878 37408 26884 37460
rect 26936 37448 26942 37460
rect 29086 37448 29092 37460
rect 26936 37420 29092 37448
rect 26936 37408 26942 37420
rect 29086 37408 29092 37420
rect 29144 37448 29150 37460
rect 29822 37448 29828 37460
rect 29144 37420 29828 37448
rect 29144 37408 29150 37420
rect 29822 37408 29828 37420
rect 29880 37408 29886 37460
rect 30101 37451 30159 37457
rect 30101 37417 30113 37451
rect 30147 37448 30159 37451
rect 30282 37448 30288 37460
rect 30147 37420 30288 37448
rect 30147 37417 30159 37420
rect 30101 37411 30159 37417
rect 30282 37408 30288 37420
rect 30340 37408 30346 37460
rect 30558 37408 30564 37460
rect 30616 37448 30622 37460
rect 31757 37451 31815 37457
rect 31757 37448 31769 37451
rect 30616 37420 31769 37448
rect 30616 37408 30622 37420
rect 10152 37352 12434 37380
rect 8757 37315 8815 37321
rect 8757 37281 8769 37315
rect 8803 37312 8815 37315
rect 9585 37315 9643 37321
rect 9585 37312 9597 37315
rect 8803 37284 9597 37312
rect 8803 37281 8815 37284
rect 8757 37275 8815 37281
rect 9585 37281 9597 37284
rect 9631 37281 9643 37315
rect 9585 37275 9643 37281
rect 8481 37247 8539 37253
rect 8481 37213 8493 37247
rect 8527 37213 8539 37247
rect 8481 37207 8539 37213
rect 8496 37176 8524 37207
rect 8662 37204 8668 37256
rect 8720 37204 8726 37256
rect 9030 37204 9036 37256
rect 9088 37204 9094 37256
rect 10152 37176 10180 37352
rect 12526 37340 12532 37392
rect 12584 37380 12590 37392
rect 12713 37383 12771 37389
rect 12713 37380 12725 37383
rect 12584 37352 12725 37380
rect 12584 37340 12590 37352
rect 12713 37349 12725 37352
rect 12759 37349 12771 37383
rect 12713 37343 12771 37349
rect 12894 37340 12900 37392
rect 12952 37380 12958 37392
rect 18874 37380 18880 37392
rect 12952 37352 18880 37380
rect 12952 37340 12958 37352
rect 18874 37340 18880 37352
rect 18932 37340 18938 37392
rect 21542 37340 21548 37392
rect 21600 37380 21606 37392
rect 21600 37352 22600 37380
rect 21600 37340 21606 37352
rect 10318 37272 10324 37324
rect 10376 37272 10382 37324
rect 11256 37284 11468 37312
rect 10965 37247 11023 37253
rect 10965 37213 10977 37247
rect 11011 37244 11023 37247
rect 11256 37244 11284 37284
rect 11011 37216 11284 37244
rect 11011 37213 11023 37216
rect 10965 37207 11023 37213
rect 11330 37204 11336 37256
rect 11388 37204 11394 37256
rect 11440 37244 11468 37284
rect 11514 37272 11520 37324
rect 11572 37312 11578 37324
rect 13633 37315 13691 37321
rect 13633 37312 13645 37315
rect 11572 37284 13645 37312
rect 11572 37272 11578 37284
rect 13633 37281 13645 37284
rect 13679 37281 13691 37315
rect 15470 37312 15476 37324
rect 13633 37275 13691 37281
rect 15212 37284 15476 37312
rect 12529 37247 12587 37253
rect 11440 37216 12434 37244
rect 8496 37148 10180 37176
rect 11146 37136 11152 37188
rect 11204 37136 11210 37188
rect 11241 37179 11299 37185
rect 11241 37145 11253 37179
rect 11287 37145 11299 37179
rect 11345 37176 11373 37204
rect 11974 37176 11980 37188
rect 11345 37148 11980 37176
rect 11241 37139 11299 37145
rect 10873 37111 10931 37117
rect 10873 37077 10885 37111
rect 10919 37108 10931 37111
rect 11256 37108 11284 37139
rect 11974 37136 11980 37148
rect 12032 37136 12038 37188
rect 10919 37080 11284 37108
rect 12406 37108 12434 37216
rect 12529 37213 12541 37247
rect 12575 37213 12587 37247
rect 12529 37207 12587 37213
rect 12989 37247 13047 37253
rect 12989 37213 13001 37247
rect 13035 37244 13047 37247
rect 13078 37244 13084 37256
rect 13035 37216 13084 37244
rect 13035 37213 13047 37216
rect 12989 37207 13047 37213
rect 12544 37176 12572 37207
rect 13078 37204 13084 37216
rect 13136 37204 13142 37256
rect 15010 37204 15016 37256
rect 15068 37204 15074 37256
rect 15212 37253 15240 37284
rect 15470 37272 15476 37284
rect 15528 37312 15534 37324
rect 16209 37315 16267 37321
rect 16209 37312 16221 37315
rect 15528 37284 15792 37312
rect 15528 37272 15534 37284
rect 15764 37256 15792 37284
rect 15948 37284 16221 37312
rect 15948 37256 15976 37284
rect 16209 37281 16221 37284
rect 16255 37312 16267 37315
rect 16482 37312 16488 37324
rect 16255 37284 16488 37312
rect 16255 37281 16267 37284
rect 16209 37275 16267 37281
rect 16482 37272 16488 37284
rect 16540 37312 16546 37324
rect 19150 37312 19156 37324
rect 16540 37284 19156 37312
rect 16540 37272 16546 37284
rect 15197 37247 15255 37253
rect 15197 37213 15209 37247
rect 15243 37213 15255 37247
rect 15197 37207 15255 37213
rect 15286 37204 15292 37256
rect 15344 37204 15350 37256
rect 15746 37204 15752 37256
rect 15804 37204 15810 37256
rect 15930 37204 15936 37256
rect 15988 37204 15994 37256
rect 16022 37204 16028 37256
rect 16080 37244 16086 37256
rect 16117 37247 16175 37253
rect 16117 37244 16129 37247
rect 16080 37216 16129 37244
rect 16080 37204 16086 37216
rect 16117 37213 16129 37216
rect 16163 37213 16175 37247
rect 16117 37207 16175 37213
rect 16574 37204 16580 37256
rect 16632 37244 16638 37256
rect 17405 37247 17463 37253
rect 17405 37244 17417 37247
rect 16632 37216 17417 37244
rect 16632 37204 16638 37216
rect 17405 37213 17417 37216
rect 17451 37213 17463 37247
rect 17405 37207 17463 37213
rect 17589 37247 17647 37253
rect 17589 37213 17601 37247
rect 17635 37213 17647 37247
rect 17589 37207 17647 37213
rect 13541 37179 13599 37185
rect 12544 37148 13124 37176
rect 12710 37108 12716 37120
rect 12406 37080 12716 37108
rect 10919 37077 10931 37080
rect 10873 37071 10931 37077
rect 12710 37068 12716 37080
rect 12768 37068 12774 37120
rect 12897 37111 12955 37117
rect 12897 37077 12909 37111
rect 12943 37108 12955 37111
rect 12986 37108 12992 37120
rect 12943 37080 12992 37108
rect 12943 37077 12955 37080
rect 12897 37071 12955 37077
rect 12986 37068 12992 37080
rect 13044 37068 13050 37120
rect 13096 37117 13124 37148
rect 13541 37145 13553 37179
rect 13587 37176 13599 37179
rect 13630 37176 13636 37188
rect 13587 37148 13636 37176
rect 13587 37145 13599 37148
rect 13541 37139 13599 37145
rect 13630 37136 13636 37148
rect 13688 37136 13694 37188
rect 15105 37179 15163 37185
rect 15105 37176 15117 37179
rect 15028 37148 15117 37176
rect 15028 37120 15056 37148
rect 15105 37145 15117 37148
rect 15151 37145 15163 37179
rect 15105 37139 15163 37145
rect 15654 37136 15660 37188
rect 15712 37176 15718 37188
rect 17218 37176 17224 37188
rect 15712 37148 17224 37176
rect 15712 37136 15718 37148
rect 17218 37136 17224 37148
rect 17276 37136 17282 37188
rect 13081 37111 13139 37117
rect 13081 37077 13093 37111
rect 13127 37077 13139 37111
rect 13081 37071 13139 37077
rect 13170 37068 13176 37120
rect 13228 37108 13234 37120
rect 13449 37111 13507 37117
rect 13449 37108 13461 37111
rect 13228 37080 13461 37108
rect 13228 37068 13234 37080
rect 13449 37077 13461 37080
rect 13495 37108 13507 37111
rect 14274 37108 14280 37120
rect 13495 37080 14280 37108
rect 13495 37077 13507 37080
rect 13449 37071 13507 37077
rect 14274 37068 14280 37080
rect 14332 37068 14338 37120
rect 15010 37068 15016 37120
rect 15068 37068 15074 37120
rect 15378 37068 15384 37120
rect 15436 37108 15442 37120
rect 17604 37108 17632 37207
rect 18138 37204 18144 37256
rect 18196 37244 18202 37256
rect 18708 37253 18736 37284
rect 19150 37272 19156 37284
rect 19208 37272 19214 37324
rect 22186 37272 22192 37324
rect 22244 37312 22250 37324
rect 22572 37312 22600 37352
rect 22833 37315 22891 37321
rect 22833 37312 22845 37315
rect 22244 37284 22508 37312
rect 22572 37284 22845 37312
rect 22244 37272 22250 37284
rect 18509 37247 18567 37253
rect 18509 37244 18521 37247
rect 18196 37216 18521 37244
rect 18196 37204 18202 37216
rect 18509 37213 18521 37216
rect 18555 37213 18567 37247
rect 18509 37207 18567 37213
rect 18693 37247 18751 37253
rect 18693 37213 18705 37247
rect 18739 37213 18751 37247
rect 19426 37244 19432 37256
rect 18693 37207 18751 37213
rect 18800 37216 19432 37244
rect 17770 37136 17776 37188
rect 17828 37136 17834 37188
rect 18049 37179 18107 37185
rect 18049 37176 18061 37179
rect 17972 37148 18061 37176
rect 17972 37120 18000 37148
rect 18049 37145 18061 37148
rect 18095 37145 18107 37179
rect 18049 37139 18107 37145
rect 15436 37080 17632 37108
rect 15436 37068 15442 37080
rect 17954 37068 17960 37120
rect 18012 37068 18018 37120
rect 18156 37108 18184 37204
rect 18265 37179 18323 37185
rect 18265 37145 18277 37179
rect 18311 37176 18323 37179
rect 18800 37176 18828 37216
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 20441 37247 20499 37253
rect 20441 37213 20453 37247
rect 20487 37244 20499 37247
rect 20530 37244 20536 37256
rect 20487 37216 20536 37244
rect 20487 37213 20499 37216
rect 20441 37207 20499 37213
rect 20530 37204 20536 37216
rect 20588 37204 20594 37256
rect 22480 37253 22508 37284
rect 22833 37281 22845 37284
rect 22879 37281 22891 37315
rect 23400 37312 23428 37408
rect 24486 37340 24492 37392
rect 24544 37380 24550 37392
rect 25222 37380 25228 37392
rect 24544 37352 25228 37380
rect 24544 37340 24550 37352
rect 25222 37340 25228 37352
rect 25280 37340 25286 37392
rect 25498 37340 25504 37392
rect 25556 37380 25562 37392
rect 26789 37383 26847 37389
rect 25556 37352 26740 37380
rect 25556 37340 25562 37352
rect 25958 37312 25964 37324
rect 23400 37284 25964 37312
rect 22833 37275 22891 37281
rect 25958 37272 25964 37284
rect 26016 37272 26022 37324
rect 20625 37247 20683 37253
rect 20625 37213 20637 37247
rect 20671 37213 20683 37247
rect 21913 37247 21971 37253
rect 21913 37244 21925 37247
rect 20625 37207 20683 37213
rect 21008 37216 21925 37244
rect 20640 37176 20668 37207
rect 21008 37188 21036 37216
rect 21913 37213 21925 37216
rect 21959 37213 21971 37247
rect 21913 37207 21971 37213
rect 22005 37247 22063 37253
rect 22005 37213 22017 37247
rect 22051 37244 22063 37247
rect 22373 37247 22431 37253
rect 22373 37244 22385 37247
rect 22051 37216 22385 37244
rect 22051 37213 22063 37216
rect 22005 37207 22063 37213
rect 22373 37213 22385 37216
rect 22419 37213 22431 37247
rect 22373 37207 22431 37213
rect 22465 37247 22523 37253
rect 22465 37213 22477 37247
rect 22511 37213 22523 37247
rect 22465 37207 22523 37213
rect 22557 37247 22615 37253
rect 22557 37213 22569 37247
rect 22603 37244 22615 37247
rect 22603 37216 22876 37244
rect 22603 37213 22615 37216
rect 22557 37207 22615 37213
rect 20990 37176 20996 37188
rect 18311 37148 18828 37176
rect 18892 37148 20996 37176
rect 18311 37145 18323 37148
rect 18265 37139 18323 37145
rect 18892 37120 18920 37148
rect 20990 37136 20996 37148
rect 21048 37136 21054 37188
rect 22738 37185 22744 37188
rect 22695 37179 22744 37185
rect 22695 37145 22707 37179
rect 22741 37145 22744 37179
rect 22695 37139 22744 37145
rect 22738 37136 22744 37139
rect 22796 37136 22802 37188
rect 22848 37176 22876 37216
rect 23014 37204 23020 37256
rect 23072 37204 23078 37256
rect 23106 37204 23112 37256
rect 23164 37204 23170 37256
rect 23201 37247 23259 37253
rect 23201 37213 23213 37247
rect 23247 37213 23259 37247
rect 23201 37207 23259 37213
rect 23293 37247 23351 37253
rect 23293 37213 23305 37247
rect 23339 37244 23351 37247
rect 23382 37244 23388 37256
rect 23339 37216 23388 37244
rect 23339 37213 23351 37216
rect 23293 37207 23351 37213
rect 23124 37176 23152 37204
rect 22848 37148 23152 37176
rect 23216 37176 23244 37207
rect 23382 37204 23388 37216
rect 23440 37204 23446 37256
rect 23474 37204 23480 37256
rect 23532 37244 23538 37256
rect 23532 37216 24992 37244
rect 23532 37204 23538 37216
rect 23658 37176 23664 37188
rect 23216 37148 23664 37176
rect 23658 37136 23664 37148
rect 23716 37136 23722 37188
rect 24964 37176 24992 37216
rect 25038 37204 25044 37256
rect 25096 37244 25102 37256
rect 25409 37247 25467 37253
rect 25409 37244 25421 37247
rect 25096 37216 25421 37244
rect 25096 37204 25102 37216
rect 25409 37213 25421 37216
rect 25455 37213 25467 37247
rect 25409 37207 25467 37213
rect 25590 37204 25596 37256
rect 25648 37204 25654 37256
rect 25682 37204 25688 37256
rect 25740 37204 25746 37256
rect 25774 37204 25780 37256
rect 25832 37204 25838 37256
rect 26237 37247 26295 37253
rect 26237 37244 26249 37247
rect 25884 37216 26249 37244
rect 25884 37176 25912 37216
rect 26237 37213 26249 37216
rect 26283 37213 26295 37247
rect 26237 37207 26295 37213
rect 26326 37204 26332 37256
rect 26384 37244 26390 37256
rect 26605 37247 26663 37253
rect 26605 37244 26617 37247
rect 26384 37216 26617 37244
rect 26384 37204 26390 37216
rect 26605 37213 26617 37216
rect 26651 37213 26663 37247
rect 26712 37244 26740 37352
rect 26789 37349 26801 37383
rect 26835 37380 26847 37383
rect 26970 37380 26976 37392
rect 26835 37352 26976 37380
rect 26835 37349 26847 37352
rect 26789 37343 26847 37349
rect 26970 37340 26976 37352
rect 27028 37340 27034 37392
rect 30024 37352 30328 37380
rect 26988 37312 27016 37340
rect 26896 37284 27016 37312
rect 26896 37253 26924 37284
rect 27614 37272 27620 37324
rect 27672 37312 27678 37324
rect 28718 37312 28724 37324
rect 27672 37284 28724 37312
rect 27672 37272 27678 37284
rect 28718 37272 28724 37284
rect 28776 37312 28782 37324
rect 30024 37312 30052 37352
rect 28776 37284 30052 37312
rect 28776 37272 28782 37284
rect 30098 37272 30104 37324
rect 30156 37312 30162 37324
rect 30300 37321 30328 37352
rect 30466 37340 30472 37392
rect 30524 37380 30530 37392
rect 31018 37380 31024 37392
rect 30524 37352 31024 37380
rect 30524 37340 30530 37352
rect 31018 37340 31024 37352
rect 31076 37340 31082 37392
rect 30285 37315 30343 37321
rect 30156 37284 30236 37312
rect 30156 37272 30162 37284
rect 26881 37247 26939 37253
rect 26712 37216 26832 37244
rect 26605 37207 26663 37213
rect 24964 37148 25912 37176
rect 26418 37136 26424 37188
rect 26476 37136 26482 37188
rect 26510 37136 26516 37188
rect 26568 37136 26574 37188
rect 18417 37111 18475 37117
rect 18417 37108 18429 37111
rect 18156 37080 18429 37108
rect 18417 37077 18429 37080
rect 18463 37077 18475 37111
rect 18417 37071 18475 37077
rect 18598 37068 18604 37120
rect 18656 37068 18662 37120
rect 18874 37068 18880 37120
rect 18932 37068 18938 37120
rect 20530 37068 20536 37120
rect 20588 37068 20594 37120
rect 22189 37111 22247 37117
rect 22189 37077 22201 37111
rect 22235 37108 22247 37111
rect 23382 37108 23388 37120
rect 22235 37080 23388 37108
rect 22235 37077 22247 37080
rect 22189 37071 22247 37077
rect 23382 37068 23388 37080
rect 23440 37068 23446 37120
rect 24394 37068 24400 37120
rect 24452 37108 24458 37120
rect 25406 37108 25412 37120
rect 24452 37080 25412 37108
rect 24452 37068 24458 37080
rect 25406 37068 25412 37080
rect 25464 37068 25470 37120
rect 26804 37108 26832 37216
rect 26881 37213 26893 37247
rect 26927 37213 26939 37247
rect 26881 37207 26939 37213
rect 26970 37204 26976 37256
rect 27028 37244 27034 37256
rect 27387 37247 27445 37253
rect 27028 37216 27073 37244
rect 27028 37204 27034 37216
rect 27387 37213 27399 37247
rect 27433 37244 27445 37247
rect 27522 37244 27528 37256
rect 27433 37216 27528 37244
rect 27433 37213 27445 37216
rect 27387 37207 27445 37213
rect 27522 37204 27528 37216
rect 27580 37204 27586 37256
rect 28258 37204 28264 37256
rect 28316 37244 28322 37256
rect 28534 37244 28540 37256
rect 28316 37216 28540 37244
rect 28316 37204 28322 37216
rect 28534 37204 28540 37216
rect 28592 37204 28598 37256
rect 28626 37204 28632 37256
rect 28684 37244 28690 37256
rect 28684 37216 29040 37244
rect 28684 37204 28690 37216
rect 29012 37188 29040 37216
rect 29362 37204 29368 37256
rect 29420 37244 29426 37256
rect 29549 37247 29607 37253
rect 29549 37244 29561 37247
rect 29420 37216 29561 37244
rect 29420 37204 29426 37216
rect 29549 37213 29561 37216
rect 29595 37213 29607 37247
rect 29549 37207 29607 37213
rect 29917 37247 29975 37253
rect 29917 37213 29929 37247
rect 29963 37244 29975 37247
rect 30006 37244 30012 37256
rect 29963 37216 30012 37244
rect 29963 37213 29975 37216
rect 29917 37207 29975 37213
rect 30006 37204 30012 37216
rect 30064 37204 30070 37256
rect 30208 37244 30236 37284
rect 30285 37281 30297 37315
rect 30331 37281 30343 37315
rect 31202 37312 31208 37324
rect 30285 37275 30343 37281
rect 30576 37284 31208 37312
rect 30469 37247 30527 37253
rect 30469 37244 30481 37247
rect 30208 37216 30481 37244
rect 30469 37213 30481 37216
rect 30515 37213 30527 37247
rect 30469 37207 30527 37213
rect 27157 37179 27215 37185
rect 27157 37145 27169 37179
rect 27203 37145 27215 37179
rect 27157 37139 27215 37145
rect 27249 37179 27307 37185
rect 27249 37145 27261 37179
rect 27295 37145 27307 37179
rect 27249 37139 27307 37145
rect 27172 37108 27200 37139
rect 26804 37080 27200 37108
rect 27264 37108 27292 37139
rect 27982 37136 27988 37188
rect 28040 37176 28046 37188
rect 28718 37176 28724 37188
rect 28040 37148 28724 37176
rect 28040 37136 28046 37148
rect 28718 37136 28724 37148
rect 28776 37136 28782 37188
rect 28994 37136 29000 37188
rect 29052 37136 29058 37188
rect 29730 37136 29736 37188
rect 29788 37136 29794 37188
rect 29825 37179 29883 37185
rect 29825 37145 29837 37179
rect 29871 37176 29883 37179
rect 30098 37176 30104 37188
rect 29871 37148 30104 37176
rect 29871 37145 29883 37148
rect 29825 37139 29883 37145
rect 30098 37136 30104 37148
rect 30156 37136 30162 37188
rect 30190 37136 30196 37188
rect 30248 37136 30254 37188
rect 27338 37108 27344 37120
rect 27264 37080 27344 37108
rect 27338 37068 27344 37080
rect 27396 37068 27402 37120
rect 27525 37111 27583 37117
rect 27525 37077 27537 37111
rect 27571 37108 27583 37111
rect 30576 37108 30604 37284
rect 31202 37272 31208 37284
rect 31260 37272 31266 37324
rect 30650 37204 30656 37256
rect 30708 37204 30714 37256
rect 30834 37204 30840 37256
rect 30892 37204 30898 37256
rect 30926 37204 30932 37256
rect 30984 37204 30990 37256
rect 31317 37253 31345 37420
rect 31757 37417 31769 37420
rect 31803 37417 31815 37451
rect 31757 37411 31815 37417
rect 32125 37451 32183 37457
rect 32125 37417 32137 37451
rect 32171 37417 32183 37451
rect 32125 37411 32183 37417
rect 31302 37247 31360 37253
rect 31302 37213 31314 37247
rect 31348 37213 31360 37247
rect 32140 37244 32168 37411
rect 31302 37207 31360 37213
rect 31496 37216 32168 37244
rect 30668 37176 30696 37204
rect 31113 37179 31171 37185
rect 31113 37176 31125 37179
rect 30668 37148 31125 37176
rect 31113 37145 31125 37148
rect 31159 37145 31171 37179
rect 31113 37139 31171 37145
rect 31202 37136 31208 37188
rect 31260 37136 31266 37188
rect 31496 37176 31524 37216
rect 32306 37204 32312 37256
rect 32364 37204 32370 37256
rect 32398 37204 32404 37256
rect 32456 37204 32462 37256
rect 33134 37204 33140 37256
rect 33192 37244 33198 37256
rect 33597 37247 33655 37253
rect 33597 37244 33609 37247
rect 33192 37216 33609 37244
rect 33192 37204 33198 37216
rect 33597 37213 33609 37216
rect 33643 37213 33655 37247
rect 33597 37207 33655 37213
rect 37550 37204 37556 37256
rect 37608 37244 37614 37256
rect 40773 37247 40831 37253
rect 40773 37244 40785 37247
rect 37608 37216 40785 37244
rect 37608 37204 37614 37216
rect 40773 37213 40785 37216
rect 40819 37213 40831 37247
rect 40773 37207 40831 37213
rect 31312 37148 31524 37176
rect 27571 37080 30604 37108
rect 30653 37111 30711 37117
rect 27571 37077 27583 37080
rect 27525 37071 27583 37077
rect 30653 37077 30665 37111
rect 30699 37108 30711 37111
rect 31312 37108 31340 37148
rect 31570 37136 31576 37188
rect 31628 37176 31634 37188
rect 31665 37179 31723 37185
rect 31665 37176 31677 37179
rect 31628 37148 31677 37176
rect 31628 37136 31634 37148
rect 31665 37145 31677 37148
rect 31711 37145 31723 37179
rect 31665 37139 31723 37145
rect 32122 37136 32128 37188
rect 32180 37136 32186 37188
rect 30699 37080 31340 37108
rect 30699 37077 30711 37080
rect 30653 37071 30711 37077
rect 31478 37068 31484 37120
rect 31536 37068 31542 37120
rect 32582 37068 32588 37120
rect 32640 37068 32646 37120
rect 33410 37068 33416 37120
rect 33468 37068 33474 37120
rect 40954 37068 40960 37120
rect 41012 37068 41018 37120
rect 1104 37018 41400 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 41400 37018
rect 1104 36944 41400 36966
rect 8662 36864 8668 36916
rect 8720 36904 8726 36916
rect 9306 36904 9312 36916
rect 8720 36876 9312 36904
rect 8720 36864 8726 36876
rect 9306 36864 9312 36876
rect 9364 36904 9370 36916
rect 11514 36904 11520 36916
rect 9364 36876 11520 36904
rect 9364 36864 9370 36876
rect 11514 36864 11520 36876
rect 11572 36864 11578 36916
rect 11716 36876 11928 36904
rect 8570 36836 8576 36848
rect 8036 36808 8576 36836
rect 8036 36777 8064 36808
rect 8570 36796 8576 36808
rect 8628 36796 8634 36848
rect 8754 36796 8760 36848
rect 8812 36796 8818 36848
rect 11146 36836 11152 36848
rect 10612 36808 11152 36836
rect 8021 36771 8079 36777
rect 8021 36737 8033 36771
rect 8067 36737 8079 36771
rect 8021 36731 8079 36737
rect 9766 36728 9772 36780
rect 9824 36768 9830 36780
rect 10612 36777 10640 36808
rect 11146 36796 11152 36808
rect 11204 36836 11210 36848
rect 11716 36836 11744 36876
rect 11204 36808 11744 36836
rect 11900 36836 11928 36876
rect 12066 36864 12072 36916
rect 12124 36864 12130 36916
rect 13354 36904 13360 36916
rect 12176 36876 13360 36904
rect 12176 36836 12204 36876
rect 13354 36864 13360 36876
rect 13412 36864 13418 36916
rect 13446 36864 13452 36916
rect 13504 36904 13510 36916
rect 13504 36876 13676 36904
rect 13504 36864 13510 36876
rect 11900 36808 12204 36836
rect 11204 36796 11210 36808
rect 9861 36771 9919 36777
rect 9861 36768 9873 36771
rect 9824 36740 9873 36768
rect 9824 36728 9830 36740
rect 9861 36737 9873 36740
rect 9907 36737 9919 36771
rect 9861 36731 9919 36737
rect 10597 36771 10655 36777
rect 10597 36737 10609 36771
rect 10643 36737 10655 36771
rect 10597 36731 10655 36737
rect 10778 36728 10784 36780
rect 10836 36728 10842 36780
rect 10873 36771 10931 36777
rect 10873 36737 10885 36771
rect 10919 36737 10931 36771
rect 10873 36731 10931 36737
rect 10965 36771 11023 36777
rect 10965 36737 10977 36771
rect 11011 36768 11023 36771
rect 11330 36768 11336 36780
rect 11011 36740 11336 36768
rect 11011 36737 11023 36740
rect 10965 36731 11023 36737
rect 8297 36703 8355 36709
rect 8297 36669 8309 36703
rect 8343 36700 8355 36703
rect 10888 36700 10916 36731
rect 11330 36728 11336 36740
rect 11388 36728 11394 36780
rect 11422 36728 11428 36780
rect 11480 36728 11486 36780
rect 11514 36728 11520 36780
rect 11572 36728 11578 36780
rect 11716 36777 11744 36808
rect 12526 36796 12532 36848
rect 12584 36796 12590 36848
rect 11701 36771 11759 36777
rect 11701 36737 11713 36771
rect 11747 36737 11759 36771
rect 11701 36731 11759 36737
rect 11790 36728 11796 36780
rect 11848 36728 11854 36780
rect 11885 36771 11943 36777
rect 11885 36737 11897 36771
rect 11931 36768 11943 36771
rect 11974 36768 11980 36780
rect 11931 36740 11980 36768
rect 11931 36737 11943 36740
rect 11885 36731 11943 36737
rect 11974 36728 11980 36740
rect 12032 36728 12038 36780
rect 13648 36754 13676 36876
rect 15194 36864 15200 36916
rect 15252 36904 15258 36916
rect 16206 36904 16212 36916
rect 15252 36876 16212 36904
rect 15252 36864 15258 36876
rect 16206 36864 16212 36876
rect 16264 36864 16270 36916
rect 17865 36907 17923 36913
rect 17865 36873 17877 36907
rect 17911 36904 17923 36907
rect 18506 36904 18512 36916
rect 17911 36876 18512 36904
rect 17911 36873 17923 36876
rect 17865 36867 17923 36873
rect 18506 36864 18512 36876
rect 18564 36864 18570 36916
rect 18598 36864 18604 36916
rect 18656 36904 18662 36916
rect 19153 36907 19211 36913
rect 19153 36904 19165 36907
rect 18656 36876 19165 36904
rect 18656 36864 18662 36876
rect 19153 36873 19165 36876
rect 19199 36873 19211 36907
rect 22554 36904 22560 36916
rect 19153 36867 19211 36873
rect 19904 36876 22560 36904
rect 19904 36848 19932 36876
rect 14274 36796 14280 36848
rect 14332 36796 14338 36848
rect 15746 36796 15752 36848
rect 15804 36796 15810 36848
rect 16390 36836 16396 36848
rect 16040 36808 16396 36836
rect 15378 36728 15384 36780
rect 15436 36728 15442 36780
rect 15565 36771 15623 36777
rect 15565 36737 15577 36771
rect 15611 36768 15623 36771
rect 16040 36768 16068 36808
rect 16390 36796 16396 36808
rect 16448 36836 16454 36848
rect 17678 36836 17684 36848
rect 16448 36808 17684 36836
rect 16448 36796 16454 36808
rect 15611 36740 16068 36768
rect 16117 36771 16175 36777
rect 15611 36737 15623 36740
rect 15565 36731 15623 36737
rect 16117 36737 16129 36771
rect 16163 36768 16175 36771
rect 16482 36768 16488 36780
rect 16163 36740 16488 36768
rect 16163 36737 16175 36740
rect 16117 36731 16175 36737
rect 16482 36728 16488 36740
rect 16540 36728 16546 36780
rect 16574 36728 16580 36780
rect 16632 36768 16638 36780
rect 16669 36771 16727 36777
rect 16669 36768 16681 36771
rect 16632 36740 16681 36768
rect 16632 36728 16638 36740
rect 16669 36737 16681 36740
rect 16715 36737 16727 36771
rect 16669 36731 16727 36737
rect 16758 36728 16764 36780
rect 16816 36768 16822 36780
rect 17604 36777 17632 36808
rect 17678 36796 17684 36808
rect 17736 36796 17742 36848
rect 18046 36796 18052 36848
rect 18104 36796 18110 36848
rect 19242 36836 19248 36848
rect 18052 36793 18110 36796
rect 16853 36771 16911 36777
rect 16853 36768 16865 36771
rect 16816 36740 16865 36768
rect 16816 36728 16822 36740
rect 16853 36737 16865 36740
rect 16899 36737 16911 36771
rect 16853 36731 16911 36737
rect 17129 36771 17187 36777
rect 17129 36737 17141 36771
rect 17175 36737 17187 36771
rect 17129 36731 17187 36737
rect 17589 36771 17647 36777
rect 17589 36737 17601 36771
rect 17635 36737 17647 36771
rect 18052 36759 18064 36793
rect 18098 36759 18110 36793
rect 18340 36808 19248 36836
rect 18052 36753 18110 36759
rect 17589 36731 17647 36737
rect 8343 36672 9996 36700
rect 8343 36669 8355 36672
rect 8297 36663 8355 36669
rect 9766 36524 9772 36576
rect 9824 36524 9830 36576
rect 9968 36564 9996 36672
rect 10060 36672 10916 36700
rect 11440 36700 11468 36728
rect 12253 36703 12311 36709
rect 12253 36700 12265 36703
rect 11440 36672 12265 36700
rect 10060 36644 10088 36672
rect 12253 36669 12265 36672
rect 12299 36669 12311 36703
rect 15396 36700 15424 36728
rect 16298 36700 16304 36712
rect 15396 36672 16304 36700
rect 12253 36663 12311 36669
rect 16298 36660 16304 36672
rect 16356 36660 16362 36712
rect 17144 36700 17172 36731
rect 18138 36728 18144 36780
rect 18196 36728 18202 36780
rect 18340 36777 18368 36808
rect 19242 36796 19248 36808
rect 19300 36796 19306 36848
rect 19886 36796 19892 36848
rect 19944 36796 19950 36848
rect 20806 36836 20812 36848
rect 20180 36808 20812 36836
rect 18325 36771 18383 36777
rect 18325 36737 18337 36771
rect 18371 36737 18383 36771
rect 18325 36731 18383 36737
rect 18417 36771 18475 36777
rect 18417 36737 18429 36771
rect 18463 36737 18475 36771
rect 18417 36731 18475 36737
rect 16684 36672 17172 36700
rect 17681 36703 17739 36709
rect 10042 36592 10048 36644
rect 10100 36592 10106 36644
rect 16684 36576 16712 36672
rect 17681 36669 17693 36703
rect 17727 36700 17739 36703
rect 17954 36700 17960 36712
rect 17727 36672 17960 36700
rect 17727 36669 17739 36672
rect 17681 36663 17739 36669
rect 17954 36660 17960 36672
rect 18012 36700 18018 36712
rect 18432 36700 18460 36731
rect 18506 36728 18512 36780
rect 18564 36728 18570 36780
rect 19058 36728 19064 36780
rect 19116 36728 19122 36780
rect 19150 36728 19156 36780
rect 19208 36768 19214 36780
rect 20180 36777 20208 36808
rect 20806 36796 20812 36808
rect 20864 36796 20870 36848
rect 20990 36796 20996 36848
rect 21048 36836 21054 36848
rect 21545 36839 21603 36845
rect 21048 36808 21496 36836
rect 21048 36796 21054 36808
rect 20165 36774 20223 36777
rect 20088 36771 20223 36774
rect 20088 36768 20177 36771
rect 19208 36746 20177 36768
rect 19208 36740 20116 36746
rect 19208 36728 19214 36740
rect 20165 36737 20177 36746
rect 20211 36737 20223 36771
rect 20165 36731 20223 36737
rect 20349 36771 20407 36777
rect 20349 36737 20361 36771
rect 20395 36768 20407 36771
rect 20438 36768 20444 36780
rect 20395 36740 20444 36768
rect 20395 36737 20407 36740
rect 20349 36731 20407 36737
rect 20438 36728 20444 36740
rect 20496 36768 20502 36780
rect 21266 36768 21272 36780
rect 20496 36740 21272 36768
rect 20496 36728 20502 36740
rect 21266 36728 21272 36740
rect 21324 36728 21330 36780
rect 21358 36728 21364 36780
rect 21416 36728 21422 36780
rect 21468 36777 21496 36808
rect 21545 36805 21557 36839
rect 21591 36836 21603 36839
rect 21591 36808 22232 36836
rect 21591 36805 21603 36808
rect 21545 36799 21603 36805
rect 21453 36771 21511 36777
rect 21453 36737 21465 36771
rect 21499 36737 21511 36771
rect 21453 36731 21511 36737
rect 21637 36771 21695 36777
rect 21637 36737 21649 36771
rect 21683 36737 21695 36771
rect 21637 36731 21695 36737
rect 18012 36672 18460 36700
rect 19245 36703 19303 36709
rect 18012 36660 18018 36672
rect 19245 36669 19257 36703
rect 19291 36669 19303 36703
rect 19245 36663 19303 36669
rect 16758 36592 16764 36644
rect 16816 36632 16822 36644
rect 18230 36632 18236 36644
rect 16816 36604 18236 36632
rect 16816 36592 16822 36604
rect 18230 36592 18236 36604
rect 18288 36592 18294 36644
rect 18874 36592 18880 36644
rect 18932 36632 18938 36644
rect 18969 36635 19027 36641
rect 18969 36632 18981 36635
rect 18932 36604 18981 36632
rect 18932 36592 18938 36604
rect 18969 36601 18981 36604
rect 19015 36601 19027 36635
rect 18969 36595 19027 36601
rect 19058 36592 19064 36644
rect 19116 36632 19122 36644
rect 19260 36632 19288 36663
rect 19518 36660 19524 36712
rect 19576 36660 19582 36712
rect 19889 36703 19947 36709
rect 19889 36669 19901 36703
rect 19935 36700 19947 36703
rect 19978 36700 19984 36712
rect 19935 36672 19984 36700
rect 19935 36669 19947 36672
rect 19889 36663 19947 36669
rect 19978 36660 19984 36672
rect 20036 36660 20042 36712
rect 20073 36703 20131 36709
rect 20073 36669 20085 36703
rect 20119 36669 20131 36703
rect 20073 36663 20131 36669
rect 20257 36703 20315 36709
rect 20257 36669 20269 36703
rect 20303 36700 20315 36703
rect 20303 36672 20484 36700
rect 20303 36669 20315 36672
rect 20257 36663 20315 36669
rect 20088 36632 20116 36663
rect 20346 36632 20352 36644
rect 19116 36604 19288 36632
rect 19352 36604 19564 36632
rect 20088 36604 20352 36632
rect 19116 36592 19122 36604
rect 11149 36567 11207 36573
rect 11149 36564 11161 36567
rect 9968 36536 11161 36564
rect 11149 36533 11161 36536
rect 11195 36533 11207 36567
rect 11149 36527 11207 36533
rect 11514 36524 11520 36576
rect 11572 36564 11578 36576
rect 15010 36564 15016 36576
rect 11572 36536 15016 36564
rect 11572 36524 11578 36536
rect 15010 36524 15016 36536
rect 15068 36524 15074 36576
rect 16666 36524 16672 36576
rect 16724 36524 16730 36576
rect 17405 36567 17463 36573
rect 17405 36533 17417 36567
rect 17451 36564 17463 36567
rect 17954 36564 17960 36576
rect 17451 36536 17960 36564
rect 17451 36533 17463 36536
rect 17405 36527 17463 36533
rect 17954 36524 17960 36536
rect 18012 36524 18018 36576
rect 18693 36567 18751 36573
rect 18693 36533 18705 36567
rect 18739 36564 18751 36567
rect 18782 36564 18788 36576
rect 18739 36536 18788 36564
rect 18739 36533 18751 36536
rect 18693 36527 18751 36533
rect 18782 36524 18788 36536
rect 18840 36524 18846 36576
rect 19150 36524 19156 36576
rect 19208 36564 19214 36576
rect 19352 36564 19380 36604
rect 19208 36536 19380 36564
rect 19208 36524 19214 36536
rect 19426 36524 19432 36576
rect 19484 36524 19490 36576
rect 19536 36564 19564 36604
rect 20346 36592 20352 36604
rect 20404 36592 20410 36644
rect 20162 36564 20168 36576
rect 19536 36536 20168 36564
rect 20162 36524 20168 36536
rect 20220 36564 20226 36576
rect 20456 36564 20484 36672
rect 20622 36660 20628 36712
rect 20680 36660 20686 36712
rect 20990 36660 20996 36712
rect 21048 36660 21054 36712
rect 21085 36703 21143 36709
rect 21085 36669 21097 36703
rect 21131 36700 21143 36703
rect 21376 36700 21404 36728
rect 21131 36672 21404 36700
rect 21131 36669 21143 36672
rect 21085 36663 21143 36669
rect 21542 36660 21548 36712
rect 21600 36700 21606 36712
rect 21652 36700 21680 36731
rect 22204 36712 22232 36808
rect 22285 36777 22313 36876
rect 22554 36864 22560 36876
rect 22612 36904 22618 36916
rect 22612 36876 23980 36904
rect 22612 36864 22618 36876
rect 23198 36796 23204 36848
rect 23256 36836 23262 36848
rect 23952 36845 23980 36876
rect 26602 36864 26608 36916
rect 26660 36904 26666 36916
rect 27338 36904 27344 36916
rect 26660 36876 27344 36904
rect 26660 36864 26666 36876
rect 27338 36864 27344 36876
rect 27396 36864 27402 36916
rect 27822 36876 28028 36904
rect 23845 36839 23903 36845
rect 23845 36836 23857 36839
rect 23256 36808 23857 36836
rect 23256 36796 23262 36808
rect 23845 36805 23857 36808
rect 23891 36805 23903 36839
rect 23845 36799 23903 36805
rect 23937 36839 23995 36845
rect 23937 36805 23949 36839
rect 23983 36805 23995 36839
rect 23937 36799 23995 36805
rect 24075 36839 24133 36845
rect 24075 36805 24087 36839
rect 24121 36836 24133 36839
rect 24210 36836 24216 36848
rect 24121 36808 24216 36836
rect 24121 36805 24133 36808
rect 24075 36799 24133 36805
rect 24210 36796 24216 36808
rect 24268 36796 24274 36848
rect 24670 36836 24676 36848
rect 24596 36808 24676 36836
rect 22281 36771 22339 36777
rect 22281 36737 22293 36771
rect 22327 36737 22339 36771
rect 22281 36731 22339 36737
rect 22738 36728 22744 36780
rect 22796 36728 22802 36780
rect 22830 36728 22836 36780
rect 22888 36728 22894 36780
rect 22925 36771 22983 36777
rect 22925 36737 22937 36771
rect 22971 36737 22983 36771
rect 22925 36731 22983 36737
rect 21600 36672 21680 36700
rect 21600 36660 21606 36672
rect 21910 36660 21916 36712
rect 21968 36660 21974 36712
rect 22094 36660 22100 36712
rect 22152 36660 22158 36712
rect 22186 36660 22192 36712
rect 22244 36660 22250 36712
rect 22373 36703 22431 36709
rect 22373 36669 22385 36703
rect 22419 36669 22431 36703
rect 22373 36663 22431 36669
rect 21269 36635 21327 36641
rect 21269 36601 21281 36635
rect 21315 36632 21327 36635
rect 22388 36632 22416 36663
rect 22940 36632 22968 36731
rect 23474 36728 23480 36780
rect 23532 36728 23538 36780
rect 23753 36771 23811 36777
rect 23753 36737 23765 36771
rect 23799 36768 23811 36771
rect 23799 36740 23980 36768
rect 24302 36750 24308 36802
rect 24360 36750 24366 36802
rect 24489 36774 24547 36777
rect 24596 36774 24624 36808
rect 24670 36796 24676 36808
rect 24728 36796 24734 36848
rect 25590 36796 25596 36848
rect 25648 36836 25654 36848
rect 25685 36839 25743 36845
rect 25685 36836 25697 36839
rect 25648 36808 25697 36836
rect 25648 36796 25654 36808
rect 25685 36805 25697 36808
rect 25731 36805 25743 36839
rect 25685 36799 25743 36805
rect 25958 36796 25964 36848
rect 26016 36836 26022 36848
rect 27822 36836 27850 36876
rect 26016 36808 27850 36836
rect 27893 36839 27951 36845
rect 26016 36796 26022 36808
rect 27893 36805 27905 36839
rect 27939 36805 27951 36839
rect 27893 36799 27951 36805
rect 28000 36836 28028 36876
rect 28258 36864 28264 36916
rect 28316 36904 28322 36916
rect 28810 36904 28816 36916
rect 28316 36876 28816 36904
rect 28316 36864 28322 36876
rect 28810 36864 28816 36876
rect 28868 36864 28874 36916
rect 29822 36864 29828 36916
rect 29880 36904 29886 36916
rect 30926 36904 30932 36916
rect 29880 36876 30932 36904
rect 29880 36864 29886 36876
rect 30926 36864 30932 36876
rect 30984 36864 30990 36916
rect 31478 36864 31484 36916
rect 31536 36864 31542 36916
rect 31941 36907 31999 36913
rect 31588 36876 31892 36904
rect 28902 36836 28908 36848
rect 28000 36808 28908 36836
rect 24489 36771 24624 36774
rect 23799 36737 23811 36740
rect 23753 36731 23811 36737
rect 23017 36703 23075 36709
rect 23017 36669 23029 36703
rect 23063 36700 23075 36703
rect 23492 36700 23520 36728
rect 23063 36672 23520 36700
rect 23063 36669 23075 36672
rect 23017 36663 23075 36669
rect 21315 36604 22416 36632
rect 22480 36604 22968 36632
rect 23952 36632 23980 36740
rect 24210 36660 24216 36712
rect 24268 36660 24274 36712
rect 24320 36709 24348 36750
rect 24489 36737 24501 36771
rect 24535 36746 24624 36771
rect 24535 36737 24547 36746
rect 24489 36731 24547 36737
rect 24946 36728 24952 36780
rect 25004 36728 25010 36780
rect 25406 36728 25412 36780
rect 25464 36728 25470 36780
rect 25498 36728 25504 36780
rect 25556 36728 25562 36780
rect 25774 36728 25780 36780
rect 25832 36728 25838 36780
rect 25874 36771 25932 36777
rect 25874 36737 25886 36771
rect 25920 36737 25932 36771
rect 25874 36731 25932 36737
rect 24305 36703 24363 36709
rect 24305 36669 24317 36703
rect 24351 36669 24363 36703
rect 24964 36700 24992 36728
rect 25517 36700 25545 36728
rect 24964 36672 25545 36700
rect 25884 36700 25912 36731
rect 26786 36700 26792 36712
rect 25884 36672 26792 36700
rect 24305 36663 24363 36669
rect 24670 36632 24676 36644
rect 23952 36604 24676 36632
rect 21315 36601 21327 36604
rect 21269 36595 21327 36601
rect 22480 36564 22508 36604
rect 24670 36592 24676 36604
rect 24728 36592 24734 36644
rect 25222 36592 25228 36644
rect 25280 36632 25286 36644
rect 25884 36632 25912 36672
rect 26786 36660 26792 36672
rect 26844 36660 26850 36712
rect 25280 36604 25912 36632
rect 26053 36635 26111 36641
rect 25280 36592 25286 36604
rect 26053 36601 26065 36635
rect 26099 36632 26111 36635
rect 27908 36632 27936 36799
rect 28000 36768 28028 36808
rect 28902 36796 28908 36808
rect 28960 36796 28966 36848
rect 28994 36796 29000 36848
rect 29052 36836 29058 36848
rect 31205 36839 31263 36845
rect 31205 36836 31217 36839
rect 29052 36808 31217 36836
rect 29052 36796 29058 36808
rect 31205 36805 31217 36808
rect 31251 36805 31263 36839
rect 31205 36799 31263 36805
rect 28169 36771 28227 36777
rect 28169 36768 28181 36771
rect 28000 36740 28181 36768
rect 28169 36737 28181 36740
rect 28215 36737 28227 36771
rect 28169 36731 28227 36737
rect 28442 36728 28448 36780
rect 28500 36768 28506 36780
rect 28500 36740 28764 36768
rect 28500 36728 28506 36740
rect 27982 36660 27988 36712
rect 28040 36660 28046 36712
rect 28736 36700 28764 36740
rect 28810 36728 28816 36780
rect 28868 36728 28874 36780
rect 30926 36728 30932 36780
rect 30984 36768 30990 36780
rect 31496 36777 31524 36864
rect 31588 36848 31616 36876
rect 31570 36796 31576 36848
rect 31628 36796 31634 36848
rect 31662 36796 31668 36848
rect 31720 36836 31726 36848
rect 31864 36836 31892 36876
rect 31941 36873 31953 36907
rect 31987 36904 31999 36907
rect 32214 36904 32220 36916
rect 31987 36876 32220 36904
rect 31987 36873 31999 36876
rect 31941 36867 31999 36873
rect 32214 36864 32220 36876
rect 32272 36864 32278 36916
rect 32398 36864 32404 36916
rect 32456 36904 32462 36916
rect 32493 36907 32551 36913
rect 32493 36904 32505 36907
rect 32456 36876 32505 36904
rect 32456 36864 32462 36876
rect 32493 36873 32505 36876
rect 32539 36873 32551 36907
rect 32493 36867 32551 36873
rect 32582 36864 32588 36916
rect 32640 36864 32646 36916
rect 33410 36864 33416 36916
rect 33468 36904 33474 36916
rect 33468 36876 34100 36904
rect 33468 36864 33474 36876
rect 32030 36836 32036 36848
rect 31720 36808 31800 36836
rect 31864 36808 32036 36836
rect 31720 36796 31726 36808
rect 31772 36777 31800 36808
rect 32030 36796 32036 36808
rect 32088 36836 32094 36848
rect 32088 36808 32260 36836
rect 32088 36796 32094 36808
rect 32232 36777 32260 36808
rect 31021 36771 31079 36777
rect 31021 36768 31033 36771
rect 30984 36740 31033 36768
rect 30984 36728 30990 36740
rect 31021 36737 31033 36740
rect 31067 36737 31079 36771
rect 31021 36731 31079 36737
rect 31481 36771 31539 36777
rect 31481 36737 31493 36771
rect 31527 36737 31539 36771
rect 31481 36731 31539 36737
rect 31757 36771 31815 36777
rect 31757 36737 31769 36771
rect 31803 36737 31815 36771
rect 31757 36731 31815 36737
rect 32125 36771 32183 36777
rect 32125 36737 32137 36771
rect 32171 36737 32183 36771
rect 32125 36731 32183 36737
rect 32217 36771 32275 36777
rect 32217 36737 32229 36771
rect 32263 36737 32275 36771
rect 32600 36768 32628 36864
rect 34072 36845 34100 36876
rect 34057 36839 34115 36845
rect 34057 36805 34069 36839
rect 34103 36805 34115 36839
rect 34057 36799 34115 36805
rect 34606 36796 34612 36848
rect 34664 36796 34670 36848
rect 33229 36771 33287 36777
rect 33229 36768 33241 36771
rect 32600 36740 33241 36768
rect 32217 36731 32275 36737
rect 33229 36737 33241 36740
rect 33275 36737 33287 36771
rect 33229 36731 33287 36737
rect 28902 36700 28908 36712
rect 28736 36672 28908 36700
rect 28902 36660 28908 36672
rect 28960 36660 28966 36712
rect 31036 36700 31064 36731
rect 31573 36703 31631 36709
rect 31573 36700 31585 36703
rect 31036 36672 31585 36700
rect 31573 36669 31585 36672
rect 31619 36669 31631 36703
rect 31573 36663 31631 36669
rect 26099 36604 28856 36632
rect 26099 36601 26111 36604
rect 26053 36595 26111 36601
rect 20220 36536 22508 36564
rect 20220 36524 20226 36536
rect 22554 36524 22560 36576
rect 22612 36524 22618 36576
rect 23569 36567 23627 36573
rect 23569 36533 23581 36567
rect 23615 36564 23627 36567
rect 25958 36564 25964 36576
rect 23615 36536 25964 36564
rect 23615 36533 23627 36536
rect 23569 36527 23627 36533
rect 25958 36524 25964 36536
rect 26016 36524 26022 36576
rect 28169 36567 28227 36573
rect 28169 36533 28181 36567
rect 28215 36564 28227 36567
rect 28258 36564 28264 36576
rect 28215 36536 28264 36564
rect 28215 36533 28227 36536
rect 28169 36527 28227 36533
rect 28258 36524 28264 36536
rect 28316 36524 28322 36576
rect 28350 36524 28356 36576
rect 28408 36524 28414 36576
rect 28828 36573 28856 36604
rect 31386 36592 31392 36644
rect 31444 36632 31450 36644
rect 32140 36632 32168 36731
rect 33594 36728 33600 36780
rect 33652 36768 33658 36780
rect 33781 36771 33839 36777
rect 33781 36768 33793 36771
rect 33652 36740 33793 36768
rect 33652 36728 33658 36740
rect 33781 36737 33793 36740
rect 33827 36737 33839 36771
rect 33781 36731 33839 36737
rect 31444 36604 32168 36632
rect 31444 36592 31450 36604
rect 28813 36567 28871 36573
rect 28813 36533 28825 36567
rect 28859 36533 28871 36567
rect 28813 36527 28871 36533
rect 29181 36567 29239 36573
rect 29181 36533 29193 36567
rect 29227 36564 29239 36567
rect 31478 36564 31484 36576
rect 29227 36536 31484 36564
rect 29227 36533 29239 36536
rect 29181 36527 29239 36533
rect 31478 36524 31484 36536
rect 31536 36524 31542 36576
rect 31938 36524 31944 36576
rect 31996 36564 32002 36576
rect 32125 36567 32183 36573
rect 32125 36564 32137 36567
rect 31996 36536 32137 36564
rect 31996 36524 32002 36536
rect 32125 36533 32137 36536
rect 32171 36533 32183 36567
rect 32125 36527 32183 36533
rect 33045 36567 33103 36573
rect 33045 36533 33057 36567
rect 33091 36564 33103 36567
rect 33226 36564 33232 36576
rect 33091 36536 33232 36564
rect 33091 36533 33103 36536
rect 33045 36527 33103 36533
rect 33226 36524 33232 36536
rect 33284 36524 33290 36576
rect 35526 36524 35532 36576
rect 35584 36524 35590 36576
rect 1104 36474 41400 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 41400 36474
rect 1104 36400 41400 36422
rect 6720 36363 6778 36369
rect 6720 36329 6732 36363
rect 6766 36360 6778 36363
rect 12066 36360 12072 36372
rect 6766 36332 12072 36360
rect 6766 36329 6778 36332
rect 6720 36323 6778 36329
rect 12066 36320 12072 36332
rect 12124 36320 12130 36372
rect 16301 36363 16359 36369
rect 16301 36329 16313 36363
rect 16347 36329 16359 36363
rect 16301 36323 16359 36329
rect 12710 36252 12716 36304
rect 12768 36292 12774 36304
rect 16316 36292 16344 36323
rect 16482 36320 16488 36372
rect 16540 36320 16546 36372
rect 16942 36360 16948 36372
rect 16592 36332 16948 36360
rect 16592 36292 16620 36332
rect 16942 36320 16948 36332
rect 17000 36360 17006 36372
rect 19150 36360 19156 36372
rect 17000 36332 19156 36360
rect 17000 36320 17006 36332
rect 19150 36320 19156 36332
rect 19208 36320 19214 36372
rect 19260 36332 19380 36360
rect 12768 36264 16252 36292
rect 16316 36264 16620 36292
rect 17696 36264 18552 36292
rect 12768 36252 12774 36264
rect 6822 36224 6828 36236
rect 6472 36196 6828 36224
rect 5994 36116 6000 36168
rect 6052 36156 6058 36168
rect 6472 36165 6500 36196
rect 6822 36184 6828 36196
rect 6880 36184 6886 36236
rect 11422 36184 11428 36236
rect 11480 36184 11486 36236
rect 16224 36224 16252 36264
rect 17586 36224 17592 36236
rect 16224 36196 17592 36224
rect 17586 36184 17592 36196
rect 17644 36184 17650 36236
rect 6457 36159 6515 36165
rect 6457 36156 6469 36159
rect 6052 36128 6469 36156
rect 6052 36116 6058 36128
rect 6457 36125 6469 36128
rect 6503 36125 6515 36159
rect 8754 36156 8760 36168
rect 6457 36119 6515 36125
rect 8128 36128 8760 36156
rect 1489 36091 1547 36097
rect 1489 36057 1501 36091
rect 1535 36088 1547 36091
rect 4798 36088 4804 36100
rect 1535 36060 4804 36088
rect 1535 36057 1547 36060
rect 1489 36051 1547 36057
rect 4798 36048 4804 36060
rect 4856 36048 4862 36100
rect 7116 36060 7222 36088
rect 7116 36032 7144 36060
rect 934 35980 940 36032
rect 992 36020 998 36032
rect 1581 36023 1639 36029
rect 1581 36020 1593 36023
rect 992 35992 1593 36020
rect 992 35980 998 35992
rect 1581 35989 1593 35992
rect 1627 35989 1639 36023
rect 1581 35983 1639 35989
rect 7098 35980 7104 36032
rect 7156 36020 7162 36032
rect 8128 36020 8156 36128
rect 8754 36116 8760 36128
rect 8812 36116 8818 36168
rect 9306 36116 9312 36168
rect 9364 36156 9370 36168
rect 10042 36156 10048 36168
rect 9364 36128 10048 36156
rect 9364 36116 9370 36128
rect 10042 36116 10048 36128
rect 10100 36116 10106 36168
rect 11701 36159 11759 36165
rect 11701 36125 11713 36159
rect 11747 36156 11759 36159
rect 15838 36156 15844 36168
rect 11747 36128 15844 36156
rect 11747 36125 11759 36128
rect 11701 36119 11759 36125
rect 15838 36116 15844 36128
rect 15896 36156 15902 36168
rect 17696 36156 17724 36264
rect 17957 36227 18015 36233
rect 17957 36193 17969 36227
rect 18003 36224 18015 36227
rect 18138 36224 18144 36236
rect 18003 36196 18144 36224
rect 18003 36193 18015 36196
rect 17957 36187 18015 36193
rect 18138 36184 18144 36196
rect 18196 36224 18202 36236
rect 18414 36224 18420 36236
rect 18196 36196 18420 36224
rect 18196 36184 18202 36196
rect 18414 36184 18420 36196
rect 18472 36184 18478 36236
rect 18524 36224 18552 36264
rect 18874 36252 18880 36304
rect 18932 36292 18938 36304
rect 19260 36292 19288 36332
rect 18932 36264 19288 36292
rect 18932 36252 18938 36264
rect 19242 36224 19248 36236
rect 18524 36196 19248 36224
rect 19242 36184 19248 36196
rect 19300 36184 19306 36236
rect 19352 36224 19380 36332
rect 19426 36320 19432 36372
rect 19484 36360 19490 36372
rect 19886 36360 19892 36372
rect 19484 36332 19892 36360
rect 19484 36320 19490 36332
rect 19886 36320 19892 36332
rect 19944 36320 19950 36372
rect 20162 36320 20168 36372
rect 20220 36320 20226 36372
rect 20438 36360 20444 36372
rect 20272 36332 20444 36360
rect 19981 36295 20039 36301
rect 19981 36261 19993 36295
rect 20027 36292 20039 36295
rect 20272 36292 20300 36332
rect 20438 36320 20444 36332
rect 20496 36320 20502 36372
rect 20622 36320 20628 36372
rect 20680 36320 20686 36372
rect 22186 36320 22192 36372
rect 22244 36360 22250 36372
rect 22244 36332 23336 36360
rect 22244 36320 22250 36332
rect 23308 36304 23336 36332
rect 24394 36320 24400 36372
rect 24452 36360 24458 36372
rect 24857 36363 24915 36369
rect 24857 36360 24869 36363
rect 24452 36332 24869 36360
rect 24452 36320 24458 36332
rect 24857 36329 24869 36332
rect 24903 36329 24915 36363
rect 24857 36323 24915 36329
rect 25038 36320 25044 36372
rect 25096 36320 25102 36372
rect 25406 36320 25412 36372
rect 25464 36360 25470 36372
rect 26694 36360 26700 36372
rect 25464 36332 26700 36360
rect 25464 36320 25470 36332
rect 26694 36320 26700 36332
rect 26752 36320 26758 36372
rect 26896 36332 27109 36360
rect 20027 36264 20300 36292
rect 20027 36261 20039 36264
rect 19981 36255 20039 36261
rect 20346 36252 20352 36304
rect 20404 36292 20410 36304
rect 22922 36292 22928 36304
rect 20404 36264 22928 36292
rect 20404 36252 20410 36264
rect 22922 36252 22928 36264
rect 22980 36252 22986 36304
rect 23290 36252 23296 36304
rect 23348 36252 23354 36304
rect 23658 36252 23664 36304
rect 23716 36252 23722 36304
rect 20257 36227 20315 36233
rect 20257 36224 20269 36227
rect 19352 36196 20269 36224
rect 20257 36193 20269 36196
rect 20303 36193 20315 36227
rect 21085 36227 21143 36233
rect 21085 36224 21097 36227
rect 20257 36187 20315 36193
rect 20364 36196 21097 36224
rect 15896 36128 17724 36156
rect 15896 36116 15902 36128
rect 17770 36116 17776 36168
rect 17828 36156 17834 36168
rect 19426 36156 19432 36168
rect 17828 36128 19432 36156
rect 17828 36116 17834 36128
rect 19426 36116 19432 36128
rect 19484 36116 19490 36168
rect 19797 36159 19855 36165
rect 19797 36125 19809 36159
rect 19843 36156 19855 36159
rect 20364 36156 20392 36196
rect 21085 36193 21097 36196
rect 21131 36193 21143 36227
rect 23676 36224 23704 36252
rect 21085 36187 21143 36193
rect 23584 36196 23704 36224
rect 23584 36168 23612 36196
rect 23842 36184 23848 36236
rect 23900 36184 23906 36236
rect 24854 36184 24860 36236
rect 24912 36184 24918 36236
rect 25056 36224 25084 36320
rect 26896 36292 26924 36332
rect 25884 36264 26924 36292
rect 25056 36196 25544 36224
rect 19843 36128 20392 36156
rect 19843 36125 19855 36128
rect 19797 36119 19855 36125
rect 20438 36116 20444 36168
rect 20496 36116 20502 36168
rect 20530 36116 20536 36168
rect 20588 36116 20594 36168
rect 20806 36116 20812 36168
rect 20864 36156 20870 36168
rect 20901 36159 20959 36165
rect 20901 36156 20913 36159
rect 20864 36128 20913 36156
rect 20864 36116 20870 36128
rect 20901 36125 20913 36128
rect 20947 36125 20959 36159
rect 20901 36119 20959 36125
rect 22186 36116 22192 36168
rect 22244 36156 22250 36168
rect 22281 36159 22339 36165
rect 22281 36156 22293 36159
rect 22244 36128 22293 36156
rect 22244 36116 22250 36128
rect 22281 36125 22293 36128
rect 22327 36125 22339 36159
rect 22281 36119 22339 36125
rect 22465 36159 22523 36165
rect 22465 36125 22477 36159
rect 22511 36156 22523 36159
rect 22554 36156 22560 36168
rect 22511 36128 22560 36156
rect 22511 36125 22523 36128
rect 22465 36119 22523 36125
rect 22554 36116 22560 36128
rect 22612 36116 22618 36168
rect 22646 36116 22652 36168
rect 22704 36116 22710 36168
rect 22738 36116 22744 36168
rect 22796 36116 22802 36168
rect 23566 36116 23572 36168
rect 23624 36116 23630 36168
rect 23658 36116 23664 36168
rect 23716 36156 23722 36168
rect 23860 36156 23888 36184
rect 23716 36128 23888 36156
rect 23716 36116 23722 36128
rect 23934 36116 23940 36168
rect 23992 36116 23998 36168
rect 24075 36159 24133 36165
rect 24075 36125 24087 36159
rect 24121 36156 24133 36159
rect 24670 36156 24676 36168
rect 24121 36128 24676 36156
rect 24121 36125 24133 36128
rect 24075 36119 24133 36125
rect 24670 36116 24676 36128
rect 24728 36116 24734 36168
rect 24872 36156 24900 36184
rect 25406 36165 25412 36168
rect 25041 36159 25099 36165
rect 25041 36156 25053 36159
rect 24872 36128 25053 36156
rect 25041 36125 25053 36128
rect 25087 36125 25099 36159
rect 25041 36119 25099 36125
rect 25363 36159 25412 36165
rect 25363 36125 25375 36159
rect 25409 36125 25412 36159
rect 25363 36119 25412 36125
rect 25406 36116 25412 36119
rect 25464 36116 25470 36168
rect 25516 36165 25544 36196
rect 25501 36159 25559 36165
rect 25501 36125 25513 36159
rect 25547 36125 25559 36159
rect 25501 36119 25559 36125
rect 25590 36116 25596 36168
rect 25648 36116 25654 36168
rect 8846 36088 8852 36100
rect 8220 36060 8852 36088
rect 8220 36029 8248 36060
rect 8846 36048 8852 36060
rect 8904 36088 8910 36100
rect 9033 36091 9091 36097
rect 9033 36088 9045 36091
rect 8904 36060 9045 36088
rect 8904 36048 8910 36060
rect 9033 36057 9045 36060
rect 9079 36088 9091 36091
rect 10502 36088 10508 36100
rect 9079 36060 10508 36088
rect 9079 36057 9091 36060
rect 9033 36051 9091 36057
rect 10502 36048 10508 36060
rect 10560 36048 10566 36100
rect 10686 36048 10692 36100
rect 10744 36048 10750 36100
rect 11330 36048 11336 36100
rect 11388 36088 11394 36100
rect 11977 36091 12035 36097
rect 11977 36088 11989 36091
rect 11388 36060 11989 36088
rect 11388 36048 11394 36060
rect 11977 36057 11989 36060
rect 12023 36088 12035 36091
rect 12250 36088 12256 36100
rect 12023 36060 12256 36088
rect 12023 36057 12035 36060
rect 11977 36051 12035 36057
rect 12250 36048 12256 36060
rect 12308 36048 12314 36100
rect 12342 36048 12348 36100
rect 12400 36088 12406 36100
rect 14182 36088 14188 36100
rect 12400 36060 14188 36088
rect 12400 36048 12406 36060
rect 14182 36048 14188 36060
rect 14240 36048 14246 36100
rect 15010 36048 15016 36100
rect 15068 36048 15074 36100
rect 16117 36091 16175 36097
rect 16117 36057 16129 36091
rect 16163 36088 16175 36091
rect 16666 36088 16672 36100
rect 16163 36060 16672 36088
rect 16163 36057 16175 36060
rect 16117 36051 16175 36057
rect 16666 36048 16672 36060
rect 16724 36048 16730 36100
rect 17681 36091 17739 36097
rect 17681 36057 17693 36091
rect 17727 36088 17739 36091
rect 17954 36088 17960 36100
rect 17727 36060 17960 36088
rect 17727 36057 17739 36060
rect 17681 36051 17739 36057
rect 17954 36048 17960 36060
rect 18012 36088 18018 36100
rect 19058 36088 19064 36100
rect 18012 36060 19064 36088
rect 18012 36048 18018 36060
rect 19058 36048 19064 36060
rect 19116 36048 19122 36100
rect 19242 36048 19248 36100
rect 19300 36048 19306 36100
rect 20165 36091 20223 36097
rect 20165 36057 20177 36091
rect 20211 36088 20223 36091
rect 20548 36088 20576 36116
rect 20211 36060 20576 36088
rect 20211 36057 20223 36060
rect 20165 36051 20223 36057
rect 20622 36048 20628 36100
rect 20680 36088 20686 36100
rect 20717 36091 20775 36097
rect 20717 36088 20729 36091
rect 20680 36060 20729 36088
rect 20680 36048 20686 36060
rect 20717 36057 20729 36060
rect 20763 36057 20775 36091
rect 20717 36051 20775 36057
rect 23842 36048 23848 36100
rect 23900 36048 23906 36100
rect 24946 36088 24952 36100
rect 24136 36060 24952 36088
rect 7156 35992 8156 36020
rect 8205 36023 8263 36029
rect 7156 35980 7162 35992
rect 8205 35989 8217 36023
rect 8251 35989 8263 36023
rect 8205 35983 8263 35989
rect 9122 35980 9128 36032
rect 9180 36020 9186 36032
rect 11790 36020 11796 36032
rect 9180 35992 11796 36020
rect 9180 35980 9186 35992
rect 11790 35980 11796 35992
rect 11848 36020 11854 36032
rect 12802 36020 12808 36032
rect 11848 35992 12808 36020
rect 11848 35980 11854 35992
rect 12802 35980 12808 35992
rect 12860 35980 12866 36032
rect 15028 36020 15056 36048
rect 16317 36023 16375 36029
rect 16317 36020 16329 36023
rect 15028 35992 16329 36020
rect 16317 35989 16329 35992
rect 16363 35989 16375 36023
rect 16317 35983 16375 35989
rect 18690 35980 18696 36032
rect 18748 36020 18754 36032
rect 19429 36023 19487 36029
rect 19429 36020 19441 36023
rect 18748 35992 19441 36020
rect 18748 35980 18754 35992
rect 19429 35989 19441 35992
rect 19475 35989 19487 36023
rect 19429 35983 19487 35989
rect 19613 36023 19671 36029
rect 19613 35989 19625 36023
rect 19659 36020 19671 36023
rect 24136 36020 24164 36060
rect 24946 36048 24952 36060
rect 25004 36048 25010 36100
rect 25130 36048 25136 36100
rect 25188 36048 25194 36100
rect 25222 36048 25228 36100
rect 25280 36048 25286 36100
rect 25608 36088 25636 36116
rect 25884 36088 25912 36264
rect 26970 36252 26976 36304
rect 27028 36252 27034 36304
rect 26694 36224 26700 36236
rect 26124 36196 26700 36224
rect 25958 36116 25964 36168
rect 26016 36116 26022 36168
rect 26124 36165 26152 36196
rect 26694 36184 26700 36196
rect 26752 36184 26758 36236
rect 26109 36159 26167 36165
rect 26109 36125 26121 36159
rect 26155 36125 26167 36159
rect 26109 36119 26167 36125
rect 26467 36159 26525 36165
rect 26467 36125 26479 36159
rect 26513 36156 26525 36159
rect 26786 36156 26792 36168
rect 26513 36128 26792 36156
rect 26513 36125 26525 36128
rect 26467 36119 26525 36125
rect 26786 36116 26792 36128
rect 26844 36116 26850 36168
rect 26988 36156 27016 36252
rect 27081 36224 27109 36332
rect 27614 36320 27620 36372
rect 27672 36360 27678 36372
rect 28077 36363 28135 36369
rect 28077 36360 28089 36363
rect 27672 36332 28089 36360
rect 27672 36320 27678 36332
rect 28077 36329 28089 36332
rect 28123 36329 28135 36363
rect 28077 36323 28135 36329
rect 28718 36320 28724 36372
rect 28776 36360 28782 36372
rect 29362 36360 29368 36372
rect 28776 36332 29368 36360
rect 28776 36320 28782 36332
rect 29362 36320 29368 36332
rect 29420 36320 29426 36372
rect 31202 36320 31208 36372
rect 31260 36320 31266 36372
rect 32122 36320 32128 36372
rect 32180 36320 32186 36372
rect 27157 36295 27215 36301
rect 27157 36261 27169 36295
rect 27203 36292 27215 36295
rect 27890 36292 27896 36304
rect 27203 36264 27896 36292
rect 27203 36261 27215 36264
rect 27157 36255 27215 36261
rect 27890 36252 27896 36264
rect 27948 36252 27954 36304
rect 28350 36292 28356 36304
rect 28000 36264 28356 36292
rect 27081 36196 27476 36224
rect 27448 36165 27476 36196
rect 27632 36196 27936 36224
rect 27632 36165 27660 36196
rect 27908 36168 27936 36196
rect 27341 36159 27399 36165
rect 27341 36156 27353 36159
rect 26988 36128 27353 36156
rect 27341 36125 27353 36128
rect 27387 36125 27399 36159
rect 27341 36119 27399 36125
rect 27433 36159 27491 36165
rect 27433 36125 27445 36159
rect 27479 36125 27491 36159
rect 27433 36119 27491 36125
rect 27617 36159 27675 36165
rect 27617 36125 27629 36159
rect 27663 36125 27675 36159
rect 27617 36119 27675 36125
rect 27706 36116 27712 36168
rect 27764 36116 27770 36168
rect 27890 36116 27896 36168
rect 27948 36116 27954 36168
rect 28000 36156 28028 36264
rect 28350 36252 28356 36264
rect 28408 36252 28414 36304
rect 28442 36252 28448 36304
rect 28500 36292 28506 36304
rect 31938 36292 31944 36304
rect 28500 36264 31944 36292
rect 28500 36252 28506 36264
rect 31938 36252 31944 36264
rect 31996 36252 32002 36304
rect 28261 36227 28319 36233
rect 28261 36193 28273 36227
rect 28307 36224 28319 36227
rect 28718 36224 28724 36236
rect 28307 36196 28724 36224
rect 28307 36193 28319 36196
rect 28261 36187 28319 36193
rect 28644 36165 28672 36196
rect 28718 36184 28724 36196
rect 28776 36184 28782 36236
rect 28997 36227 29055 36233
rect 28997 36193 29009 36227
rect 29043 36224 29055 36227
rect 31294 36224 31300 36236
rect 29043 36196 31300 36224
rect 29043 36193 29055 36196
rect 28997 36187 29055 36193
rect 31294 36184 31300 36196
rect 31352 36184 31358 36236
rect 31386 36184 31392 36236
rect 31444 36184 31450 36236
rect 28077 36159 28135 36165
rect 28077 36156 28089 36159
rect 28000 36128 28089 36156
rect 28077 36125 28089 36128
rect 28123 36125 28135 36159
rect 28077 36119 28135 36125
rect 28353 36159 28411 36165
rect 28353 36125 28365 36159
rect 28399 36125 28411 36159
rect 28353 36119 28411 36125
rect 28629 36159 28687 36165
rect 28629 36125 28641 36159
rect 28675 36156 28687 36159
rect 31312 36156 31340 36184
rect 31481 36159 31539 36165
rect 31481 36156 31493 36159
rect 28675 36128 28709 36156
rect 31312 36128 31493 36156
rect 28675 36125 28687 36128
rect 28629 36119 28687 36125
rect 31481 36125 31493 36128
rect 31527 36125 31539 36159
rect 31481 36119 31539 36125
rect 26237 36091 26295 36097
rect 26237 36088 26249 36091
rect 25608 36060 26249 36088
rect 26237 36057 26249 36060
rect 26283 36057 26295 36091
rect 26237 36051 26295 36057
rect 26329 36091 26387 36097
rect 26329 36057 26341 36091
rect 26375 36088 26387 36091
rect 26970 36088 26976 36100
rect 26375 36060 26976 36088
rect 26375 36057 26387 36060
rect 26329 36051 26387 36057
rect 26970 36048 26976 36060
rect 27028 36048 27034 36100
rect 19659 35992 24164 36020
rect 24213 36023 24271 36029
rect 19659 35989 19671 35992
rect 19613 35983 19671 35989
rect 24213 35989 24225 36023
rect 24259 36020 24271 36023
rect 26142 36020 26148 36032
rect 24259 35992 26148 36020
rect 24259 35989 24271 35992
rect 24213 35983 24271 35989
rect 26142 35980 26148 35992
rect 26200 35980 26206 36032
rect 26605 36023 26663 36029
rect 26605 35989 26617 36023
rect 26651 36020 26663 36023
rect 27246 36020 27252 36032
rect 26651 35992 27252 36020
rect 26651 35989 26663 35992
rect 26605 35983 26663 35989
rect 27246 35980 27252 35992
rect 27304 36020 27310 36032
rect 28368 36020 28396 36119
rect 28718 36048 28724 36100
rect 28776 36088 28782 36100
rect 28813 36091 28871 36097
rect 28813 36088 28825 36091
rect 28776 36060 28825 36088
rect 28776 36048 28782 36060
rect 28813 36057 28825 36060
rect 28859 36057 28871 36091
rect 28813 36051 28871 36057
rect 29914 36048 29920 36100
rect 29972 36088 29978 36100
rect 31205 36091 31263 36097
rect 31205 36088 31217 36091
rect 29972 36060 31217 36088
rect 29972 36048 29978 36060
rect 31205 36057 31217 36060
rect 31251 36057 31263 36091
rect 32140 36088 32168 36320
rect 33594 36184 33600 36236
rect 33652 36224 33658 36236
rect 34241 36227 34299 36233
rect 34241 36224 34253 36227
rect 33652 36196 34253 36224
rect 33652 36184 33658 36196
rect 34241 36193 34253 36196
rect 34287 36193 34299 36227
rect 34241 36187 34299 36193
rect 31205 36051 31263 36057
rect 31312 36060 32168 36088
rect 33505 36091 33563 36097
rect 27304 35992 28396 36020
rect 28537 36023 28595 36029
rect 27304 35980 27310 35992
rect 28537 35989 28549 36023
rect 28583 36020 28595 36023
rect 31312 36020 31340 36060
rect 33505 36057 33517 36091
rect 33551 36088 33563 36091
rect 37274 36088 37280 36100
rect 33551 36060 37280 36088
rect 33551 36057 33563 36060
rect 33505 36051 33563 36057
rect 37274 36048 37280 36060
rect 37332 36048 37338 36100
rect 28583 35992 31340 36020
rect 31665 36023 31723 36029
rect 28583 35989 28595 35992
rect 28537 35983 28595 35989
rect 31665 35989 31677 36023
rect 31711 36020 31723 36023
rect 32490 36020 32496 36032
rect 31711 35992 32496 36020
rect 31711 35989 31723 35992
rect 31665 35983 31723 35989
rect 32490 35980 32496 35992
rect 32548 35980 32554 36032
rect 1104 35930 41400 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 41400 35930
rect 1104 35856 41400 35878
rect 9033 35819 9091 35825
rect 9033 35785 9045 35819
rect 9079 35785 9091 35819
rect 9033 35779 9091 35785
rect 7098 35708 7104 35760
rect 7156 35708 7162 35760
rect 8938 35640 8944 35692
rect 8996 35640 9002 35692
rect 9048 35680 9076 35779
rect 9490 35776 9496 35828
rect 9548 35816 9554 35828
rect 10226 35816 10232 35828
rect 9548 35788 9720 35816
rect 9548 35776 9554 35788
rect 9692 35757 9720 35788
rect 10157 35788 10232 35816
rect 9309 35751 9367 35757
rect 9309 35717 9321 35751
rect 9355 35748 9367 35751
rect 9666 35751 9724 35757
rect 9666 35748 9678 35751
rect 9355 35720 9678 35748
rect 9355 35717 9367 35720
rect 9309 35711 9367 35717
rect 9666 35717 9678 35720
rect 9712 35717 9724 35751
rect 9666 35711 9724 35717
rect 9493 35683 9551 35689
rect 9048 35652 9444 35680
rect 5994 35572 6000 35624
rect 6052 35612 6058 35624
rect 6365 35615 6423 35621
rect 6365 35612 6377 35615
rect 6052 35584 6377 35612
rect 6052 35572 6058 35584
rect 6365 35581 6377 35584
rect 6411 35581 6423 35615
rect 6365 35575 6423 35581
rect 6730 35572 6736 35624
rect 6788 35572 6794 35624
rect 9030 35572 9036 35624
rect 9088 35612 9094 35624
rect 9125 35615 9183 35621
rect 9125 35612 9137 35615
rect 9088 35584 9137 35612
rect 9088 35572 9094 35584
rect 9125 35581 9137 35584
rect 9171 35581 9183 35615
rect 9416 35612 9444 35652
rect 9493 35649 9505 35683
rect 9539 35680 9551 35683
rect 10157 35680 10185 35788
rect 10226 35776 10232 35788
rect 10284 35776 10290 35828
rect 10965 35819 11023 35825
rect 10965 35785 10977 35819
rect 11011 35785 11023 35819
rect 10965 35779 11023 35785
rect 10980 35748 11008 35779
rect 12342 35776 12348 35828
rect 12400 35776 12406 35828
rect 13081 35819 13139 35825
rect 13081 35785 13093 35819
rect 13127 35816 13139 35819
rect 13998 35816 14004 35828
rect 13127 35788 14004 35816
rect 13127 35785 13139 35788
rect 13081 35779 13139 35785
rect 13998 35776 14004 35788
rect 14056 35776 14062 35828
rect 15194 35776 15200 35828
rect 15252 35816 15258 35828
rect 22738 35816 22744 35828
rect 15252 35788 22744 35816
rect 15252 35776 15258 35788
rect 22738 35776 22744 35788
rect 22796 35776 22802 35828
rect 23014 35776 23020 35828
rect 23072 35776 23078 35828
rect 23566 35776 23572 35828
rect 23624 35816 23630 35828
rect 24305 35819 24363 35825
rect 24305 35816 24317 35819
rect 23624 35788 24317 35816
rect 23624 35776 23630 35788
rect 24305 35785 24317 35788
rect 24351 35785 24363 35819
rect 24305 35779 24363 35785
rect 24412 35788 25636 35816
rect 12360 35748 12388 35776
rect 10244 35720 11008 35748
rect 11992 35720 12388 35748
rect 10244 35689 10272 35720
rect 9539 35652 10185 35680
rect 10229 35683 10287 35689
rect 9539 35649 9551 35652
rect 9493 35643 9551 35649
rect 10229 35649 10241 35683
rect 10275 35649 10287 35683
rect 10229 35643 10287 35649
rect 10689 35683 10747 35689
rect 10689 35649 10701 35683
rect 10735 35649 10747 35683
rect 10689 35643 10747 35649
rect 10134 35612 10140 35624
rect 9416 35584 10140 35612
rect 9125 35575 9183 35581
rect 10134 35572 10140 35584
rect 10192 35572 10198 35624
rect 10704 35612 10732 35643
rect 10778 35640 10784 35692
rect 10836 35680 10842 35692
rect 11992 35689 12020 35720
rect 12802 35708 12808 35760
rect 12860 35711 12866 35760
rect 12860 35708 12873 35711
rect 12986 35708 12992 35760
rect 13044 35748 13050 35760
rect 21542 35748 21548 35760
rect 13044 35720 21548 35748
rect 13044 35708 13050 35720
rect 21542 35708 21548 35720
rect 21600 35708 21606 35760
rect 23032 35748 23060 35776
rect 22204 35720 23060 35748
rect 23477 35751 23535 35757
rect 12815 35705 12873 35708
rect 11977 35683 12035 35689
rect 11977 35680 11989 35683
rect 10836 35652 11989 35680
rect 10836 35640 10842 35652
rect 11977 35649 11989 35652
rect 12023 35649 12035 35683
rect 12815 35671 12827 35705
rect 12861 35671 12873 35705
rect 12815 35665 12873 35671
rect 19705 35683 19763 35689
rect 11977 35643 12035 35649
rect 19705 35649 19717 35683
rect 19751 35680 19763 35683
rect 19886 35680 19892 35692
rect 19751 35652 19892 35680
rect 19751 35649 19763 35652
rect 19705 35643 19763 35649
rect 19886 35640 19892 35652
rect 19944 35640 19950 35692
rect 21266 35640 21272 35692
rect 21324 35680 21330 35692
rect 21726 35680 21732 35692
rect 21324 35652 21732 35680
rect 21324 35640 21330 35652
rect 21726 35640 21732 35652
rect 21784 35680 21790 35692
rect 22204 35680 22232 35720
rect 23477 35717 23489 35751
rect 23523 35748 23535 35751
rect 23934 35748 23940 35760
rect 23523 35720 23940 35748
rect 23523 35717 23535 35720
rect 23477 35711 23535 35717
rect 23934 35708 23940 35720
rect 23992 35708 23998 35760
rect 21784 35652 22232 35680
rect 21784 35640 21790 35652
rect 22278 35640 22284 35692
rect 22336 35680 22342 35692
rect 22649 35683 22707 35689
rect 22649 35680 22661 35683
rect 22336 35652 22661 35680
rect 22336 35640 22342 35652
rect 22649 35649 22661 35652
rect 22695 35649 22707 35683
rect 22649 35643 22707 35649
rect 22922 35640 22928 35692
rect 22980 35680 22986 35692
rect 23109 35683 23167 35689
rect 23109 35680 23121 35683
rect 22980 35652 23121 35680
rect 22980 35640 22986 35652
rect 23109 35649 23121 35652
rect 23155 35649 23167 35683
rect 23109 35643 23167 35649
rect 23201 35683 23259 35689
rect 23201 35649 23213 35683
rect 23247 35649 23259 35683
rect 23201 35643 23259 35649
rect 11793 35615 11851 35621
rect 11793 35612 11805 35615
rect 10704 35584 11805 35612
rect 8018 35504 8024 35556
rect 8076 35544 8082 35556
rect 8159 35547 8217 35553
rect 8159 35544 8171 35547
rect 8076 35516 8171 35544
rect 8076 35504 8082 35516
rect 8159 35513 8171 35516
rect 8205 35544 8217 35547
rect 10704 35544 10732 35584
rect 11793 35581 11805 35584
rect 11839 35581 11851 35615
rect 11793 35575 11851 35581
rect 13081 35615 13139 35621
rect 13081 35581 13093 35615
rect 13127 35581 13139 35615
rect 13081 35575 13139 35581
rect 8205 35516 10732 35544
rect 8205 35513 8217 35516
rect 8159 35507 8217 35513
rect 10870 35504 10876 35556
rect 10928 35544 10934 35556
rect 11698 35544 11704 35556
rect 10928 35516 11704 35544
rect 10928 35504 10934 35516
rect 11698 35504 11704 35516
rect 11756 35504 11762 35556
rect 11882 35504 11888 35556
rect 11940 35544 11946 35556
rect 12897 35547 12955 35553
rect 12897 35544 12909 35547
rect 11940 35516 12909 35544
rect 11940 35504 11946 35516
rect 12897 35513 12909 35516
rect 12943 35544 12955 35547
rect 12986 35544 12992 35556
rect 12943 35516 12992 35544
rect 12943 35513 12955 35516
rect 12897 35507 12955 35513
rect 12986 35504 12992 35516
rect 13044 35504 13050 35556
rect 9217 35479 9275 35485
rect 9217 35445 9229 35479
rect 9263 35476 9275 35479
rect 9306 35476 9312 35488
rect 9263 35448 9312 35476
rect 9263 35445 9275 35448
rect 9217 35439 9275 35445
rect 9306 35436 9312 35448
rect 9364 35436 9370 35488
rect 9858 35436 9864 35488
rect 9916 35436 9922 35488
rect 10042 35436 10048 35488
rect 10100 35436 10106 35488
rect 10226 35436 10232 35488
rect 10284 35476 10290 35488
rect 11606 35476 11612 35488
rect 10284 35448 11612 35476
rect 10284 35436 10290 35448
rect 11606 35436 11612 35448
rect 11664 35436 11670 35488
rect 12161 35479 12219 35485
rect 12161 35445 12173 35479
rect 12207 35476 12219 35479
rect 12618 35476 12624 35488
rect 12207 35448 12624 35476
rect 12207 35445 12219 35448
rect 12161 35439 12219 35445
rect 12618 35436 12624 35448
rect 12676 35436 12682 35488
rect 12710 35436 12716 35488
rect 12768 35476 12774 35488
rect 13096 35476 13124 35575
rect 14734 35572 14740 35624
rect 14792 35612 14798 35624
rect 19981 35615 20039 35621
rect 19981 35612 19993 35615
rect 14792 35584 19993 35612
rect 14792 35572 14798 35584
rect 19981 35581 19993 35584
rect 20027 35612 20039 35615
rect 20622 35612 20628 35624
rect 20027 35584 20628 35612
rect 20027 35581 20039 35584
rect 19981 35575 20039 35581
rect 20622 35572 20628 35584
rect 20680 35572 20686 35624
rect 22370 35572 22376 35624
rect 22428 35572 22434 35624
rect 22833 35615 22891 35621
rect 22833 35581 22845 35615
rect 22879 35612 22891 35615
rect 23216 35612 23244 35643
rect 23290 35640 23296 35692
rect 23348 35640 23354 35692
rect 23382 35640 23388 35692
rect 23440 35680 23446 35692
rect 23569 35683 23627 35689
rect 23569 35680 23581 35683
rect 23440 35652 23581 35680
rect 23440 35640 23446 35652
rect 23569 35649 23581 35652
rect 23615 35649 23627 35683
rect 23569 35643 23627 35649
rect 23658 35640 23664 35692
rect 23716 35689 23722 35692
rect 23716 35683 23765 35689
rect 23716 35649 23719 35683
rect 23753 35680 23765 35683
rect 24412 35680 24440 35788
rect 25608 35760 25636 35788
rect 25866 35776 25872 35828
rect 25924 35776 25930 35828
rect 25958 35776 25964 35828
rect 26016 35816 26022 35828
rect 26016 35788 26648 35816
rect 26016 35776 26022 35788
rect 24581 35751 24639 35757
rect 24581 35717 24593 35751
rect 24627 35748 24639 35751
rect 24627 35720 25176 35748
rect 24627 35717 24639 35720
rect 24581 35711 24639 35717
rect 25148 35692 25176 35720
rect 25590 35708 25596 35760
rect 25648 35708 25654 35760
rect 25976 35720 26372 35748
rect 23753 35652 24440 35680
rect 23753 35649 23765 35652
rect 23716 35643 23765 35649
rect 23716 35640 23722 35643
rect 24486 35640 24492 35692
rect 24544 35640 24550 35692
rect 24670 35640 24676 35692
rect 24728 35640 24734 35692
rect 24791 35683 24849 35689
rect 24791 35649 24803 35683
rect 24837 35649 24849 35683
rect 24791 35643 24849 35649
rect 24949 35683 25007 35689
rect 24949 35649 24961 35683
rect 24995 35680 25007 35683
rect 25038 35680 25044 35692
rect 24995 35652 25044 35680
rect 24995 35649 25007 35652
rect 24949 35643 25007 35649
rect 23934 35612 23940 35624
rect 22879 35584 23940 35612
rect 22879 35581 22891 35584
rect 22833 35575 22891 35581
rect 23934 35572 23940 35584
rect 23992 35572 23998 35624
rect 24578 35572 24584 35624
rect 24636 35612 24642 35624
rect 24806 35612 24834 35643
rect 25038 35640 25044 35652
rect 25096 35640 25102 35692
rect 25130 35640 25136 35692
rect 25188 35640 25194 35692
rect 24636 35584 24834 35612
rect 24636 35572 24642 35584
rect 13906 35504 13912 35556
rect 13964 35544 13970 35556
rect 14826 35544 14832 35556
rect 13964 35516 14832 35544
rect 13964 35504 13970 35516
rect 14826 35504 14832 35516
rect 14884 35504 14890 35556
rect 19521 35547 19579 35553
rect 19521 35513 19533 35547
rect 19567 35544 19579 35547
rect 25976 35544 26004 35720
rect 26344 35692 26372 35720
rect 26234 35689 26240 35692
rect 26053 35683 26111 35689
rect 26053 35649 26065 35683
rect 26099 35649 26111 35683
rect 26053 35643 26111 35649
rect 26191 35683 26240 35689
rect 26191 35649 26203 35683
rect 26237 35649 26240 35683
rect 26191 35643 26240 35649
rect 26068 35612 26096 35643
rect 26234 35640 26240 35643
rect 26292 35640 26298 35692
rect 26326 35640 26332 35692
rect 26384 35640 26390 35692
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35649 26479 35683
rect 26421 35643 26479 35649
rect 26436 35612 26464 35643
rect 26620 35612 26648 35788
rect 27338 35776 27344 35828
rect 27396 35776 27402 35828
rect 27709 35819 27767 35825
rect 27709 35785 27721 35819
rect 27755 35816 27767 35819
rect 28718 35816 28724 35828
rect 27755 35788 28724 35816
rect 27755 35785 27767 35788
rect 27709 35779 27767 35785
rect 28718 35776 28724 35788
rect 28776 35776 28782 35828
rect 30285 35819 30343 35825
rect 30285 35785 30297 35819
rect 30331 35816 30343 35819
rect 31202 35816 31208 35828
rect 30331 35788 31208 35816
rect 30331 35785 30343 35788
rect 30285 35779 30343 35785
rect 31202 35776 31208 35788
rect 31260 35776 31266 35828
rect 33594 35776 33600 35828
rect 33652 35776 33658 35828
rect 26896 35720 27292 35748
rect 26896 35692 26924 35720
rect 26786 35640 26792 35692
rect 26844 35640 26850 35692
rect 26878 35640 26884 35692
rect 26936 35640 26942 35692
rect 27062 35640 27068 35692
rect 27120 35640 27126 35692
rect 27158 35683 27216 35689
rect 27158 35649 27170 35683
rect 27204 35649 27216 35683
rect 27158 35643 27216 35649
rect 26068 35584 26280 35612
rect 26436 35584 26648 35612
rect 26804 35612 26832 35640
rect 27173 35612 27201 35643
rect 26804 35584 27201 35612
rect 27264 35612 27292 35720
rect 27356 35689 27384 35776
rect 27586 35720 30006 35748
rect 27586 35692 27614 35720
rect 29978 35692 30006 35720
rect 30650 35708 30656 35760
rect 30708 35748 30714 35760
rect 30708 35720 30880 35748
rect 30708 35708 30714 35720
rect 27341 35683 27399 35689
rect 27341 35649 27353 35683
rect 27387 35649 27399 35683
rect 27341 35643 27399 35649
rect 27430 35640 27436 35692
rect 27488 35640 27494 35692
rect 27522 35640 27528 35692
rect 27580 35680 27614 35692
rect 27801 35683 27859 35689
rect 27580 35652 27625 35680
rect 27580 35643 27588 35652
rect 27801 35649 27813 35683
rect 27847 35649 27859 35683
rect 27801 35643 27859 35649
rect 27985 35683 28043 35689
rect 27985 35649 27997 35683
rect 28031 35649 28043 35683
rect 27985 35643 28043 35649
rect 27580 35640 27586 35643
rect 27816 35612 27844 35643
rect 28000 35612 28028 35643
rect 28074 35640 28080 35692
rect 28132 35640 28138 35692
rect 28169 35683 28227 35689
rect 28169 35649 28181 35683
rect 28215 35680 28227 35683
rect 28442 35680 28448 35692
rect 28215 35652 28448 35680
rect 28215 35649 28227 35652
rect 28169 35643 28227 35649
rect 28442 35640 28448 35652
rect 28500 35640 28506 35692
rect 29638 35689 29644 35692
rect 29457 35683 29515 35689
rect 29457 35649 29469 35683
rect 29503 35649 29515 35683
rect 29457 35643 29515 35649
rect 29605 35683 29644 35689
rect 29605 35649 29617 35683
rect 29605 35643 29644 35649
rect 27264 35584 27844 35612
rect 27908 35584 28488 35612
rect 26252 35556 26280 35584
rect 19567 35516 26004 35544
rect 19567 35513 19579 35516
rect 19521 35507 19579 35513
rect 26234 35504 26240 35556
rect 26292 35504 26298 35556
rect 26418 35504 26424 35556
rect 26476 35544 26482 35556
rect 27908 35544 27936 35584
rect 28353 35547 28411 35553
rect 28353 35544 28365 35547
rect 26476 35516 27936 35544
rect 28000 35516 28365 35544
rect 26476 35504 26482 35516
rect 12768 35448 13124 35476
rect 12768 35436 12774 35448
rect 13354 35436 13360 35488
rect 13412 35476 13418 35488
rect 15010 35476 15016 35488
rect 13412 35448 15016 35476
rect 13412 35436 13418 35448
rect 15010 35436 15016 35448
rect 15068 35436 15074 35488
rect 19058 35436 19064 35488
rect 19116 35476 19122 35488
rect 19886 35476 19892 35488
rect 19116 35448 19892 35476
rect 19116 35436 19122 35448
rect 19886 35436 19892 35448
rect 19944 35436 19950 35488
rect 22738 35436 22744 35488
rect 22796 35436 22802 35488
rect 23845 35479 23903 35485
rect 23845 35445 23857 35479
rect 23891 35476 23903 35479
rect 27614 35476 27620 35488
rect 23891 35448 27620 35476
rect 23891 35445 23903 35448
rect 23845 35439 23903 35445
rect 27614 35436 27620 35448
rect 27672 35436 27678 35488
rect 27890 35436 27896 35488
rect 27948 35476 27954 35488
rect 28000 35476 28028 35516
rect 28353 35513 28365 35516
rect 28399 35513 28411 35547
rect 28460 35544 28488 35584
rect 28626 35572 28632 35624
rect 28684 35612 28690 35624
rect 29472 35612 29500 35643
rect 29638 35640 29644 35643
rect 29696 35640 29702 35692
rect 29730 35640 29736 35692
rect 29788 35640 29794 35692
rect 29822 35640 29828 35692
rect 29880 35640 29886 35692
rect 29978 35689 30012 35692
rect 29963 35683 30012 35689
rect 29963 35649 29975 35683
rect 30009 35649 30012 35683
rect 29963 35643 30012 35649
rect 30006 35640 30012 35643
rect 30064 35640 30070 35692
rect 30742 35640 30748 35692
rect 30800 35640 30806 35692
rect 30852 35689 30880 35720
rect 33226 35708 33232 35760
rect 33284 35708 33290 35760
rect 33612 35748 33640 35776
rect 33336 35720 33640 35748
rect 30837 35683 30895 35689
rect 30837 35649 30849 35683
rect 30883 35649 30895 35683
rect 30837 35643 30895 35649
rect 31021 35683 31079 35689
rect 31021 35649 31033 35683
rect 31067 35680 31079 35683
rect 31110 35680 31116 35692
rect 31067 35652 31116 35680
rect 31067 35649 31079 35652
rect 31021 35643 31079 35649
rect 31110 35640 31116 35652
rect 31168 35640 31174 35692
rect 32490 35640 32496 35692
rect 32548 35640 32554 35692
rect 28684 35584 29500 35612
rect 29656 35612 29684 35640
rect 30282 35612 30288 35624
rect 29656 35584 30288 35612
rect 28684 35572 28690 35584
rect 30282 35572 30288 35584
rect 30340 35572 30346 35624
rect 30374 35572 30380 35624
rect 30432 35612 30438 35624
rect 30653 35615 30711 35621
rect 30653 35612 30665 35615
rect 30432 35584 30665 35612
rect 30432 35572 30438 35584
rect 30653 35581 30665 35584
rect 30699 35581 30711 35615
rect 30653 35575 30711 35581
rect 30101 35547 30159 35553
rect 28460 35516 29684 35544
rect 28353 35507 28411 35513
rect 29656 35488 29684 35516
rect 30101 35513 30113 35547
rect 30147 35544 30159 35547
rect 30760 35544 30788 35640
rect 33244 35612 33272 35708
rect 33336 35692 33364 35720
rect 34606 35708 34612 35760
rect 34664 35708 34670 35760
rect 33318 35640 33324 35692
rect 33376 35640 33382 35692
rect 33597 35615 33655 35621
rect 33597 35612 33609 35615
rect 33244 35584 33609 35612
rect 33597 35581 33609 35584
rect 33643 35581 33655 35615
rect 33597 35575 33655 35581
rect 30147 35516 30788 35544
rect 30147 35513 30159 35516
rect 30101 35507 30159 35513
rect 31478 35504 31484 35556
rect 31536 35544 31542 35556
rect 35069 35547 35127 35553
rect 31536 35516 33456 35544
rect 31536 35504 31542 35516
rect 27948 35448 28028 35476
rect 27948 35436 27954 35448
rect 29638 35436 29644 35488
rect 29696 35436 29702 35488
rect 29914 35436 29920 35488
rect 29972 35476 29978 35488
rect 30190 35476 30196 35488
rect 29972 35448 30196 35476
rect 29972 35436 29978 35448
rect 30190 35436 30196 35448
rect 30248 35476 30254 35488
rect 30561 35479 30619 35485
rect 30561 35476 30573 35479
rect 30248 35448 30573 35476
rect 30248 35436 30254 35448
rect 30561 35445 30573 35448
rect 30607 35445 30619 35479
rect 30561 35439 30619 35445
rect 30834 35436 30840 35488
rect 30892 35476 30898 35488
rect 32214 35476 32220 35488
rect 30892 35448 32220 35476
rect 30892 35436 30898 35448
rect 32214 35436 32220 35448
rect 32272 35436 32278 35488
rect 32306 35436 32312 35488
rect 32364 35436 32370 35488
rect 33428 35476 33456 35516
rect 35069 35513 35081 35547
rect 35115 35513 35127 35547
rect 35069 35507 35127 35513
rect 35084 35476 35112 35507
rect 33428 35448 35112 35476
rect 1104 35386 41400 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 41400 35386
rect 1104 35312 41400 35334
rect 6730 35232 6736 35284
rect 6788 35232 6794 35284
rect 8018 35232 8024 35284
rect 8076 35232 8082 35284
rect 9214 35232 9220 35284
rect 9272 35272 9278 35284
rect 9858 35272 9864 35284
rect 9272 35244 9864 35272
rect 9272 35232 9278 35244
rect 9858 35232 9864 35244
rect 9916 35232 9922 35284
rect 10045 35275 10103 35281
rect 10045 35241 10057 35275
rect 10091 35272 10103 35275
rect 10226 35272 10232 35284
rect 10091 35244 10232 35272
rect 10091 35241 10103 35244
rect 10045 35235 10103 35241
rect 10226 35232 10232 35244
rect 10284 35232 10290 35284
rect 10413 35275 10471 35281
rect 10413 35241 10425 35275
rect 10459 35241 10471 35275
rect 13170 35272 13176 35284
rect 10413 35235 10471 35241
rect 10628 35244 13176 35272
rect 8036 35145 8064 35232
rect 8662 35204 8668 35216
rect 8312 35176 8668 35204
rect 8021 35139 8079 35145
rect 8021 35105 8033 35139
rect 8067 35105 8079 35139
rect 8021 35099 8079 35105
rect 6917 35071 6975 35077
rect 6917 35037 6929 35071
rect 6963 35068 6975 35071
rect 7745 35071 7803 35077
rect 6963 35040 7420 35068
rect 6963 35037 6975 35040
rect 6917 35031 6975 35037
rect 7392 34941 7420 35040
rect 7745 35037 7757 35071
rect 7791 35068 7803 35071
rect 8312 35068 8340 35176
rect 8662 35164 8668 35176
rect 8720 35164 8726 35216
rect 9582 35204 9588 35216
rect 8772 35176 9588 35204
rect 8772 35136 8800 35176
rect 9582 35164 9588 35176
rect 9640 35164 9646 35216
rect 9677 35207 9735 35213
rect 9677 35173 9689 35207
rect 9723 35204 9735 35207
rect 10318 35204 10324 35216
rect 9723 35176 10324 35204
rect 9723 35173 9735 35176
rect 9677 35167 9735 35173
rect 10318 35164 10324 35176
rect 10376 35164 10382 35216
rect 8404 35108 8800 35136
rect 8404 35077 8432 35108
rect 9490 35096 9496 35148
rect 9548 35136 9554 35148
rect 9953 35139 10011 35145
rect 9953 35136 9965 35139
rect 9548 35108 9965 35136
rect 9548 35096 9554 35108
rect 9953 35105 9965 35108
rect 9999 35136 10011 35139
rect 10428 35136 10456 35235
rect 9999 35108 10456 35136
rect 9999 35105 10011 35108
rect 9953 35099 10011 35105
rect 10502 35096 10508 35148
rect 10560 35096 10566 35148
rect 7791 35040 8340 35068
rect 8389 35071 8447 35077
rect 7791 35037 7803 35040
rect 7745 35031 7803 35037
rect 8389 35037 8401 35071
rect 8435 35037 8447 35071
rect 8389 35031 8447 35037
rect 8662 35028 8668 35080
rect 8720 35028 8726 35080
rect 9861 35071 9919 35077
rect 9861 35037 9873 35071
rect 9907 35068 9919 35071
rect 10226 35068 10232 35080
rect 9907 35040 10232 35068
rect 9907 35037 9919 35040
rect 9861 35031 9919 35037
rect 10226 35028 10232 35040
rect 10284 35068 10290 35080
rect 10413 35071 10471 35077
rect 10413 35068 10425 35071
rect 10284 35040 10425 35068
rect 10284 35028 10290 35040
rect 10413 35037 10425 35040
rect 10459 35068 10471 35071
rect 10628 35068 10656 35244
rect 13170 35232 13176 35244
rect 13228 35232 13234 35284
rect 13262 35232 13268 35284
rect 13320 35272 13326 35284
rect 22465 35275 22523 35281
rect 13320 35244 16160 35272
rect 13320 35232 13326 35244
rect 10873 35207 10931 35213
rect 10873 35173 10885 35207
rect 10919 35173 10931 35207
rect 10873 35167 10931 35173
rect 10888 35136 10916 35167
rect 12158 35164 12164 35216
rect 12216 35164 12222 35216
rect 12268 35176 15332 35204
rect 10888 35108 11376 35136
rect 10459 35040 10656 35068
rect 10689 35071 10747 35077
rect 10459 35037 10471 35040
rect 10413 35031 10471 35037
rect 10689 35037 10701 35071
rect 10735 35068 10747 35071
rect 10870 35068 10876 35080
rect 10735 35040 10876 35068
rect 10735 35037 10747 35040
rect 10689 35031 10747 35037
rect 10870 35028 10876 35040
rect 10928 35028 10934 35080
rect 11348 35077 11376 35108
rect 11698 35096 11704 35148
rect 11756 35096 11762 35148
rect 11790 35096 11796 35148
rect 11848 35136 11854 35148
rect 12176 35136 12204 35164
rect 11848 35108 12204 35136
rect 11848 35096 11854 35108
rect 11241 35071 11299 35077
rect 11241 35037 11253 35071
rect 11287 35037 11299 35071
rect 11241 35031 11299 35037
rect 11333 35071 11391 35077
rect 11333 35037 11345 35071
rect 11379 35037 11391 35071
rect 11333 35031 11391 35037
rect 8573 35003 8631 35009
rect 8573 34969 8585 35003
rect 8619 34969 8631 35003
rect 8573 34963 8631 34969
rect 7377 34935 7435 34941
rect 7377 34901 7389 34935
rect 7423 34901 7435 34935
rect 7377 34895 7435 34901
rect 7837 34935 7895 34941
rect 7837 34901 7849 34935
rect 7883 34932 7895 34935
rect 8205 34935 8263 34941
rect 8205 34932 8217 34935
rect 7883 34904 8217 34932
rect 7883 34901 7895 34904
rect 7837 34895 7895 34901
rect 8205 34901 8217 34904
rect 8251 34901 8263 34935
rect 8588 34932 8616 34963
rect 9398 34960 9404 35012
rect 9456 34960 9462 35012
rect 9508 34972 10364 35000
rect 9508 34932 9536 34972
rect 8588 34904 9536 34932
rect 8205 34895 8263 34901
rect 9582 34892 9588 34944
rect 9640 34932 9646 34944
rect 10229 34935 10287 34941
rect 10229 34932 10241 34935
rect 9640 34904 10241 34932
rect 9640 34892 9646 34904
rect 10229 34901 10241 34904
rect 10275 34901 10287 34935
rect 10336 34932 10364 34972
rect 10778 34960 10784 35012
rect 10836 34960 10842 35012
rect 11256 35000 11284 35031
rect 11514 35028 11520 35080
rect 11572 35028 11578 35080
rect 11609 35071 11667 35077
rect 11609 35037 11621 35071
rect 11655 35068 11667 35071
rect 11716 35068 11744 35096
rect 11655 35040 11744 35068
rect 11655 35037 11667 35040
rect 11609 35031 11667 35037
rect 11882 35028 11888 35080
rect 11940 35028 11946 35080
rect 11977 35071 12035 35077
rect 11977 35037 11989 35071
rect 12023 35068 12035 35071
rect 12066 35068 12072 35080
rect 12023 35040 12072 35068
rect 12023 35037 12035 35040
rect 11977 35031 12035 35037
rect 12066 35028 12072 35040
rect 12124 35028 12130 35080
rect 12176 35077 12204 35108
rect 12268 35077 12296 35176
rect 13998 35096 14004 35148
rect 14056 35136 14062 35148
rect 14056 35108 15148 35136
rect 14056 35096 14062 35108
rect 12161 35071 12219 35077
rect 12161 35037 12173 35071
rect 12207 35037 12219 35071
rect 12161 35031 12219 35037
rect 12253 35071 12311 35077
rect 12253 35037 12265 35071
rect 12299 35037 12311 35071
rect 12253 35031 12311 35037
rect 11701 35003 11759 35009
rect 11701 35000 11713 35003
rect 11256 34972 11713 35000
rect 11701 34969 11713 34972
rect 11747 34969 11759 35003
rect 11701 34963 11759 34969
rect 10796 34932 10824 34960
rect 10336 34904 10824 34932
rect 10229 34895 10287 34901
rect 11054 34892 11060 34944
rect 11112 34892 11118 34944
rect 11514 34892 11520 34944
rect 11572 34932 11578 34944
rect 11900 34932 11928 35028
rect 12268 35000 12296 35031
rect 12618 35028 12624 35080
rect 12676 35068 12682 35080
rect 13262 35068 13268 35080
rect 12676 35040 13268 35068
rect 12676 35028 12682 35040
rect 13262 35028 13268 35040
rect 13320 35028 13326 35080
rect 13906 35068 13912 35080
rect 13464 35040 13912 35068
rect 12084 34972 12296 35000
rect 12084 34944 12112 34972
rect 12802 34960 12808 35012
rect 12860 35000 12866 35012
rect 12897 35003 12955 35009
rect 12897 35000 12909 35003
rect 12860 34972 12909 35000
rect 12860 34960 12866 34972
rect 12897 34969 12909 34972
rect 12943 35000 12955 35003
rect 13170 35000 13176 35012
rect 12943 34972 13176 35000
rect 12943 34969 12955 34972
rect 12897 34963 12955 34969
rect 13170 34960 13176 34972
rect 13228 34960 13234 35012
rect 13464 35009 13492 35040
rect 13906 35028 13912 35040
rect 13964 35028 13970 35080
rect 14090 35028 14096 35080
rect 14148 35028 14154 35080
rect 14274 35028 14280 35080
rect 14332 35068 14338 35080
rect 14737 35071 14795 35077
rect 14737 35068 14749 35071
rect 14332 35040 14749 35068
rect 14332 35028 14338 35040
rect 14737 35037 14749 35040
rect 14783 35037 14795 35071
rect 14737 35031 14795 35037
rect 14826 35028 14832 35080
rect 14884 35068 14890 35080
rect 14921 35071 14979 35077
rect 14921 35068 14933 35071
rect 14884 35040 14933 35068
rect 14884 35028 14890 35040
rect 14921 35037 14933 35040
rect 14967 35037 14979 35071
rect 14921 35031 14979 35037
rect 15010 35028 15016 35080
rect 15068 35028 15074 35080
rect 15120 35077 15148 35108
rect 15304 35077 15332 35176
rect 15930 35164 15936 35216
rect 15988 35164 15994 35216
rect 15105 35071 15163 35077
rect 15105 35037 15117 35071
rect 15151 35037 15163 35071
rect 15105 35031 15163 35037
rect 15289 35071 15347 35077
rect 15289 35037 15301 35071
rect 15335 35037 15347 35071
rect 15289 35031 15347 35037
rect 15378 35028 15384 35080
rect 15436 35028 15442 35080
rect 16132 35077 16160 35244
rect 22465 35241 22477 35275
rect 22511 35272 22523 35275
rect 22738 35272 22744 35284
rect 22511 35244 22744 35272
rect 22511 35241 22523 35244
rect 22465 35235 22523 35241
rect 22738 35232 22744 35244
rect 22796 35232 22802 35284
rect 22922 35232 22928 35284
rect 22980 35232 22986 35284
rect 23934 35232 23940 35284
rect 23992 35272 23998 35284
rect 25133 35275 25191 35281
rect 25133 35272 25145 35275
rect 23992 35244 25145 35272
rect 23992 35232 23998 35244
rect 25133 35241 25145 35244
rect 25179 35241 25191 35275
rect 26786 35272 26792 35284
rect 25133 35235 25191 35241
rect 26620 35244 26792 35272
rect 16482 35204 16488 35216
rect 16280 35176 16488 35204
rect 16280 35077 16308 35176
rect 16482 35164 16488 35176
rect 16540 35164 16546 35216
rect 16666 35164 16672 35216
rect 16724 35204 16730 35216
rect 16724 35176 17724 35204
rect 16724 35164 16730 35176
rect 17586 35136 17592 35148
rect 16500 35108 17592 35136
rect 16500 35077 16528 35108
rect 17586 35096 17592 35108
rect 17644 35096 17650 35148
rect 17696 35136 17724 35176
rect 18138 35164 18144 35216
rect 18196 35204 18202 35216
rect 18196 35176 22324 35204
rect 18196 35164 18202 35176
rect 17696 35108 22232 35136
rect 15801 35071 15859 35077
rect 15801 35037 15813 35071
rect 15847 35068 15859 35071
rect 16117 35071 16175 35077
rect 15847 35040 15976 35068
rect 15847 35037 15859 35040
rect 15801 35031 15859 35037
rect 13449 35003 13507 35009
rect 13449 34969 13461 35003
rect 13495 34969 13507 35003
rect 13449 34963 13507 34969
rect 13630 34960 13636 35012
rect 13688 34960 13694 35012
rect 13722 34960 13728 35012
rect 13780 35000 13786 35012
rect 14185 35003 14243 35009
rect 14185 35000 14197 35003
rect 13780 34972 14197 35000
rect 13780 34960 13786 34972
rect 14185 34969 14197 34972
rect 14231 34969 14243 35003
rect 14185 34963 14243 34969
rect 15197 35003 15255 35009
rect 15197 34969 15209 35003
rect 15243 35000 15255 35003
rect 15565 35003 15623 35009
rect 15565 35000 15577 35003
rect 15243 34972 15577 35000
rect 15243 34969 15255 34972
rect 15197 34963 15255 34969
rect 15565 34969 15577 34972
rect 15611 34969 15623 35003
rect 15565 34963 15623 34969
rect 15657 35003 15715 35009
rect 15657 34969 15669 35003
rect 15703 34969 15715 35003
rect 15657 34963 15715 34969
rect 11572 34904 11928 34932
rect 11572 34892 11578 34904
rect 12066 34892 12072 34944
rect 12124 34892 12130 34944
rect 13817 34935 13875 34941
rect 13817 34901 13829 34935
rect 13863 34932 13875 34935
rect 14090 34932 14096 34944
rect 13863 34904 14096 34932
rect 13863 34901 13875 34904
rect 13817 34895 13875 34901
rect 14090 34892 14096 34904
rect 14148 34892 14154 34944
rect 14550 34892 14556 34944
rect 14608 34892 14614 34944
rect 15672 34932 15700 34963
rect 15746 34932 15752 34944
rect 15672 34904 15752 34932
rect 15746 34892 15752 34904
rect 15804 34892 15810 34944
rect 15948 34932 15976 35040
rect 16117 35037 16129 35071
rect 16163 35037 16175 35071
rect 16117 35031 16175 35037
rect 16265 35071 16323 35077
rect 16265 35037 16277 35071
rect 16311 35037 16323 35071
rect 16265 35031 16323 35037
rect 16485 35071 16543 35077
rect 16485 35037 16497 35071
rect 16531 35037 16543 35071
rect 16485 35031 16543 35037
rect 16623 35071 16681 35077
rect 16623 35037 16635 35071
rect 16669 35068 16681 35071
rect 17034 35068 17040 35080
rect 16669 35040 17040 35068
rect 16669 35037 16681 35040
rect 16623 35031 16681 35037
rect 17034 35028 17040 35040
rect 17092 35028 17098 35080
rect 17604 35068 17632 35096
rect 20254 35068 20260 35080
rect 17604 35040 20260 35068
rect 20254 35028 20260 35040
rect 20312 35028 20318 35080
rect 16022 34960 16028 35012
rect 16080 35000 16086 35012
rect 16393 35003 16451 35009
rect 16393 35000 16405 35003
rect 16080 34972 16405 35000
rect 16080 34960 16086 34972
rect 16393 34969 16405 34972
rect 16439 34969 16451 35003
rect 21450 35000 21456 35012
rect 16393 34963 16451 34969
rect 16684 34972 21456 35000
rect 16684 34932 16712 34972
rect 21450 34960 21456 34972
rect 21508 34960 21514 35012
rect 15948 34904 16712 34932
rect 16758 34892 16764 34944
rect 16816 34892 16822 34944
rect 18506 34892 18512 34944
rect 18564 34932 18570 34944
rect 20898 34932 20904 34944
rect 18564 34904 20904 34932
rect 18564 34892 18570 34904
rect 20898 34892 20904 34904
rect 20956 34892 20962 34944
rect 22204 34932 22232 35108
rect 22296 35077 22324 35176
rect 22373 35139 22431 35145
rect 22373 35105 22385 35139
rect 22419 35105 22431 35139
rect 22940 35136 22968 35232
rect 24578 35164 24584 35216
rect 24636 35204 24642 35216
rect 26620 35204 26648 35244
rect 26786 35232 26792 35244
rect 26844 35232 26850 35284
rect 27433 35275 27491 35281
rect 27433 35241 27445 35275
rect 27479 35272 27491 35275
rect 27706 35272 27712 35284
rect 27479 35244 27712 35272
rect 27479 35241 27491 35244
rect 27433 35235 27491 35241
rect 27706 35232 27712 35244
rect 27764 35232 27770 35284
rect 28629 35275 28687 35281
rect 28629 35241 28641 35275
rect 28675 35272 28687 35275
rect 28810 35272 28816 35284
rect 28675 35244 28816 35272
rect 28675 35241 28687 35244
rect 28629 35235 28687 35241
rect 28810 35232 28816 35244
rect 28868 35232 28874 35284
rect 28994 35232 29000 35284
rect 29052 35272 29058 35284
rect 30374 35272 30380 35284
rect 29052 35244 30380 35272
rect 29052 35232 29058 35244
rect 30374 35232 30380 35244
rect 30432 35232 30438 35284
rect 31110 35272 31116 35284
rect 30852 35244 31116 35272
rect 24636 35176 26648 35204
rect 24636 35164 24642 35176
rect 26694 35164 26700 35216
rect 26752 35204 26758 35216
rect 27614 35204 27620 35216
rect 26752 35176 27620 35204
rect 26752 35164 26758 35176
rect 27614 35164 27620 35176
rect 27672 35164 27678 35216
rect 28902 35164 28908 35216
rect 28960 35204 28966 35216
rect 30101 35207 30159 35213
rect 28960 35176 29960 35204
rect 28960 35164 28966 35176
rect 26878 35136 26884 35148
rect 22940 35108 26884 35136
rect 22373 35099 22431 35105
rect 22281 35071 22339 35077
rect 22281 35037 22293 35071
rect 22327 35037 22339 35071
rect 22388 35068 22416 35099
rect 23198 35068 23204 35080
rect 22388 35040 23204 35068
rect 22281 35031 22339 35037
rect 23198 35028 23204 35040
rect 23256 35028 23262 35080
rect 24486 35028 24492 35080
rect 24544 35068 24550 35080
rect 24964 35077 24992 35108
rect 26878 35096 26884 35108
rect 26936 35096 26942 35148
rect 27798 35096 27804 35148
rect 27856 35096 27862 35148
rect 27893 35139 27951 35145
rect 27893 35105 27905 35139
rect 27939 35136 27951 35139
rect 28350 35136 28356 35148
rect 27939 35108 28356 35136
rect 27939 35105 27951 35108
rect 27893 35099 27951 35105
rect 28350 35096 28356 35108
rect 28408 35096 28414 35148
rect 28736 35108 29040 35136
rect 24581 35071 24639 35077
rect 24581 35068 24593 35071
rect 24544 35040 24593 35068
rect 24544 35028 24550 35040
rect 24581 35037 24593 35040
rect 24627 35037 24639 35071
rect 24581 35031 24639 35037
rect 24949 35071 25007 35077
rect 24949 35037 24961 35071
rect 24995 35037 25007 35071
rect 24949 35031 25007 35037
rect 25038 35028 25044 35080
rect 25096 35068 25102 35080
rect 25225 35071 25283 35077
rect 25225 35068 25237 35071
rect 25096 35040 25237 35068
rect 25096 35028 25102 35040
rect 25225 35037 25237 35040
rect 25271 35037 25283 35071
rect 25225 35031 25283 35037
rect 25406 35028 25412 35080
rect 25464 35028 25470 35080
rect 25590 35028 25596 35080
rect 25648 35068 25654 35080
rect 25866 35068 25872 35080
rect 25648 35040 25872 35068
rect 25648 35028 25654 35040
rect 25866 35028 25872 35040
rect 25924 35068 25930 35080
rect 26234 35068 26240 35080
rect 25924 35040 26240 35068
rect 25924 35028 25930 35040
rect 26234 35028 26240 35040
rect 26292 35028 26298 35080
rect 27522 35028 27528 35080
rect 27580 35068 27586 35080
rect 27617 35071 27675 35077
rect 27617 35068 27629 35071
rect 27580 35040 27629 35068
rect 27580 35028 27586 35040
rect 27617 35037 27629 35040
rect 27663 35037 27675 35071
rect 27617 35031 27675 35037
rect 27709 35071 27767 35077
rect 27709 35037 27721 35071
rect 27755 35068 27767 35071
rect 28736 35068 28764 35108
rect 27755 35040 28764 35068
rect 27755 35037 27767 35040
rect 27709 35031 27767 35037
rect 22554 34960 22560 35012
rect 22612 34960 22618 35012
rect 24765 35003 24823 35009
rect 24765 34969 24777 35003
rect 24811 34969 24823 35003
rect 24765 34963 24823 34969
rect 24857 35003 24915 35009
rect 24857 34969 24869 35003
rect 24903 35000 24915 35003
rect 25056 35000 25084 35028
rect 28368 35012 28396 35040
rect 28810 35028 28816 35080
rect 28868 35028 28874 35080
rect 29012 35077 29040 35108
rect 28997 35071 29055 35077
rect 28997 35037 29009 35071
rect 29043 35037 29055 35071
rect 28997 35031 29055 35037
rect 29270 35028 29276 35080
rect 29328 35028 29334 35080
rect 29362 35028 29368 35080
rect 29420 35078 29426 35080
rect 29420 35077 29592 35078
rect 29420 35071 29607 35077
rect 29420 35050 29561 35071
rect 29420 35028 29426 35050
rect 29549 35037 29561 35050
rect 29595 35037 29607 35071
rect 29549 35031 29607 35037
rect 29638 35028 29644 35080
rect 29696 35068 29702 35080
rect 29932 35077 29960 35176
rect 30101 35173 30113 35207
rect 30147 35204 30159 35207
rect 30466 35204 30472 35216
rect 30147 35176 30472 35204
rect 30147 35173 30159 35176
rect 30101 35167 30159 35173
rect 30466 35164 30472 35176
rect 30524 35164 30530 35216
rect 30852 35136 30880 35244
rect 31110 35232 31116 35244
rect 31168 35272 31174 35284
rect 31168 35244 31754 35272
rect 31168 35232 31174 35244
rect 30926 35164 30932 35216
rect 30984 35164 30990 35216
rect 31021 35207 31079 35213
rect 31021 35173 31033 35207
rect 31067 35204 31079 35207
rect 31570 35204 31576 35216
rect 31067 35176 31576 35204
rect 31067 35173 31079 35176
rect 31021 35167 31079 35173
rect 31570 35164 31576 35176
rect 31628 35164 31634 35216
rect 31726 35204 31754 35244
rect 32306 35232 32312 35284
rect 32364 35272 32370 35284
rect 32658 35275 32716 35281
rect 32658 35272 32670 35275
rect 32364 35244 32670 35272
rect 32364 35232 32370 35244
rect 32658 35241 32670 35244
rect 32704 35241 32716 35275
rect 32658 35235 32716 35241
rect 31726 35176 31800 35204
rect 30760 35108 30880 35136
rect 30944 35136 30972 35164
rect 30944 35108 31248 35136
rect 29733 35071 29791 35077
rect 29733 35068 29745 35071
rect 29696 35040 29745 35068
rect 29696 35028 29702 35040
rect 29733 35037 29745 35040
rect 29779 35037 29791 35071
rect 29733 35031 29791 35037
rect 29917 35071 29975 35077
rect 29917 35037 29929 35071
rect 29963 35037 29975 35071
rect 29917 35031 29975 35037
rect 30374 35028 30380 35080
rect 30432 35077 30438 35080
rect 30432 35068 30442 35077
rect 30525 35071 30583 35077
rect 30432 35040 30477 35068
rect 30432 35031 30442 35040
rect 30525 35037 30537 35071
rect 30571 35068 30583 35071
rect 30760 35068 30788 35108
rect 30571 35040 30788 35068
rect 30842 35071 30900 35077
rect 30571 35037 30583 35040
rect 30525 35031 30583 35037
rect 30842 35037 30854 35071
rect 30888 35037 30900 35071
rect 30842 35031 30900 35037
rect 30432 35028 30438 35031
rect 24903 34972 25084 35000
rect 25501 35003 25559 35009
rect 24903 34969 24915 34972
rect 24857 34963 24915 34969
rect 25501 34969 25513 35003
rect 25547 34969 25559 35003
rect 27982 35000 27988 35012
rect 25501 34963 25559 34969
rect 25608 34972 27988 35000
rect 23290 34932 23296 34944
rect 22204 34904 23296 34932
rect 23290 34892 23296 34904
rect 23348 34892 23354 34944
rect 24780 34932 24808 34963
rect 24946 34932 24952 34944
rect 24780 34904 24952 34932
rect 24946 34892 24952 34904
rect 25004 34892 25010 34944
rect 25038 34892 25044 34944
rect 25096 34932 25102 34944
rect 25516 34932 25544 34963
rect 25608 34944 25636 34972
rect 27982 34960 27988 34972
rect 28040 34960 28046 35012
rect 28350 34960 28356 35012
rect 28408 34960 28414 35012
rect 28718 34960 28724 35012
rect 28776 35000 28782 35012
rect 28905 35003 28963 35009
rect 28905 35000 28917 35003
rect 28776 34972 28917 35000
rect 28776 34960 28782 34972
rect 28905 34969 28917 34972
rect 28951 34969 28963 35003
rect 29135 35003 29193 35009
rect 29135 35000 29147 35003
rect 28905 34963 28963 34969
rect 29130 34969 29147 35000
rect 29181 34969 29193 35003
rect 29130 34963 29193 34969
rect 29825 35003 29883 35009
rect 29825 34969 29837 35003
rect 29871 35000 29883 35003
rect 30653 35003 30711 35009
rect 30653 35000 30665 35003
rect 29871 34972 30052 35000
rect 29871 34969 29883 34972
rect 29825 34963 29883 34969
rect 29130 34944 29158 34963
rect 25096 34904 25544 34932
rect 25096 34892 25102 34904
rect 25590 34892 25596 34944
rect 25648 34892 25654 34944
rect 25777 34935 25835 34941
rect 25777 34901 25789 34935
rect 25823 34932 25835 34935
rect 28810 34932 28816 34944
rect 25823 34904 28816 34932
rect 25823 34901 25835 34904
rect 25777 34895 25835 34901
rect 28810 34892 28816 34904
rect 28868 34892 28874 34944
rect 29086 34892 29092 34944
rect 29144 34904 29158 34944
rect 30024 34932 30052 34972
rect 30392 34972 30665 35000
rect 30392 34944 30420 34972
rect 30653 34969 30665 34972
rect 30699 34969 30711 35003
rect 30653 34963 30711 34969
rect 30745 35003 30803 35009
rect 30745 34969 30757 35003
rect 30791 34969 30803 35003
rect 30745 34963 30803 34969
rect 30190 34932 30196 34944
rect 30024 34904 30196 34932
rect 29144 34892 29150 34904
rect 30190 34892 30196 34904
rect 30248 34892 30254 34944
rect 30374 34892 30380 34944
rect 30432 34892 30438 34944
rect 30466 34892 30472 34944
rect 30524 34932 30530 34944
rect 30760 34932 30788 34963
rect 30857 34944 30885 35031
rect 31110 35028 31116 35080
rect 31168 35028 31174 35080
rect 31220 35077 31248 35108
rect 31386 35096 31392 35148
rect 31444 35096 31450 35148
rect 31772 35136 31800 35176
rect 32401 35139 32459 35145
rect 31772 35108 31984 35136
rect 31205 35071 31263 35077
rect 31205 35037 31217 35071
rect 31251 35037 31263 35071
rect 31205 35031 31263 35037
rect 31294 35028 31300 35080
rect 31352 35028 31358 35080
rect 31404 35068 31432 35096
rect 31670 35071 31728 35077
rect 31670 35068 31682 35071
rect 31404 35040 31682 35068
rect 31670 35037 31682 35040
rect 31716 35037 31728 35071
rect 31670 35031 31728 35037
rect 31846 35028 31852 35080
rect 31904 35028 31910 35080
rect 31956 35077 31984 35108
rect 32401 35105 32413 35139
rect 32447 35136 32459 35139
rect 33318 35136 33324 35148
rect 32447 35108 33324 35136
rect 32447 35105 32459 35108
rect 32401 35099 32459 35105
rect 33318 35096 33324 35108
rect 33376 35096 33382 35148
rect 34514 35096 34520 35148
rect 34572 35136 34578 35148
rect 34882 35136 34888 35148
rect 34572 35108 34888 35136
rect 34572 35096 34578 35108
rect 34882 35096 34888 35108
rect 34940 35096 34946 35148
rect 31941 35071 31999 35077
rect 31941 35037 31953 35071
rect 31987 35037 31999 35071
rect 31941 35031 31999 35037
rect 32030 35028 32036 35080
rect 32088 35068 32094 35080
rect 32125 35071 32183 35077
rect 32125 35068 32137 35071
rect 32088 35040 32137 35068
rect 32088 35028 32094 35040
rect 32125 35037 32137 35040
rect 32171 35037 32183 35071
rect 34606 35068 34612 35080
rect 33810 35040 34612 35068
rect 32125 35031 32183 35037
rect 34606 35028 34612 35040
rect 34664 35028 34670 35080
rect 34790 35028 34796 35080
rect 34848 35028 34854 35080
rect 31128 35000 31156 35028
rect 31481 35003 31539 35009
rect 31481 35000 31493 35003
rect 31128 34972 31493 35000
rect 31481 34969 31493 34972
rect 31527 34969 31539 35003
rect 31481 34963 31539 34969
rect 31570 34960 31576 35012
rect 31628 34960 31634 35012
rect 30524 34904 30788 34932
rect 30524 34892 30530 34904
rect 30834 34892 30840 34944
rect 30892 34892 30898 34944
rect 31864 34941 31892 35028
rect 31849 34935 31907 34941
rect 31849 34901 31861 34935
rect 31895 34901 31907 34935
rect 31849 34895 31907 34901
rect 32030 34892 32036 34944
rect 32088 34892 32094 34944
rect 32398 34892 32404 34944
rect 32456 34932 32462 34944
rect 34149 34935 34207 34941
rect 34149 34932 34161 34935
rect 32456 34904 34161 34932
rect 32456 34892 32462 34904
rect 34149 34901 34161 34904
rect 34195 34901 34207 34935
rect 34149 34895 34207 34901
rect 34606 34892 34612 34944
rect 34664 34932 34670 34944
rect 34885 34935 34943 34941
rect 34885 34932 34897 34935
rect 34664 34904 34897 34932
rect 34664 34892 34670 34904
rect 34885 34901 34897 34904
rect 34931 34901 34943 34935
rect 34885 34895 34943 34901
rect 1104 34842 41400 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 41400 34842
rect 1104 34768 41400 34790
rect 9398 34688 9404 34740
rect 9456 34728 9462 34740
rect 10229 34731 10287 34737
rect 10229 34728 10241 34731
rect 9456 34700 10241 34728
rect 9456 34688 9462 34700
rect 10229 34697 10241 34700
rect 10275 34697 10287 34731
rect 10229 34691 10287 34697
rect 13081 34731 13139 34737
rect 13081 34697 13093 34731
rect 13127 34728 13139 34731
rect 13127 34700 13860 34728
rect 13127 34697 13139 34700
rect 13081 34691 13139 34697
rect 5534 34620 5540 34672
rect 5592 34660 5598 34672
rect 6641 34663 6699 34669
rect 6641 34660 6653 34663
rect 5592 34632 6653 34660
rect 5592 34620 5598 34632
rect 6641 34629 6653 34632
rect 6687 34660 6699 34663
rect 6822 34660 6828 34672
rect 6687 34632 6828 34660
rect 6687 34629 6699 34632
rect 6641 34623 6699 34629
rect 6822 34620 6828 34632
rect 6880 34620 6886 34672
rect 9214 34620 9220 34672
rect 9272 34660 9278 34672
rect 9309 34663 9367 34669
rect 9309 34660 9321 34663
rect 9272 34632 9321 34660
rect 9272 34620 9278 34632
rect 9309 34629 9321 34632
rect 9355 34629 9367 34663
rect 9861 34663 9919 34669
rect 9861 34660 9873 34663
rect 9309 34623 9367 34629
rect 9508 34632 9873 34660
rect 9508 34601 9536 34632
rect 9861 34629 9873 34632
rect 9907 34660 9919 34663
rect 11790 34660 11796 34672
rect 9907 34632 11796 34660
rect 9907 34629 9919 34632
rect 9861 34623 9919 34629
rect 11790 34620 11796 34632
rect 11848 34620 11854 34672
rect 13170 34620 13176 34672
rect 13228 34660 13234 34672
rect 13228 34632 13584 34660
rect 13228 34620 13234 34632
rect 9493 34595 9551 34601
rect 9493 34561 9505 34595
rect 9539 34561 9551 34595
rect 9493 34555 9551 34561
rect 9585 34595 9643 34601
rect 9585 34561 9597 34595
rect 9631 34561 9643 34595
rect 9585 34555 9643 34561
rect 10045 34595 10103 34601
rect 10045 34561 10057 34595
rect 10091 34561 10103 34595
rect 10045 34555 10103 34561
rect 5994 34484 6000 34536
rect 6052 34524 6058 34536
rect 7377 34527 7435 34533
rect 7377 34524 7389 34527
rect 6052 34496 7389 34524
rect 6052 34484 6058 34496
rect 7377 34493 7389 34496
rect 7423 34493 7435 34527
rect 7377 34487 7435 34493
rect 9306 34484 9312 34536
rect 9364 34524 9370 34536
rect 9600 34524 9628 34555
rect 10060 34524 10088 34555
rect 10134 34552 10140 34604
rect 10192 34592 10198 34604
rect 11882 34592 11888 34604
rect 10192 34564 11888 34592
rect 10192 34552 10198 34564
rect 11882 34552 11888 34564
rect 11940 34552 11946 34604
rect 12621 34595 12679 34601
rect 12621 34561 12633 34595
rect 12667 34592 12679 34595
rect 12710 34592 12716 34604
rect 12667 34564 12716 34592
rect 12667 34561 12679 34564
rect 12621 34555 12679 34561
rect 12710 34552 12716 34564
rect 12768 34552 12774 34604
rect 13354 34592 13360 34604
rect 12820 34564 13360 34592
rect 9364 34496 9628 34524
rect 9876 34496 10088 34524
rect 9364 34484 9370 34496
rect 9876 34456 9904 34496
rect 11422 34484 11428 34536
rect 11480 34524 11486 34536
rect 12820 34524 12848 34564
rect 13354 34552 13360 34564
rect 13412 34552 13418 34604
rect 13556 34601 13584 34632
rect 13449 34595 13507 34601
rect 13449 34561 13461 34595
rect 13495 34561 13507 34595
rect 13449 34555 13507 34561
rect 13541 34595 13599 34601
rect 13541 34561 13553 34595
rect 13587 34561 13599 34595
rect 13541 34555 13599 34561
rect 11480 34496 12848 34524
rect 11480 34484 11486 34496
rect 9324 34428 9904 34456
rect 9030 34348 9036 34400
rect 9088 34388 9094 34400
rect 9324 34397 9352 34428
rect 10042 34416 10048 34468
rect 10100 34416 10106 34468
rect 13464 34456 13492 34555
rect 13722 34552 13728 34604
rect 13780 34552 13786 34604
rect 13832 34601 13860 34700
rect 13998 34688 14004 34740
rect 14056 34688 14062 34740
rect 14461 34731 14519 34737
rect 14461 34697 14473 34731
rect 14507 34697 14519 34731
rect 17770 34728 17776 34740
rect 14461 34691 14519 34697
rect 15948 34700 17776 34728
rect 14016 34660 14044 34688
rect 14093 34663 14151 34669
rect 14093 34660 14105 34663
rect 14016 34632 14105 34660
rect 14093 34629 14105 34632
rect 14139 34629 14151 34663
rect 14093 34623 14151 34629
rect 13817 34595 13875 34601
rect 13817 34561 13829 34595
rect 13863 34561 13875 34595
rect 13817 34555 13875 34561
rect 13965 34595 14023 34601
rect 13965 34561 13977 34595
rect 14011 34561 14023 34595
rect 13965 34555 14023 34561
rect 14185 34595 14243 34601
rect 14185 34561 14197 34595
rect 14231 34561 14243 34595
rect 14185 34555 14243 34561
rect 14282 34595 14340 34601
rect 14282 34561 14294 34595
rect 14328 34592 14340 34595
rect 14476 34592 14504 34691
rect 14553 34595 14611 34601
rect 14553 34592 14565 34595
rect 14328 34564 14412 34592
rect 14476 34564 14565 34592
rect 14328 34561 14340 34564
rect 14282 34555 14340 34561
rect 13980 34524 14008 34555
rect 14090 34524 14096 34536
rect 13980 34496 14096 34524
rect 14090 34484 14096 34496
rect 14148 34484 14154 34536
rect 14200 34524 14228 34555
rect 14200 34496 14320 34524
rect 14182 34456 14188 34468
rect 13464 34428 14188 34456
rect 14182 34416 14188 34428
rect 14240 34416 14246 34468
rect 9309 34391 9367 34397
rect 9309 34388 9321 34391
rect 9088 34360 9321 34388
rect 9088 34348 9094 34360
rect 9309 34357 9321 34360
rect 9355 34357 9367 34391
rect 9309 34351 9367 34357
rect 9398 34348 9404 34400
rect 9456 34388 9462 34400
rect 9674 34388 9680 34400
rect 9456 34360 9680 34388
rect 9456 34348 9462 34360
rect 9674 34348 9680 34360
rect 9732 34348 9738 34400
rect 9769 34391 9827 34397
rect 9769 34357 9781 34391
rect 9815 34388 9827 34391
rect 10060 34388 10088 34416
rect 9815 34360 10088 34388
rect 9815 34357 9827 34360
rect 9769 34351 9827 34357
rect 12618 34348 12624 34400
rect 12676 34388 12682 34400
rect 12713 34391 12771 34397
rect 12713 34388 12725 34391
rect 12676 34360 12725 34388
rect 12676 34348 12682 34360
rect 12713 34357 12725 34360
rect 12759 34357 12771 34391
rect 12713 34351 12771 34357
rect 13446 34348 13452 34400
rect 13504 34388 13510 34400
rect 14292 34388 14320 34496
rect 14384 34456 14412 34564
rect 14553 34561 14565 34564
rect 14599 34561 14611 34595
rect 14553 34555 14611 34561
rect 14737 34595 14795 34601
rect 14737 34561 14749 34595
rect 14783 34592 14795 34595
rect 15948 34592 15976 34700
rect 17770 34688 17776 34700
rect 17828 34688 17834 34740
rect 18877 34731 18935 34737
rect 18877 34697 18889 34731
rect 18923 34697 18935 34731
rect 18877 34691 18935 34697
rect 16022 34620 16028 34672
rect 16080 34620 16086 34672
rect 18892 34660 18920 34691
rect 19150 34688 19156 34740
rect 19208 34688 19214 34740
rect 21450 34688 21456 34740
rect 21508 34688 21514 34740
rect 22189 34731 22247 34737
rect 22189 34697 22201 34731
rect 22235 34728 22247 34731
rect 22370 34728 22376 34740
rect 22235 34700 22376 34728
rect 22235 34697 22247 34700
rect 22189 34691 22247 34697
rect 22370 34688 22376 34700
rect 22428 34688 22434 34740
rect 26050 34688 26056 34740
rect 26108 34688 26114 34740
rect 26878 34688 26884 34740
rect 26936 34728 26942 34740
rect 27985 34731 28043 34737
rect 26936 34700 27476 34728
rect 26936 34688 26942 34700
rect 19168 34660 19196 34688
rect 17144 34632 17448 34660
rect 14783 34564 15976 34592
rect 14783 34561 14795 34564
rect 14737 34555 14795 34561
rect 14458 34484 14464 34536
rect 14516 34524 14522 34536
rect 14752 34524 14780 34555
rect 14516 34496 14780 34524
rect 14516 34484 14522 34496
rect 14826 34484 14832 34536
rect 14884 34524 14890 34536
rect 16040 34524 16068 34620
rect 17144 34604 17172 34632
rect 16758 34552 16764 34604
rect 16816 34592 16822 34604
rect 16945 34595 17003 34601
rect 16945 34592 16957 34595
rect 16816 34564 16957 34592
rect 16816 34552 16822 34564
rect 16945 34561 16957 34564
rect 16991 34561 17003 34595
rect 16945 34555 17003 34561
rect 17126 34552 17132 34604
rect 17184 34552 17190 34604
rect 17218 34552 17224 34604
rect 17276 34552 17282 34604
rect 17420 34601 17448 34632
rect 17512 34632 18920 34660
rect 19076 34632 19196 34660
rect 20993 34663 21051 34669
rect 17512 34601 17540 34632
rect 17405 34595 17463 34601
rect 17405 34561 17417 34595
rect 17451 34561 17463 34595
rect 17405 34555 17463 34561
rect 17497 34595 17555 34601
rect 17497 34561 17509 34595
rect 17543 34561 17555 34595
rect 17497 34555 17555 34561
rect 14884 34496 16068 34524
rect 17037 34527 17095 34533
rect 14884 34484 14890 34496
rect 17037 34493 17049 34527
rect 17083 34524 17095 34527
rect 17512 34524 17540 34555
rect 17586 34552 17592 34604
rect 17644 34592 17650 34604
rect 17773 34595 17831 34601
rect 17644 34564 17689 34592
rect 17644 34552 17650 34564
rect 17773 34561 17785 34595
rect 17819 34561 17831 34595
rect 17773 34555 17831 34561
rect 17083 34496 17540 34524
rect 17083 34493 17095 34496
rect 17037 34487 17095 34493
rect 17678 34484 17684 34536
rect 17736 34524 17742 34536
rect 17788 34524 17816 34555
rect 17862 34552 17868 34604
rect 17920 34552 17926 34604
rect 18046 34601 18052 34604
rect 18003 34595 18052 34601
rect 18003 34561 18015 34595
rect 18049 34561 18052 34595
rect 18003 34555 18052 34561
rect 18046 34552 18052 34555
rect 18104 34552 18110 34604
rect 18325 34595 18383 34601
rect 18325 34561 18337 34595
rect 18371 34561 18383 34595
rect 18325 34555 18383 34561
rect 18340 34524 18368 34555
rect 18506 34552 18512 34604
rect 18564 34552 18570 34604
rect 18598 34552 18604 34604
rect 18656 34552 18662 34604
rect 18693 34595 18751 34601
rect 18693 34561 18705 34595
rect 18739 34592 18751 34595
rect 19076 34592 19104 34632
rect 20993 34629 21005 34663
rect 21039 34660 21051 34663
rect 22465 34663 22523 34669
rect 21039 34632 22140 34660
rect 21039 34629 21051 34632
rect 20993 34623 21051 34629
rect 22112 34604 22140 34632
rect 22465 34629 22477 34663
rect 22511 34660 22523 34663
rect 22554 34660 22560 34672
rect 22511 34632 22560 34660
rect 22511 34629 22523 34632
rect 22465 34623 22523 34629
rect 22554 34620 22560 34632
rect 22612 34660 22618 34672
rect 22612 34632 27108 34660
rect 22612 34620 22618 34632
rect 18739 34564 19104 34592
rect 19153 34595 19211 34601
rect 18739 34561 18751 34564
rect 18693 34555 18751 34561
rect 19153 34561 19165 34595
rect 19199 34561 19211 34595
rect 19153 34555 19211 34561
rect 21269 34595 21327 34601
rect 21269 34561 21281 34595
rect 21315 34592 21327 34595
rect 21634 34592 21640 34604
rect 21315 34564 21640 34592
rect 21315 34561 21327 34564
rect 21269 34555 21327 34561
rect 19168 34524 19196 34555
rect 21634 34552 21640 34564
rect 21692 34552 21698 34604
rect 22094 34552 22100 34604
rect 22152 34552 22158 34604
rect 22189 34595 22247 34601
rect 22189 34561 22201 34595
rect 22235 34592 22247 34595
rect 22646 34592 22652 34604
rect 22235 34564 22652 34592
rect 22235 34561 22247 34564
rect 22189 34555 22247 34561
rect 22646 34552 22652 34564
rect 22704 34592 22710 34604
rect 25961 34595 26019 34601
rect 25961 34592 25973 34595
rect 22704 34564 25973 34592
rect 22704 34552 22710 34564
rect 25961 34561 25973 34564
rect 26007 34592 26019 34595
rect 26050 34592 26056 34604
rect 26007 34564 26056 34592
rect 26007 34561 26019 34564
rect 25961 34555 26019 34561
rect 26050 34552 26056 34564
rect 26108 34552 26114 34604
rect 26145 34595 26203 34601
rect 26145 34561 26157 34595
rect 26191 34561 26203 34595
rect 26145 34555 26203 34561
rect 26150 34554 26188 34555
rect 17736 34496 17816 34524
rect 18067 34496 19196 34524
rect 19429 34527 19487 34533
rect 17736 34484 17742 34496
rect 15194 34456 15200 34468
rect 14384 34428 15200 34456
rect 15194 34416 15200 34428
rect 15252 34416 15258 34468
rect 18067 34456 18095 34496
rect 19429 34493 19441 34527
rect 19475 34524 19487 34527
rect 20806 34524 20812 34536
rect 19475 34496 20812 34524
rect 19475 34493 19487 34496
rect 19429 34487 19487 34493
rect 20806 34484 20812 34496
rect 20864 34484 20870 34536
rect 21177 34527 21235 34533
rect 21177 34493 21189 34527
rect 21223 34524 21235 34527
rect 25222 34524 25228 34536
rect 21223 34496 25228 34524
rect 21223 34493 21235 34496
rect 21177 34487 21235 34493
rect 25222 34484 25228 34496
rect 25280 34524 25286 34536
rect 25590 34524 25596 34536
rect 25280 34496 25596 34524
rect 25280 34484 25286 34496
rect 25590 34484 25596 34496
rect 25648 34484 25654 34536
rect 26150 34524 26178 34554
rect 27080 34536 27108 34632
rect 27448 34601 27476 34700
rect 27985 34697 27997 34731
rect 28031 34728 28043 34731
rect 28258 34728 28264 34740
rect 28031 34700 28264 34728
rect 28031 34697 28043 34700
rect 27985 34691 28043 34697
rect 28258 34688 28264 34700
rect 28316 34688 28322 34740
rect 29825 34731 29883 34737
rect 29825 34697 29837 34731
rect 29871 34728 29883 34731
rect 29914 34728 29920 34740
rect 29871 34700 29920 34728
rect 29871 34697 29883 34700
rect 29825 34691 29883 34697
rect 29914 34688 29920 34700
rect 29972 34688 29978 34740
rect 30282 34728 30288 34740
rect 30024 34700 30288 34728
rect 27614 34620 27620 34672
rect 27672 34620 27678 34672
rect 29549 34663 29607 34669
rect 29549 34660 29561 34663
rect 29104 34632 29561 34660
rect 29104 34604 29132 34632
rect 29549 34629 29561 34632
rect 29595 34629 29607 34663
rect 29549 34623 29607 34629
rect 27433 34595 27491 34601
rect 27433 34561 27445 34595
rect 27479 34561 27491 34595
rect 27433 34555 27491 34561
rect 27706 34552 27712 34604
rect 27764 34552 27770 34604
rect 27801 34595 27859 34601
rect 27801 34561 27813 34595
rect 27847 34592 27859 34595
rect 28442 34592 28448 34604
rect 27847 34564 28448 34592
rect 27847 34561 27859 34564
rect 27801 34555 27859 34561
rect 28442 34552 28448 34564
rect 28500 34552 28506 34604
rect 29086 34552 29092 34604
rect 29144 34552 29150 34604
rect 29273 34595 29331 34601
rect 29273 34561 29285 34595
rect 29319 34592 29331 34595
rect 29362 34592 29368 34604
rect 29319 34564 29368 34592
rect 29319 34561 29331 34564
rect 29273 34555 29331 34561
rect 29362 34552 29368 34564
rect 29420 34552 29426 34604
rect 29457 34595 29515 34601
rect 29457 34561 29469 34595
rect 29503 34592 29515 34595
rect 29641 34595 29699 34601
rect 29503 34564 29592 34592
rect 29503 34561 29515 34564
rect 29457 34555 29515 34561
rect 26150 34496 26280 34524
rect 26252 34468 26280 34496
rect 27062 34484 27068 34536
rect 27120 34484 27126 34536
rect 28460 34524 28488 34552
rect 29564 34524 29592 34564
rect 29641 34561 29653 34595
rect 29687 34592 29699 34595
rect 29914 34592 29920 34604
rect 29687 34564 29920 34592
rect 29687 34561 29699 34564
rect 29641 34555 29699 34561
rect 29914 34552 29920 34564
rect 29972 34552 29978 34604
rect 30024 34601 30052 34700
rect 30282 34688 30288 34700
rect 30340 34688 30346 34740
rect 30561 34731 30619 34737
rect 30561 34697 30573 34731
rect 30607 34728 30619 34731
rect 30650 34728 30656 34740
rect 30607 34700 30656 34728
rect 30607 34697 30619 34700
rect 30561 34691 30619 34697
rect 30650 34688 30656 34700
rect 30708 34688 30714 34740
rect 30834 34688 30840 34740
rect 30892 34728 30898 34740
rect 31294 34728 31300 34740
rect 30892 34700 31300 34728
rect 30892 34688 30898 34700
rect 31294 34688 31300 34700
rect 31352 34688 31358 34740
rect 35069 34731 35127 34737
rect 35069 34728 35081 34731
rect 31404 34700 32352 34728
rect 30193 34663 30251 34669
rect 30193 34629 30205 34663
rect 30239 34660 30251 34663
rect 30742 34660 30748 34672
rect 30239 34632 30748 34660
rect 30239 34629 30251 34632
rect 30193 34623 30251 34629
rect 30742 34620 30748 34632
rect 30800 34620 30806 34672
rect 30009 34595 30067 34601
rect 30009 34561 30021 34595
rect 30055 34561 30067 34595
rect 30009 34555 30067 34561
rect 30282 34552 30288 34604
rect 30340 34552 30346 34604
rect 30377 34595 30435 34601
rect 30377 34561 30389 34595
rect 30423 34592 30435 34595
rect 30653 34595 30711 34601
rect 30653 34592 30665 34595
rect 30423 34564 30665 34592
rect 30423 34561 30435 34564
rect 30377 34555 30435 34561
rect 30653 34561 30665 34564
rect 30699 34561 30711 34595
rect 31404 34592 31432 34700
rect 31846 34660 31852 34672
rect 31680 34632 31852 34660
rect 31680 34601 31708 34632
rect 31846 34620 31852 34632
rect 31904 34620 31910 34672
rect 32214 34620 32220 34672
rect 32272 34620 32278 34672
rect 32324 34604 32352 34700
rect 34900 34700 35081 34728
rect 34900 34660 34928 34700
rect 35069 34697 35081 34700
rect 35115 34697 35127 34731
rect 35069 34691 35127 34697
rect 33888 34632 34928 34660
rect 35084 34632 35664 34660
rect 31481 34595 31539 34601
rect 31481 34592 31493 34595
rect 31404 34564 31493 34592
rect 30653 34555 30711 34561
rect 31481 34561 31493 34564
rect 31527 34561 31539 34595
rect 31481 34555 31539 34561
rect 31665 34595 31723 34601
rect 31665 34561 31677 34595
rect 31711 34561 31723 34595
rect 31665 34555 31723 34561
rect 31757 34595 31815 34601
rect 31757 34561 31769 34595
rect 31803 34592 31815 34595
rect 32030 34592 32036 34604
rect 31803 34564 32036 34592
rect 31803 34561 31815 34564
rect 31757 34555 31815 34561
rect 29730 34524 29736 34536
rect 28460 34496 28994 34524
rect 29564 34496 29736 34524
rect 17052 34428 18095 34456
rect 17052 34400 17080 34428
rect 18138 34416 18144 34468
rect 18196 34416 18202 34468
rect 19337 34459 19395 34465
rect 19337 34425 19349 34459
rect 19383 34456 19395 34459
rect 21910 34456 21916 34468
rect 19383 34428 21916 34456
rect 19383 34425 19395 34428
rect 19337 34419 19395 34425
rect 21910 34416 21916 34428
rect 21968 34416 21974 34468
rect 22278 34416 22284 34468
rect 22336 34456 22342 34468
rect 24210 34456 24216 34468
rect 22336 34428 24216 34456
rect 22336 34416 22342 34428
rect 24210 34416 24216 34428
rect 24268 34416 24274 34468
rect 26234 34416 26240 34468
rect 26292 34416 26298 34468
rect 28966 34456 28994 34496
rect 29730 34484 29736 34496
rect 29788 34484 29794 34536
rect 30392 34524 30420 34555
rect 32030 34552 32036 34564
rect 32088 34552 32094 34604
rect 32125 34595 32183 34601
rect 32125 34561 32137 34595
rect 32171 34561 32183 34595
rect 32125 34555 32183 34561
rect 30300 34496 30420 34524
rect 31297 34527 31355 34533
rect 30300 34456 30328 34496
rect 31297 34493 31309 34527
rect 31343 34524 31355 34527
rect 32140 34524 32168 34555
rect 32306 34552 32312 34604
rect 32364 34552 32370 34604
rect 33888 34601 33916 34632
rect 33873 34595 33931 34601
rect 33873 34561 33885 34595
rect 33919 34561 33931 34595
rect 33873 34555 33931 34561
rect 34425 34595 34483 34601
rect 34425 34561 34437 34595
rect 34471 34592 34483 34595
rect 34514 34592 34520 34604
rect 34471 34564 34520 34592
rect 34471 34561 34483 34564
rect 34425 34555 34483 34561
rect 34514 34552 34520 34564
rect 34572 34552 34578 34604
rect 34606 34552 34612 34604
rect 34664 34552 34670 34604
rect 34698 34552 34704 34604
rect 34756 34552 34762 34604
rect 34790 34552 34796 34604
rect 34848 34552 34854 34604
rect 34882 34552 34888 34604
rect 34940 34592 34946 34604
rect 35084 34592 35112 34632
rect 34940 34564 35112 34592
rect 35161 34595 35219 34601
rect 34940 34552 34946 34564
rect 35161 34561 35173 34595
rect 35207 34561 35219 34595
rect 35161 34555 35219 34561
rect 34057 34527 34115 34533
rect 34057 34524 34069 34527
rect 31343 34496 32168 34524
rect 32232 34496 34069 34524
rect 31343 34493 31355 34496
rect 31297 34487 31355 34493
rect 28966 34428 30328 34456
rect 31202 34416 31208 34468
rect 31260 34456 31266 34468
rect 31573 34459 31631 34465
rect 31573 34456 31585 34459
rect 31260 34428 31585 34456
rect 31260 34416 31266 34428
rect 31573 34425 31585 34428
rect 31619 34425 31631 34459
rect 32232 34456 32260 34496
rect 34057 34493 34069 34496
rect 34103 34493 34115 34527
rect 34624 34524 34652 34552
rect 34057 34487 34115 34493
rect 34532 34496 34652 34524
rect 34808 34524 34836 34552
rect 35176 34524 35204 34555
rect 35526 34552 35532 34604
rect 35584 34552 35590 34604
rect 35636 34601 35664 34632
rect 35621 34595 35679 34601
rect 35621 34561 35633 34595
rect 35667 34561 35679 34595
rect 35621 34555 35679 34561
rect 34808 34496 35204 34524
rect 31573 34419 31631 34425
rect 31726 34428 32260 34456
rect 13504 34360 14320 34388
rect 13504 34348 13510 34360
rect 14550 34348 14556 34400
rect 14608 34348 14614 34400
rect 14642 34348 14648 34400
rect 14700 34388 14706 34400
rect 14921 34391 14979 34397
rect 14921 34388 14933 34391
rect 14700 34360 14933 34388
rect 14700 34348 14706 34360
rect 14921 34357 14933 34360
rect 14967 34357 14979 34391
rect 14921 34351 14979 34357
rect 16666 34348 16672 34400
rect 16724 34348 16730 34400
rect 17034 34348 17040 34400
rect 17092 34348 17098 34400
rect 17129 34391 17187 34397
rect 17129 34357 17141 34391
rect 17175 34388 17187 34391
rect 17954 34388 17960 34400
rect 17175 34360 17960 34388
rect 17175 34357 17187 34360
rect 17129 34351 17187 34357
rect 17954 34348 17960 34360
rect 18012 34348 18018 34400
rect 18966 34348 18972 34400
rect 19024 34348 19030 34400
rect 19518 34348 19524 34400
rect 19576 34388 19582 34400
rect 20070 34388 20076 34400
rect 19576 34360 20076 34388
rect 19576 34348 19582 34360
rect 20070 34348 20076 34360
rect 20128 34388 20134 34400
rect 21174 34388 21180 34400
rect 20128 34360 21180 34388
rect 20128 34348 20134 34360
rect 21174 34348 21180 34360
rect 21232 34348 21238 34400
rect 21269 34391 21327 34397
rect 21269 34357 21281 34391
rect 21315 34388 21327 34391
rect 26326 34388 26332 34400
rect 21315 34360 26332 34388
rect 21315 34357 21327 34360
rect 21269 34351 21327 34357
rect 26326 34348 26332 34360
rect 26384 34348 26390 34400
rect 26418 34348 26424 34400
rect 26476 34388 26482 34400
rect 31726 34388 31754 34428
rect 26476 34360 31754 34388
rect 26476 34348 26482 34360
rect 34422 34348 34428 34400
rect 34480 34388 34486 34400
rect 34532 34397 34560 34496
rect 34606 34416 34612 34468
rect 34664 34456 34670 34468
rect 35805 34459 35863 34465
rect 35805 34456 35817 34459
rect 34664 34428 35817 34456
rect 34664 34416 34670 34428
rect 35805 34425 35817 34428
rect 35851 34425 35863 34459
rect 35805 34419 35863 34425
rect 34517 34391 34575 34397
rect 34517 34388 34529 34391
rect 34480 34360 34529 34388
rect 34480 34348 34486 34360
rect 34517 34357 34529 34360
rect 34563 34357 34575 34391
rect 34517 34351 34575 34357
rect 34698 34348 34704 34400
rect 34756 34388 34762 34400
rect 35342 34388 35348 34400
rect 34756 34360 35348 34388
rect 34756 34348 34762 34360
rect 35342 34348 35348 34360
rect 35400 34348 35406 34400
rect 1104 34298 41400 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 41400 34298
rect 1104 34224 41400 34246
rect 9674 34144 9680 34196
rect 9732 34184 9738 34196
rect 14090 34184 14096 34196
rect 9732 34156 12296 34184
rect 9732 34144 9738 34156
rect 7926 34076 7932 34128
rect 7984 34076 7990 34128
rect 8754 34076 8760 34128
rect 8812 34116 8818 34128
rect 9398 34116 9404 34128
rect 8812 34088 9404 34116
rect 8812 34076 8818 34088
rect 9398 34076 9404 34088
rect 9456 34076 9462 34128
rect 10226 34116 10232 34128
rect 9646 34088 10232 34116
rect 9401 33983 9459 33989
rect 9401 33949 9413 33983
rect 9447 33949 9459 33983
rect 9401 33943 9459 33949
rect 9549 33983 9607 33989
rect 9549 33949 9561 33983
rect 9595 33980 9607 33983
rect 9646 33980 9674 34088
rect 10226 34076 10232 34088
rect 10284 34116 10290 34128
rect 10778 34116 10784 34128
rect 10284 34088 10784 34116
rect 10284 34076 10290 34088
rect 10778 34076 10784 34088
rect 10836 34076 10842 34128
rect 11146 34076 11152 34128
rect 11204 34076 11210 34128
rect 12066 34116 12072 34128
rect 11716 34088 12072 34116
rect 9950 34048 9956 34060
rect 9784 34020 9956 34048
rect 9784 33989 9812 34020
rect 9950 34008 9956 34020
rect 10008 34008 10014 34060
rect 11716 34057 11744 34088
rect 12066 34076 12072 34088
rect 12124 34076 12130 34128
rect 11701 34051 11759 34057
rect 11701 34048 11713 34051
rect 10520 34020 11713 34048
rect 10520 33992 10548 34020
rect 11701 34017 11713 34020
rect 11747 34017 11759 34051
rect 11701 34011 11759 34017
rect 11793 34051 11851 34057
rect 11793 34017 11805 34051
rect 11839 34048 11851 34051
rect 11882 34048 11888 34060
rect 11839 34020 11888 34048
rect 11839 34017 11851 34020
rect 11793 34011 11851 34017
rect 11882 34008 11888 34020
rect 11940 34008 11946 34060
rect 9595 33952 9674 33980
rect 9769 33983 9827 33989
rect 9595 33949 9607 33952
rect 9549 33943 9607 33949
rect 9769 33949 9781 33983
rect 9815 33949 9827 33983
rect 9769 33943 9827 33949
rect 7561 33915 7619 33921
rect 7561 33881 7573 33915
rect 7607 33912 7619 33915
rect 8202 33912 8208 33924
rect 7607 33884 8208 33912
rect 7607 33881 7619 33884
rect 7561 33875 7619 33881
rect 8202 33872 8208 33884
rect 8260 33872 8266 33924
rect 9416 33912 9444 33943
rect 9858 33940 9864 33992
rect 9916 33989 9922 33992
rect 9916 33980 9924 33989
rect 9916 33952 9961 33980
rect 9916 33943 9924 33952
rect 9916 33940 9922 33943
rect 10502 33940 10508 33992
rect 10560 33940 10566 33992
rect 10870 33940 10876 33992
rect 10928 33940 10934 33992
rect 11330 33983 11388 33989
rect 11330 33949 11342 33983
rect 11376 33980 11388 33983
rect 11606 33980 11612 33992
rect 11376 33952 11612 33980
rect 11376 33949 11388 33952
rect 11330 33943 11388 33949
rect 11606 33940 11612 33952
rect 11664 33940 11670 33992
rect 12268 33980 12296 34156
rect 13556 34156 14096 34184
rect 12342 34076 12348 34128
rect 12400 34116 12406 34128
rect 13556 34125 13584 34156
rect 14090 34144 14096 34156
rect 14148 34184 14154 34196
rect 14734 34184 14740 34196
rect 14148 34156 14740 34184
rect 14148 34144 14154 34156
rect 14734 34144 14740 34156
rect 14792 34144 14798 34196
rect 17034 34144 17040 34196
rect 17092 34144 17098 34196
rect 18598 34144 18604 34196
rect 18656 34184 18662 34196
rect 20809 34187 20867 34193
rect 20809 34184 20821 34187
rect 18656 34156 19564 34184
rect 18656 34144 18662 34156
rect 13541 34119 13599 34125
rect 13541 34116 13553 34119
rect 12400 34088 13553 34116
rect 12400 34076 12406 34088
rect 13541 34085 13553 34088
rect 13587 34085 13599 34119
rect 13541 34079 13599 34085
rect 16868 34088 19288 34116
rect 12713 33983 12771 33989
rect 12713 33980 12725 33983
rect 12268 33952 12725 33980
rect 12713 33949 12725 33952
rect 12759 33980 12771 33983
rect 12986 33980 12992 33992
rect 12759 33952 12992 33980
rect 12759 33949 12771 33952
rect 12713 33943 12771 33949
rect 12986 33940 12992 33952
rect 13044 33940 13050 33992
rect 15289 33983 15347 33989
rect 15289 33980 15301 33983
rect 13096 33952 15301 33980
rect 9677 33915 9735 33921
rect 9416 33884 9536 33912
rect 9508 33856 9536 33884
rect 9677 33881 9689 33915
rect 9723 33912 9735 33915
rect 10318 33912 10324 33924
rect 9723 33884 10324 33912
rect 9723 33881 9735 33884
rect 9677 33875 9735 33881
rect 10318 33872 10324 33884
rect 10376 33872 10382 33924
rect 10888 33912 10916 33940
rect 10888 33884 11744 33912
rect 8018 33804 8024 33856
rect 8076 33804 8082 33856
rect 9490 33804 9496 33856
rect 9548 33804 9554 33856
rect 9950 33804 9956 33856
rect 10008 33844 10014 33856
rect 10045 33847 10103 33853
rect 10045 33844 10057 33847
rect 10008 33816 10057 33844
rect 10008 33804 10014 33816
rect 10045 33813 10057 33816
rect 10091 33813 10103 33847
rect 10045 33807 10103 33813
rect 11054 33804 11060 33856
rect 11112 33844 11118 33856
rect 11333 33847 11391 33853
rect 11333 33844 11345 33847
rect 11112 33816 11345 33844
rect 11112 33804 11118 33816
rect 11333 33813 11345 33816
rect 11379 33813 11391 33847
rect 11716 33844 11744 33884
rect 11882 33872 11888 33924
rect 11940 33912 11946 33924
rect 11977 33915 12035 33921
rect 11977 33912 11989 33915
rect 11940 33884 11989 33912
rect 11940 33872 11946 33884
rect 11977 33881 11989 33884
rect 12023 33912 12035 33915
rect 13096 33912 13124 33952
rect 15289 33949 15301 33952
rect 15335 33980 15347 33983
rect 15470 33980 15476 33992
rect 15335 33952 15476 33980
rect 15335 33949 15347 33952
rect 15289 33943 15347 33949
rect 15470 33940 15476 33952
rect 15528 33940 15534 33992
rect 16868 33989 16896 34088
rect 18966 34008 18972 34060
rect 19024 34008 19030 34060
rect 16853 33983 16911 33989
rect 16853 33980 16865 33983
rect 16224 33952 16865 33980
rect 16224 33924 16252 33952
rect 16853 33949 16865 33952
rect 16899 33949 16911 33983
rect 16853 33943 16911 33949
rect 17034 33940 17040 33992
rect 17092 33980 17098 33992
rect 17589 33983 17647 33989
rect 17589 33980 17601 33983
rect 17092 33952 17601 33980
rect 17092 33940 17098 33952
rect 17589 33949 17601 33952
rect 17635 33949 17647 33983
rect 17589 33943 17647 33949
rect 18417 33983 18475 33989
rect 18417 33949 18429 33983
rect 18463 33949 18475 33983
rect 18417 33943 18475 33949
rect 18509 33983 18567 33989
rect 18509 33949 18521 33983
rect 18555 33980 18567 33983
rect 18693 33983 18751 33989
rect 18555 33952 18644 33980
rect 18555 33949 18567 33952
rect 18509 33943 18567 33949
rect 12023 33884 13124 33912
rect 13265 33915 13323 33921
rect 12023 33881 12035 33884
rect 11977 33875 12035 33881
rect 13265 33881 13277 33915
rect 13311 33912 13323 33915
rect 13814 33912 13820 33924
rect 13311 33884 13820 33912
rect 13311 33881 13323 33884
rect 13265 33875 13323 33881
rect 13814 33872 13820 33884
rect 13872 33872 13878 33924
rect 14093 33915 14151 33921
rect 14093 33881 14105 33915
rect 14139 33912 14151 33915
rect 14182 33912 14188 33924
rect 14139 33884 14188 33912
rect 14139 33881 14151 33884
rect 14093 33875 14151 33881
rect 14182 33872 14188 33884
rect 14240 33872 14246 33924
rect 14277 33915 14335 33921
rect 14277 33881 14289 33915
rect 14323 33912 14335 33915
rect 14366 33912 14372 33924
rect 14323 33884 14372 33912
rect 14323 33881 14335 33884
rect 14277 33875 14335 33881
rect 14366 33872 14372 33884
rect 14424 33912 14430 33924
rect 15565 33915 15623 33921
rect 14424 33884 15516 33912
rect 14424 33872 14430 33884
rect 12066 33844 12072 33856
rect 11716 33816 12072 33844
rect 11333 33807 11391 33813
rect 12066 33804 12072 33816
rect 12124 33804 12130 33856
rect 12710 33804 12716 33856
rect 12768 33844 12774 33856
rect 12805 33847 12863 33853
rect 12805 33844 12817 33847
rect 12768 33816 12817 33844
rect 12768 33804 12774 33816
rect 12805 33813 12817 33816
rect 12851 33813 12863 33847
rect 12805 33807 12863 33813
rect 13630 33804 13636 33856
rect 13688 33844 13694 33856
rect 13998 33844 14004 33856
rect 13688 33816 14004 33844
rect 13688 33804 13694 33816
rect 13998 33804 14004 33816
rect 14056 33844 14062 33856
rect 14461 33847 14519 33853
rect 14461 33844 14473 33847
rect 14056 33816 14473 33844
rect 14056 33804 14062 33816
rect 14461 33813 14473 33816
rect 14507 33813 14519 33847
rect 15488 33844 15516 33884
rect 15565 33881 15577 33915
rect 15611 33912 15623 33915
rect 15746 33912 15752 33924
rect 15611 33884 15752 33912
rect 15611 33881 15623 33884
rect 15565 33875 15623 33881
rect 15746 33872 15752 33884
rect 15804 33872 15810 33924
rect 16114 33872 16120 33924
rect 16172 33872 16178 33924
rect 16206 33872 16212 33924
rect 16264 33872 16270 33924
rect 16669 33915 16727 33921
rect 16669 33881 16681 33915
rect 16715 33912 16727 33915
rect 16758 33912 16764 33924
rect 16715 33884 16764 33912
rect 16715 33881 16727 33884
rect 16669 33875 16727 33881
rect 16758 33872 16764 33884
rect 16816 33872 16822 33924
rect 18233 33915 18291 33921
rect 18233 33912 18245 33915
rect 16960 33884 18245 33912
rect 16132 33844 16160 33872
rect 15488 33816 16160 33844
rect 14461 33807 14519 33813
rect 16574 33804 16580 33856
rect 16632 33844 16638 33856
rect 16960 33844 16988 33884
rect 18233 33881 18245 33884
rect 18279 33881 18291 33915
rect 18432 33912 18460 33943
rect 18432 33884 18552 33912
rect 18233 33875 18291 33881
rect 18524 33856 18552 33884
rect 18616 33856 18644 33952
rect 18693 33949 18705 33983
rect 18739 33949 18751 33983
rect 18693 33943 18751 33949
rect 18785 33983 18843 33989
rect 18785 33949 18797 33983
rect 18831 33980 18843 33983
rect 18984 33980 19012 34008
rect 19260 33992 19288 34088
rect 19426 34008 19432 34060
rect 19484 34008 19490 34060
rect 18831 33952 19012 33980
rect 18831 33949 18843 33952
rect 18785 33943 18843 33949
rect 18708 33856 18736 33943
rect 19242 33940 19248 33992
rect 19300 33940 19306 33992
rect 19444 33921 19472 34008
rect 19536 33989 19564 34156
rect 20272 34156 20821 34184
rect 20272 34048 20300 34156
rect 20809 34153 20821 34156
rect 20855 34153 20867 34187
rect 20809 34147 20867 34153
rect 21634 34144 21640 34196
rect 21692 34184 21698 34196
rect 21729 34187 21787 34193
rect 21729 34184 21741 34187
rect 21692 34156 21741 34184
rect 21692 34144 21698 34156
rect 21729 34153 21741 34156
rect 21775 34153 21787 34187
rect 21729 34147 21787 34153
rect 22922 34144 22928 34196
rect 22980 34184 22986 34196
rect 23382 34184 23388 34196
rect 22980 34156 23388 34184
rect 22980 34144 22986 34156
rect 23382 34144 23388 34156
rect 23440 34144 23446 34196
rect 24302 34144 24308 34196
rect 24360 34184 24366 34196
rect 25038 34184 25044 34196
rect 24360 34156 25044 34184
rect 24360 34144 24366 34156
rect 25038 34144 25044 34156
rect 25096 34144 25102 34196
rect 25130 34144 25136 34196
rect 25188 34184 25194 34196
rect 25317 34187 25375 34193
rect 25317 34184 25329 34187
rect 25188 34156 25329 34184
rect 25188 34144 25194 34156
rect 25317 34153 25329 34156
rect 25363 34153 25375 34187
rect 30650 34184 30656 34196
rect 25317 34147 25375 34153
rect 28966 34156 30656 34184
rect 21450 34116 21456 34128
rect 21284 34088 21456 34116
rect 20088 34020 20300 34048
rect 19521 33983 19579 33989
rect 19521 33949 19533 33983
rect 19567 33949 19579 33983
rect 19521 33943 19579 33949
rect 19429 33915 19487 33921
rect 19429 33881 19441 33915
rect 19475 33881 19487 33915
rect 19536 33912 19564 33943
rect 19610 33940 19616 33992
rect 19668 33940 19674 33992
rect 20088 33989 20116 34020
rect 20714 34008 20720 34060
rect 20772 34048 20778 34060
rect 21284 34057 21312 34088
rect 21450 34076 21456 34088
rect 21508 34116 21514 34128
rect 28442 34116 28448 34128
rect 21508 34088 23612 34116
rect 21508 34076 21514 34088
rect 23584 34060 23612 34088
rect 25332 34088 28448 34116
rect 21269 34051 21327 34057
rect 20772 34020 21036 34048
rect 20772 34008 20778 34020
rect 20073 33983 20131 33989
rect 20073 33949 20085 33983
rect 20119 33949 20131 33983
rect 20073 33943 20131 33949
rect 20162 33940 20168 33992
rect 20220 33980 20226 33992
rect 21008 33989 21036 34020
rect 21269 34017 21281 34051
rect 21315 34017 21327 34051
rect 21269 34011 21327 34017
rect 21744 34020 22324 34048
rect 20579 33983 20637 33989
rect 20220 33952 20265 33980
rect 20220 33940 20226 33952
rect 20579 33949 20591 33983
rect 20625 33980 20637 33983
rect 20993 33983 21051 33989
rect 20625 33952 20944 33980
rect 20625 33949 20637 33952
rect 20579 33943 20637 33949
rect 19536 33884 20300 33912
rect 19429 33875 19487 33881
rect 16632 33816 16988 33844
rect 16632 33804 16638 33816
rect 17034 33804 17040 33856
rect 17092 33844 17098 33856
rect 17678 33844 17684 33856
rect 17092 33816 17684 33844
rect 17092 33804 17098 33816
rect 17678 33804 17684 33816
rect 17736 33804 17742 33856
rect 18506 33804 18512 33856
rect 18564 33804 18570 33856
rect 18598 33804 18604 33856
rect 18656 33804 18662 33856
rect 18690 33804 18696 33856
rect 18748 33844 18754 33856
rect 19797 33847 19855 33853
rect 19797 33844 19809 33847
rect 18748 33816 19809 33844
rect 18748 33804 18754 33816
rect 19797 33813 19809 33816
rect 19843 33813 19855 33847
rect 19797 33807 19855 33813
rect 19978 33804 19984 33856
rect 20036 33844 20042 33856
rect 20162 33844 20168 33856
rect 20036 33816 20168 33844
rect 20036 33804 20042 33816
rect 20162 33804 20168 33816
rect 20220 33804 20226 33856
rect 20272 33844 20300 33884
rect 20346 33872 20352 33924
rect 20404 33872 20410 33924
rect 20441 33915 20499 33921
rect 20441 33881 20453 33915
rect 20487 33881 20499 33915
rect 20916 33912 20944 33952
rect 20993 33949 21005 33983
rect 21039 33949 21051 33983
rect 20993 33943 21051 33949
rect 21174 33940 21180 33992
rect 21232 33940 21238 33992
rect 21744 33989 21772 34020
rect 22296 33992 22324 34020
rect 23290 34008 23296 34060
rect 23348 34048 23354 34060
rect 23348 34020 23520 34048
rect 23348 34008 23354 34020
rect 21729 33983 21787 33989
rect 21729 33949 21741 33983
rect 21775 33949 21787 33983
rect 21729 33943 21787 33949
rect 21913 33983 21971 33989
rect 21913 33949 21925 33983
rect 21959 33980 21971 33983
rect 22094 33980 22100 33992
rect 21959 33952 22100 33980
rect 21959 33949 21971 33952
rect 21913 33943 21971 33949
rect 22094 33940 22100 33952
rect 22152 33940 22158 33992
rect 22278 33940 22284 33992
rect 22336 33940 22342 33992
rect 22830 33940 22836 33992
rect 22888 33940 22894 33992
rect 22925 33983 22983 33989
rect 22925 33949 22937 33983
rect 22971 33949 22983 33983
rect 22925 33943 22983 33949
rect 23109 33983 23167 33989
rect 23109 33949 23121 33983
rect 23155 33980 23167 33983
rect 23382 33980 23388 33992
rect 23155 33952 23388 33980
rect 23155 33949 23167 33952
rect 23109 33943 23167 33949
rect 22646 33912 22652 33924
rect 20916 33884 22652 33912
rect 20441 33875 20499 33881
rect 20456 33844 20484 33875
rect 22646 33872 22652 33884
rect 22704 33912 22710 33924
rect 22848 33912 22876 33940
rect 22704 33884 22876 33912
rect 22940 33912 22968 33943
rect 23382 33940 23388 33952
rect 23440 33940 23446 33992
rect 23492 33980 23520 34020
rect 23566 34008 23572 34060
rect 23624 34008 23630 34060
rect 24412 34020 25176 34048
rect 24412 33980 24440 34020
rect 25148 33989 25176 34020
rect 24949 33983 25007 33989
rect 24949 33980 24961 33983
rect 23492 33952 24440 33980
rect 24504 33952 24961 33980
rect 23934 33912 23940 33924
rect 22940 33884 23940 33912
rect 22704 33872 22710 33884
rect 23934 33872 23940 33884
rect 23992 33912 23998 33924
rect 24118 33912 24124 33924
rect 23992 33884 24124 33912
rect 23992 33872 23998 33884
rect 24118 33872 24124 33884
rect 24176 33872 24182 33924
rect 20272 33816 20484 33844
rect 20714 33804 20720 33856
rect 20772 33804 20778 33856
rect 23014 33804 23020 33856
rect 23072 33844 23078 33856
rect 24504 33844 24532 33952
rect 24949 33949 24961 33952
rect 24995 33949 25007 33983
rect 24949 33943 25007 33949
rect 25133 33983 25191 33989
rect 25133 33949 25145 33983
rect 25179 33949 25191 33983
rect 25133 33943 25191 33949
rect 24964 33912 24992 33943
rect 25332 33912 25360 34088
rect 28442 34076 28448 34088
rect 28500 34116 28506 34128
rect 28966 34116 28994 34156
rect 30650 34144 30656 34156
rect 30708 34144 30714 34196
rect 31570 34144 31576 34196
rect 31628 34184 31634 34196
rect 31757 34187 31815 34193
rect 31757 34184 31769 34187
rect 31628 34156 31769 34184
rect 31628 34144 31634 34156
rect 31757 34153 31769 34156
rect 31803 34153 31815 34187
rect 31757 34147 31815 34153
rect 34238 34144 34244 34196
rect 34296 34144 34302 34196
rect 34330 34144 34336 34196
rect 34388 34144 34394 34196
rect 35161 34187 35219 34193
rect 35161 34153 35173 34187
rect 35207 34184 35219 34187
rect 35342 34184 35348 34196
rect 35207 34156 35348 34184
rect 35207 34153 35219 34156
rect 35161 34147 35219 34153
rect 35342 34144 35348 34156
rect 35400 34144 35406 34196
rect 28500 34088 28994 34116
rect 28500 34076 28506 34088
rect 27614 34048 27620 34060
rect 25608 34020 27620 34048
rect 25409 33983 25467 33989
rect 25409 33949 25421 33983
rect 25455 33949 25467 33983
rect 25409 33943 25467 33949
rect 24964 33884 25360 33912
rect 25424 33912 25452 33943
rect 25498 33940 25504 33992
rect 25556 33980 25562 33992
rect 25608 33989 25636 34020
rect 27614 34008 27620 34020
rect 27672 34008 27678 34060
rect 30190 34008 30196 34060
rect 30248 34048 30254 34060
rect 33689 34051 33747 34057
rect 33689 34048 33701 34051
rect 30248 34020 33701 34048
rect 30248 34008 30254 34020
rect 33689 34017 33701 34020
rect 33735 34017 33747 34051
rect 34348 34048 34376 34144
rect 34514 34076 34520 34128
rect 34572 34116 34578 34128
rect 34572 34088 35020 34116
rect 34572 34076 34578 34088
rect 34992 34048 35020 34088
rect 35069 34051 35127 34057
rect 35069 34048 35081 34051
rect 34348 34020 34744 34048
rect 34992 34020 35081 34048
rect 33689 34011 33747 34017
rect 34716 33992 34744 34020
rect 35069 34017 35081 34020
rect 35115 34048 35127 34051
rect 35526 34048 35532 34060
rect 35115 34020 35532 34048
rect 35115 34017 35127 34020
rect 35069 34011 35127 34017
rect 35526 34008 35532 34020
rect 35584 34008 35590 34060
rect 25593 33983 25651 33989
rect 25593 33980 25605 33983
rect 25556 33952 25605 33980
rect 25556 33940 25562 33952
rect 25593 33949 25605 33952
rect 25639 33949 25651 33983
rect 25593 33943 25651 33949
rect 26326 33940 26332 33992
rect 26384 33980 26390 33992
rect 28718 33980 28724 33992
rect 26384 33952 28724 33980
rect 26384 33940 26390 33952
rect 28718 33940 28724 33952
rect 28776 33980 28782 33992
rect 30098 33980 30104 33992
rect 28776 33952 30104 33980
rect 28776 33940 28782 33952
rect 30098 33940 30104 33952
rect 30156 33940 30162 33992
rect 31757 33983 31815 33989
rect 31757 33949 31769 33983
rect 31803 33980 31815 33983
rect 31941 33983 31999 33989
rect 31803 33952 31837 33980
rect 31803 33949 31815 33952
rect 31757 33943 31815 33949
rect 31941 33949 31953 33983
rect 31987 33980 31999 33983
rect 32306 33980 32312 33992
rect 31987 33952 32312 33980
rect 31987 33949 31999 33952
rect 31941 33943 31999 33949
rect 26234 33912 26240 33924
rect 25424 33884 26240 33912
rect 26234 33872 26240 33884
rect 26292 33912 26298 33924
rect 26694 33912 26700 33924
rect 26292 33884 26700 33912
rect 26292 33872 26298 33884
rect 26694 33872 26700 33884
rect 26752 33872 26758 33924
rect 27522 33872 27528 33924
rect 27580 33912 27586 33924
rect 28258 33912 28264 33924
rect 27580 33884 28264 33912
rect 27580 33872 27586 33884
rect 28258 33872 28264 33884
rect 28316 33912 28322 33924
rect 31772 33912 31800 33943
rect 31846 33912 31852 33924
rect 28316 33884 31852 33912
rect 28316 33872 28322 33884
rect 31846 33872 31852 33884
rect 31904 33872 31910 33924
rect 23072 33816 24532 33844
rect 23072 33804 23078 33816
rect 24578 33804 24584 33856
rect 24636 33844 24642 33856
rect 25501 33847 25559 33853
rect 25501 33844 25513 33847
rect 24636 33816 25513 33844
rect 24636 33804 24642 33816
rect 25501 33813 25513 33816
rect 25547 33813 25559 33847
rect 25501 33807 25559 33813
rect 27062 33804 27068 33856
rect 27120 33844 27126 33856
rect 31956 33844 31984 33943
rect 32306 33940 32312 33952
rect 32364 33940 32370 33992
rect 33505 33983 33563 33989
rect 33505 33949 33517 33983
rect 33551 33949 33563 33983
rect 34606 33980 34612 33992
rect 33505 33943 33563 33949
rect 34348 33952 34612 33980
rect 27120 33816 31984 33844
rect 33520 33844 33548 33943
rect 34149 33915 34207 33921
rect 34149 33881 34161 33915
rect 34195 33912 34207 33915
rect 34348 33912 34376 33952
rect 34606 33940 34612 33952
rect 34664 33940 34670 33992
rect 34698 33940 34704 33992
rect 34756 33940 34762 33992
rect 34790 33940 34796 33992
rect 34848 33940 34854 33992
rect 35161 33983 35219 33989
rect 35161 33980 35173 33983
rect 35084 33952 35173 33980
rect 34195 33884 34376 33912
rect 34808 33912 34836 33940
rect 35084 33912 35112 33952
rect 35161 33949 35173 33952
rect 35207 33949 35219 33983
rect 35161 33943 35219 33949
rect 34808 33884 35112 33912
rect 34195 33881 34207 33884
rect 34149 33875 34207 33881
rect 35345 33847 35403 33853
rect 35345 33844 35357 33847
rect 33520 33816 35357 33844
rect 27120 33804 27126 33816
rect 35345 33813 35357 33816
rect 35391 33813 35403 33847
rect 35345 33807 35403 33813
rect 1104 33754 41400 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 41400 33754
rect 1104 33680 41400 33702
rect 8018 33600 8024 33652
rect 8076 33600 8082 33652
rect 9582 33600 9588 33652
rect 9640 33600 9646 33652
rect 11330 33600 11336 33652
rect 11388 33640 11394 33652
rect 11882 33640 11888 33652
rect 11388 33612 11888 33640
rect 11388 33600 11394 33612
rect 11882 33600 11888 33612
rect 11940 33600 11946 33652
rect 12618 33600 12624 33652
rect 12676 33600 12682 33652
rect 13449 33643 13507 33649
rect 13449 33609 13461 33643
rect 13495 33640 13507 33643
rect 14366 33640 14372 33652
rect 13495 33612 14372 33640
rect 13495 33609 13507 33612
rect 13449 33603 13507 33609
rect 14366 33600 14372 33612
rect 14424 33600 14430 33652
rect 16666 33640 16672 33652
rect 15948 33612 16672 33640
rect 7098 33532 7104 33584
rect 7156 33532 7162 33584
rect 8036 33572 8064 33600
rect 8757 33575 8815 33581
rect 8757 33572 8769 33575
rect 8036 33544 8769 33572
rect 8757 33541 8769 33544
rect 8803 33541 8815 33575
rect 10137 33575 10195 33581
rect 10137 33572 10149 33575
rect 8757 33535 8815 33541
rect 9600 33544 10149 33572
rect 8202 33464 8208 33516
rect 8260 33464 8266 33516
rect 9490 33513 9496 33516
rect 9447 33507 9496 33513
rect 9447 33473 9459 33507
rect 9493 33473 9496 33507
rect 9447 33467 9496 33473
rect 9490 33464 9496 33467
rect 9548 33504 9554 33516
rect 9600 33504 9628 33544
rect 10137 33541 10149 33544
rect 10183 33541 10195 33575
rect 12066 33572 12072 33584
rect 10137 33535 10195 33541
rect 11440 33544 12072 33572
rect 9548 33476 9628 33504
rect 9677 33507 9735 33513
rect 9548 33464 9554 33476
rect 9677 33473 9689 33507
rect 9723 33504 9735 33507
rect 9858 33504 9864 33516
rect 9723 33476 9864 33504
rect 9723 33473 9735 33476
rect 9677 33467 9735 33473
rect 5994 33396 6000 33448
rect 6052 33436 6058 33448
rect 6365 33439 6423 33445
rect 6365 33436 6377 33439
rect 6052 33408 6377 33436
rect 6052 33396 6058 33408
rect 6365 33405 6377 33408
rect 6411 33405 6423 33439
rect 6365 33399 6423 33405
rect 6730 33396 6736 33448
rect 6788 33396 6794 33448
rect 9033 33439 9091 33445
rect 9033 33405 9045 33439
rect 9079 33436 9091 33439
rect 9214 33436 9220 33448
rect 9079 33408 9220 33436
rect 9079 33405 9091 33408
rect 9033 33399 9091 33405
rect 9214 33396 9220 33408
rect 9272 33436 9278 33448
rect 9692 33436 9720 33467
rect 9858 33464 9864 33476
rect 9916 33464 9922 33516
rect 9953 33507 10011 33513
rect 9953 33473 9965 33507
rect 9999 33504 10011 33507
rect 11440 33504 11468 33544
rect 12066 33532 12072 33544
rect 12124 33532 12130 33584
rect 12636 33572 12664 33600
rect 15948 33581 15976 33612
rect 16666 33600 16672 33612
rect 16724 33600 16730 33652
rect 17678 33600 17684 33652
rect 17736 33640 17742 33652
rect 18414 33640 18420 33652
rect 17736 33612 18420 33640
rect 17736 33600 17742 33612
rect 18414 33600 18420 33612
rect 18472 33600 18478 33652
rect 18877 33643 18935 33649
rect 18877 33609 18889 33643
rect 18923 33640 18935 33643
rect 19978 33640 19984 33652
rect 18923 33612 19984 33640
rect 18923 33609 18935 33612
rect 18877 33603 18935 33609
rect 13173 33575 13231 33581
rect 13173 33572 13185 33575
rect 12636 33544 13185 33572
rect 13173 33541 13185 33544
rect 13219 33541 13231 33575
rect 15933 33575 15991 33581
rect 13173 33535 13231 33541
rect 13648 33544 14228 33572
rect 9999 33476 11468 33504
rect 9999 33473 10011 33476
rect 9953 33467 10011 33473
rect 11514 33464 11520 33516
rect 11572 33464 11578 33516
rect 11606 33464 11612 33516
rect 11664 33504 11670 33516
rect 12621 33507 12679 33513
rect 11664 33476 12572 33504
rect 11664 33464 11670 33476
rect 12544 33448 12572 33476
rect 12621 33473 12633 33507
rect 12667 33504 12679 33507
rect 13648 33504 13676 33544
rect 14200 33516 14228 33544
rect 15488 33544 15792 33572
rect 12667 33476 13676 33504
rect 12667 33473 12679 33476
rect 12621 33467 12679 33473
rect 13906 33464 13912 33516
rect 13964 33504 13970 33516
rect 14001 33507 14059 33513
rect 14001 33504 14013 33507
rect 13964 33476 14013 33504
rect 13964 33464 13970 33476
rect 14001 33473 14013 33476
rect 14047 33473 14059 33507
rect 14001 33467 14059 33473
rect 14182 33464 14188 33516
rect 14240 33464 14246 33516
rect 15010 33464 15016 33516
rect 15068 33464 15074 33516
rect 15488 33513 15516 33544
rect 15473 33507 15531 33513
rect 15473 33473 15485 33507
rect 15519 33473 15531 33507
rect 15473 33467 15531 33473
rect 15657 33507 15715 33513
rect 15657 33473 15669 33507
rect 15703 33473 15715 33507
rect 15657 33467 15715 33473
rect 9272 33408 9720 33436
rect 9769 33439 9827 33445
rect 9272 33396 9278 33408
rect 9769 33405 9781 33439
rect 9815 33436 9827 33439
rect 11330 33436 11336 33448
rect 9815 33408 11336 33436
rect 9815 33405 9827 33408
rect 9769 33399 9827 33405
rect 9876 33380 9904 33408
rect 11330 33396 11336 33408
rect 11388 33396 11394 33448
rect 11793 33439 11851 33445
rect 11793 33405 11805 33439
rect 11839 33405 11851 33439
rect 11793 33399 11851 33405
rect 9858 33328 9864 33380
rect 9916 33328 9922 33380
rect 11808 33368 11836 33399
rect 12526 33396 12532 33448
rect 12584 33396 12590 33448
rect 12713 33439 12771 33445
rect 12713 33405 12725 33439
rect 12759 33436 12771 33439
rect 13538 33436 13544 33448
rect 12759 33408 13544 33436
rect 12759 33405 12771 33408
rect 12713 33399 12771 33405
rect 13538 33396 13544 33408
rect 13596 33396 13602 33448
rect 14093 33439 14151 33445
rect 14093 33405 14105 33439
rect 14139 33436 14151 33439
rect 15028 33436 15056 33464
rect 14139 33408 15056 33436
rect 14139 33405 14151 33408
rect 14093 33399 14151 33405
rect 11624 33340 11836 33368
rect 12989 33371 13047 33377
rect 9030 33260 9036 33312
rect 9088 33300 9094 33312
rect 9217 33303 9275 33309
rect 9217 33300 9229 33303
rect 9088 33272 9229 33300
rect 9088 33260 9094 33272
rect 9217 33269 9229 33272
rect 9263 33300 9275 33303
rect 11054 33300 11060 33312
rect 9263 33272 11060 33300
rect 9263 33269 9275 33272
rect 9217 33263 9275 33269
rect 11054 33260 11060 33272
rect 11112 33300 11118 33312
rect 11624 33300 11652 33340
rect 12989 33337 13001 33371
rect 13035 33368 13047 33371
rect 14550 33368 14556 33380
rect 13035 33340 14556 33368
rect 13035 33337 13047 33340
rect 12989 33331 13047 33337
rect 14550 33328 14556 33340
rect 14608 33328 14614 33380
rect 15672 33368 15700 33467
rect 15764 33436 15792 33544
rect 15933 33541 15945 33575
rect 15979 33541 15991 33575
rect 16390 33572 16396 33584
rect 15933 33535 15991 33541
rect 16224 33544 16396 33572
rect 16224 33513 16252 33544
rect 16390 33532 16396 33544
rect 16448 33532 16454 33584
rect 18892 33572 18920 33603
rect 19978 33600 19984 33612
rect 20036 33600 20042 33652
rect 21358 33640 21364 33652
rect 20272 33612 21364 33640
rect 19058 33572 19064 33584
rect 17328 33544 19064 33572
rect 17328 33516 17356 33544
rect 19058 33532 19064 33544
rect 19116 33532 19122 33584
rect 19242 33532 19248 33584
rect 19300 33572 19306 33584
rect 20162 33572 20168 33584
rect 19300 33544 20168 33572
rect 19300 33532 19306 33544
rect 20162 33532 20168 33544
rect 20220 33532 20226 33584
rect 16209 33507 16267 33513
rect 16209 33473 16221 33507
rect 16255 33473 16267 33507
rect 16209 33467 16267 33473
rect 17310 33464 17316 33516
rect 17368 33464 17374 33516
rect 18690 33464 18696 33516
rect 18748 33464 18754 33516
rect 18969 33507 19027 33513
rect 18969 33473 18981 33507
rect 19015 33504 19027 33507
rect 20272 33504 20300 33612
rect 21358 33600 21364 33612
rect 21416 33600 21422 33652
rect 22738 33600 22744 33652
rect 22796 33640 22802 33652
rect 22796 33612 23244 33640
rect 22796 33600 22802 33612
rect 23216 33584 23244 33612
rect 23474 33600 23480 33652
rect 23532 33600 23538 33652
rect 23937 33643 23995 33649
rect 23937 33609 23949 33643
rect 23983 33640 23995 33643
rect 24026 33640 24032 33652
rect 23983 33612 24032 33640
rect 23983 33609 23995 33612
rect 23937 33603 23995 33609
rect 24026 33600 24032 33612
rect 24084 33600 24090 33652
rect 24136 33612 26464 33640
rect 20346 33532 20352 33584
rect 20404 33572 20410 33584
rect 21726 33572 21732 33584
rect 20404 33544 20852 33572
rect 20404 33532 20410 33544
rect 19015 33476 20300 33504
rect 19015 33473 19027 33476
rect 18969 33467 19027 33473
rect 16117 33439 16175 33445
rect 16117 33436 16129 33439
rect 15764 33408 16129 33436
rect 16117 33405 16129 33408
rect 16163 33436 16175 33439
rect 18233 33439 18291 33445
rect 18233 33436 18245 33439
rect 16163 33408 18245 33436
rect 16163 33405 16175 33408
rect 16117 33399 16175 33405
rect 18233 33405 18245 33408
rect 18279 33405 18291 33439
rect 18233 33399 18291 33405
rect 18506 33396 18512 33448
rect 18564 33436 18570 33448
rect 18984 33436 19012 33467
rect 20530 33464 20536 33516
rect 20588 33504 20594 33516
rect 20625 33507 20683 33513
rect 20625 33504 20637 33507
rect 20588 33476 20637 33504
rect 20588 33464 20594 33476
rect 20625 33473 20637 33476
rect 20671 33473 20683 33507
rect 20625 33467 20683 33473
rect 20714 33464 20720 33516
rect 20772 33464 20778 33516
rect 18564 33408 19012 33436
rect 18564 33396 18570 33408
rect 20732 33368 20760 33464
rect 20824 33445 20852 33544
rect 21652 33544 21732 33572
rect 20898 33464 20904 33516
rect 20956 33464 20962 33516
rect 21082 33464 21088 33516
rect 21140 33504 21146 33516
rect 21652 33504 21680 33544
rect 21726 33532 21732 33544
rect 21784 33572 21790 33584
rect 21913 33575 21971 33581
rect 21913 33572 21925 33575
rect 21784 33544 21925 33572
rect 21784 33532 21790 33544
rect 21913 33541 21925 33544
rect 21959 33541 21971 33575
rect 21913 33535 21971 33541
rect 23014 33532 23020 33584
rect 23072 33532 23078 33584
rect 23198 33532 23204 33584
rect 23256 33572 23262 33584
rect 24136 33572 24164 33612
rect 23256 33544 24164 33572
rect 23256 33532 23262 33544
rect 21140 33476 21680 33504
rect 21821 33507 21879 33513
rect 21140 33464 21146 33476
rect 21821 33473 21833 33507
rect 21867 33473 21879 33507
rect 21821 33467 21879 33473
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33504 22063 33507
rect 22094 33504 22100 33516
rect 22051 33476 22100 33504
rect 22051 33473 22063 33476
rect 22005 33467 22063 33473
rect 20809 33439 20867 33445
rect 20809 33405 20821 33439
rect 20855 33436 20867 33439
rect 21542 33436 21548 33448
rect 20855 33408 21548 33436
rect 20855 33405 20867 33408
rect 20809 33399 20867 33405
rect 21542 33396 21548 33408
rect 21600 33396 21606 33448
rect 21836 33436 21864 33467
rect 22094 33464 22100 33476
rect 22152 33464 22158 33516
rect 22189 33507 22247 33513
rect 22189 33473 22201 33507
rect 22235 33504 22247 33507
rect 22373 33507 22431 33513
rect 22235 33476 22324 33504
rect 22235 33473 22247 33476
rect 22189 33467 22247 33473
rect 22296 33448 22324 33476
rect 22373 33473 22385 33507
rect 22419 33473 22431 33507
rect 22373 33467 22431 33473
rect 22278 33436 22284 33448
rect 21836 33408 22284 33436
rect 22278 33396 22284 33408
rect 22336 33396 22342 33448
rect 22388 33436 22416 33467
rect 22554 33464 22560 33516
rect 22612 33464 22618 33516
rect 22833 33507 22891 33513
rect 22833 33473 22845 33507
rect 22879 33504 22891 33507
rect 23106 33504 23112 33516
rect 22879 33476 23112 33504
rect 22879 33473 22891 33476
rect 22833 33467 22891 33473
rect 23106 33464 23112 33476
rect 23164 33464 23170 33516
rect 23768 33513 23796 33544
rect 24302 33532 24308 33584
rect 24360 33532 24366 33584
rect 25424 33544 25912 33572
rect 23569 33507 23627 33513
rect 23569 33473 23581 33507
rect 23615 33473 23627 33507
rect 23569 33467 23627 33473
rect 23753 33507 23811 33513
rect 23753 33473 23765 33507
rect 23799 33473 23811 33507
rect 23753 33467 23811 33473
rect 23845 33507 23903 33513
rect 23845 33473 23857 33507
rect 23891 33504 23903 33507
rect 23934 33504 23940 33516
rect 23891 33476 23940 33504
rect 23891 33473 23903 33476
rect 23845 33467 23903 33473
rect 23382 33436 23388 33448
rect 22388 33408 23388 33436
rect 23382 33396 23388 33408
rect 23440 33436 23446 33448
rect 23584 33436 23612 33467
rect 23934 33464 23940 33476
rect 23992 33464 23998 33516
rect 24029 33507 24087 33513
rect 24029 33473 24041 33507
rect 24075 33473 24087 33507
rect 24029 33467 24087 33473
rect 24044 33436 24072 33467
rect 24210 33464 24216 33516
rect 24268 33464 24274 33516
rect 23440 33408 23888 33436
rect 23440 33396 23446 33408
rect 15672 33340 20760 33368
rect 16224 33312 16252 33340
rect 21266 33328 21272 33380
rect 21324 33328 21330 33380
rect 21634 33328 21640 33380
rect 21692 33368 21698 33380
rect 22373 33371 22431 33377
rect 22373 33368 22385 33371
rect 21692 33340 22385 33368
rect 21692 33328 21698 33340
rect 22373 33337 22385 33340
rect 22419 33337 22431 33371
rect 22373 33331 22431 33337
rect 22833 33371 22891 33377
rect 22833 33337 22845 33371
rect 22879 33337 22891 33371
rect 22833 33331 22891 33337
rect 11112 33272 11652 33300
rect 11112 33260 11118 33272
rect 11698 33260 11704 33312
rect 11756 33260 11762 33312
rect 12342 33260 12348 33312
rect 12400 33300 12406 33312
rect 12621 33303 12679 33309
rect 12621 33300 12633 33303
rect 12400 33272 12633 33300
rect 12400 33260 12406 33272
rect 12621 33269 12633 33272
rect 12667 33269 12679 33303
rect 12621 33263 12679 33269
rect 13998 33260 14004 33312
rect 14056 33260 14062 33312
rect 14366 33260 14372 33312
rect 14424 33260 14430 33312
rect 15286 33260 15292 33312
rect 15344 33300 15350 33312
rect 15841 33303 15899 33309
rect 15841 33300 15853 33303
rect 15344 33272 15853 33300
rect 15344 33260 15350 33272
rect 15841 33269 15853 33272
rect 15887 33269 15899 33303
rect 15841 33263 15899 33269
rect 16206 33260 16212 33312
rect 16264 33260 16270 33312
rect 16298 33260 16304 33312
rect 16356 33300 16362 33312
rect 16393 33303 16451 33309
rect 16393 33300 16405 33303
rect 16356 33272 16405 33300
rect 16356 33260 16362 33272
rect 16393 33269 16405 33272
rect 16439 33269 16451 33303
rect 16393 33263 16451 33269
rect 18506 33260 18512 33312
rect 18564 33260 18570 33312
rect 18601 33303 18659 33309
rect 18601 33269 18613 33303
rect 18647 33300 18659 33303
rect 18966 33300 18972 33312
rect 18647 33272 18972 33300
rect 18647 33269 18659 33272
rect 18601 33263 18659 33269
rect 18966 33260 18972 33272
rect 19024 33260 19030 33312
rect 20806 33260 20812 33312
rect 20864 33260 20870 33312
rect 21082 33260 21088 33312
rect 21140 33260 21146 33312
rect 21284 33300 21312 33328
rect 22848 33300 22876 33331
rect 23014 33328 23020 33380
rect 23072 33368 23078 33380
rect 23290 33368 23296 33380
rect 23072 33340 23296 33368
rect 23072 33328 23078 33340
rect 23290 33328 23296 33340
rect 23348 33328 23354 33380
rect 23569 33371 23627 33377
rect 23569 33337 23581 33371
rect 23615 33368 23627 33371
rect 23750 33368 23756 33380
rect 23615 33340 23756 33368
rect 23615 33337 23627 33340
rect 23569 33331 23627 33337
rect 21284 33272 22876 33300
rect 22922 33260 22928 33312
rect 22980 33300 22986 33312
rect 23584 33300 23612 33331
rect 23750 33328 23756 33340
rect 23808 33328 23814 33380
rect 22980 33272 23612 33300
rect 23860 33300 23888 33408
rect 23952 33408 24072 33436
rect 24320 33436 24348 33532
rect 24394 33464 24400 33516
rect 24452 33464 24458 33516
rect 24489 33513 24547 33519
rect 24489 33479 24501 33513
rect 24535 33479 24547 33513
rect 24489 33473 24547 33479
rect 24504 33436 24532 33473
rect 24854 33464 24860 33516
rect 24912 33504 24918 33516
rect 24949 33507 25007 33513
rect 24949 33504 24961 33507
rect 24912 33476 24961 33504
rect 24912 33464 24918 33476
rect 24949 33473 24961 33476
rect 24995 33473 25007 33507
rect 24949 33467 25007 33473
rect 25130 33464 25136 33516
rect 25188 33464 25194 33516
rect 25314 33464 25320 33516
rect 25372 33464 25378 33516
rect 24320 33408 24532 33436
rect 23952 33380 23980 33408
rect 24578 33396 24584 33448
rect 24636 33396 24642 33448
rect 23934 33328 23940 33380
rect 23992 33368 23998 33380
rect 25424 33368 25452 33544
rect 25590 33464 25596 33516
rect 25648 33504 25654 33516
rect 25774 33504 25780 33516
rect 25648 33476 25780 33504
rect 25648 33464 25654 33476
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 25884 33513 25912 33544
rect 26234 33532 26240 33584
rect 26292 33532 26298 33584
rect 26436 33516 26464 33612
rect 26602 33600 26608 33652
rect 26660 33640 26666 33652
rect 26697 33643 26755 33649
rect 26697 33640 26709 33643
rect 26660 33612 26709 33640
rect 26660 33600 26666 33612
rect 26697 33609 26709 33612
rect 26743 33609 26755 33643
rect 26697 33603 26755 33609
rect 26786 33600 26792 33652
rect 26844 33640 26850 33652
rect 27065 33643 27123 33649
rect 27065 33640 27077 33643
rect 26844 33612 27077 33640
rect 26844 33600 26850 33612
rect 27065 33609 27077 33612
rect 27111 33640 27123 33643
rect 27154 33640 27160 33652
rect 27111 33612 27160 33640
rect 27111 33609 27123 33612
rect 27065 33603 27123 33609
rect 27154 33600 27160 33612
rect 27212 33600 27218 33652
rect 28166 33600 28172 33652
rect 28224 33600 28230 33652
rect 29365 33643 29423 33649
rect 29365 33640 29377 33643
rect 28276 33612 29377 33640
rect 26878 33532 26884 33584
rect 26936 33572 26942 33584
rect 28276 33572 28304 33612
rect 29365 33609 29377 33612
rect 29411 33609 29423 33643
rect 29365 33603 29423 33609
rect 34701 33643 34759 33649
rect 34701 33609 34713 33643
rect 34747 33609 34759 33643
rect 34701 33603 34759 33609
rect 26936 33544 28304 33572
rect 28368 33544 31616 33572
rect 26936 33532 26942 33544
rect 25869 33507 25927 33513
rect 25869 33473 25881 33507
rect 25915 33473 25927 33507
rect 25869 33467 25927 33473
rect 25501 33439 25559 33445
rect 25501 33405 25513 33439
rect 25547 33436 25559 33439
rect 25682 33436 25688 33448
rect 25547 33408 25688 33436
rect 25547 33405 25559 33408
rect 25501 33399 25559 33405
rect 25682 33396 25688 33408
rect 25740 33396 25746 33448
rect 25884 33436 25912 33467
rect 25958 33464 25964 33516
rect 26016 33504 26022 33516
rect 26053 33507 26111 33513
rect 26053 33504 26065 33507
rect 26016 33476 26065 33504
rect 26016 33464 26022 33476
rect 26053 33473 26065 33476
rect 26099 33473 26111 33507
rect 26053 33467 26111 33473
rect 26418 33464 26424 33516
rect 26476 33504 26482 33516
rect 26605 33507 26663 33513
rect 26605 33504 26617 33507
rect 26476 33476 26617 33504
rect 26476 33464 26482 33476
rect 26605 33473 26617 33476
rect 26651 33473 26663 33507
rect 26605 33467 26663 33473
rect 26789 33507 26847 33513
rect 26789 33473 26801 33507
rect 26835 33473 26847 33507
rect 26789 33467 26847 33473
rect 26804 33436 26832 33467
rect 27062 33464 27068 33516
rect 27120 33464 27126 33516
rect 27154 33464 27160 33516
rect 27212 33464 27218 33516
rect 27433 33507 27491 33513
rect 27433 33473 27445 33507
rect 27479 33504 27491 33507
rect 27522 33504 27528 33516
rect 27479 33476 27528 33504
rect 27479 33473 27491 33476
rect 27433 33467 27491 33473
rect 27522 33464 27528 33476
rect 27580 33464 27586 33516
rect 27617 33507 27675 33513
rect 27617 33473 27629 33507
rect 27663 33473 27675 33507
rect 27617 33467 27675 33473
rect 27632 33436 27660 33467
rect 27982 33464 27988 33516
rect 28040 33504 28046 33516
rect 28077 33507 28135 33513
rect 28077 33504 28089 33507
rect 28040 33476 28089 33504
rect 28040 33464 28046 33476
rect 28077 33473 28089 33476
rect 28123 33473 28135 33507
rect 28077 33467 28135 33473
rect 28258 33464 28264 33516
rect 28316 33464 28322 33516
rect 27798 33436 27804 33448
rect 25884 33408 27804 33436
rect 27798 33396 27804 33408
rect 27856 33396 27862 33448
rect 23992 33340 25452 33368
rect 25608 33340 26648 33368
rect 23992 33328 23998 33340
rect 24394 33300 24400 33312
rect 23860 33272 24400 33300
rect 22980 33260 22986 33272
rect 24394 33260 24400 33272
rect 24452 33260 24458 33312
rect 24486 33260 24492 33312
rect 24544 33260 24550 33312
rect 24854 33260 24860 33312
rect 24912 33260 24918 33312
rect 24946 33260 24952 33312
rect 25004 33300 25010 33312
rect 25314 33300 25320 33312
rect 25004 33272 25320 33300
rect 25004 33260 25010 33272
rect 25314 33260 25320 33272
rect 25372 33260 25378 33312
rect 25608 33309 25636 33340
rect 26620 33312 26648 33340
rect 27154 33328 27160 33380
rect 27212 33368 27218 33380
rect 28368 33368 28396 33544
rect 28534 33464 28540 33516
rect 28592 33504 28598 33516
rect 28902 33504 28908 33516
rect 28592 33476 28908 33504
rect 28592 33464 28598 33476
rect 28902 33464 28908 33476
rect 28960 33464 28966 33516
rect 29221 33507 29279 33513
rect 29221 33473 29233 33507
rect 29267 33504 29279 33507
rect 29537 33507 29595 33513
rect 29267 33476 29500 33504
rect 29267 33473 29279 33476
rect 29221 33467 29279 33473
rect 28997 33439 29055 33445
rect 28997 33405 29009 33439
rect 29043 33405 29055 33439
rect 29472 33436 29500 33476
rect 29537 33473 29549 33507
rect 29583 33504 29595 33507
rect 29656 33504 29684 33544
rect 29583 33476 29684 33504
rect 29733 33507 29791 33513
rect 29583 33473 29595 33476
rect 29537 33467 29595 33473
rect 29733 33473 29745 33507
rect 29779 33504 29791 33507
rect 30006 33504 30012 33516
rect 29779 33476 30012 33504
rect 29779 33473 29791 33476
rect 29733 33467 29791 33473
rect 30006 33464 30012 33476
rect 30064 33464 30070 33516
rect 30282 33464 30288 33516
rect 30340 33464 30346 33516
rect 31389 33507 31447 33513
rect 31389 33473 31401 33507
rect 31435 33504 31447 33507
rect 31478 33504 31484 33516
rect 31435 33476 31484 33504
rect 31435 33473 31447 33476
rect 31389 33467 31447 33473
rect 31478 33464 31484 33476
rect 31536 33464 31542 33516
rect 31588 33504 31616 33544
rect 31846 33532 31852 33584
rect 31904 33572 31910 33584
rect 33410 33572 33416 33584
rect 31904 33544 33416 33572
rect 31904 33532 31910 33544
rect 33410 33532 33416 33544
rect 33468 33572 33474 33584
rect 34716 33572 34744 33603
rect 33468 33544 34744 33572
rect 35161 33575 35219 33581
rect 33468 33532 33474 33544
rect 35161 33541 35173 33575
rect 35207 33572 35219 33575
rect 35342 33572 35348 33584
rect 35207 33544 35348 33572
rect 35207 33541 35219 33544
rect 35161 33535 35219 33541
rect 35342 33532 35348 33544
rect 35400 33532 35406 33584
rect 34238 33504 34244 33516
rect 31588 33476 34244 33504
rect 34238 33464 34244 33476
rect 34296 33464 34302 33516
rect 34606 33464 34612 33516
rect 34664 33464 34670 33516
rect 35437 33507 35495 33513
rect 35437 33473 35449 33507
rect 35483 33504 35495 33507
rect 35526 33504 35532 33516
rect 35483 33476 35532 33504
rect 35483 33473 35495 33476
rect 35437 33467 35495 33473
rect 35526 33464 35532 33476
rect 35584 33464 35590 33516
rect 30300 33436 30328 33464
rect 29472 33408 30328 33436
rect 28997 33399 29055 33405
rect 27212 33340 28396 33368
rect 29012 33368 29040 33399
rect 30650 33396 30656 33448
rect 30708 33436 30714 33448
rect 31570 33436 31576 33448
rect 30708 33408 31576 33436
rect 30708 33396 30714 33408
rect 31570 33396 31576 33408
rect 31628 33396 31634 33448
rect 29270 33368 29276 33380
rect 29012 33340 29276 33368
rect 27212 33328 27218 33340
rect 29270 33328 29276 33340
rect 29328 33328 29334 33380
rect 25593 33303 25651 33309
rect 25593 33269 25605 33303
rect 25639 33269 25651 33303
rect 25593 33263 25651 33269
rect 25774 33260 25780 33312
rect 25832 33260 25838 33312
rect 26602 33260 26608 33312
rect 26660 33260 26666 33312
rect 27430 33260 27436 33312
rect 27488 33300 27494 33312
rect 28626 33300 28632 33312
rect 27488 33272 28632 33300
rect 27488 33260 27494 33272
rect 28626 33260 28632 33272
rect 28684 33260 28690 33312
rect 29181 33303 29239 33309
rect 29181 33269 29193 33303
rect 29227 33300 29239 33303
rect 29546 33300 29552 33312
rect 29227 33272 29552 33300
rect 29227 33269 29239 33272
rect 29181 33263 29239 33269
rect 29546 33260 29552 33272
rect 29604 33260 29610 33312
rect 34790 33260 34796 33312
rect 34848 33300 34854 33312
rect 35253 33303 35311 33309
rect 35253 33300 35265 33303
rect 34848 33272 35265 33300
rect 34848 33260 34854 33272
rect 35253 33269 35265 33272
rect 35299 33269 35311 33303
rect 35253 33263 35311 33269
rect 35618 33260 35624 33312
rect 35676 33260 35682 33312
rect 1104 33210 41400 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 41400 33210
rect 1104 33136 41400 33158
rect 5537 33099 5595 33105
rect 5537 33065 5549 33099
rect 5583 33096 5595 33099
rect 6730 33096 6736 33108
rect 5583 33068 6736 33096
rect 5583 33065 5595 33068
rect 5537 33059 5595 33065
rect 6730 33056 6736 33068
rect 6788 33056 6794 33108
rect 8113 33099 8171 33105
rect 8113 33065 8125 33099
rect 8159 33096 8171 33099
rect 8294 33096 8300 33108
rect 8159 33068 8300 33096
rect 8159 33065 8171 33068
rect 8113 33059 8171 33065
rect 8294 33056 8300 33068
rect 8352 33056 8358 33108
rect 13538 33096 13544 33108
rect 13101 33068 13544 33096
rect 6825 33031 6883 33037
rect 6825 33028 6837 33031
rect 5920 33000 6837 33028
rect 5920 32904 5948 33000
rect 6825 32997 6837 33000
rect 6871 32997 6883 33031
rect 13101 33028 13129 33068
rect 13538 33056 13544 33068
rect 13596 33056 13602 33108
rect 13630 33056 13636 33108
rect 13688 33056 13694 33108
rect 13906 33056 13912 33108
rect 13964 33056 13970 33108
rect 14090 33056 14096 33108
rect 14148 33056 14154 33108
rect 15470 33056 15476 33108
rect 15528 33096 15534 33108
rect 17402 33096 17408 33108
rect 15528 33068 17408 33096
rect 15528 33056 15534 33068
rect 17402 33056 17408 33068
rect 17460 33056 17466 33108
rect 17862 33056 17868 33108
rect 17920 33096 17926 33108
rect 18230 33096 18236 33108
rect 17920 33068 18236 33096
rect 17920 33056 17926 33068
rect 18230 33056 18236 33068
rect 18288 33056 18294 33108
rect 18506 33056 18512 33108
rect 18564 33096 18570 33108
rect 18601 33099 18659 33105
rect 18601 33096 18613 33099
rect 18564 33068 18613 33096
rect 18564 33056 18570 33068
rect 18601 33065 18613 33068
rect 18647 33065 18659 33099
rect 18601 33059 18659 33065
rect 21174 33056 21180 33108
rect 21232 33096 21238 33108
rect 21545 33099 21603 33105
rect 21545 33096 21557 33099
rect 21232 33068 21557 33096
rect 21232 33056 21238 33068
rect 21545 33065 21557 33068
rect 21591 33065 21603 33099
rect 21545 33059 21603 33065
rect 6825 32991 6883 32997
rect 8220 33000 13129 33028
rect 13173 33031 13231 33037
rect 5997 32963 6055 32969
rect 5997 32929 6009 32963
rect 6043 32960 6055 32963
rect 7650 32960 7656 32972
rect 6043 32932 7656 32960
rect 6043 32929 6055 32932
rect 5997 32923 6055 32929
rect 7650 32920 7656 32932
rect 7708 32920 7714 32972
rect 5721 32895 5779 32901
rect 5721 32861 5733 32895
rect 5767 32861 5779 32895
rect 5721 32855 5779 32861
rect 5813 32895 5871 32901
rect 5813 32861 5825 32895
rect 5859 32892 5871 32895
rect 5902 32892 5908 32904
rect 5859 32864 5908 32892
rect 5859 32861 5871 32864
rect 5813 32855 5871 32861
rect 5736 32824 5764 32855
rect 5902 32852 5908 32864
rect 5960 32852 5966 32904
rect 6086 32852 6092 32904
rect 6144 32852 6150 32904
rect 6270 32852 6276 32904
rect 6328 32892 6334 32904
rect 8220 32892 8248 33000
rect 13173 32997 13185 33031
rect 13219 33028 13231 33031
rect 13924 33028 13952 33056
rect 13219 33000 13952 33028
rect 14108 33028 14136 33056
rect 14108 33000 14233 33028
rect 13219 32997 13231 33000
rect 13173 32991 13231 32997
rect 8478 32920 8484 32972
rect 8536 32960 8542 32972
rect 8665 32963 8723 32969
rect 8665 32960 8677 32963
rect 8536 32932 8677 32960
rect 8536 32920 8542 32932
rect 8665 32929 8677 32932
rect 8711 32960 8723 32963
rect 8754 32960 8760 32972
rect 8711 32932 8760 32960
rect 8711 32929 8723 32932
rect 8665 32923 8723 32929
rect 8754 32920 8760 32932
rect 8812 32920 8818 32972
rect 13265 32963 13323 32969
rect 13265 32929 13277 32963
rect 13311 32960 13323 32963
rect 14205 32960 14233 33000
rect 15378 32988 15384 33040
rect 15436 33028 15442 33040
rect 15436 33000 18368 33028
rect 15436 32988 15442 33000
rect 18340 32960 18368 33000
rect 20254 32988 20260 33040
rect 20312 33028 20318 33040
rect 21560 33028 21588 33059
rect 21634 33056 21640 33108
rect 21692 33096 21698 33108
rect 22922 33096 22928 33108
rect 21692 33068 22928 33096
rect 21692 33056 21698 33068
rect 22922 33056 22928 33068
rect 22980 33056 22986 33108
rect 23658 33056 23664 33108
rect 23716 33096 23722 33108
rect 27522 33096 27528 33108
rect 23716 33068 24716 33096
rect 23716 33056 23722 33068
rect 24578 33028 24584 33040
rect 20312 33000 21404 33028
rect 21560 33000 24584 33028
rect 20312 32988 20318 33000
rect 21376 32960 21404 33000
rect 24578 32988 24584 33000
rect 24636 32988 24642 33040
rect 24688 33037 24716 33068
rect 24872 33068 27528 33096
rect 24673 33031 24731 33037
rect 24673 32997 24685 33031
rect 24719 32997 24731 33031
rect 24673 32991 24731 32997
rect 13311 32932 14136 32960
rect 14205 32932 14284 32960
rect 13311 32929 13323 32932
rect 13265 32923 13323 32929
rect 6328 32864 8248 32892
rect 6328 32852 6334 32864
rect 8386 32852 8392 32904
rect 8444 32852 8450 32904
rect 11422 32852 11428 32904
rect 11480 32852 11486 32904
rect 13449 32895 13507 32901
rect 11716 32864 13124 32892
rect 6454 32824 6460 32836
rect 5736 32796 6460 32824
rect 6454 32784 6460 32796
rect 6512 32784 6518 32836
rect 7834 32784 7840 32836
rect 7892 32824 7898 32836
rect 8202 32824 8208 32836
rect 7892 32796 8208 32824
rect 7892 32784 7898 32796
rect 8202 32784 8208 32796
rect 8260 32784 8266 32836
rect 8018 32716 8024 32768
rect 8076 32756 8082 32768
rect 8404 32756 8432 32852
rect 8570 32784 8576 32836
rect 8628 32824 8634 32836
rect 8846 32824 8852 32836
rect 8628 32796 8852 32824
rect 8628 32784 8634 32796
rect 8846 32784 8852 32796
rect 8904 32824 8910 32836
rect 11716 32824 11744 32864
rect 8904 32796 11744 32824
rect 12805 32827 12863 32833
rect 8904 32784 8910 32796
rect 12805 32793 12817 32827
rect 12851 32824 12863 32827
rect 12894 32824 12900 32836
rect 12851 32796 12900 32824
rect 12851 32793 12863 32796
rect 12805 32787 12863 32793
rect 12894 32784 12900 32796
rect 12952 32784 12958 32836
rect 12989 32827 13047 32833
rect 12989 32793 13001 32827
rect 13035 32793 13047 32827
rect 13096 32824 13124 32864
rect 13449 32861 13461 32895
rect 13495 32892 13507 32895
rect 13630 32892 13636 32904
rect 13495 32864 13636 32892
rect 13495 32861 13507 32864
rect 13449 32855 13507 32861
rect 13630 32852 13636 32864
rect 13688 32852 13694 32904
rect 14108 32901 14136 32932
rect 14256 32901 14284 32932
rect 18340 32932 20852 32960
rect 13725 32895 13783 32901
rect 13725 32861 13737 32895
rect 13771 32861 13783 32895
rect 13725 32855 13783 32861
rect 14093 32895 14151 32901
rect 14093 32861 14105 32895
rect 14139 32861 14151 32895
rect 14093 32855 14151 32861
rect 14241 32895 14299 32901
rect 14241 32861 14253 32895
rect 14287 32861 14299 32895
rect 14241 32855 14299 32861
rect 13740 32824 13768 32855
rect 14366 32852 14372 32904
rect 14424 32852 14430 32904
rect 14550 32852 14556 32904
rect 14608 32901 14614 32904
rect 14608 32892 14616 32901
rect 14608 32864 14653 32892
rect 14608 32855 14616 32864
rect 14608 32852 14614 32855
rect 15194 32852 15200 32904
rect 15252 32852 15258 32904
rect 16022 32852 16028 32904
rect 16080 32852 16086 32904
rect 16114 32852 16120 32904
rect 16172 32852 16178 32904
rect 16206 32852 16212 32904
rect 16264 32892 16270 32904
rect 16301 32895 16359 32901
rect 16301 32892 16313 32895
rect 16264 32864 16313 32892
rect 16264 32852 16270 32864
rect 16301 32861 16313 32864
rect 16347 32861 16359 32895
rect 16301 32855 16359 32861
rect 16393 32895 16451 32901
rect 16393 32861 16405 32895
rect 16439 32861 16451 32895
rect 16393 32855 16451 32861
rect 14461 32827 14519 32833
rect 14461 32824 14473 32827
rect 13096 32796 13768 32824
rect 13832 32796 14473 32824
rect 12989 32787 13047 32793
rect 8076 32728 8432 32756
rect 8076 32716 8082 32728
rect 8938 32716 8944 32768
rect 8996 32756 9002 32768
rect 10042 32756 10048 32768
rect 8996 32728 10048 32756
rect 8996 32716 9002 32728
rect 10042 32716 10048 32728
rect 10100 32716 10106 32768
rect 11701 32759 11759 32765
rect 11701 32725 11713 32759
rect 11747 32756 11759 32759
rect 11790 32756 11796 32768
rect 11747 32728 11796 32756
rect 11747 32725 11759 32728
rect 11701 32719 11759 32725
rect 11790 32716 11796 32728
rect 11848 32716 11854 32768
rect 12158 32716 12164 32768
rect 12216 32756 12222 32768
rect 12434 32756 12440 32768
rect 12216 32728 12440 32756
rect 12216 32716 12222 32728
rect 12434 32716 12440 32728
rect 12492 32716 12498 32768
rect 13004 32756 13032 32787
rect 13832 32768 13860 32796
rect 14461 32793 14473 32796
rect 14507 32824 14519 32827
rect 14918 32824 14924 32836
rect 14507 32796 14924 32824
rect 14507 32793 14519 32796
rect 14461 32787 14519 32793
rect 14918 32784 14924 32796
rect 14976 32824 14982 32836
rect 15212 32824 15240 32852
rect 14976 32796 15240 32824
rect 14976 32784 14982 32796
rect 15930 32784 15936 32836
rect 15988 32824 15994 32836
rect 16408 32824 16436 32855
rect 17034 32852 17040 32904
rect 17092 32892 17098 32904
rect 17678 32892 17684 32904
rect 17092 32864 17684 32892
rect 17092 32852 17098 32864
rect 17678 32852 17684 32864
rect 17736 32892 17742 32904
rect 18340 32901 18368 32932
rect 18049 32895 18107 32901
rect 18049 32892 18061 32895
rect 17736 32864 18061 32892
rect 17736 32852 17742 32864
rect 18049 32861 18061 32864
rect 18095 32861 18107 32895
rect 18049 32855 18107 32861
rect 18233 32895 18291 32901
rect 18233 32861 18245 32895
rect 18279 32861 18291 32895
rect 18233 32855 18291 32861
rect 18325 32895 18383 32901
rect 18325 32861 18337 32895
rect 18371 32861 18383 32895
rect 18325 32855 18383 32861
rect 18248 32824 18276 32855
rect 18414 32852 18420 32904
rect 18472 32892 18478 32904
rect 18966 32892 18972 32904
rect 18472 32864 18972 32892
rect 18472 32852 18478 32864
rect 18966 32852 18972 32864
rect 19024 32852 19030 32904
rect 19518 32852 19524 32904
rect 19576 32852 19582 32904
rect 15988 32796 16436 32824
rect 16868 32796 18276 32824
rect 15988 32784 15994 32796
rect 13354 32756 13360 32768
rect 13004 32728 13360 32756
rect 13354 32716 13360 32728
rect 13412 32716 13418 32768
rect 13814 32716 13820 32768
rect 13872 32716 13878 32768
rect 14366 32716 14372 32768
rect 14424 32756 14430 32768
rect 14737 32759 14795 32765
rect 14737 32756 14749 32759
rect 14424 32728 14749 32756
rect 14424 32716 14430 32728
rect 14737 32725 14749 32728
rect 14783 32725 14795 32759
rect 14737 32719 14795 32725
rect 15654 32716 15660 32768
rect 15712 32756 15718 32768
rect 15841 32759 15899 32765
rect 15841 32756 15853 32759
rect 15712 32728 15853 32756
rect 15712 32716 15718 32728
rect 15841 32725 15853 32728
rect 15887 32725 15899 32759
rect 15841 32719 15899 32725
rect 16022 32716 16028 32768
rect 16080 32756 16086 32768
rect 16868 32756 16896 32796
rect 16080 32728 16896 32756
rect 16080 32716 16086 32728
rect 16942 32716 16948 32768
rect 17000 32756 17006 32768
rect 17862 32756 17868 32768
rect 17000 32728 17868 32756
rect 17000 32716 17006 32728
rect 17862 32716 17868 32728
rect 17920 32716 17926 32768
rect 18248 32756 18276 32796
rect 18690 32784 18696 32836
rect 18748 32824 18754 32836
rect 19536 32824 19564 32852
rect 18748 32796 19564 32824
rect 18748 32784 18754 32796
rect 20714 32784 20720 32836
rect 20772 32784 20778 32836
rect 20824 32824 20852 32932
rect 21376 32932 24520 32960
rect 21376 32901 21404 32932
rect 21361 32895 21419 32901
rect 21361 32861 21373 32895
rect 21407 32861 21419 32895
rect 21361 32855 21419 32861
rect 21450 32852 21456 32904
rect 21508 32852 21514 32904
rect 21726 32852 21732 32904
rect 21784 32892 21790 32904
rect 22002 32892 22008 32904
rect 21784 32864 22008 32892
rect 21784 32852 21790 32864
rect 22002 32852 22008 32864
rect 22060 32852 22066 32904
rect 22554 32852 22560 32904
rect 22612 32892 22618 32904
rect 24302 32892 24308 32904
rect 22612 32864 24308 32892
rect 22612 32852 22618 32864
rect 24302 32852 24308 32864
rect 24360 32892 24366 32904
rect 24397 32895 24455 32901
rect 24397 32892 24409 32895
rect 24360 32864 24409 32892
rect 24360 32852 24366 32864
rect 24397 32861 24409 32864
rect 24443 32861 24455 32895
rect 24397 32855 24455 32861
rect 20824 32796 21864 32824
rect 20732 32756 20760 32784
rect 18248 32728 20760 32756
rect 21726 32716 21732 32768
rect 21784 32716 21790 32768
rect 21836 32756 21864 32796
rect 22830 32756 22836 32768
rect 21836 32728 22836 32756
rect 22830 32716 22836 32728
rect 22888 32716 22894 32768
rect 24492 32756 24520 32932
rect 24578 32852 24584 32904
rect 24636 32892 24642 32904
rect 24673 32895 24731 32901
rect 24673 32892 24685 32895
rect 24636 32864 24685 32892
rect 24636 32852 24642 32864
rect 24673 32861 24685 32864
rect 24719 32892 24731 32895
rect 24872 32892 24900 33068
rect 27522 33056 27528 33068
rect 27580 33056 27586 33108
rect 27617 33099 27675 33105
rect 27617 33065 27629 33099
rect 27663 33096 27675 33099
rect 28166 33096 28172 33108
rect 27663 33068 28172 33096
rect 27663 33065 27675 33068
rect 27617 33059 27675 33065
rect 28166 33056 28172 33068
rect 28224 33056 28230 33108
rect 28534 33056 28540 33108
rect 28592 33096 28598 33108
rect 30190 33096 30196 33108
rect 28592 33068 30196 33096
rect 28592 33056 28598 33068
rect 30190 33056 30196 33068
rect 30248 33056 30254 33108
rect 30374 33056 30380 33108
rect 30432 33096 30438 33108
rect 31202 33096 31208 33108
rect 30432 33068 31208 33096
rect 30432 33056 30438 33068
rect 31202 33056 31208 33068
rect 31260 33096 31266 33108
rect 31260 33068 31754 33096
rect 31260 33056 31266 33068
rect 27706 33028 27712 33040
rect 25424 33000 27712 33028
rect 24719 32864 24900 32892
rect 24719 32861 24731 32864
rect 24673 32855 24731 32861
rect 24946 32852 24952 32904
rect 25004 32852 25010 32904
rect 25038 32852 25044 32904
rect 25096 32892 25102 32904
rect 25225 32895 25283 32901
rect 25225 32892 25237 32895
rect 25096 32864 25237 32892
rect 25096 32852 25102 32864
rect 25225 32861 25237 32864
rect 25271 32861 25283 32895
rect 25225 32855 25283 32861
rect 25314 32852 25320 32904
rect 25372 32852 25378 32904
rect 25424 32901 25452 33000
rect 27706 32988 27712 33000
rect 27764 33028 27770 33040
rect 27764 33000 28028 33028
rect 27764 32988 27770 33000
rect 27246 32920 27252 32972
rect 27304 32920 27310 32972
rect 27338 32920 27344 32972
rect 27396 32960 27402 32972
rect 27396 32932 27568 32960
rect 27396 32920 27402 32932
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32861 25467 32895
rect 26050 32892 26056 32904
rect 25409 32855 25467 32861
rect 25516 32864 26056 32892
rect 24964 32824 24992 32852
rect 25424 32824 25452 32855
rect 24964 32796 25452 32824
rect 25516 32756 25544 32864
rect 26050 32852 26056 32864
rect 26108 32852 26114 32904
rect 26234 32852 26240 32904
rect 26292 32892 26298 32904
rect 27433 32895 27491 32901
rect 27433 32892 27445 32895
rect 26292 32864 27445 32892
rect 26292 32852 26298 32864
rect 27433 32861 27445 32864
rect 27479 32861 27491 32895
rect 27540 32892 27568 32932
rect 27614 32920 27620 32972
rect 27672 32960 27678 32972
rect 28000 32969 28028 33000
rect 30006 32988 30012 33040
rect 30064 33028 30070 33040
rect 31297 33031 31355 33037
rect 31297 33028 31309 33031
rect 30064 33000 31309 33028
rect 30064 32988 30070 33000
rect 31297 32997 31309 33000
rect 31343 32997 31355 33031
rect 31726 33028 31754 33068
rect 34606 33056 34612 33108
rect 34664 33056 34670 33108
rect 35253 33099 35311 33105
rect 35253 33065 35265 33099
rect 35299 33096 35311 33099
rect 35618 33096 35624 33108
rect 35299 33068 35624 33096
rect 35299 33065 35311 33068
rect 35253 33059 35311 33065
rect 35618 33056 35624 33068
rect 35676 33056 35682 33108
rect 34624 33028 34652 33056
rect 35437 33031 35495 33037
rect 35437 33028 35449 33031
rect 31726 33000 34100 33028
rect 34624 33000 35449 33028
rect 31297 32991 31355 32997
rect 27985 32963 28043 32969
rect 27672 32932 27844 32960
rect 27672 32920 27678 32932
rect 27816 32901 27844 32932
rect 27985 32929 27997 32963
rect 28031 32929 28043 32963
rect 28166 32960 28172 32972
rect 27985 32923 28043 32929
rect 28092 32932 28172 32960
rect 27709 32895 27767 32901
rect 27709 32892 27721 32895
rect 27540 32864 27721 32892
rect 27433 32855 27491 32861
rect 27709 32861 27721 32864
rect 27755 32861 27767 32895
rect 27709 32855 27767 32861
rect 27801 32895 27859 32901
rect 27801 32861 27813 32895
rect 27847 32892 27859 32895
rect 28092 32892 28120 32932
rect 28166 32920 28172 32932
rect 28224 32960 28230 32972
rect 28537 32963 28595 32969
rect 28537 32960 28549 32963
rect 28224 32932 28549 32960
rect 28224 32920 28230 32932
rect 28537 32929 28549 32932
rect 28583 32929 28595 32963
rect 28537 32923 28595 32929
rect 27847 32864 28120 32892
rect 28353 32895 28411 32901
rect 27847 32861 27859 32864
rect 27801 32855 27859 32861
rect 28353 32861 28365 32895
rect 28399 32892 28411 32895
rect 29362 32892 29368 32904
rect 28399 32864 29368 32892
rect 28399 32861 28411 32864
rect 28353 32855 28411 32861
rect 29362 32852 29368 32864
rect 29420 32892 29426 32904
rect 30024 32901 30052 32988
rect 34072 32972 34100 33000
rect 35437 32997 35449 33000
rect 35483 32997 35495 33031
rect 35437 32991 35495 32997
rect 30098 32920 30104 32972
rect 30156 32960 30162 32972
rect 30469 32963 30527 32969
rect 30469 32960 30481 32963
rect 30156 32932 30481 32960
rect 30156 32920 30162 32932
rect 30469 32929 30481 32932
rect 30515 32960 30527 32963
rect 30515 32932 31892 32960
rect 30515 32929 30527 32932
rect 30469 32923 30527 32929
rect 31864 32904 31892 32932
rect 34054 32920 34060 32972
rect 34112 32920 34118 32972
rect 34514 32920 34520 32972
rect 34572 32920 34578 32972
rect 34790 32920 34796 32972
rect 34848 32920 34854 32972
rect 30009 32895 30067 32901
rect 30009 32892 30021 32895
rect 29420 32864 30021 32892
rect 29420 32852 29426 32864
rect 30009 32861 30021 32864
rect 30055 32861 30067 32895
rect 30009 32855 30067 32861
rect 30190 32852 30196 32904
rect 30248 32852 30254 32904
rect 30745 32895 30803 32901
rect 30745 32861 30757 32895
rect 30791 32892 30803 32895
rect 31021 32895 31079 32901
rect 31021 32892 31033 32895
rect 30791 32864 31033 32892
rect 30791 32861 30803 32864
rect 30745 32855 30803 32861
rect 31021 32861 31033 32864
rect 31067 32892 31079 32895
rect 31386 32892 31392 32904
rect 31067 32864 31392 32892
rect 31067 32861 31079 32864
rect 31021 32855 31079 32861
rect 31386 32852 31392 32864
rect 31444 32852 31450 32904
rect 31665 32895 31723 32901
rect 31665 32861 31677 32895
rect 31711 32861 31723 32895
rect 31665 32855 31723 32861
rect 30374 32824 30380 32836
rect 25608 32796 30380 32824
rect 25608 32768 25636 32796
rect 30374 32784 30380 32796
rect 30432 32784 30438 32836
rect 30561 32827 30619 32833
rect 30561 32793 30573 32827
rect 30607 32824 30619 32827
rect 30834 32824 30840 32836
rect 30607 32796 30840 32824
rect 30607 32793 30619 32796
rect 30561 32787 30619 32793
rect 30834 32784 30840 32796
rect 30892 32784 30898 32836
rect 30926 32784 30932 32836
rect 30984 32784 30990 32836
rect 31680 32824 31708 32855
rect 31846 32852 31852 32904
rect 31904 32852 31910 32904
rect 32033 32895 32091 32901
rect 32033 32861 32045 32895
rect 32079 32892 32091 32895
rect 32398 32892 32404 32904
rect 32079 32864 32404 32892
rect 32079 32861 32091 32864
rect 32033 32855 32091 32861
rect 32398 32852 32404 32864
rect 32456 32852 32462 32904
rect 33873 32895 33931 32901
rect 33873 32861 33885 32895
rect 33919 32892 33931 32895
rect 34330 32892 34336 32904
rect 33919 32864 34336 32892
rect 33919 32861 33931 32864
rect 33873 32855 33931 32861
rect 34330 32852 34336 32864
rect 34388 32852 34394 32904
rect 34532 32892 34560 32920
rect 34882 32892 34888 32904
rect 34532 32864 34888 32892
rect 32309 32827 32367 32833
rect 32309 32824 32321 32827
rect 31680 32796 32321 32824
rect 24492 32728 25544 32756
rect 25590 32716 25596 32768
rect 25648 32716 25654 32768
rect 25958 32716 25964 32768
rect 26016 32756 26022 32768
rect 27154 32756 27160 32768
rect 26016 32728 27160 32756
rect 26016 32716 26022 32728
rect 27154 32716 27160 32728
rect 27212 32716 27218 32768
rect 28994 32716 29000 32768
rect 29052 32756 29058 32768
rect 29822 32756 29828 32768
rect 29052 32728 29828 32756
rect 29052 32716 29058 32728
rect 29822 32716 29828 32728
rect 29880 32756 29886 32768
rect 30098 32756 30104 32768
rect 29880 32728 30104 32756
rect 29880 32716 29886 32728
rect 30098 32716 30104 32728
rect 30156 32716 30162 32768
rect 30190 32716 30196 32768
rect 30248 32756 30254 32768
rect 31726 32756 31754 32796
rect 32309 32793 32321 32796
rect 32355 32793 32367 32827
rect 32309 32787 32367 32793
rect 32858 32784 32864 32836
rect 32916 32784 32922 32836
rect 32950 32784 32956 32836
rect 33008 32824 33014 32836
rect 33597 32827 33655 32833
rect 33597 32824 33609 32827
rect 33008 32796 33609 32824
rect 33008 32784 33014 32796
rect 33597 32793 33609 32796
rect 33643 32793 33655 32827
rect 33597 32787 33655 32793
rect 33778 32784 33784 32836
rect 33836 32824 33842 32836
rect 34532 32824 34560 32864
rect 34882 32852 34888 32864
rect 34940 32852 34946 32904
rect 35253 32895 35311 32901
rect 35253 32861 35265 32895
rect 35299 32892 35311 32895
rect 35529 32895 35587 32901
rect 35529 32892 35541 32895
rect 35299 32864 35541 32892
rect 35299 32861 35311 32864
rect 35253 32855 35311 32861
rect 35529 32861 35541 32864
rect 35575 32861 35587 32895
rect 35529 32855 35587 32861
rect 33836 32796 34560 32824
rect 33836 32784 33842 32796
rect 34698 32784 34704 32836
rect 34756 32824 34762 32836
rect 35268 32824 35296 32855
rect 39114 32852 39120 32904
rect 39172 32892 39178 32904
rect 40773 32895 40831 32901
rect 40773 32892 40785 32895
rect 39172 32864 40785 32892
rect 39172 32852 39178 32864
rect 40773 32861 40785 32864
rect 40819 32861 40831 32895
rect 40773 32855 40831 32861
rect 34756 32796 35296 32824
rect 34756 32784 34762 32796
rect 30248 32728 31754 32756
rect 30248 32716 30254 32728
rect 34974 32716 34980 32768
rect 35032 32756 35038 32768
rect 35713 32759 35771 32765
rect 35713 32756 35725 32759
rect 35032 32728 35725 32756
rect 35032 32716 35038 32728
rect 35713 32725 35725 32728
rect 35759 32725 35771 32759
rect 35713 32719 35771 32725
rect 40954 32716 40960 32768
rect 41012 32716 41018 32768
rect 1104 32666 41400 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 41400 32666
rect 1104 32592 41400 32614
rect 5626 32552 5632 32564
rect 1504 32524 5632 32552
rect 1504 32493 1532 32524
rect 5626 32512 5632 32524
rect 5684 32512 5690 32564
rect 6089 32555 6147 32561
rect 6089 32521 6101 32555
rect 6135 32552 6147 32555
rect 6270 32552 6276 32564
rect 6135 32524 6276 32552
rect 6135 32521 6147 32524
rect 6089 32515 6147 32521
rect 6270 32512 6276 32524
rect 6328 32512 6334 32564
rect 6454 32512 6460 32564
rect 6512 32512 6518 32564
rect 8478 32552 8484 32564
rect 7760 32524 8484 32552
rect 1489 32487 1547 32493
rect 1489 32453 1501 32487
rect 1535 32453 1547 32487
rect 7098 32484 7104 32496
rect 5842 32456 7104 32484
rect 1489 32447 1547 32453
rect 7098 32444 7104 32456
rect 7156 32444 7162 32496
rect 6362 32376 6368 32428
rect 6420 32376 6426 32428
rect 7760 32425 7788 32524
rect 8478 32512 8484 32524
rect 8536 32512 8542 32564
rect 8662 32512 8668 32564
rect 8720 32552 8726 32564
rect 9033 32555 9091 32561
rect 9033 32552 9045 32555
rect 8720 32524 9045 32552
rect 8720 32512 8726 32524
rect 9033 32521 9045 32524
rect 9079 32521 9091 32555
rect 9033 32515 9091 32521
rect 9306 32512 9312 32564
rect 9364 32552 9370 32564
rect 10594 32552 10600 32564
rect 9364 32524 10600 32552
rect 9364 32512 9370 32524
rect 10594 32512 10600 32524
rect 10652 32512 10658 32564
rect 12526 32552 12532 32564
rect 12452 32524 12532 32552
rect 10505 32487 10563 32493
rect 7944 32456 8248 32484
rect 7944 32425 7972 32456
rect 8220 32428 8248 32456
rect 8680 32456 9628 32484
rect 7745 32419 7803 32425
rect 7745 32385 7757 32419
rect 7791 32385 7803 32419
rect 7745 32379 7803 32385
rect 7929 32419 7987 32425
rect 7929 32385 7941 32419
rect 7975 32385 7987 32419
rect 7929 32379 7987 32385
rect 8113 32419 8171 32425
rect 8113 32385 8125 32419
rect 8159 32385 8171 32419
rect 8113 32379 8171 32385
rect 4341 32351 4399 32357
rect 4341 32317 4353 32351
rect 4387 32317 4399 32351
rect 4341 32311 4399 32317
rect 4617 32351 4675 32357
rect 4617 32317 4629 32351
rect 4663 32348 4675 32351
rect 6178 32348 6184 32360
rect 4663 32320 6184 32348
rect 4663 32317 4675 32320
rect 4617 32311 4675 32317
rect 934 32172 940 32224
rect 992 32212 998 32224
rect 1581 32215 1639 32221
rect 1581 32212 1593 32215
rect 992 32184 1593 32212
rect 992 32172 998 32184
rect 1581 32181 1593 32184
rect 1627 32181 1639 32215
rect 4356 32212 4384 32311
rect 6178 32308 6184 32320
rect 6236 32308 6242 32360
rect 7837 32351 7895 32357
rect 7837 32317 7849 32351
rect 7883 32348 7895 32351
rect 8128 32348 8156 32379
rect 8202 32376 8208 32428
rect 8260 32376 8266 32428
rect 8297 32419 8355 32425
rect 8297 32385 8309 32419
rect 8343 32416 8355 32419
rect 8343 32388 8524 32416
rect 8343 32385 8355 32388
rect 8297 32379 8355 32385
rect 7883 32320 8156 32348
rect 7883 32317 7895 32320
rect 7837 32311 7895 32317
rect 8128 32224 8156 32320
rect 8496 32224 8524 32388
rect 8570 32376 8576 32428
rect 8628 32376 8634 32428
rect 8680 32348 8708 32456
rect 9600 32425 9628 32456
rect 10505 32453 10517 32487
rect 10551 32484 10563 32487
rect 10551 32456 12020 32484
rect 10551 32453 10563 32456
rect 10505 32447 10563 32453
rect 8757 32419 8815 32425
rect 8757 32385 8769 32419
rect 8803 32416 8815 32419
rect 9125 32419 9183 32425
rect 9125 32416 9137 32419
rect 8803 32388 9137 32416
rect 8803 32385 8815 32388
rect 8757 32379 8815 32385
rect 9125 32385 9137 32388
rect 9171 32385 9183 32419
rect 9125 32379 9183 32385
rect 9309 32419 9367 32425
rect 9309 32385 9321 32419
rect 9355 32385 9367 32419
rect 9309 32379 9367 32385
rect 9585 32419 9643 32425
rect 9585 32385 9597 32419
rect 9631 32416 9643 32419
rect 10689 32419 10747 32425
rect 10689 32416 10701 32419
rect 9631 32388 10701 32416
rect 9631 32385 9643 32388
rect 9585 32379 9643 32385
rect 10689 32385 10701 32388
rect 10735 32385 10747 32419
rect 10689 32379 10747 32385
rect 10781 32419 10839 32425
rect 10781 32385 10793 32419
rect 10827 32385 10839 32419
rect 10781 32379 10839 32385
rect 8588 32320 8708 32348
rect 8588 32292 8616 32320
rect 9030 32308 9036 32360
rect 9088 32308 9094 32360
rect 9324 32348 9352 32379
rect 10134 32348 10140 32360
rect 9232 32320 10140 32348
rect 8570 32240 8576 32292
rect 8628 32240 8634 32292
rect 9122 32240 9128 32292
rect 9180 32280 9186 32292
rect 9232 32280 9260 32320
rect 10134 32308 10140 32320
rect 10192 32308 10198 32360
rect 10594 32308 10600 32360
rect 10652 32348 10658 32360
rect 10796 32348 10824 32379
rect 10870 32376 10876 32428
rect 10928 32416 10934 32428
rect 10965 32419 11023 32425
rect 10965 32416 10977 32419
rect 10928 32388 10977 32416
rect 10928 32376 10934 32388
rect 10965 32385 10977 32388
rect 11011 32385 11023 32419
rect 10965 32379 11023 32385
rect 11054 32376 11060 32428
rect 11112 32376 11118 32428
rect 11606 32376 11612 32428
rect 11664 32416 11670 32428
rect 11701 32419 11759 32425
rect 11701 32416 11713 32419
rect 11664 32388 11713 32416
rect 11664 32376 11670 32388
rect 11701 32385 11713 32388
rect 11747 32385 11759 32419
rect 11701 32379 11759 32385
rect 11882 32376 11888 32428
rect 11940 32376 11946 32428
rect 11992 32425 12020 32456
rect 11977 32419 12035 32425
rect 11977 32385 11989 32419
rect 12023 32385 12035 32419
rect 11977 32379 12035 32385
rect 12158 32376 12164 32428
rect 12216 32376 12222 32428
rect 10652 32320 10824 32348
rect 10652 32308 10658 32320
rect 11146 32308 11152 32360
rect 11204 32348 11210 32360
rect 11624 32348 11652 32376
rect 12176 32348 12204 32376
rect 11204 32320 11652 32348
rect 11716 32320 12204 32348
rect 12452 32348 12480 32524
rect 12526 32512 12532 32524
rect 12584 32512 12590 32564
rect 12894 32512 12900 32564
rect 12952 32512 12958 32564
rect 14369 32555 14427 32561
rect 14369 32521 14381 32555
rect 14415 32552 14427 32555
rect 15841 32555 15899 32561
rect 14415 32524 14780 32552
rect 14415 32521 14427 32524
rect 14369 32515 14427 32521
rect 12912 32484 12940 32512
rect 13265 32487 13323 32493
rect 12544 32456 13032 32484
rect 12544 32428 12572 32456
rect 12526 32376 12532 32428
rect 12584 32376 12590 32428
rect 12621 32419 12679 32425
rect 12621 32385 12633 32419
rect 12667 32385 12679 32419
rect 12621 32379 12679 32385
rect 12713 32419 12771 32425
rect 12713 32385 12725 32419
rect 12759 32385 12771 32419
rect 12713 32379 12771 32385
rect 12636 32348 12664 32379
rect 12452 32320 12664 32348
rect 12728 32348 12756 32379
rect 12894 32376 12900 32428
rect 12952 32376 12958 32428
rect 13004 32416 13032 32456
rect 13265 32453 13277 32487
rect 13311 32484 13323 32487
rect 13538 32484 13544 32496
rect 13311 32456 13544 32484
rect 13311 32453 13323 32456
rect 13265 32447 13323 32453
rect 13538 32444 13544 32456
rect 13596 32444 13602 32496
rect 13633 32487 13691 32493
rect 13633 32453 13645 32487
rect 13679 32484 13691 32487
rect 14001 32487 14059 32493
rect 14001 32484 14013 32487
rect 13679 32456 14013 32484
rect 13679 32453 13691 32456
rect 13633 32447 13691 32453
rect 14001 32453 14013 32456
rect 14047 32453 14059 32487
rect 14550 32484 14556 32496
rect 14001 32447 14059 32453
rect 14108 32456 14556 32484
rect 13449 32419 13507 32425
rect 13449 32416 13461 32419
rect 13004 32388 13461 32416
rect 13449 32385 13461 32388
rect 13495 32385 13507 32419
rect 13725 32419 13783 32425
rect 13725 32416 13737 32419
rect 13449 32379 13507 32385
rect 13556 32388 13737 32416
rect 12728 32320 13216 32348
rect 11204 32308 11210 32320
rect 9180 32252 9260 32280
rect 9180 32240 9186 32252
rect 9306 32240 9312 32292
rect 9364 32280 9370 32292
rect 9401 32283 9459 32289
rect 9401 32280 9413 32283
rect 9364 32252 9413 32280
rect 9364 32240 9370 32252
rect 9401 32249 9413 32252
rect 9447 32249 9459 32283
rect 9401 32243 9459 32249
rect 9490 32240 9496 32292
rect 9548 32280 9554 32292
rect 11716 32280 11744 32320
rect 9548 32252 11744 32280
rect 9548 32240 9554 32252
rect 11882 32240 11888 32292
rect 11940 32280 11946 32292
rect 12452 32280 12480 32320
rect 13188 32292 13216 32320
rect 11940 32252 12480 32280
rect 11940 32240 11946 32252
rect 13170 32240 13176 32292
rect 13228 32240 13234 32292
rect 13464 32280 13492 32379
rect 13556 32360 13584 32388
rect 13725 32385 13737 32388
rect 13771 32385 13783 32419
rect 13725 32379 13783 32385
rect 13814 32376 13820 32428
rect 13872 32416 13878 32428
rect 14108 32425 14136 32456
rect 14550 32444 14556 32456
rect 14608 32444 14614 32496
rect 14752 32493 14780 32524
rect 15841 32521 15853 32555
rect 15887 32552 15899 32555
rect 15930 32552 15936 32564
rect 15887 32524 15936 32552
rect 15887 32521 15899 32524
rect 15841 32515 15899 32521
rect 15930 32512 15936 32524
rect 15988 32512 15994 32564
rect 16390 32512 16396 32564
rect 16448 32512 16454 32564
rect 17310 32512 17316 32564
rect 17368 32512 17374 32564
rect 17954 32512 17960 32564
rect 18012 32552 18018 32564
rect 18509 32555 18567 32561
rect 18509 32552 18521 32555
rect 18012 32524 18521 32552
rect 18012 32512 18018 32524
rect 18509 32521 18521 32524
rect 18555 32552 18567 32555
rect 18555 32524 18920 32552
rect 18555 32521 18567 32524
rect 18509 32515 18567 32521
rect 14737 32487 14795 32493
rect 14737 32453 14749 32487
rect 14783 32453 14795 32487
rect 16408 32484 16436 32512
rect 16669 32487 16727 32493
rect 16669 32484 16681 32487
rect 14737 32447 14795 32453
rect 15028 32456 16681 32484
rect 14093 32419 14151 32425
rect 13872 32388 13917 32416
rect 13872 32376 13878 32388
rect 14093 32385 14105 32419
rect 14139 32385 14151 32419
rect 14093 32379 14151 32385
rect 14182 32376 14188 32428
rect 14240 32425 14246 32428
rect 15028 32425 15056 32456
rect 16669 32453 16681 32456
rect 16715 32453 16727 32487
rect 17328 32484 17356 32512
rect 17328 32456 18000 32484
rect 16669 32447 16727 32453
rect 14240 32379 14248 32425
rect 15013 32419 15071 32425
rect 14384 32388 14964 32416
rect 14240 32376 14246 32379
rect 13538 32308 13544 32360
rect 13596 32308 13602 32360
rect 13814 32280 13820 32292
rect 13464 32252 13820 32280
rect 13814 32240 13820 32252
rect 13872 32240 13878 32292
rect 14090 32240 14096 32292
rect 14148 32280 14154 32292
rect 14384 32280 14412 32388
rect 14826 32308 14832 32360
rect 14884 32308 14890 32360
rect 14936 32348 14964 32388
rect 15013 32385 15025 32419
rect 15059 32385 15071 32419
rect 15013 32379 15071 32385
rect 15289 32419 15347 32425
rect 15289 32385 15301 32419
rect 15335 32416 15347 32419
rect 15378 32416 15384 32428
rect 15335 32388 15384 32416
rect 15335 32385 15347 32388
rect 15289 32379 15347 32385
rect 15378 32376 15384 32388
rect 15436 32376 15442 32428
rect 15473 32419 15531 32425
rect 15473 32385 15485 32419
rect 15519 32385 15531 32419
rect 15473 32379 15531 32385
rect 15488 32348 15516 32379
rect 15562 32376 15568 32428
rect 15620 32376 15626 32428
rect 15657 32419 15715 32425
rect 15657 32385 15669 32419
rect 15703 32416 15715 32419
rect 16022 32416 16028 32428
rect 15703 32388 16028 32416
rect 15703 32385 15715 32388
rect 15657 32379 15715 32385
rect 16022 32376 16028 32388
rect 16080 32376 16086 32428
rect 16117 32419 16175 32425
rect 16117 32385 16129 32419
rect 16163 32385 16175 32419
rect 16117 32379 16175 32385
rect 16209 32419 16267 32425
rect 16209 32385 16221 32419
rect 16255 32416 16267 32419
rect 16298 32416 16304 32428
rect 16255 32388 16304 32416
rect 16255 32385 16267 32388
rect 16209 32379 16267 32385
rect 16132 32348 16160 32379
rect 14936 32320 15516 32348
rect 16040 32320 16160 32348
rect 14148 32252 14412 32280
rect 15028 32252 15332 32280
rect 14148 32240 14154 32252
rect 4614 32212 4620 32224
rect 4356 32184 4620 32212
rect 1581 32175 1639 32181
rect 4614 32172 4620 32184
rect 4672 32212 4678 32224
rect 5994 32212 6000 32224
rect 4672 32184 6000 32212
rect 4672 32172 4678 32184
rect 5994 32172 6000 32184
rect 6052 32172 6058 32224
rect 8110 32172 8116 32224
rect 8168 32172 8174 32224
rect 8478 32172 8484 32224
rect 8536 32212 8542 32224
rect 10410 32212 10416 32224
rect 8536 32184 10416 32212
rect 8536 32172 8542 32184
rect 10410 32172 10416 32184
rect 10468 32172 10474 32224
rect 10778 32172 10784 32224
rect 10836 32212 10842 32224
rect 11054 32212 11060 32224
rect 10836 32184 11060 32212
rect 10836 32172 10842 32184
rect 11054 32172 11060 32184
rect 11112 32172 11118 32224
rect 11514 32172 11520 32224
rect 11572 32172 11578 32224
rect 12250 32172 12256 32224
rect 12308 32172 12314 32224
rect 15028 32221 15056 32252
rect 15304 32224 15332 32252
rect 15013 32215 15071 32221
rect 15013 32181 15025 32215
rect 15059 32181 15071 32215
rect 15013 32175 15071 32181
rect 15194 32172 15200 32224
rect 15252 32172 15258 32224
rect 15286 32172 15292 32224
rect 15344 32172 15350 32224
rect 15930 32172 15936 32224
rect 15988 32172 15994 32224
rect 16040 32212 16068 32320
rect 16114 32240 16120 32292
rect 16172 32280 16178 32292
rect 16224 32280 16252 32379
rect 16298 32376 16304 32388
rect 16356 32376 16362 32428
rect 16390 32376 16396 32428
rect 16448 32376 16454 32428
rect 16485 32419 16543 32425
rect 16485 32385 16497 32419
rect 16531 32416 16543 32419
rect 16850 32416 16856 32428
rect 16531 32388 16856 32416
rect 16531 32385 16543 32388
rect 16485 32379 16543 32385
rect 16850 32376 16856 32388
rect 16908 32416 16914 32428
rect 16945 32419 17003 32425
rect 16945 32416 16957 32419
rect 16908 32388 16957 32416
rect 16908 32376 16914 32388
rect 16945 32385 16957 32388
rect 16991 32385 17003 32419
rect 16945 32379 17003 32385
rect 17405 32419 17463 32425
rect 17405 32385 17417 32419
rect 17451 32385 17463 32419
rect 17405 32379 17463 32385
rect 17681 32419 17739 32425
rect 17681 32385 17693 32419
rect 17727 32385 17739 32419
rect 17681 32379 17739 32385
rect 16408 32348 16436 32376
rect 17037 32351 17095 32357
rect 17037 32348 17049 32351
rect 16408 32320 17049 32348
rect 17037 32317 17049 32320
rect 17083 32317 17095 32351
rect 17420 32348 17448 32379
rect 17037 32311 17095 32317
rect 17144 32320 17448 32348
rect 17144 32280 17172 32320
rect 16172 32252 16252 32280
rect 16592 32252 17172 32280
rect 16172 32240 16178 32252
rect 16592 32212 16620 32252
rect 16040 32184 16620 32212
rect 16666 32172 16672 32224
rect 16724 32212 16730 32224
rect 17129 32215 17187 32221
rect 17129 32212 17141 32215
rect 16724 32184 17141 32212
rect 16724 32172 16730 32184
rect 17129 32181 17141 32184
rect 17175 32181 17187 32215
rect 17420 32212 17448 32320
rect 17494 32308 17500 32360
rect 17552 32308 17558 32360
rect 17586 32308 17592 32360
rect 17644 32348 17650 32360
rect 17696 32348 17724 32379
rect 17862 32376 17868 32428
rect 17920 32376 17926 32428
rect 17972 32425 18000 32456
rect 18138 32444 18144 32496
rect 18196 32444 18202 32496
rect 18414 32484 18420 32496
rect 18248 32456 18420 32484
rect 18248 32425 18276 32456
rect 18414 32444 18420 32456
rect 18472 32444 18478 32496
rect 17957 32419 18015 32425
rect 17957 32385 17969 32419
rect 18003 32385 18015 32419
rect 17957 32379 18015 32385
rect 18233 32419 18291 32425
rect 18233 32385 18245 32419
rect 18279 32385 18291 32419
rect 18233 32379 18291 32385
rect 18325 32419 18383 32425
rect 18325 32385 18337 32419
rect 18371 32416 18383 32419
rect 18598 32416 18604 32428
rect 18371 32388 18604 32416
rect 18371 32385 18383 32388
rect 18325 32379 18383 32385
rect 18598 32376 18604 32388
rect 18656 32376 18662 32428
rect 18690 32348 18696 32360
rect 17644 32320 18696 32348
rect 17644 32308 17650 32320
rect 18690 32308 18696 32320
rect 18748 32308 18754 32360
rect 18892 32280 18920 32524
rect 19242 32512 19248 32564
rect 19300 32552 19306 32564
rect 20165 32555 20223 32561
rect 20165 32552 20177 32555
rect 19300 32524 20177 32552
rect 19300 32512 19306 32524
rect 20165 32521 20177 32524
rect 20211 32521 20223 32555
rect 20165 32515 20223 32521
rect 22002 32512 22008 32564
rect 22060 32512 22066 32564
rect 22094 32512 22100 32564
rect 22152 32512 22158 32564
rect 23014 32512 23020 32564
rect 23072 32552 23078 32564
rect 24210 32552 24216 32564
rect 23072 32524 24216 32552
rect 23072 32512 23078 32524
rect 24210 32512 24216 32524
rect 24268 32552 24274 32564
rect 24268 32524 26464 32552
rect 24268 32512 24274 32524
rect 19153 32487 19211 32493
rect 19153 32453 19165 32487
rect 19199 32484 19211 32487
rect 21542 32484 21548 32496
rect 19199 32456 20024 32484
rect 19199 32453 19211 32456
rect 19153 32447 19211 32453
rect 19337 32419 19395 32425
rect 19337 32385 19349 32419
rect 19383 32416 19395 32419
rect 19426 32416 19432 32428
rect 19383 32388 19432 32416
rect 19383 32385 19395 32388
rect 19337 32379 19395 32385
rect 19426 32376 19432 32388
rect 19484 32376 19490 32428
rect 19996 32425 20024 32456
rect 20456 32456 21548 32484
rect 20456 32425 20484 32456
rect 21542 32444 21548 32456
rect 21600 32444 21606 32496
rect 19705 32419 19763 32425
rect 19705 32385 19717 32419
rect 19751 32416 19763 32419
rect 19981 32419 20039 32425
rect 19751 32388 19932 32416
rect 19751 32385 19763 32388
rect 19705 32379 19763 32385
rect 19610 32308 19616 32360
rect 19668 32308 19674 32360
rect 19797 32351 19855 32357
rect 19797 32317 19809 32351
rect 19843 32317 19855 32351
rect 19904 32348 19932 32388
rect 19981 32385 19993 32419
rect 20027 32385 20039 32419
rect 20441 32419 20499 32425
rect 19981 32379 20039 32385
rect 20088 32388 20392 32416
rect 20088 32348 20116 32388
rect 19904 32320 20116 32348
rect 20257 32351 20315 32357
rect 19797 32311 19855 32317
rect 20257 32317 20269 32351
rect 20303 32317 20315 32351
rect 20364 32348 20392 32388
rect 20441 32385 20453 32419
rect 20487 32385 20499 32419
rect 20441 32379 20499 32385
rect 21174 32376 21180 32428
rect 21232 32416 21238 32428
rect 21634 32416 21640 32428
rect 21232 32388 21640 32416
rect 21232 32376 21238 32388
rect 21634 32376 21640 32388
rect 21692 32416 21698 32428
rect 21821 32419 21879 32425
rect 21821 32416 21833 32419
rect 21692 32388 21833 32416
rect 21692 32376 21698 32388
rect 21821 32385 21833 32388
rect 21867 32385 21879 32419
rect 22020 32416 22048 32512
rect 22112 32484 22140 32512
rect 23566 32484 23572 32496
rect 22112 32456 23572 32484
rect 23566 32444 23572 32456
rect 23624 32484 23630 32496
rect 24305 32487 24363 32493
rect 23624 32456 23980 32484
rect 23624 32444 23630 32456
rect 22097 32419 22155 32425
rect 22097 32416 22109 32419
rect 22020 32388 22109 32416
rect 21821 32379 21879 32385
rect 22097 32385 22109 32388
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 20364 32320 20576 32348
rect 20257 32311 20315 32317
rect 19812 32280 19840 32311
rect 18892 32252 19840 32280
rect 19886 32240 19892 32292
rect 19944 32280 19950 32292
rect 20272 32280 20300 32311
rect 20548 32292 20576 32320
rect 21266 32308 21272 32360
rect 21324 32348 21330 32360
rect 22005 32351 22063 32357
rect 22005 32348 22017 32351
rect 21324 32320 22017 32348
rect 21324 32308 21330 32320
rect 22005 32317 22017 32320
rect 22051 32348 22063 32351
rect 23845 32351 23903 32357
rect 22051 32320 22140 32348
rect 22051 32317 22063 32320
rect 22005 32311 22063 32317
rect 22112 32292 22140 32320
rect 23845 32317 23857 32351
rect 23891 32317 23903 32351
rect 23952 32348 23980 32456
rect 24305 32453 24317 32487
rect 24351 32484 24363 32487
rect 25130 32484 25136 32496
rect 24351 32456 25136 32484
rect 24351 32453 24363 32456
rect 24305 32447 24363 32453
rect 25130 32444 25136 32456
rect 25188 32444 25194 32496
rect 25406 32444 25412 32496
rect 25464 32484 25470 32496
rect 25958 32484 25964 32496
rect 25464 32456 25964 32484
rect 25464 32444 25470 32456
rect 25958 32444 25964 32456
rect 26016 32444 26022 32496
rect 26436 32428 26464 32524
rect 27338 32512 27344 32564
rect 27396 32512 27402 32564
rect 28810 32512 28816 32564
rect 28868 32552 28874 32564
rect 28905 32555 28963 32561
rect 28905 32552 28917 32555
rect 28868 32524 28917 32552
rect 28868 32512 28874 32524
rect 28905 32521 28917 32524
rect 28951 32552 28963 32555
rect 29086 32552 29092 32564
rect 28951 32524 29092 32552
rect 28951 32521 28963 32524
rect 28905 32515 28963 32521
rect 29086 32512 29092 32524
rect 29144 32512 29150 32564
rect 29546 32512 29552 32564
rect 29604 32552 29610 32564
rect 30193 32555 30251 32561
rect 30193 32552 30205 32555
rect 29604 32524 30205 32552
rect 29604 32512 29610 32524
rect 30193 32521 30205 32524
rect 30239 32552 30251 32555
rect 30282 32552 30288 32564
rect 30239 32524 30288 32552
rect 30239 32521 30251 32524
rect 30193 32515 30251 32521
rect 30282 32512 30288 32524
rect 30340 32512 30346 32564
rect 31202 32552 31208 32564
rect 30392 32524 31208 32552
rect 27062 32444 27068 32496
rect 27120 32484 27126 32496
rect 30392 32484 30420 32524
rect 31202 32512 31208 32524
rect 31260 32512 31266 32564
rect 32398 32512 32404 32564
rect 32456 32512 32462 32564
rect 32858 32512 32864 32564
rect 32916 32552 32922 32564
rect 33965 32555 34023 32561
rect 33965 32552 33977 32555
rect 32916 32524 33977 32552
rect 32916 32512 32922 32524
rect 33965 32521 33977 32524
rect 34011 32521 34023 32555
rect 33965 32515 34023 32521
rect 34330 32512 34336 32564
rect 34388 32552 34394 32564
rect 34793 32555 34851 32561
rect 34793 32552 34805 32555
rect 34388 32524 34805 32552
rect 34388 32512 34394 32524
rect 34793 32521 34805 32524
rect 34839 32521 34851 32555
rect 34793 32515 34851 32521
rect 34882 32512 34888 32564
rect 34940 32552 34946 32564
rect 34940 32524 35112 32552
rect 34940 32512 34946 32524
rect 27120 32456 30420 32484
rect 27120 32444 27126 32456
rect 24029 32419 24087 32425
rect 24029 32385 24041 32419
rect 24075 32416 24087 32419
rect 24210 32416 24216 32428
rect 24075 32388 24216 32416
rect 24075 32385 24087 32388
rect 24029 32379 24087 32385
rect 24210 32376 24216 32388
rect 24268 32416 24274 32428
rect 24762 32416 24768 32428
rect 24268 32388 24768 32416
rect 24268 32376 24274 32388
rect 24762 32376 24768 32388
rect 24820 32416 24826 32428
rect 24820 32388 26372 32416
rect 24820 32376 24826 32388
rect 24397 32351 24455 32357
rect 24397 32348 24409 32351
rect 23952 32320 24409 32348
rect 23845 32311 23903 32317
rect 24397 32317 24409 32320
rect 24443 32348 24455 32351
rect 24946 32348 24952 32360
rect 24443 32320 24952 32348
rect 24443 32317 24455 32320
rect 24397 32311 24455 32317
rect 19944 32252 20300 32280
rect 19944 32240 19950 32252
rect 20530 32240 20536 32292
rect 20588 32280 20594 32292
rect 20625 32283 20683 32289
rect 20625 32280 20637 32283
rect 20588 32252 20637 32280
rect 20588 32240 20594 32252
rect 20625 32249 20637 32252
rect 20671 32249 20683 32283
rect 20625 32243 20683 32249
rect 22094 32240 22100 32292
rect 22152 32240 22158 32292
rect 23860 32280 23888 32311
rect 24946 32308 24952 32320
rect 25004 32308 25010 32360
rect 26344 32348 26372 32388
rect 26418 32376 26424 32428
rect 26476 32376 26482 32428
rect 27154 32376 27160 32428
rect 27212 32376 27218 32428
rect 27356 32425 27384 32456
rect 27341 32419 27399 32425
rect 27341 32385 27353 32419
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 27525 32419 27583 32425
rect 27525 32385 27537 32419
rect 27571 32385 27583 32419
rect 27525 32379 27583 32385
rect 27540 32348 27568 32379
rect 27706 32376 27712 32428
rect 27764 32376 27770 32428
rect 27982 32376 27988 32428
rect 28040 32416 28046 32428
rect 28801 32419 28859 32425
rect 28801 32416 28813 32419
rect 28040 32388 28813 32416
rect 28040 32376 28046 32388
rect 28801 32385 28813 32388
rect 28847 32416 28859 32419
rect 28902 32416 28908 32428
rect 28847 32388 28908 32416
rect 28847 32385 28859 32388
rect 28801 32379 28859 32385
rect 28902 32376 28908 32388
rect 28960 32376 28966 32428
rect 29012 32425 29040 32456
rect 30834 32444 30840 32496
rect 30892 32484 30898 32496
rect 32416 32484 32444 32512
rect 30892 32456 32444 32484
rect 33428 32456 34560 32484
rect 30892 32444 30898 32456
rect 28997 32419 29055 32425
rect 28997 32385 29009 32419
rect 29043 32416 29055 32419
rect 29086 32416 29092 32428
rect 29043 32388 29092 32416
rect 29043 32385 29055 32388
rect 28997 32379 29055 32385
rect 29086 32376 29092 32388
rect 29144 32376 29150 32428
rect 30098 32376 30104 32428
rect 30156 32376 30162 32428
rect 30285 32419 30343 32425
rect 30285 32385 30297 32419
rect 30331 32416 30343 32419
rect 30926 32416 30932 32428
rect 30331 32388 30932 32416
rect 30331 32385 30343 32388
rect 30285 32379 30343 32385
rect 30926 32376 30932 32388
rect 30984 32376 30990 32428
rect 31036 32425 31064 32456
rect 31021 32419 31079 32425
rect 31021 32385 31033 32419
rect 31067 32385 31079 32419
rect 31021 32379 31079 32385
rect 31570 32376 31576 32428
rect 31628 32416 31634 32428
rect 31665 32419 31723 32425
rect 31665 32416 31677 32419
rect 31628 32388 31677 32416
rect 31628 32376 31634 32388
rect 31665 32385 31677 32388
rect 31711 32385 31723 32419
rect 31665 32379 31723 32385
rect 32674 32376 32680 32428
rect 32732 32376 32738 32428
rect 33428 32425 33456 32456
rect 34532 32428 34560 32456
rect 33413 32419 33471 32425
rect 33413 32385 33425 32419
rect 33459 32385 33471 32419
rect 33413 32379 33471 32385
rect 33778 32376 33784 32428
rect 33836 32376 33842 32428
rect 34241 32419 34299 32425
rect 34241 32416 34253 32419
rect 34072 32388 34253 32416
rect 28534 32348 28540 32360
rect 26344 32320 28540 32348
rect 28534 32308 28540 32320
rect 28592 32308 28598 32360
rect 28626 32308 28632 32360
rect 28684 32348 28690 32360
rect 30190 32348 30196 32360
rect 28684 32320 30196 32348
rect 28684 32308 28690 32320
rect 30190 32308 30196 32320
rect 30248 32348 30254 32360
rect 30377 32351 30435 32357
rect 30377 32348 30389 32351
rect 30248 32320 30389 32348
rect 30248 32308 30254 32320
rect 30377 32317 30389 32320
rect 30423 32317 30435 32351
rect 31110 32348 31116 32360
rect 30377 32311 30435 32317
rect 30484 32320 31116 32348
rect 24302 32280 24308 32292
rect 22204 32252 23796 32280
rect 23860 32252 24308 32280
rect 18690 32212 18696 32224
rect 17420 32184 18696 32212
rect 17129 32175 17187 32181
rect 18690 32172 18696 32184
rect 18748 32172 18754 32224
rect 19521 32215 19579 32221
rect 19521 32181 19533 32215
rect 19567 32212 19579 32215
rect 19702 32212 19708 32224
rect 19567 32184 19708 32212
rect 19567 32181 19579 32184
rect 19521 32175 19579 32181
rect 19702 32172 19708 32184
rect 19760 32172 19766 32224
rect 19981 32215 20039 32221
rect 19981 32181 19993 32215
rect 20027 32212 20039 32215
rect 20898 32212 20904 32224
rect 20027 32184 20904 32212
rect 20027 32181 20039 32184
rect 19981 32175 20039 32181
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 21910 32172 21916 32224
rect 21968 32212 21974 32224
rect 22204 32212 22232 32252
rect 21968 32184 22232 32212
rect 21968 32172 21974 32184
rect 22278 32172 22284 32224
rect 22336 32172 22342 32224
rect 22830 32172 22836 32224
rect 22888 32212 22894 32224
rect 23198 32212 23204 32224
rect 22888 32184 23204 32212
rect 22888 32172 22894 32184
rect 23198 32172 23204 32184
rect 23256 32172 23262 32224
rect 23768 32212 23796 32252
rect 24302 32240 24308 32252
rect 24360 32280 24366 32292
rect 25038 32280 25044 32292
rect 24360 32252 25044 32280
rect 24360 32240 24366 32252
rect 25038 32240 25044 32252
rect 25096 32240 25102 32292
rect 27430 32240 27436 32292
rect 27488 32280 27494 32292
rect 30484 32280 30512 32320
rect 31110 32308 31116 32320
rect 31168 32308 31174 32360
rect 32858 32308 32864 32360
rect 32916 32308 32922 32360
rect 33321 32351 33379 32357
rect 33321 32317 33333 32351
rect 33367 32348 33379 32351
rect 34072 32348 34100 32388
rect 34241 32385 34253 32388
rect 34287 32416 34299 32419
rect 34422 32416 34428 32428
rect 34287 32388 34428 32416
rect 34287 32385 34299 32388
rect 34241 32379 34299 32385
rect 34422 32376 34428 32388
rect 34480 32376 34486 32428
rect 34514 32376 34520 32428
rect 34572 32416 34578 32428
rect 34609 32419 34667 32425
rect 34609 32416 34621 32419
rect 34572 32388 34621 32416
rect 34572 32376 34578 32388
rect 34609 32385 34621 32388
rect 34655 32416 34667 32419
rect 34974 32416 34980 32428
rect 34655 32388 34980 32416
rect 34655 32385 34667 32388
rect 34609 32379 34667 32385
rect 34974 32376 34980 32388
rect 35032 32376 35038 32428
rect 35084 32425 35112 32524
rect 37274 32444 37280 32496
rect 37332 32484 37338 32496
rect 37369 32487 37427 32493
rect 37369 32484 37381 32487
rect 37332 32456 37381 32484
rect 37332 32444 37338 32456
rect 37369 32453 37381 32456
rect 37415 32453 37427 32487
rect 37369 32447 37427 32453
rect 35069 32419 35127 32425
rect 35069 32385 35081 32419
rect 35115 32385 35127 32419
rect 35069 32379 35127 32385
rect 35437 32419 35495 32425
rect 35437 32385 35449 32419
rect 35483 32385 35495 32419
rect 37384 32416 37412 32447
rect 37642 32444 37648 32496
rect 37700 32484 37706 32496
rect 38102 32484 38108 32496
rect 37700 32456 38108 32484
rect 37700 32444 37706 32456
rect 38102 32444 38108 32456
rect 38160 32444 38166 32496
rect 37734 32416 37740 32428
rect 37384 32388 37740 32416
rect 35437 32379 35495 32385
rect 33367 32320 34100 32348
rect 34149 32351 34207 32357
rect 33367 32317 33379 32320
rect 33321 32311 33379 32317
rect 34149 32317 34161 32351
rect 34195 32348 34207 32351
rect 34790 32348 34796 32360
rect 34195 32320 34796 32348
rect 34195 32317 34207 32320
rect 34149 32311 34207 32317
rect 27488 32252 30512 32280
rect 27488 32240 27494 32252
rect 30650 32240 30656 32292
rect 30708 32240 30714 32292
rect 31297 32283 31355 32289
rect 31297 32280 31309 32283
rect 30760 32252 31309 32280
rect 25314 32212 25320 32224
rect 23768 32184 25320 32212
rect 25314 32172 25320 32184
rect 25372 32172 25378 32224
rect 26050 32172 26056 32224
rect 26108 32212 26114 32224
rect 27338 32212 27344 32224
rect 26108 32184 27344 32212
rect 26108 32172 26114 32184
rect 27338 32172 27344 32184
rect 27396 32172 27402 32224
rect 27522 32172 27528 32224
rect 27580 32172 27586 32224
rect 29178 32172 29184 32224
rect 29236 32212 29242 32224
rect 30006 32212 30012 32224
rect 29236 32184 30012 32212
rect 29236 32172 29242 32184
rect 30006 32172 30012 32184
rect 30064 32172 30070 32224
rect 30282 32172 30288 32224
rect 30340 32212 30346 32224
rect 30760 32212 30788 32252
rect 31297 32249 31309 32252
rect 31343 32249 31355 32283
rect 31297 32243 31355 32249
rect 30340 32184 30788 32212
rect 30340 32172 30346 32184
rect 30834 32172 30840 32224
rect 30892 32172 30898 32224
rect 33502 32172 33508 32224
rect 33560 32212 33566 32224
rect 33781 32215 33839 32221
rect 33781 32212 33793 32215
rect 33560 32184 33793 32212
rect 33560 32172 33566 32184
rect 33781 32181 33793 32184
rect 33827 32212 33839 32215
rect 34164 32212 34192 32311
rect 34790 32308 34796 32320
rect 34848 32348 34854 32360
rect 35452 32348 35480 32379
rect 37734 32376 37740 32388
rect 37792 32376 37798 32428
rect 35526 32348 35532 32360
rect 34848 32320 35532 32348
rect 34848 32308 34854 32320
rect 35526 32308 35532 32320
rect 35584 32308 35590 32360
rect 35618 32308 35624 32360
rect 35676 32308 35682 32360
rect 37642 32308 37648 32360
rect 37700 32348 37706 32360
rect 38562 32348 38568 32360
rect 37700 32320 38568 32348
rect 37700 32308 37706 32320
rect 38562 32308 38568 32320
rect 38620 32308 38626 32360
rect 34698 32240 34704 32292
rect 34756 32280 34762 32292
rect 35636 32280 35664 32308
rect 34756 32252 35664 32280
rect 34756 32240 34762 32252
rect 33827 32184 34192 32212
rect 34609 32215 34667 32221
rect 33827 32181 33839 32184
rect 33781 32175 33839 32181
rect 34609 32181 34621 32215
rect 34655 32212 34667 32215
rect 34882 32212 34888 32224
rect 34655 32184 34888 32212
rect 34655 32181 34667 32184
rect 34609 32175 34667 32181
rect 34882 32172 34888 32184
rect 34940 32172 34946 32224
rect 35452 32221 35480 32252
rect 35437 32215 35495 32221
rect 35437 32181 35449 32215
rect 35483 32181 35495 32215
rect 35437 32175 35495 32181
rect 35618 32172 35624 32224
rect 35676 32172 35682 32224
rect 1104 32122 41400 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 41400 32122
rect 1104 32048 41400 32070
rect 5902 31968 5908 32020
rect 5960 31968 5966 32020
rect 6178 31968 6184 32020
rect 6236 31968 6242 32020
rect 7926 31968 7932 32020
rect 7984 31968 7990 32020
rect 8478 32008 8484 32020
rect 8220 31980 8484 32008
rect 5629 31807 5687 31813
rect 5629 31773 5641 31807
rect 5675 31804 5687 31807
rect 5718 31804 5724 31816
rect 5675 31776 5724 31804
rect 5675 31773 5687 31776
rect 5629 31767 5687 31773
rect 5718 31764 5724 31776
rect 5776 31764 5782 31816
rect 5920 31813 5948 31968
rect 5905 31807 5963 31813
rect 5905 31773 5917 31807
rect 5951 31773 5963 31807
rect 5905 31767 5963 31773
rect 5994 31764 6000 31816
rect 6052 31764 6058 31816
rect 8110 31764 8116 31816
rect 8168 31764 8174 31816
rect 8220 31813 8248 31980
rect 8478 31968 8484 31980
rect 8536 31968 8542 32020
rect 8754 31968 8760 32020
rect 8812 32008 8818 32020
rect 9033 32011 9091 32017
rect 9033 32008 9045 32011
rect 8812 31980 9045 32008
rect 8812 31968 8818 31980
rect 9033 31977 9045 31980
rect 9079 31977 9091 32011
rect 9674 32008 9680 32020
rect 9033 31971 9091 31977
rect 9140 31980 9680 32008
rect 9140 31952 9168 31980
rect 9674 31968 9680 31980
rect 9732 31968 9738 32020
rect 9766 31968 9772 32020
rect 9824 32008 9830 32020
rect 10597 32011 10655 32017
rect 10597 32008 10609 32011
rect 9824 31980 10609 32008
rect 9824 31968 9830 31980
rect 10597 31977 10609 31980
rect 10643 31977 10655 32011
rect 10597 31971 10655 31977
rect 12250 31968 12256 32020
rect 12308 31968 12314 32020
rect 12342 31968 12348 32020
rect 12400 32008 12406 32020
rect 14090 32008 14096 32020
rect 12400 31980 14096 32008
rect 12400 31968 12406 31980
rect 14090 31968 14096 31980
rect 14148 31968 14154 32020
rect 14274 32008 14280 32020
rect 14200 31980 14280 32008
rect 9122 31940 9128 31952
rect 8312 31912 9128 31940
rect 8312 31813 8340 31912
rect 9122 31900 9128 31912
rect 9180 31900 9186 31952
rect 10226 31940 10232 31952
rect 9784 31912 10232 31940
rect 8573 31875 8631 31881
rect 8573 31841 8585 31875
rect 8619 31872 8631 31875
rect 8938 31872 8944 31884
rect 8619 31844 8944 31872
rect 8619 31841 8631 31844
rect 8573 31835 8631 31841
rect 8938 31832 8944 31844
rect 8996 31832 9002 31884
rect 9677 31875 9735 31881
rect 9677 31841 9689 31875
rect 9723 31841 9735 31875
rect 9677 31835 9735 31841
rect 8205 31807 8263 31813
rect 8205 31773 8217 31807
rect 8251 31773 8263 31807
rect 8205 31767 8263 31773
rect 8297 31807 8355 31813
rect 8297 31773 8309 31807
rect 8343 31773 8355 31807
rect 9217 31807 9275 31813
rect 9217 31804 9229 31807
rect 8297 31767 8355 31773
rect 9048 31776 9229 31804
rect 9048 31748 9076 31776
rect 9217 31773 9229 31776
rect 9263 31773 9275 31807
rect 9217 31767 9275 31773
rect 9309 31807 9367 31813
rect 9309 31773 9321 31807
rect 9355 31798 9367 31807
rect 9478 31807 9536 31813
rect 9355 31773 9444 31798
rect 9309 31770 9444 31773
rect 9309 31767 9367 31770
rect 5810 31696 5816 31748
rect 5868 31736 5874 31748
rect 8478 31745 8484 31748
rect 8435 31739 8484 31745
rect 5868 31708 6408 31736
rect 5868 31696 5874 31708
rect 6380 31680 6408 31708
rect 8435 31705 8447 31739
rect 8481 31705 8484 31739
rect 8435 31699 8484 31705
rect 8478 31696 8484 31699
rect 8536 31696 8542 31748
rect 9030 31696 9036 31748
rect 9088 31696 9094 31748
rect 6362 31628 6368 31680
rect 6420 31628 6426 31680
rect 8570 31628 8576 31680
rect 8628 31668 8634 31680
rect 8846 31668 8852 31680
rect 8628 31640 8852 31668
rect 8628 31628 8634 31640
rect 8846 31628 8852 31640
rect 8904 31628 8910 31680
rect 9214 31628 9220 31680
rect 9272 31668 9278 31680
rect 9416 31668 9444 31770
rect 9478 31773 9490 31807
rect 9524 31773 9536 31807
rect 9478 31767 9536 31773
rect 9272 31640 9444 31668
rect 9508 31668 9536 31767
rect 9595 31785 9653 31791
rect 9595 31751 9607 31785
rect 9641 31782 9653 31785
rect 9692 31782 9720 31835
rect 9641 31754 9720 31782
rect 9784 31804 9812 31912
rect 10226 31900 10232 31912
rect 10284 31940 10290 31952
rect 10284 31912 10548 31940
rect 10284 31900 10290 31912
rect 10042 31832 10048 31884
rect 10100 31832 10106 31884
rect 10321 31875 10379 31881
rect 10321 31841 10333 31875
rect 10367 31872 10379 31875
rect 10410 31872 10416 31884
rect 10367 31844 10416 31872
rect 10367 31841 10379 31844
rect 10321 31835 10379 31841
rect 10410 31832 10416 31844
rect 10468 31832 10474 31884
rect 10520 31872 10548 31912
rect 10778 31900 10784 31952
rect 10836 31900 10842 31952
rect 11882 31872 11888 31884
rect 10520 31844 11888 31872
rect 11882 31832 11888 31844
rect 11940 31832 11946 31884
rect 9861 31807 9919 31813
rect 9861 31804 9873 31807
rect 9784 31776 9873 31804
rect 9861 31773 9873 31776
rect 9907 31773 9919 31807
rect 10060 31804 10088 31832
rect 9861 31767 9919 31773
rect 9968 31776 10088 31804
rect 10183 31807 10241 31813
rect 9641 31751 9653 31754
rect 9595 31745 9653 31751
rect 9968 31745 9996 31776
rect 10183 31773 10195 31807
rect 10229 31773 10241 31807
rect 12268 31804 12296 31968
rect 13817 31943 13875 31949
rect 13817 31940 13829 31943
rect 12729 31912 13829 31940
rect 12729 31813 12757 31912
rect 13817 31909 13829 31912
rect 13863 31940 13875 31943
rect 14200 31940 14228 31980
rect 14274 31968 14280 31980
rect 14332 32008 14338 32020
rect 15010 32008 15016 32020
rect 14332 31980 15016 32008
rect 14332 31968 14338 31980
rect 15010 31968 15016 31980
rect 15068 31968 15074 32020
rect 15930 31968 15936 32020
rect 15988 31968 15994 32020
rect 16666 31968 16672 32020
rect 16724 31968 16730 32020
rect 18417 32011 18475 32017
rect 16776 31980 18368 32008
rect 16776 31940 16804 31980
rect 13863 31912 14228 31940
rect 14256 31912 16804 31940
rect 13863 31909 13875 31912
rect 13817 31903 13875 31909
rect 13078 31872 13084 31884
rect 12820 31844 13084 31872
rect 12820 31813 12848 31844
rect 13078 31832 13084 31844
rect 13136 31872 13142 31884
rect 13449 31875 13507 31881
rect 13136 31844 13308 31872
rect 13136 31832 13142 31844
rect 12437 31807 12495 31813
rect 12437 31804 12449 31807
rect 12268 31776 12449 31804
rect 10183 31767 10241 31773
rect 12437 31773 12449 31776
rect 12483 31773 12495 31807
rect 9953 31739 10011 31745
rect 9953 31705 9965 31739
rect 9999 31705 10011 31739
rect 9953 31699 10011 31705
rect 10042 31696 10048 31748
rect 10100 31696 10106 31748
rect 9582 31668 9588 31680
rect 9508 31640 9588 31668
rect 9272 31628 9278 31640
rect 9582 31628 9588 31640
rect 9640 31628 9646 31680
rect 9766 31628 9772 31680
rect 9824 31668 9830 31680
rect 10198 31668 10226 31767
rect 10520 31748 10640 31770
rect 12437 31767 12495 31773
rect 12530 31807 12588 31813
rect 12530 31773 12542 31807
rect 12576 31804 12588 31807
rect 12713 31807 12771 31813
rect 12576 31776 12609 31804
rect 12576 31773 12588 31776
rect 12530 31767 12588 31773
rect 12713 31773 12725 31807
rect 12759 31773 12771 31807
rect 12713 31767 12771 31773
rect 12805 31807 12863 31813
rect 12805 31773 12817 31807
rect 12851 31773 12863 31807
rect 12805 31767 12863 31773
rect 10413 31739 10471 31745
rect 10413 31705 10425 31739
rect 10459 31736 10471 31739
rect 10502 31736 10508 31748
rect 10459 31708 10508 31736
rect 10459 31705 10471 31708
rect 10413 31699 10471 31705
rect 10502 31696 10508 31708
rect 10560 31742 10640 31748
rect 10560 31696 10566 31742
rect 10612 31736 10640 31742
rect 11606 31736 11612 31748
rect 10612 31708 11612 31736
rect 11606 31696 11612 31708
rect 11664 31696 11670 31748
rect 12544 31736 12572 31767
rect 12894 31764 12900 31816
rect 12952 31813 12958 31816
rect 12952 31804 12960 31813
rect 12952 31776 12997 31804
rect 12952 31767 12960 31776
rect 12952 31764 12958 31767
rect 12544 31708 13216 31736
rect 13188 31680 13216 31708
rect 9824 31640 10226 31668
rect 10623 31671 10681 31677
rect 9824 31628 9830 31640
rect 10623 31637 10635 31671
rect 10669 31668 10681 31671
rect 10962 31668 10968 31680
rect 10669 31640 10968 31668
rect 10669 31637 10681 31640
rect 10623 31631 10681 31637
rect 10962 31628 10968 31640
rect 11020 31628 11026 31680
rect 12618 31628 12624 31680
rect 12676 31668 12682 31680
rect 13081 31671 13139 31677
rect 13081 31668 13093 31671
rect 12676 31640 13093 31668
rect 12676 31628 12682 31640
rect 13081 31637 13093 31640
rect 13127 31637 13139 31671
rect 13081 31631 13139 31637
rect 13170 31628 13176 31680
rect 13228 31628 13234 31680
rect 13280 31668 13308 31844
rect 13449 31841 13461 31875
rect 13495 31872 13507 31875
rect 13538 31872 13544 31884
rect 13495 31844 13544 31872
rect 13495 31841 13507 31844
rect 13449 31835 13507 31841
rect 13538 31832 13544 31844
rect 13596 31872 13602 31884
rect 13596 31844 13860 31872
rect 13596 31832 13602 31844
rect 13633 31807 13691 31813
rect 13633 31773 13645 31807
rect 13679 31804 13691 31807
rect 13832 31804 13860 31844
rect 13906 31832 13912 31884
rect 13964 31832 13970 31884
rect 14090 31804 14096 31816
rect 13679 31776 13713 31804
rect 13832 31776 14096 31804
rect 13679 31773 13691 31776
rect 13633 31767 13691 31773
rect 13446 31696 13452 31748
rect 13504 31736 13510 31748
rect 13648 31736 13676 31767
rect 14090 31764 14096 31776
rect 14148 31764 14154 31816
rect 13504 31708 13676 31736
rect 13504 31696 13510 31708
rect 14256 31668 14284 31912
rect 17034 31900 17040 31952
rect 17092 31900 17098 31952
rect 17862 31900 17868 31952
rect 17920 31900 17926 31952
rect 18230 31900 18236 31952
rect 18288 31900 18294 31952
rect 18340 31940 18368 31980
rect 18417 31977 18429 32011
rect 18463 32008 18475 32011
rect 19242 32008 19248 32020
rect 18463 31980 19248 32008
rect 18463 31977 18475 31980
rect 18417 31971 18475 31977
rect 19242 31968 19248 31980
rect 19300 31968 19306 32020
rect 20806 31968 20812 32020
rect 20864 31968 20870 32020
rect 21082 31968 21088 32020
rect 21140 32008 21146 32020
rect 21177 32011 21235 32017
rect 21177 32008 21189 32011
rect 21140 31980 21189 32008
rect 21140 31968 21146 31980
rect 21177 31977 21189 31980
rect 21223 31977 21235 32011
rect 21177 31971 21235 31977
rect 21266 31968 21272 32020
rect 21324 31968 21330 32020
rect 21358 31968 21364 32020
rect 21416 32008 21422 32020
rect 21637 32011 21695 32017
rect 21637 32008 21649 32011
rect 21416 31980 21649 32008
rect 21416 31968 21422 31980
rect 21637 31977 21649 31980
rect 21683 32008 21695 32011
rect 22189 32011 22247 32017
rect 22189 32008 22201 32011
rect 21683 31980 22201 32008
rect 21683 31977 21695 31980
rect 21637 31971 21695 31977
rect 22189 31977 22201 31980
rect 22235 31977 22247 32011
rect 22189 31971 22247 31977
rect 22285 31980 26453 32008
rect 19886 31940 19892 31952
rect 18340 31912 19892 31940
rect 19886 31900 19892 31912
rect 19944 31900 19950 31952
rect 20990 31940 20996 31952
rect 20824 31912 20996 31940
rect 15841 31875 15899 31881
rect 15841 31841 15853 31875
rect 15887 31872 15899 31875
rect 16574 31872 16580 31884
rect 15887 31844 16580 31872
rect 15887 31841 15899 31844
rect 15841 31835 15899 31841
rect 16574 31832 16580 31844
rect 16632 31832 16638 31884
rect 17402 31872 17408 31884
rect 16868 31844 17408 31872
rect 15654 31764 15660 31816
rect 15712 31764 15718 31816
rect 15930 31764 15936 31816
rect 15988 31764 15994 31816
rect 16114 31764 16120 31816
rect 16172 31804 16178 31816
rect 16868 31813 16896 31844
rect 17402 31832 17408 31844
rect 17460 31832 17466 31884
rect 17880 31872 17908 31900
rect 18248 31872 18276 31900
rect 20824 31884 20852 31912
rect 20990 31900 20996 31912
rect 21048 31900 21054 31952
rect 22097 31943 22155 31949
rect 22097 31940 22109 31943
rect 21560 31912 22109 31940
rect 17880 31844 18092 31872
rect 18248 31844 18552 31872
rect 16853 31807 16911 31813
rect 16853 31804 16865 31807
rect 16172 31776 16865 31804
rect 16172 31764 16178 31776
rect 16853 31773 16865 31776
rect 16899 31773 16911 31807
rect 16853 31767 16911 31773
rect 17126 31764 17132 31816
rect 17184 31764 17190 31816
rect 17954 31764 17960 31816
rect 18012 31764 18018 31816
rect 18064 31804 18092 31844
rect 18233 31807 18291 31813
rect 18233 31804 18245 31807
rect 18064 31776 18245 31804
rect 18233 31773 18245 31776
rect 18279 31773 18291 31807
rect 18233 31767 18291 31773
rect 18322 31764 18328 31816
rect 18380 31764 18386 31816
rect 18524 31813 18552 31844
rect 20806 31832 20812 31884
rect 20864 31832 20870 31884
rect 21008 31844 21496 31872
rect 18509 31807 18567 31813
rect 18509 31773 18521 31807
rect 18555 31773 18567 31807
rect 18509 31767 18567 31773
rect 15838 31696 15844 31748
rect 15896 31736 15902 31748
rect 16574 31736 16580 31748
rect 15896 31708 16580 31736
rect 15896 31696 15902 31708
rect 16574 31696 16580 31708
rect 16632 31696 16638 31748
rect 13280 31640 14284 31668
rect 15010 31628 15016 31680
rect 15068 31668 15074 31680
rect 15930 31668 15936 31680
rect 15068 31640 15936 31668
rect 15068 31628 15074 31640
rect 15930 31628 15936 31640
rect 15988 31628 15994 31680
rect 16022 31628 16028 31680
rect 16080 31668 16086 31680
rect 16117 31671 16175 31677
rect 16117 31668 16129 31671
rect 16080 31640 16129 31668
rect 16080 31628 16086 31640
rect 16117 31637 16129 31640
rect 16163 31637 16175 31671
rect 17144 31668 17172 31764
rect 18524 31736 18552 31767
rect 18690 31764 18696 31816
rect 18748 31804 18754 31816
rect 21008 31804 21036 31844
rect 18748 31776 21036 31804
rect 21085 31807 21143 31813
rect 18748 31764 18754 31776
rect 21085 31773 21097 31807
rect 21131 31773 21143 31807
rect 21266 31804 21272 31816
rect 21085 31767 21143 31773
rect 21192 31776 21272 31804
rect 21100 31736 21128 31767
rect 21192 31748 21220 31776
rect 21266 31764 21272 31776
rect 21324 31764 21330 31816
rect 21358 31764 21364 31816
rect 21416 31764 21422 31816
rect 18524 31708 21128 31736
rect 21174 31696 21180 31748
rect 21232 31696 21238 31748
rect 21468 31736 21496 31844
rect 21560 31813 21588 31912
rect 22097 31909 22109 31912
rect 22143 31909 22155 31943
rect 22097 31903 22155 31909
rect 21726 31832 21732 31884
rect 21784 31832 21790 31884
rect 22285 31872 22313 31980
rect 22462 31900 22468 31952
rect 22520 31900 22526 31952
rect 22646 31900 22652 31952
rect 22704 31940 22710 31952
rect 22830 31940 22836 31952
rect 22704 31912 22836 31940
rect 22704 31900 22710 31912
rect 22830 31900 22836 31912
rect 22888 31900 22894 31952
rect 24394 31900 24400 31952
rect 24452 31940 24458 31952
rect 24578 31940 24584 31952
rect 24452 31912 24584 31940
rect 24452 31900 24458 31912
rect 24578 31900 24584 31912
rect 24636 31900 24642 31952
rect 24670 31900 24676 31952
rect 24728 31940 24734 31952
rect 25222 31940 25228 31952
rect 24728 31912 25228 31940
rect 24728 31900 24734 31912
rect 25222 31900 25228 31912
rect 25280 31900 25286 31952
rect 25774 31900 25780 31952
rect 25832 31940 25838 31952
rect 25961 31943 26019 31949
rect 25961 31940 25973 31943
rect 25832 31912 25973 31940
rect 25832 31900 25838 31912
rect 25961 31909 25973 31912
rect 26007 31909 26019 31943
rect 25961 31903 26019 31909
rect 26234 31900 26240 31952
rect 26292 31900 26298 31952
rect 26326 31900 26332 31952
rect 26384 31900 26390 31952
rect 26425 31940 26453 31980
rect 26510 31968 26516 32020
rect 26568 32008 26574 32020
rect 27801 32011 27859 32017
rect 27801 32008 27813 32011
rect 26568 31980 27813 32008
rect 26568 31968 26574 31980
rect 27801 31977 27813 31980
rect 27847 32008 27859 32011
rect 27847 31980 28304 32008
rect 27847 31977 27859 31980
rect 27801 31971 27859 31977
rect 28169 31943 28227 31949
rect 28169 31940 28181 31943
rect 26425 31912 28181 31940
rect 28169 31909 28181 31912
rect 28215 31909 28227 31943
rect 28276 31940 28304 31980
rect 28718 31968 28724 32020
rect 28776 32008 28782 32020
rect 28776 31980 29316 32008
rect 28776 31968 28782 31980
rect 29288 31952 29316 31980
rect 29730 31968 29736 32020
rect 29788 31968 29794 32020
rect 30006 31968 30012 32020
rect 30064 32008 30070 32020
rect 30834 32008 30840 32020
rect 30064 31980 30840 32008
rect 30064 31968 30070 31980
rect 30834 31968 30840 31980
rect 30892 31968 30898 32020
rect 30926 31968 30932 32020
rect 30984 31968 30990 32020
rect 31294 31968 31300 32020
rect 31352 32008 31358 32020
rect 31849 32011 31907 32017
rect 31849 32008 31861 32011
rect 31352 31980 31861 32008
rect 31352 31968 31358 31980
rect 31849 31977 31861 31980
rect 31895 31977 31907 32011
rect 31849 31971 31907 31977
rect 32674 31968 32680 32020
rect 32732 31968 32738 32020
rect 33778 31968 33784 32020
rect 33836 31968 33842 32020
rect 35618 31968 35624 32020
rect 35676 31968 35682 32020
rect 28994 31940 29000 31952
rect 28276 31912 29000 31940
rect 28169 31903 28227 31909
rect 28994 31900 29000 31912
rect 29052 31900 29058 31952
rect 29086 31900 29092 31952
rect 29144 31940 29150 31952
rect 29144 31912 29217 31940
rect 29144 31900 29150 31912
rect 22480 31872 22508 31900
rect 26252 31872 26280 31900
rect 27893 31875 27951 31881
rect 21836 31844 22313 31872
rect 22388 31844 22508 31872
rect 24504 31844 26004 31872
rect 26252 31844 26464 31872
rect 21545 31807 21603 31813
rect 21545 31773 21557 31807
rect 21591 31773 21603 31807
rect 21545 31767 21603 31773
rect 21634 31764 21640 31816
rect 21692 31764 21698 31816
rect 21836 31736 21864 31844
rect 21910 31764 21916 31816
rect 21968 31764 21974 31816
rect 22189 31807 22247 31813
rect 22189 31773 22201 31807
rect 22235 31804 22247 31807
rect 22388 31804 22416 31844
rect 22235 31776 22416 31804
rect 22465 31807 22523 31813
rect 22235 31773 22247 31776
rect 22189 31767 22247 31773
rect 22465 31773 22477 31807
rect 22511 31804 22523 31807
rect 23014 31804 23020 31816
rect 22511 31776 23020 31804
rect 22511 31773 22523 31776
rect 22465 31767 22523 31773
rect 23014 31764 23020 31776
rect 23072 31764 23078 31816
rect 24504 31813 24532 31844
rect 25976 31816 26004 31844
rect 24489 31807 24547 31813
rect 24489 31773 24501 31807
rect 24535 31773 24547 31807
rect 24489 31767 24547 31773
rect 24946 31764 24952 31816
rect 25004 31764 25010 31816
rect 25038 31764 25044 31816
rect 25096 31804 25102 31816
rect 25096 31776 25176 31804
rect 25096 31764 25102 31776
rect 21468 31708 21864 31736
rect 22370 31696 22376 31748
rect 22428 31736 22434 31748
rect 24964 31736 24992 31764
rect 25148 31745 25176 31776
rect 25314 31764 25320 31816
rect 25372 31764 25378 31816
rect 25958 31764 25964 31816
rect 26016 31764 26022 31816
rect 26050 31764 26056 31816
rect 26108 31804 26114 31816
rect 26436 31813 26464 31844
rect 27893 31841 27905 31875
rect 27939 31872 27951 31875
rect 28074 31872 28080 31884
rect 27939 31844 28080 31872
rect 27939 31841 27951 31844
rect 27893 31835 27951 31841
rect 28074 31832 28080 31844
rect 28132 31832 28138 31884
rect 28810 31832 28816 31884
rect 28868 31872 28874 31884
rect 28868 31844 29040 31872
rect 28868 31832 28874 31844
rect 26145 31807 26203 31813
rect 26145 31804 26157 31807
rect 26108 31776 26157 31804
rect 26108 31764 26114 31776
rect 26145 31773 26157 31776
rect 26191 31773 26203 31807
rect 26145 31767 26203 31773
rect 26237 31807 26295 31813
rect 26237 31773 26249 31807
rect 26283 31773 26295 31807
rect 26237 31767 26295 31773
rect 26421 31807 26479 31813
rect 26421 31773 26433 31807
rect 26467 31773 26479 31807
rect 26421 31767 26479 31773
rect 22428 31708 24992 31736
rect 25133 31739 25191 31745
rect 22428 31696 22434 31708
rect 25133 31705 25145 31739
rect 25179 31705 25191 31739
rect 25332 31736 25360 31764
rect 26252 31736 26280 31767
rect 27246 31764 27252 31816
rect 27304 31804 27310 31816
rect 27801 31807 27859 31813
rect 27801 31804 27813 31807
rect 27304 31776 27813 31804
rect 27304 31764 27310 31776
rect 27801 31773 27813 31776
rect 27847 31804 27859 31807
rect 27982 31804 27988 31816
rect 27847 31776 27988 31804
rect 27847 31773 27859 31776
rect 27801 31767 27859 31773
rect 27982 31764 27988 31776
rect 28040 31764 28046 31816
rect 26602 31736 26608 31748
rect 25332 31708 26608 31736
rect 25133 31699 25191 31705
rect 26602 31696 26608 31708
rect 26660 31696 26666 31748
rect 18782 31668 18788 31680
rect 17144 31640 18788 31668
rect 16117 31631 16175 31637
rect 18782 31628 18788 31640
rect 18840 31668 18846 31680
rect 19610 31668 19616 31680
rect 18840 31640 19616 31668
rect 18840 31628 18846 31640
rect 19610 31628 19616 31640
rect 19668 31668 19674 31680
rect 22002 31668 22008 31680
rect 19668 31640 22008 31668
rect 19668 31628 19674 31640
rect 22002 31628 22008 31640
rect 22060 31628 22066 31680
rect 23106 31628 23112 31680
rect 23164 31668 23170 31680
rect 25590 31668 25596 31680
rect 23164 31640 25596 31668
rect 23164 31628 23170 31640
rect 25590 31628 25596 31640
rect 25648 31628 25654 31680
rect 26142 31628 26148 31680
rect 26200 31668 26206 31680
rect 26510 31668 26516 31680
rect 26200 31640 26516 31668
rect 26200 31628 26206 31640
rect 26510 31628 26516 31640
rect 26568 31668 26574 31680
rect 26970 31668 26976 31680
rect 26568 31640 26976 31668
rect 26568 31628 26574 31640
rect 26970 31628 26976 31640
rect 27028 31628 27034 31680
rect 27246 31628 27252 31680
rect 27304 31668 27310 31680
rect 27522 31668 27528 31680
rect 27304 31640 27528 31668
rect 27304 31628 27310 31640
rect 27522 31628 27528 31640
rect 27580 31628 27586 31680
rect 28092 31668 28120 31832
rect 28258 31764 28264 31816
rect 28316 31804 28322 31816
rect 28537 31807 28595 31813
rect 28537 31804 28549 31807
rect 28316 31776 28549 31804
rect 28316 31764 28322 31776
rect 28537 31773 28549 31776
rect 28583 31773 28595 31807
rect 28537 31767 28595 31773
rect 28721 31807 28779 31813
rect 28721 31773 28733 31807
rect 28767 31773 28779 31807
rect 28721 31767 28779 31773
rect 28736 31736 28764 31767
rect 28902 31764 28908 31816
rect 28960 31764 28966 31816
rect 29012 31813 29040 31844
rect 28997 31807 29055 31813
rect 28997 31773 29009 31807
rect 29043 31773 29055 31807
rect 28997 31767 29055 31773
rect 29086 31764 29092 31816
rect 29144 31764 29150 31816
rect 29189 31813 29217 31912
rect 29270 31900 29276 31952
rect 29328 31900 29334 31952
rect 29748 31940 29776 31968
rect 29914 31940 29920 31952
rect 29748 31912 29920 31940
rect 29914 31900 29920 31912
rect 29972 31940 29978 31952
rect 29972 31912 30604 31940
rect 29972 31900 29978 31912
rect 29288 31872 29316 31900
rect 30576 31881 30604 31912
rect 30561 31875 30619 31881
rect 29288 31844 30328 31872
rect 30300 31816 30328 31844
rect 30561 31841 30573 31875
rect 30607 31841 30619 31875
rect 30561 31835 30619 31841
rect 29189 31807 29263 31813
rect 29189 31776 29217 31807
rect 29205 31773 29217 31776
rect 29251 31773 29263 31807
rect 29205 31767 29263 31773
rect 29362 31764 29368 31816
rect 29420 31764 29426 31816
rect 30282 31764 30288 31816
rect 30340 31764 30346 31816
rect 30374 31764 30380 31816
rect 30432 31804 30438 31816
rect 30944 31813 30972 31968
rect 31110 31900 31116 31952
rect 31168 31940 31174 31952
rect 32692 31940 32720 31968
rect 33965 31943 34023 31949
rect 33965 31940 33977 31943
rect 31168 31912 31892 31940
rect 32692 31912 33977 31940
rect 31168 31900 31174 31912
rect 31312 31844 31800 31872
rect 30469 31807 30527 31813
rect 30469 31804 30481 31807
rect 30432 31776 30481 31804
rect 30432 31764 30438 31776
rect 30469 31773 30481 31776
rect 30515 31773 30527 31807
rect 30469 31767 30527 31773
rect 30929 31807 30987 31813
rect 30929 31773 30941 31807
rect 30975 31804 30987 31807
rect 30975 31776 31156 31804
rect 30975 31773 30987 31776
rect 30929 31767 30987 31773
rect 29098 31736 29126 31764
rect 28736 31708 29126 31736
rect 31128 31736 31156 31776
rect 31312 31736 31340 31844
rect 31772 31813 31800 31844
rect 31389 31807 31447 31813
rect 31389 31773 31401 31807
rect 31435 31804 31447 31807
rect 31757 31807 31815 31813
rect 31435 31776 31708 31804
rect 31435 31773 31447 31776
rect 31389 31767 31447 31773
rect 31128 31708 31340 31736
rect 31680 31736 31708 31776
rect 31757 31773 31769 31807
rect 31803 31773 31815 31807
rect 31757 31767 31815 31773
rect 31864 31804 31892 31912
rect 33965 31909 33977 31912
rect 34011 31909 34023 31943
rect 33965 31903 34023 31909
rect 33594 31832 33600 31884
rect 33652 31872 33658 31884
rect 33689 31875 33747 31881
rect 33689 31872 33701 31875
rect 33652 31844 33701 31872
rect 33652 31832 33658 31844
rect 33689 31841 33701 31844
rect 33735 31872 33747 31875
rect 34422 31872 34428 31884
rect 33735 31844 34428 31872
rect 33735 31841 33747 31844
rect 33689 31835 33747 31841
rect 34422 31832 34428 31844
rect 34480 31832 34486 31884
rect 34885 31875 34943 31881
rect 34885 31872 34897 31875
rect 34624 31844 34897 31872
rect 33321 31807 33379 31813
rect 31864 31776 33272 31804
rect 31864 31736 31892 31776
rect 31680 31708 31892 31736
rect 33244 31736 33272 31776
rect 33321 31773 33333 31807
rect 33367 31804 33379 31807
rect 33502 31804 33508 31816
rect 33367 31776 33508 31804
rect 33367 31773 33379 31776
rect 33321 31767 33379 31773
rect 33502 31764 33508 31776
rect 33560 31764 33566 31816
rect 33781 31807 33839 31813
rect 33781 31773 33793 31807
rect 33827 31804 33839 31807
rect 34514 31804 34520 31816
rect 33827 31776 34520 31804
rect 33827 31773 33839 31776
rect 33781 31767 33839 31773
rect 34514 31764 34520 31776
rect 34572 31764 34578 31816
rect 34624 31736 34652 31844
rect 34885 31841 34897 31844
rect 34931 31841 34943 31875
rect 34885 31835 34943 31841
rect 34701 31807 34759 31813
rect 34701 31773 34713 31807
rect 34747 31804 34759 31807
rect 35636 31804 35664 31968
rect 34747 31776 35664 31804
rect 34747 31773 34759 31776
rect 34701 31767 34759 31773
rect 33244 31708 34652 31736
rect 28629 31671 28687 31677
rect 28629 31668 28641 31671
rect 28092 31640 28641 31668
rect 28629 31637 28641 31640
rect 28675 31668 28687 31671
rect 28810 31668 28816 31680
rect 28675 31640 28816 31668
rect 28675 31637 28687 31640
rect 28629 31631 28687 31637
rect 28810 31628 28816 31640
rect 28868 31628 28874 31680
rect 29178 31628 29184 31680
rect 29236 31668 29242 31680
rect 29273 31671 29331 31677
rect 29273 31668 29285 31671
rect 29236 31640 29285 31668
rect 29236 31628 29242 31640
rect 29273 31637 29285 31640
rect 29319 31637 29331 31671
rect 29273 31631 29331 31637
rect 30926 31628 30932 31680
rect 30984 31628 30990 31680
rect 1104 31578 41400 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 41400 31578
rect 1104 31504 41400 31526
rect 6181 31467 6239 31473
rect 6181 31433 6193 31467
rect 6227 31433 6239 31467
rect 6181 31427 6239 31433
rect 6196 31396 6224 31427
rect 7650 31424 7656 31476
rect 7708 31464 7714 31476
rect 8846 31464 8852 31476
rect 7708 31436 8852 31464
rect 7708 31424 7714 31436
rect 6641 31399 6699 31405
rect 6641 31396 6653 31399
rect 5644 31368 6132 31396
rect 6196 31368 6653 31396
rect 5644 31337 5672 31368
rect 6104 31340 6132 31368
rect 6641 31365 6653 31368
rect 6687 31365 6699 31399
rect 6641 31359 6699 31365
rect 7282 31356 7288 31408
rect 7340 31356 7346 31408
rect 8018 31356 8024 31408
rect 8076 31396 8082 31408
rect 8389 31399 8447 31405
rect 8389 31396 8401 31399
rect 8076 31368 8401 31396
rect 8076 31356 8082 31368
rect 8389 31365 8401 31368
rect 8435 31365 8447 31399
rect 8389 31359 8447 31365
rect 5629 31331 5687 31337
rect 5629 31297 5641 31331
rect 5675 31297 5687 31331
rect 5629 31291 5687 31297
rect 5810 31288 5816 31340
rect 5868 31288 5874 31340
rect 5902 31288 5908 31340
rect 5960 31288 5966 31340
rect 5994 31288 6000 31340
rect 6052 31288 6058 31340
rect 6086 31288 6092 31340
rect 6144 31288 6150 31340
rect 8496 31337 8524 31436
rect 8846 31424 8852 31436
rect 8904 31424 8910 31476
rect 9214 31424 9220 31476
rect 9272 31464 9278 31476
rect 9272 31436 9720 31464
rect 9272 31424 9278 31436
rect 9398 31396 9404 31408
rect 8680 31368 9404 31396
rect 8680 31337 8708 31368
rect 9398 31356 9404 31368
rect 9456 31356 9462 31408
rect 9582 31356 9588 31408
rect 9640 31356 9646 31408
rect 8481 31331 8539 31337
rect 8481 31297 8493 31331
rect 8527 31297 8539 31331
rect 8481 31291 8539 31297
rect 8665 31331 8723 31337
rect 8665 31297 8677 31331
rect 8711 31297 8723 31331
rect 8665 31291 8723 31297
rect 8754 31288 8760 31340
rect 8812 31288 8818 31340
rect 8850 31331 8908 31337
rect 8850 31297 8862 31331
rect 8896 31297 8908 31331
rect 8850 31291 8908 31297
rect 4614 31220 4620 31272
rect 4672 31260 4678 31272
rect 6365 31263 6423 31269
rect 6365 31260 6377 31263
rect 4672 31232 6377 31260
rect 4672 31220 4678 31232
rect 6365 31229 6377 31232
rect 6411 31229 6423 31263
rect 6365 31223 6423 31229
rect 8662 31152 8668 31204
rect 8720 31192 8726 31204
rect 8864 31192 8892 31291
rect 8938 31288 8944 31340
rect 8996 31328 9002 31340
rect 9692 31337 9720 31436
rect 10042 31424 10048 31476
rect 10100 31464 10106 31476
rect 10502 31464 10508 31476
rect 10100 31436 10508 31464
rect 10100 31424 10106 31436
rect 10502 31424 10508 31436
rect 10560 31424 10566 31476
rect 13170 31464 13176 31476
rect 12406 31436 13176 31464
rect 9309 31331 9367 31337
rect 9309 31328 9321 31331
rect 8996 31300 9321 31328
rect 8996 31288 9002 31300
rect 9309 31297 9321 31300
rect 9355 31297 9367 31331
rect 9309 31291 9367 31297
rect 9493 31331 9551 31337
rect 9493 31297 9505 31331
rect 9539 31297 9551 31331
rect 9493 31291 9551 31297
rect 9677 31331 9735 31337
rect 9677 31297 9689 31331
rect 9723 31297 9735 31331
rect 12406 31328 12434 31436
rect 13170 31424 13176 31436
rect 13228 31464 13234 31476
rect 13354 31464 13360 31476
rect 13228 31436 13360 31464
rect 13228 31424 13234 31436
rect 13354 31424 13360 31436
rect 13412 31424 13418 31476
rect 13648 31436 15608 31464
rect 12989 31399 13047 31405
rect 12989 31396 13001 31399
rect 9677 31291 9735 31297
rect 9784 31300 12434 31328
rect 12544 31368 13001 31396
rect 8720 31164 8892 31192
rect 9125 31195 9183 31201
rect 8720 31152 8726 31164
rect 9125 31161 9137 31195
rect 9171 31161 9183 31195
rect 9125 31155 9183 31161
rect 6454 31084 6460 31136
rect 6512 31124 6518 31136
rect 9140 31124 9168 31155
rect 9398 31152 9404 31204
rect 9456 31192 9462 31204
rect 9508 31192 9536 31291
rect 9582 31220 9588 31272
rect 9640 31260 9646 31272
rect 9784 31260 9812 31300
rect 9640 31232 9812 31260
rect 9640 31220 9646 31232
rect 10962 31220 10968 31272
rect 11020 31260 11026 31272
rect 12544 31260 12572 31368
rect 12989 31365 13001 31368
rect 13035 31396 13047 31399
rect 13648 31396 13676 31436
rect 15580 31408 15608 31436
rect 17402 31424 17408 31476
rect 17460 31464 17466 31476
rect 17460 31436 22232 31464
rect 17460 31424 17466 31436
rect 13035 31368 13676 31396
rect 13035 31365 13047 31368
rect 12989 31359 13047 31365
rect 13814 31356 13820 31408
rect 13872 31396 13878 31408
rect 14461 31399 14519 31405
rect 14461 31396 14473 31399
rect 13872 31368 14473 31396
rect 13872 31356 13878 31368
rect 14461 31365 14473 31368
rect 14507 31396 14519 31399
rect 14507 31368 15056 31396
rect 14507 31365 14519 31368
rect 14461 31359 14519 31365
rect 12618 31288 12624 31340
rect 12676 31288 12682 31340
rect 12710 31288 12716 31340
rect 12768 31328 12774 31340
rect 12768 31300 12813 31328
rect 12768 31288 12774 31300
rect 12894 31288 12900 31340
rect 12952 31288 12958 31340
rect 13086 31331 13144 31337
rect 13086 31297 13098 31331
rect 13132 31328 13144 31331
rect 13630 31328 13636 31340
rect 13132 31300 13636 31328
rect 13132 31297 13144 31300
rect 13086 31291 13144 31297
rect 11020 31232 12572 31260
rect 11020 31220 11026 31232
rect 12250 31192 12256 31204
rect 9456 31164 12256 31192
rect 9456 31152 9462 31164
rect 12250 31152 12256 31164
rect 12308 31152 12314 31204
rect 12618 31152 12624 31204
rect 12676 31192 12682 31204
rect 13101 31192 13129 31291
rect 13630 31288 13636 31300
rect 13688 31288 13694 31340
rect 14090 31288 14096 31340
rect 14148 31288 14154 31340
rect 14274 31337 14280 31340
rect 14241 31331 14280 31337
rect 14241 31297 14253 31331
rect 14241 31291 14280 31297
rect 14274 31288 14280 31291
rect 14332 31288 14338 31340
rect 14369 31331 14427 31337
rect 14369 31297 14381 31331
rect 14415 31297 14427 31331
rect 14369 31291 14427 31297
rect 14599 31331 14657 31337
rect 14599 31297 14611 31331
rect 14645 31328 14657 31331
rect 14918 31328 14924 31340
rect 14645 31300 14924 31328
rect 14645 31297 14657 31300
rect 14599 31291 14657 31297
rect 14384 31260 14412 31291
rect 14918 31288 14924 31300
rect 14976 31288 14982 31340
rect 15028 31328 15056 31368
rect 15562 31356 15568 31408
rect 15620 31356 15626 31408
rect 15930 31356 15936 31408
rect 15988 31396 15994 31408
rect 22204 31396 22232 31436
rect 22462 31424 22468 31476
rect 22520 31464 22526 31476
rect 29089 31467 29147 31473
rect 29089 31464 29101 31467
rect 22520 31436 29101 31464
rect 22520 31424 22526 31436
rect 29089 31433 29101 31436
rect 29135 31433 29147 31467
rect 31018 31464 31024 31476
rect 29089 31427 29147 31433
rect 29840 31436 31024 31464
rect 15988 31368 22140 31396
rect 22204 31368 24520 31396
rect 15988 31356 15994 31368
rect 16114 31328 16120 31340
rect 15028 31300 16120 31328
rect 16114 31288 16120 31300
rect 16172 31288 16178 31340
rect 16298 31288 16304 31340
rect 16356 31328 16362 31340
rect 18506 31328 18512 31340
rect 16356 31300 18512 31328
rect 16356 31288 16362 31300
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 19978 31288 19984 31340
rect 20036 31328 20042 31340
rect 20441 31331 20499 31337
rect 20441 31328 20453 31331
rect 20036 31300 20453 31328
rect 20036 31288 20042 31300
rect 20441 31297 20453 31300
rect 20487 31297 20499 31331
rect 20441 31291 20499 31297
rect 20809 31331 20867 31337
rect 20809 31297 20821 31331
rect 20855 31297 20867 31331
rect 20809 31291 20867 31297
rect 16482 31260 16488 31272
rect 14384 31232 16488 31260
rect 14568 31204 14596 31232
rect 16482 31220 16488 31232
rect 16540 31260 16546 31272
rect 17402 31260 17408 31272
rect 16540 31232 17408 31260
rect 16540 31220 16546 31232
rect 17402 31220 17408 31232
rect 17460 31220 17466 31272
rect 20824 31260 20852 31291
rect 21082 31288 21088 31340
rect 21140 31288 21146 31340
rect 21174 31288 21180 31340
rect 21232 31288 21238 31340
rect 21542 31288 21548 31340
rect 21600 31288 21606 31340
rect 22005 31331 22063 31337
rect 22005 31297 22017 31331
rect 22051 31297 22063 31331
rect 22112 31328 22140 31368
rect 22270 31331 22328 31337
rect 22270 31328 22282 31331
rect 22112 31300 22282 31328
rect 22005 31291 22063 31297
rect 22270 31297 22282 31300
rect 22316 31297 22328 31331
rect 22270 31291 22328 31297
rect 21821 31263 21879 31269
rect 21821 31260 21833 31263
rect 20824 31232 21833 31260
rect 21821 31229 21833 31232
rect 21867 31229 21879 31263
rect 21821 31223 21879 31229
rect 12676 31164 13129 31192
rect 12676 31152 12682 31164
rect 14550 31152 14556 31204
rect 14608 31152 14614 31204
rect 15930 31152 15936 31204
rect 15988 31192 15994 31204
rect 20533 31195 20591 31201
rect 20533 31192 20545 31195
rect 15988 31164 20545 31192
rect 15988 31152 15994 31164
rect 20533 31161 20545 31164
rect 20579 31161 20591 31195
rect 20533 31155 20591 31161
rect 21358 31152 21364 31204
rect 21416 31192 21422 31204
rect 22020 31192 22048 31291
rect 22370 31288 22376 31340
rect 22428 31328 22434 31340
rect 23474 31328 23480 31340
rect 22428 31300 23480 31328
rect 22428 31288 22434 31300
rect 23474 31288 23480 31300
rect 23532 31288 23538 31340
rect 23753 31331 23811 31337
rect 23753 31297 23765 31331
rect 23799 31328 23811 31331
rect 23842 31328 23848 31340
rect 23799 31300 23848 31328
rect 23799 31297 23811 31300
rect 23753 31291 23811 31297
rect 23842 31288 23848 31300
rect 23900 31288 23906 31340
rect 24026 31288 24032 31340
rect 24084 31328 24090 31340
rect 24121 31331 24179 31337
rect 24121 31328 24133 31331
rect 24084 31300 24133 31328
rect 24084 31288 24090 31300
rect 24121 31297 24133 31300
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 24210 31288 24216 31340
rect 24268 31328 24274 31340
rect 24397 31331 24455 31337
rect 24397 31328 24409 31331
rect 24268 31300 24409 31328
rect 24268 31288 24274 31300
rect 24397 31297 24409 31300
rect 24443 31297 24455 31331
rect 24492 31328 24520 31368
rect 24670 31356 24676 31408
rect 24728 31396 24734 31408
rect 24949 31399 25007 31405
rect 24949 31396 24961 31399
rect 24728 31368 24961 31396
rect 24728 31356 24734 31368
rect 24949 31365 24961 31368
rect 24995 31365 25007 31399
rect 24949 31359 25007 31365
rect 25682 31356 25688 31408
rect 25740 31396 25746 31408
rect 25740 31368 25912 31396
rect 25740 31356 25746 31368
rect 24492 31300 24716 31328
rect 24397 31291 24455 31297
rect 24688 31272 24716 31300
rect 24762 31288 24768 31340
rect 24820 31331 24826 31340
rect 24820 31288 24834 31331
rect 25038 31288 25044 31340
rect 25096 31288 25102 31340
rect 25130 31288 25136 31340
rect 25188 31288 25194 31340
rect 25590 31288 25596 31340
rect 25648 31288 25654 31340
rect 25774 31288 25780 31340
rect 25832 31288 25838 31340
rect 25884 31328 25912 31368
rect 25958 31356 25964 31408
rect 26016 31396 26022 31408
rect 27154 31396 27160 31408
rect 26016 31368 27160 31396
rect 26016 31356 26022 31368
rect 26050 31328 26056 31340
rect 25884 31300 26056 31328
rect 26050 31288 26056 31300
rect 26108 31288 26114 31340
rect 26160 31337 26188 31368
rect 27154 31356 27160 31368
rect 27212 31396 27218 31408
rect 27614 31396 27620 31408
rect 27212 31368 27620 31396
rect 27212 31356 27218 31368
rect 27614 31356 27620 31368
rect 27672 31396 27678 31408
rect 27709 31399 27767 31405
rect 27709 31396 27721 31399
rect 27672 31368 27721 31396
rect 27672 31356 27678 31368
rect 27709 31365 27721 31368
rect 27755 31365 27767 31399
rect 28718 31396 28724 31408
rect 27709 31359 27767 31365
rect 28276 31368 28724 31396
rect 28276 31340 28304 31368
rect 28718 31356 28724 31368
rect 28776 31356 28782 31408
rect 29840 31396 29868 31436
rect 31018 31424 31024 31436
rect 31076 31424 31082 31476
rect 31202 31424 31208 31476
rect 31260 31464 31266 31476
rect 33965 31467 34023 31473
rect 33965 31464 33977 31467
rect 31260 31436 33977 31464
rect 31260 31424 31266 31436
rect 33965 31433 33977 31436
rect 34011 31433 34023 31467
rect 33965 31427 34023 31433
rect 31294 31396 31300 31408
rect 29012 31368 29408 31396
rect 26145 31331 26203 31337
rect 26145 31297 26157 31331
rect 26191 31297 26203 31331
rect 26145 31291 26203 31297
rect 26234 31288 26240 31340
rect 26292 31288 26298 31340
rect 26421 31331 26479 31337
rect 26421 31297 26433 31331
rect 26467 31297 26479 31331
rect 26421 31291 26479 31297
rect 22094 31220 22100 31272
rect 22152 31220 22158 31272
rect 22189 31263 22247 31269
rect 22189 31229 22201 31263
rect 22235 31260 22247 31263
rect 22554 31260 22560 31272
rect 22235 31232 22560 31260
rect 22235 31229 22247 31232
rect 22189 31223 22247 31229
rect 22554 31220 22560 31232
rect 22612 31220 22618 31272
rect 22664 31232 23796 31260
rect 22664 31192 22692 31232
rect 21416 31164 22692 31192
rect 21416 31152 21422 31164
rect 23106 31152 23112 31204
rect 23164 31192 23170 31204
rect 23382 31192 23388 31204
rect 23164 31164 23388 31192
rect 23164 31152 23170 31164
rect 23382 31152 23388 31164
rect 23440 31152 23446 31204
rect 23658 31152 23664 31204
rect 23716 31152 23722 31204
rect 23768 31192 23796 31232
rect 24670 31220 24676 31272
rect 24728 31220 24734 31272
rect 24806 31260 24834 31288
rect 26252 31260 26280 31288
rect 24806 31232 26280 31260
rect 26436 31260 26464 31291
rect 26510 31288 26516 31340
rect 26568 31328 26574 31340
rect 26605 31331 26663 31337
rect 26605 31328 26617 31331
rect 26568 31300 26617 31328
rect 26568 31288 26574 31300
rect 26605 31297 26617 31300
rect 26651 31297 26663 31331
rect 26605 31291 26663 31297
rect 26973 31331 27031 31337
rect 26973 31297 26985 31331
rect 27019 31328 27031 31331
rect 27985 31331 28043 31337
rect 27985 31328 27997 31331
rect 27019 31300 27997 31328
rect 27019 31297 27031 31300
rect 26973 31291 27031 31297
rect 27985 31297 27997 31300
rect 28031 31328 28043 31331
rect 28258 31328 28264 31340
rect 28031 31300 28264 31328
rect 28031 31297 28043 31300
rect 27985 31291 28043 31297
rect 28258 31288 28264 31300
rect 28316 31288 28322 31340
rect 28534 31288 28540 31340
rect 28592 31288 28598 31340
rect 29012 31337 29040 31368
rect 29380 31340 29408 31368
rect 29748 31368 29868 31396
rect 31036 31368 31300 31396
rect 28997 31331 29055 31337
rect 28997 31297 29009 31331
rect 29043 31297 29055 31331
rect 28997 31291 29055 31297
rect 29086 31288 29092 31340
rect 29144 31328 29150 31340
rect 29273 31331 29331 31337
rect 29273 31328 29285 31331
rect 29144 31300 29285 31328
rect 29144 31288 29150 31300
rect 29273 31297 29285 31300
rect 29319 31297 29331 31331
rect 29273 31291 29331 31297
rect 29362 31288 29368 31340
rect 29420 31328 29426 31340
rect 29641 31331 29699 31337
rect 29641 31328 29653 31331
rect 29420 31300 29653 31328
rect 29420 31288 29426 31300
rect 29641 31297 29653 31300
rect 29687 31297 29699 31331
rect 29641 31291 29699 31297
rect 26436 31232 27568 31260
rect 26234 31192 26240 31204
rect 23768 31164 26240 31192
rect 26234 31152 26240 31164
rect 26292 31152 26298 31204
rect 6512 31096 9168 31124
rect 6512 31084 6518 31096
rect 9858 31084 9864 31136
rect 9916 31084 9922 31136
rect 10042 31084 10048 31136
rect 10100 31124 10106 31136
rect 10410 31124 10416 31136
rect 10100 31096 10416 31124
rect 10100 31084 10106 31096
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10502 31084 10508 31136
rect 10560 31124 10566 31136
rect 11238 31124 11244 31136
rect 10560 31096 11244 31124
rect 10560 31084 10566 31096
rect 11238 31084 11244 31096
rect 11296 31084 11302 31136
rect 11422 31084 11428 31136
rect 11480 31124 11486 31136
rect 11790 31124 11796 31136
rect 11480 31096 11796 31124
rect 11480 31084 11486 31096
rect 11790 31084 11796 31096
rect 11848 31084 11854 31136
rect 12342 31084 12348 31136
rect 12400 31124 12406 31136
rect 13265 31127 13323 31133
rect 13265 31124 13277 31127
rect 12400 31096 13277 31124
rect 12400 31084 12406 31096
rect 13265 31093 13277 31096
rect 13311 31093 13323 31127
rect 13265 31087 13323 31093
rect 14737 31127 14795 31133
rect 14737 31093 14749 31127
rect 14783 31124 14795 31127
rect 16114 31124 16120 31136
rect 14783 31096 16120 31124
rect 14783 31093 14795 31096
rect 14737 31087 14795 31093
rect 16114 31084 16120 31096
rect 16172 31084 16178 31136
rect 19242 31084 19248 31136
rect 19300 31124 19306 31136
rect 24486 31124 24492 31136
rect 19300 31096 24492 31124
rect 19300 31084 19306 31096
rect 24486 31084 24492 31096
rect 24544 31084 24550 31136
rect 24946 31084 24952 31136
rect 25004 31124 25010 31136
rect 25130 31124 25136 31136
rect 25004 31096 25136 31124
rect 25004 31084 25010 31096
rect 25130 31084 25136 31096
rect 25188 31084 25194 31136
rect 25314 31084 25320 31136
rect 25372 31084 25378 31136
rect 25590 31084 25596 31136
rect 25648 31124 25654 31136
rect 26436 31124 26464 31232
rect 27540 31204 27568 31232
rect 28074 31220 28080 31272
rect 28132 31260 28138 31272
rect 28445 31263 28503 31269
rect 28445 31260 28457 31263
rect 28132 31232 28457 31260
rect 28132 31220 28138 31232
rect 28445 31229 28457 31232
rect 28491 31229 28503 31263
rect 28445 31223 28503 31229
rect 27522 31152 27528 31204
rect 27580 31152 27586 31204
rect 28552 31192 28580 31288
rect 28718 31220 28724 31272
rect 28776 31260 28782 31272
rect 29748 31260 29776 31368
rect 30190 31288 30196 31340
rect 30248 31288 30254 31340
rect 30834 31288 30840 31340
rect 30892 31328 30898 31340
rect 31036 31337 31064 31368
rect 31294 31356 31300 31368
rect 31352 31356 31358 31408
rect 33505 31399 33563 31405
rect 33505 31365 33517 31399
rect 33551 31396 33563 31399
rect 33594 31396 33600 31408
rect 33551 31368 33600 31396
rect 33551 31365 33563 31368
rect 33505 31359 33563 31365
rect 33594 31356 33600 31368
rect 33652 31356 33658 31408
rect 31021 31331 31079 31337
rect 31021 31328 31033 31331
rect 30892 31300 31033 31328
rect 30892 31288 30898 31300
rect 31021 31297 31033 31300
rect 31067 31297 31079 31331
rect 31021 31291 31079 31297
rect 31202 31288 31208 31340
rect 31260 31328 31266 31340
rect 32398 31328 32404 31340
rect 31260 31300 32404 31328
rect 31260 31288 31266 31300
rect 32398 31288 32404 31300
rect 32456 31288 32462 31340
rect 32766 31288 32772 31340
rect 32824 31328 32830 31340
rect 33781 31331 33839 31337
rect 33781 31328 33793 31331
rect 32824 31300 33793 31328
rect 32824 31288 32830 31300
rect 33781 31297 33793 31300
rect 33827 31297 33839 31331
rect 33781 31291 33839 31297
rect 28776 31232 29776 31260
rect 28776 31220 28782 31232
rect 29822 31220 29828 31272
rect 29880 31260 29886 31272
rect 30101 31263 30159 31269
rect 30101 31260 30113 31263
rect 29880 31232 30113 31260
rect 29880 31220 29886 31232
rect 30101 31229 30113 31232
rect 30147 31229 30159 31263
rect 31938 31260 31944 31272
rect 30101 31223 30159 31229
rect 31726 31232 31944 31260
rect 31726 31192 31754 31232
rect 31938 31220 31944 31232
rect 31996 31260 32002 31272
rect 32950 31260 32956 31272
rect 31996 31232 32956 31260
rect 31996 31220 32002 31232
rect 32950 31220 32956 31232
rect 33008 31220 33014 31272
rect 33502 31220 33508 31272
rect 33560 31260 33566 31272
rect 33597 31263 33655 31269
rect 33597 31260 33609 31263
rect 33560 31232 33609 31260
rect 33560 31220 33566 31232
rect 33597 31229 33609 31232
rect 33643 31229 33655 31263
rect 33597 31223 33655 31229
rect 28552 31164 31754 31192
rect 25648 31096 26464 31124
rect 25648 31084 25654 31096
rect 26694 31084 26700 31136
rect 26752 31124 26758 31136
rect 30098 31124 30104 31136
rect 26752 31096 30104 31124
rect 26752 31084 26758 31096
rect 30098 31084 30104 31096
rect 30156 31084 30162 31136
rect 33778 31084 33784 31136
rect 33836 31084 33842 31136
rect 1104 31034 41400 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 41400 31034
rect 1104 30960 41400 30982
rect 7282 30880 7288 30932
rect 7340 30880 7346 30932
rect 9582 30920 9588 30932
rect 7484 30892 9588 30920
rect 7300 30852 7328 30880
rect 6104 30824 7328 30852
rect 4157 30787 4215 30793
rect 4157 30753 4169 30787
rect 4203 30784 4215 30787
rect 4522 30784 4528 30796
rect 4203 30756 4528 30784
rect 4203 30753 4215 30756
rect 4157 30747 4215 30753
rect 4522 30744 4528 30756
rect 4580 30744 4586 30796
rect 5442 30676 5448 30728
rect 5500 30716 5506 30728
rect 6104 30716 6132 30824
rect 6178 30744 6184 30796
rect 6236 30784 6242 30796
rect 6236 30756 6684 30784
rect 6236 30744 6242 30756
rect 5500 30688 6132 30716
rect 5500 30676 5506 30688
rect 6270 30676 6276 30728
rect 6328 30676 6334 30728
rect 6454 30676 6460 30728
rect 6512 30676 6518 30728
rect 6656 30725 6684 30756
rect 6641 30719 6699 30725
rect 6641 30685 6653 30719
rect 6687 30685 6699 30719
rect 6641 30679 6699 30685
rect 7190 30676 7196 30728
rect 7248 30676 7254 30728
rect 4433 30651 4491 30657
rect 4433 30617 4445 30651
rect 4479 30617 4491 30651
rect 4433 30611 4491 30617
rect 4448 30580 4476 30611
rect 6178 30608 6184 30660
rect 6236 30648 6242 30660
rect 6549 30651 6607 30657
rect 6549 30648 6561 30651
rect 6236 30620 6561 30648
rect 6236 30608 6242 30620
rect 6549 30617 6561 30620
rect 6595 30648 6607 30651
rect 7484 30648 7512 30892
rect 9582 30880 9588 30892
rect 9640 30880 9646 30932
rect 9769 30923 9827 30929
rect 9769 30889 9781 30923
rect 9815 30889 9827 30923
rect 9769 30883 9827 30889
rect 10137 30923 10195 30929
rect 10137 30889 10149 30923
rect 10183 30920 10195 30923
rect 10962 30920 10968 30932
rect 10183 30892 10968 30920
rect 10183 30889 10195 30892
rect 10137 30883 10195 30889
rect 9784 30852 9812 30883
rect 10962 30880 10968 30892
rect 11020 30880 11026 30932
rect 12342 30880 12348 30932
rect 12400 30880 12406 30932
rect 12710 30880 12716 30932
rect 12768 30920 12774 30932
rect 15838 30920 15844 30932
rect 12768 30892 15844 30920
rect 12768 30880 12774 30892
rect 15838 30880 15844 30892
rect 15896 30880 15902 30932
rect 16390 30880 16396 30932
rect 16448 30920 16454 30932
rect 16485 30923 16543 30929
rect 16485 30920 16497 30923
rect 16448 30892 16497 30920
rect 16448 30880 16454 30892
rect 16485 30889 16497 30892
rect 16531 30889 16543 30923
rect 16485 30883 16543 30889
rect 16942 30880 16948 30932
rect 17000 30920 17006 30932
rect 17681 30923 17739 30929
rect 17000 30892 17633 30920
rect 17000 30880 17006 30892
rect 9784 30824 10180 30852
rect 7558 30744 7564 30796
rect 7616 30784 7622 30796
rect 9677 30787 9735 30793
rect 7616 30756 9628 30784
rect 7616 30744 7622 30756
rect 9401 30719 9459 30725
rect 9401 30716 9413 30719
rect 6595 30620 7512 30648
rect 8956 30688 9413 30716
rect 6595 30617 6607 30620
rect 6549 30611 6607 30617
rect 8956 30592 8984 30688
rect 9401 30685 9413 30688
rect 9447 30685 9459 30719
rect 9600 30716 9628 30756
rect 9677 30753 9689 30787
rect 9723 30784 9735 30787
rect 9950 30784 9956 30796
rect 9723 30756 9956 30784
rect 9723 30753 9735 30756
rect 9677 30747 9735 30753
rect 9950 30744 9956 30756
rect 10008 30744 10014 30796
rect 10152 30784 10180 30824
rect 10686 30812 10692 30864
rect 10744 30852 10750 30864
rect 10744 30824 11836 30852
rect 10744 30812 10750 30824
rect 10778 30784 10784 30796
rect 10152 30756 10784 30784
rect 10778 30744 10784 30756
rect 10836 30744 10842 30796
rect 11422 30744 11428 30796
rect 11480 30744 11486 30796
rect 10045 30719 10103 30725
rect 10045 30716 10057 30719
rect 9600 30688 10057 30716
rect 9401 30679 9459 30685
rect 10045 30685 10057 30688
rect 10091 30685 10103 30719
rect 10045 30679 10103 30685
rect 10229 30719 10287 30725
rect 10229 30685 10241 30719
rect 10275 30716 10287 30719
rect 10962 30716 10968 30728
rect 10275 30688 10968 30716
rect 10275 30685 10287 30688
rect 10229 30679 10287 30685
rect 9030 30608 9036 30660
rect 9088 30648 9094 30660
rect 9582 30648 9588 30660
rect 9088 30620 9588 30648
rect 9088 30608 9094 30620
rect 9582 30608 9588 30620
rect 9640 30608 9646 30660
rect 10060 30648 10088 30679
rect 10962 30676 10968 30688
rect 11020 30676 11026 30728
rect 11330 30676 11336 30728
rect 11388 30676 11394 30728
rect 11808 30725 11836 30824
rect 12360 30725 12388 30880
rect 15102 30852 15108 30864
rect 14292 30824 15108 30852
rect 12636 30756 13768 30784
rect 12636 30725 12664 30756
rect 13740 30728 13768 30756
rect 14292 30728 14320 30824
rect 15102 30812 15108 30824
rect 15160 30852 15166 30864
rect 17218 30852 17224 30864
rect 15160 30824 17224 30852
rect 15160 30812 15166 30824
rect 17218 30812 17224 30824
rect 17276 30812 17282 30864
rect 17605 30852 17633 30892
rect 17681 30889 17693 30923
rect 17727 30920 17739 30923
rect 18322 30920 18328 30932
rect 17727 30892 18328 30920
rect 17727 30889 17739 30892
rect 17681 30883 17739 30889
rect 18322 30880 18328 30892
rect 18380 30880 18386 30932
rect 19242 30880 19248 30932
rect 19300 30880 19306 30932
rect 22186 30880 22192 30932
rect 22244 30920 22250 30932
rect 22462 30920 22468 30932
rect 22244 30892 22468 30920
rect 22244 30880 22250 30892
rect 22462 30880 22468 30892
rect 22520 30880 22526 30932
rect 22554 30880 22560 30932
rect 22612 30920 22618 30932
rect 23106 30920 23112 30932
rect 22612 30892 23112 30920
rect 22612 30880 22618 30892
rect 23106 30880 23112 30892
rect 23164 30880 23170 30932
rect 24302 30880 24308 30932
rect 24360 30920 24366 30932
rect 24946 30920 24952 30932
rect 24360 30892 24952 30920
rect 24360 30880 24366 30892
rect 24946 30880 24952 30892
rect 25004 30920 25010 30932
rect 25590 30920 25596 30932
rect 25004 30892 25596 30920
rect 25004 30880 25010 30892
rect 25590 30880 25596 30892
rect 25648 30880 25654 30932
rect 26050 30880 26056 30932
rect 26108 30880 26114 30932
rect 26234 30880 26240 30932
rect 26292 30880 26298 30932
rect 26602 30880 26608 30932
rect 26660 30880 26666 30932
rect 27154 30880 27160 30932
rect 27212 30920 27218 30932
rect 28718 30920 28724 30932
rect 27212 30892 28724 30920
rect 27212 30880 27218 30892
rect 28718 30880 28724 30892
rect 28776 30920 28782 30932
rect 28905 30923 28963 30929
rect 28905 30920 28917 30923
rect 28776 30892 28917 30920
rect 28776 30880 28782 30892
rect 28905 30889 28917 30892
rect 28951 30889 28963 30923
rect 28905 30883 28963 30889
rect 28994 30880 29000 30932
rect 29052 30920 29058 30932
rect 29181 30923 29239 30929
rect 29181 30920 29193 30923
rect 29052 30892 29193 30920
rect 29052 30880 29058 30892
rect 29181 30889 29193 30892
rect 29227 30920 29239 30923
rect 29641 30923 29699 30929
rect 29641 30920 29653 30923
rect 29227 30892 29653 30920
rect 29227 30889 29239 30892
rect 29181 30883 29239 30889
rect 29641 30889 29653 30892
rect 29687 30889 29699 30923
rect 29641 30883 29699 30889
rect 18049 30855 18107 30861
rect 18049 30852 18061 30855
rect 17605 30824 18061 30852
rect 18049 30821 18061 30824
rect 18095 30852 18107 30855
rect 19260 30852 19288 30880
rect 18095 30824 19288 30852
rect 18095 30821 18107 30824
rect 18049 30815 18107 30821
rect 20254 30812 20260 30864
rect 20312 30852 20318 30864
rect 21266 30852 21272 30864
rect 20312 30824 21272 30852
rect 20312 30812 20318 30824
rect 21266 30812 21272 30824
rect 21324 30812 21330 30864
rect 22278 30812 22284 30864
rect 22336 30852 22342 30864
rect 22572 30852 22600 30880
rect 22336 30824 22600 30852
rect 22664 30824 24256 30852
rect 22336 30812 22342 30824
rect 14550 30744 14556 30796
rect 14608 30784 14614 30796
rect 14918 30784 14924 30796
rect 14608 30756 14924 30784
rect 14608 30744 14614 30756
rect 14918 30744 14924 30756
rect 14976 30744 14982 30796
rect 17236 30784 17264 30812
rect 15120 30756 15700 30784
rect 11793 30719 11851 30725
rect 11793 30685 11805 30719
rect 11839 30685 11851 30719
rect 11793 30679 11851 30685
rect 12345 30719 12403 30725
rect 12345 30685 12357 30719
rect 12391 30685 12403 30719
rect 12345 30679 12403 30685
rect 12621 30719 12679 30725
rect 12621 30685 12633 30719
rect 12667 30685 12679 30719
rect 12621 30679 12679 30685
rect 12802 30676 12808 30728
rect 12860 30716 12866 30728
rect 12989 30719 13047 30725
rect 12989 30716 13001 30719
rect 12860 30688 13001 30716
rect 12860 30676 12866 30688
rect 12989 30685 13001 30688
rect 13035 30685 13047 30719
rect 12989 30679 13047 30685
rect 13722 30676 13728 30728
rect 13780 30676 13786 30728
rect 14274 30676 14280 30728
rect 14332 30676 14338 30728
rect 15120 30648 15148 30756
rect 15197 30719 15255 30725
rect 15197 30685 15209 30719
rect 15243 30685 15255 30719
rect 15197 30679 15255 30685
rect 15381 30719 15439 30725
rect 15381 30685 15393 30719
rect 15427 30716 15439 30719
rect 15562 30716 15568 30728
rect 15427 30688 15568 30716
rect 15427 30685 15439 30688
rect 15381 30679 15439 30685
rect 10060 30620 15148 30648
rect 15212 30648 15240 30679
rect 15562 30676 15568 30688
rect 15620 30676 15626 30728
rect 15672 30716 15700 30756
rect 16224 30756 16712 30784
rect 17236 30756 17632 30784
rect 16224 30716 16252 30756
rect 15672 30688 16252 30716
rect 15930 30648 15936 30660
rect 15212 30620 15936 30648
rect 15930 30608 15936 30620
rect 15988 30608 15994 30660
rect 16224 30657 16252 30688
rect 16482 30676 16488 30728
rect 16540 30676 16546 30728
rect 16684 30725 16712 30756
rect 16669 30719 16727 30725
rect 16669 30685 16681 30719
rect 16715 30716 16727 30719
rect 17494 30716 17500 30728
rect 16715 30688 17500 30716
rect 16715 30685 16727 30688
rect 16669 30679 16727 30685
rect 17494 30676 17500 30688
rect 17552 30676 17558 30728
rect 17604 30716 17632 30756
rect 17678 30744 17684 30796
rect 17736 30784 17742 30796
rect 18874 30784 18880 30796
rect 17736 30756 18880 30784
rect 17736 30744 17742 30756
rect 18874 30744 18880 30756
rect 18932 30744 18938 30796
rect 22664 30784 22692 30824
rect 24228 30784 24256 30824
rect 24486 30812 24492 30864
rect 24544 30812 24550 30864
rect 26973 30855 27031 30861
rect 26973 30852 26985 30855
rect 24596 30824 26985 30852
rect 24596 30784 24624 30824
rect 26973 30821 26985 30824
rect 27019 30821 27031 30855
rect 26973 30815 27031 30821
rect 27338 30812 27344 30864
rect 27396 30852 27402 30864
rect 28629 30855 28687 30861
rect 28629 30852 28641 30855
rect 27396 30824 28641 30852
rect 27396 30812 27402 30824
rect 28629 30821 28641 30824
rect 28675 30821 28687 30855
rect 28629 30815 28687 30821
rect 29362 30812 29368 30864
rect 29420 30812 29426 30864
rect 29546 30812 29552 30864
rect 29604 30812 29610 30864
rect 25958 30784 25964 30796
rect 19444 30756 22692 30784
rect 22940 30756 24164 30784
rect 24228 30756 24624 30784
rect 24780 30756 25964 30784
rect 19444 30728 19472 30756
rect 17865 30719 17923 30725
rect 17865 30716 17877 30719
rect 17604 30688 17877 30716
rect 17865 30685 17877 30688
rect 17911 30685 17923 30719
rect 17865 30679 17923 30685
rect 18141 30719 18199 30725
rect 18141 30685 18153 30719
rect 18187 30716 18199 30719
rect 18414 30716 18420 30728
rect 18187 30688 18420 30716
rect 18187 30685 18199 30688
rect 18141 30679 18199 30685
rect 18414 30676 18420 30688
rect 18472 30676 18478 30728
rect 18690 30676 18696 30728
rect 18748 30716 18754 30728
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 18748 30688 19257 30716
rect 18748 30676 18754 30688
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19426 30676 19432 30728
rect 19484 30676 19490 30728
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 19978 30716 19984 30728
rect 19751 30688 19984 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 19978 30676 19984 30688
rect 20036 30676 20042 30728
rect 21468 30725 21496 30756
rect 21453 30719 21511 30725
rect 21453 30685 21465 30719
rect 21499 30685 21511 30719
rect 21453 30679 21511 30685
rect 21542 30676 21548 30728
rect 21600 30716 21606 30728
rect 21910 30716 21916 30728
rect 21600 30688 21916 30716
rect 21600 30676 21606 30688
rect 21910 30676 21916 30688
rect 21968 30676 21974 30728
rect 22738 30676 22744 30728
rect 22796 30676 22802 30728
rect 22940 30725 22968 30756
rect 23768 30725 23796 30756
rect 22925 30719 22983 30725
rect 22925 30685 22937 30719
rect 22971 30685 22983 30719
rect 22925 30679 22983 30685
rect 23109 30719 23167 30725
rect 23109 30685 23121 30719
rect 23155 30685 23167 30719
rect 23109 30679 23167 30685
rect 23201 30719 23259 30725
rect 23201 30685 23213 30719
rect 23247 30716 23259 30719
rect 23753 30719 23811 30725
rect 23247 30688 23337 30716
rect 23247 30685 23259 30688
rect 23201 30679 23259 30685
rect 16025 30651 16083 30657
rect 16025 30617 16037 30651
rect 16071 30617 16083 30651
rect 16025 30611 16083 30617
rect 16209 30651 16267 30657
rect 16209 30617 16221 30651
rect 16255 30617 16267 30651
rect 18230 30648 18236 30660
rect 16209 30611 16267 30617
rect 16316 30620 18236 30648
rect 6825 30583 6883 30589
rect 6825 30580 6837 30583
rect 4448 30552 6837 30580
rect 6825 30549 6837 30552
rect 6871 30549 6883 30583
rect 6825 30543 6883 30549
rect 8938 30540 8944 30592
rect 8996 30540 9002 30592
rect 9950 30540 9956 30592
rect 10008 30540 10014 30592
rect 10410 30540 10416 30592
rect 10468 30580 10474 30592
rect 11330 30580 11336 30592
rect 10468 30552 11336 30580
rect 10468 30540 10474 30552
rect 11330 30540 11336 30552
rect 11388 30540 11394 30592
rect 15010 30540 15016 30592
rect 15068 30580 15074 30592
rect 15289 30583 15347 30589
rect 15289 30580 15301 30583
rect 15068 30552 15301 30580
rect 15068 30540 15074 30552
rect 15289 30549 15301 30552
rect 15335 30549 15347 30583
rect 16040 30580 16068 30611
rect 16316 30580 16344 30620
rect 18230 30608 18236 30620
rect 18288 30608 18294 30660
rect 19794 30608 19800 30660
rect 19852 30648 19858 30660
rect 20254 30648 20260 30660
rect 19852 30620 20260 30648
rect 19852 30608 19858 30620
rect 20254 30608 20260 30620
rect 20312 30608 20318 30660
rect 22756 30648 22784 30676
rect 23014 30648 23020 30660
rect 22756 30620 23020 30648
rect 23014 30608 23020 30620
rect 23072 30648 23078 30660
rect 23124 30648 23152 30679
rect 23072 30620 23152 30648
rect 23072 30608 23078 30620
rect 16040 30552 16344 30580
rect 15289 30543 15347 30549
rect 16390 30540 16396 30592
rect 16448 30540 16454 30592
rect 17770 30540 17776 30592
rect 17828 30580 17834 30592
rect 21358 30580 21364 30592
rect 17828 30552 21364 30580
rect 17828 30540 17834 30552
rect 21358 30540 21364 30552
rect 21416 30540 21422 30592
rect 22738 30540 22744 30592
rect 22796 30540 22802 30592
rect 23309 30580 23337 30688
rect 23753 30685 23765 30719
rect 23799 30685 23811 30719
rect 23753 30679 23811 30685
rect 24026 30676 24032 30728
rect 24084 30676 24090 30728
rect 24136 30716 24164 30756
rect 24581 30719 24639 30725
rect 24581 30716 24593 30719
rect 24136 30688 24593 30716
rect 24581 30685 24593 30688
rect 24627 30716 24639 30719
rect 24780 30716 24808 30756
rect 25958 30744 25964 30756
rect 26016 30744 26022 30796
rect 26421 30787 26479 30793
rect 26421 30784 26433 30787
rect 26068 30756 26433 30784
rect 24627 30688 24808 30716
rect 24627 30685 24639 30688
rect 24581 30679 24639 30685
rect 24946 30676 24952 30728
rect 25004 30676 25010 30728
rect 25225 30719 25283 30725
rect 25225 30685 25237 30719
rect 25271 30685 25283 30719
rect 25225 30679 25283 30685
rect 24213 30651 24271 30657
rect 24213 30617 24225 30651
rect 24259 30648 24271 30651
rect 24670 30648 24676 30660
rect 24259 30620 24676 30648
rect 24259 30617 24271 30620
rect 24213 30611 24271 30617
rect 24670 30608 24676 30620
rect 24728 30608 24734 30660
rect 25240 30580 25268 30679
rect 25866 30676 25872 30728
rect 25924 30676 25930 30728
rect 26068 30725 26096 30756
rect 26421 30753 26433 30756
rect 26467 30753 26479 30787
rect 26421 30747 26479 30753
rect 26528 30756 27660 30784
rect 26528 30728 26556 30756
rect 27632 30728 27660 30756
rect 27798 30744 27804 30796
rect 27856 30744 27862 30796
rect 29089 30787 29147 30793
rect 29089 30753 29101 30787
rect 29135 30784 29147 30787
rect 29380 30784 29408 30812
rect 29135 30756 29408 30784
rect 29135 30753 29147 30756
rect 29089 30747 29147 30753
rect 26053 30719 26111 30725
rect 26053 30685 26065 30719
rect 26099 30685 26111 30719
rect 26053 30679 26111 30685
rect 26329 30719 26387 30725
rect 26329 30685 26341 30719
rect 26375 30718 26387 30719
rect 26375 30690 26453 30718
rect 26375 30685 26387 30690
rect 26329 30679 26387 30685
rect 25590 30608 25596 30660
rect 25648 30608 25654 30660
rect 26425 30648 26453 30690
rect 26510 30676 26516 30728
rect 26568 30676 26574 30728
rect 26602 30676 26608 30728
rect 26660 30676 26666 30728
rect 26694 30676 26700 30728
rect 26752 30676 26758 30728
rect 26789 30719 26847 30725
rect 26789 30685 26801 30719
rect 26835 30716 26847 30719
rect 26835 30688 27568 30716
rect 26835 30685 26847 30688
rect 26789 30679 26847 30685
rect 26712 30648 26740 30676
rect 26425 30620 26740 30648
rect 26878 30608 26884 30660
rect 26936 30648 26942 30660
rect 27157 30651 27215 30657
rect 27157 30648 27169 30651
rect 26936 30620 27169 30648
rect 26936 30608 26942 30620
rect 27157 30617 27169 30620
rect 27203 30617 27215 30651
rect 27157 30611 27215 30617
rect 27430 30608 27436 30660
rect 27488 30608 27494 30660
rect 27540 30657 27568 30688
rect 27614 30676 27620 30728
rect 27672 30676 27678 30728
rect 27706 30676 27712 30728
rect 27764 30716 27770 30728
rect 28166 30716 28172 30728
rect 27764 30688 28172 30716
rect 27764 30676 27770 30688
rect 28166 30676 28172 30688
rect 28224 30716 28230 30728
rect 28353 30719 28411 30725
rect 28353 30716 28365 30719
rect 28224 30688 28365 30716
rect 28224 30676 28230 30688
rect 28353 30685 28365 30688
rect 28399 30685 28411 30719
rect 28353 30679 28411 30685
rect 28629 30719 28687 30725
rect 28629 30685 28641 30719
rect 28675 30685 28687 30719
rect 28629 30679 28687 30685
rect 27525 30651 27583 30657
rect 27525 30617 27537 30651
rect 27571 30617 27583 30651
rect 28644 30648 28672 30679
rect 28810 30676 28816 30728
rect 28868 30676 28874 30728
rect 29181 30719 29239 30725
rect 29181 30685 29193 30719
rect 29227 30685 29239 30719
rect 29181 30679 29239 30685
rect 29196 30648 29224 30679
rect 29362 30676 29368 30728
rect 29420 30676 29426 30728
rect 29564 30725 29592 30812
rect 29638 30744 29644 30796
rect 29696 30784 29702 30796
rect 29825 30787 29883 30793
rect 29825 30784 29837 30787
rect 29696 30756 29837 30784
rect 29696 30744 29702 30756
rect 29825 30753 29837 30756
rect 29871 30753 29883 30787
rect 29825 30747 29883 30753
rect 32674 30744 32680 30796
rect 32732 30784 32738 30796
rect 33597 30787 33655 30793
rect 33597 30784 33609 30787
rect 32732 30756 33609 30784
rect 32732 30744 32738 30756
rect 33597 30753 33609 30756
rect 33643 30753 33655 30787
rect 33597 30747 33655 30753
rect 34054 30744 34060 30796
rect 34112 30784 34118 30796
rect 35529 30787 35587 30793
rect 35529 30784 35541 30787
rect 34112 30756 35541 30784
rect 34112 30744 34118 30756
rect 35529 30753 35541 30756
rect 35575 30753 35587 30787
rect 35529 30747 35587 30753
rect 29549 30719 29607 30725
rect 29549 30685 29561 30719
rect 29595 30685 29607 30719
rect 29549 30679 29607 30685
rect 31202 30676 31208 30728
rect 31260 30676 31266 30728
rect 33413 30719 33471 30725
rect 33413 30685 33425 30719
rect 33459 30716 33471 30719
rect 33502 30716 33508 30728
rect 33459 30688 33508 30716
rect 33459 30685 33471 30688
rect 33413 30679 33471 30685
rect 33502 30676 33508 30688
rect 33560 30676 33566 30728
rect 35253 30719 35311 30725
rect 35253 30685 35265 30719
rect 35299 30716 35311 30719
rect 35434 30716 35440 30728
rect 35299 30688 35440 30716
rect 35299 30685 35311 30688
rect 35253 30679 35311 30685
rect 35434 30676 35440 30688
rect 35492 30676 35498 30728
rect 31220 30648 31248 30676
rect 28644 30620 29224 30648
rect 27525 30611 27583 30617
rect 26602 30580 26608 30592
rect 23309 30552 26608 30580
rect 26602 30540 26608 30552
rect 26660 30540 26666 30592
rect 26970 30540 26976 30592
rect 27028 30580 27034 30592
rect 27249 30583 27307 30589
rect 27249 30580 27261 30583
rect 27028 30552 27261 30580
rect 27028 30540 27034 30552
rect 27249 30549 27261 30552
rect 27295 30549 27307 30583
rect 27249 30543 27307 30549
rect 27341 30583 27399 30589
rect 27341 30549 27353 30583
rect 27387 30580 27399 30583
rect 27448 30580 27476 30608
rect 27387 30552 27476 30580
rect 27540 30580 27568 30611
rect 27614 30580 27620 30592
rect 27540 30552 27620 30580
rect 27387 30549 27399 30552
rect 27341 30543 27399 30549
rect 27614 30540 27620 30552
rect 27672 30540 27678 30592
rect 29086 30540 29092 30592
rect 29144 30540 29150 30592
rect 29196 30580 29224 30620
rect 29380 30620 31248 30648
rect 29380 30580 29408 30620
rect 32766 30608 32772 30660
rect 32824 30648 32830 30660
rect 32953 30651 33011 30657
rect 32953 30648 32965 30651
rect 32824 30620 32965 30648
rect 32824 30608 32830 30620
rect 32953 30617 32965 30620
rect 32999 30648 33011 30651
rect 32999 30620 33640 30648
rect 32999 30617 33011 30620
rect 32953 30611 33011 30617
rect 29196 30552 29408 30580
rect 29454 30540 29460 30592
rect 29512 30580 29518 30592
rect 29825 30583 29883 30589
rect 29825 30580 29837 30583
rect 29512 30552 29837 30580
rect 29512 30540 29518 30552
rect 29825 30549 29837 30552
rect 29871 30549 29883 30583
rect 29825 30543 29883 30549
rect 31570 30540 31576 30592
rect 31628 30580 31634 30592
rect 33226 30580 33232 30592
rect 31628 30552 33232 30580
rect 31628 30540 31634 30552
rect 33226 30540 33232 30552
rect 33284 30540 33290 30592
rect 33612 30580 33640 30620
rect 33870 30608 33876 30660
rect 33928 30648 33934 30660
rect 34793 30651 34851 30657
rect 33928 30620 34744 30648
rect 33928 30608 33934 30620
rect 34146 30580 34152 30592
rect 33612 30552 34152 30580
rect 34146 30540 34152 30552
rect 34204 30580 34210 30592
rect 34606 30580 34612 30592
rect 34204 30552 34612 30580
rect 34204 30540 34210 30552
rect 34606 30540 34612 30552
rect 34664 30540 34670 30592
rect 34716 30580 34744 30620
rect 34793 30617 34805 30651
rect 34839 30648 34851 30651
rect 34839 30620 35480 30648
rect 34839 30617 34851 30620
rect 34793 30611 34851 30617
rect 34885 30583 34943 30589
rect 34885 30580 34897 30583
rect 34716 30552 34897 30580
rect 34885 30549 34897 30552
rect 34931 30549 34943 30583
rect 35452 30580 35480 30620
rect 35894 30580 35900 30592
rect 35452 30552 35900 30580
rect 34885 30543 34943 30549
rect 35894 30540 35900 30552
rect 35952 30540 35958 30592
rect 1104 30490 41400 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 41400 30490
rect 1104 30416 41400 30438
rect 8478 30336 8484 30388
rect 8536 30376 8542 30388
rect 8665 30379 8723 30385
rect 8665 30376 8677 30379
rect 8536 30348 8677 30376
rect 8536 30336 8542 30348
rect 8665 30345 8677 30348
rect 8711 30345 8723 30379
rect 8665 30339 8723 30345
rect 9674 30336 9680 30388
rect 9732 30376 9738 30388
rect 11054 30376 11060 30388
rect 9732 30348 11060 30376
rect 9732 30336 9738 30348
rect 11054 30336 11060 30348
rect 11112 30336 11118 30388
rect 11241 30379 11299 30385
rect 11241 30345 11253 30379
rect 11287 30376 11299 30379
rect 13998 30376 14004 30388
rect 11287 30348 14004 30376
rect 11287 30345 11299 30348
rect 11241 30339 11299 30345
rect 13998 30336 14004 30348
rect 14056 30336 14062 30388
rect 15654 30376 15660 30388
rect 14752 30348 15660 30376
rect 10873 30311 10931 30317
rect 10873 30308 10885 30311
rect 8496 30280 10885 30308
rect 7650 30200 7656 30252
rect 7708 30240 7714 30252
rect 8496 30249 8524 30280
rect 10873 30277 10885 30280
rect 10919 30277 10931 30311
rect 10873 30271 10931 30277
rect 10965 30311 11023 30317
rect 10965 30277 10977 30311
rect 11011 30308 11023 30311
rect 11072 30308 11100 30336
rect 12250 30308 12256 30320
rect 11011 30280 12256 30308
rect 11011 30277 11023 30280
rect 10965 30271 11023 30277
rect 12250 30268 12256 30280
rect 12308 30268 12314 30320
rect 13722 30268 13728 30320
rect 13780 30308 13786 30320
rect 14752 30308 14780 30348
rect 15654 30336 15660 30348
rect 15712 30336 15718 30388
rect 16025 30379 16083 30385
rect 16025 30345 16037 30379
rect 16071 30376 16083 30379
rect 16390 30376 16396 30388
rect 16071 30348 16396 30376
rect 16071 30345 16083 30348
rect 16025 30339 16083 30345
rect 15562 30308 15568 30320
rect 13780 30280 14780 30308
rect 14844 30280 15568 30308
rect 13780 30268 13786 30280
rect 8481 30243 8539 30249
rect 8481 30240 8493 30243
rect 7708 30212 8493 30240
rect 7708 30200 7714 30212
rect 8481 30209 8493 30212
rect 8527 30209 8539 30243
rect 8481 30203 8539 30209
rect 8941 30243 8999 30249
rect 8941 30209 8953 30243
rect 8987 30209 8999 30243
rect 8941 30203 8999 30209
rect 7926 30132 7932 30184
rect 7984 30172 7990 30184
rect 8754 30172 8760 30184
rect 7984 30144 8760 30172
rect 7984 30132 7990 30144
rect 8754 30132 8760 30144
rect 8812 30172 8818 30184
rect 8956 30172 8984 30203
rect 10410 30200 10416 30252
rect 10468 30240 10474 30252
rect 10597 30243 10655 30249
rect 10597 30240 10609 30243
rect 10468 30212 10609 30240
rect 10468 30200 10474 30212
rect 10597 30209 10609 30212
rect 10643 30209 10655 30243
rect 10597 30203 10655 30209
rect 10686 30200 10692 30252
rect 10744 30240 10750 30252
rect 11062 30243 11120 30249
rect 10744 30212 10789 30240
rect 10744 30200 10750 30212
rect 11062 30209 11074 30243
rect 11108 30209 11120 30243
rect 11062 30203 11120 30209
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30240 11759 30243
rect 11747 30212 11836 30240
rect 11747 30209 11759 30212
rect 11701 30203 11759 30209
rect 10502 30172 10508 30184
rect 8812 30144 8984 30172
rect 9048 30144 10508 30172
rect 8812 30132 8818 30144
rect 8846 30064 8852 30116
rect 8904 30104 8910 30116
rect 9048 30104 9076 30144
rect 10502 30132 10508 30144
rect 10560 30132 10566 30184
rect 11077 30172 11105 30203
rect 10612 30144 11105 30172
rect 10612 30116 10640 30144
rect 11514 30132 11520 30184
rect 11572 30132 11578 30184
rect 8904 30076 9076 30104
rect 8904 30064 8910 30076
rect 9582 30064 9588 30116
rect 9640 30104 9646 30116
rect 10594 30104 10600 30116
rect 9640 30076 10600 30104
rect 9640 30064 9646 30076
rect 10594 30064 10600 30076
rect 10652 30064 10658 30116
rect 11808 30104 11836 30212
rect 11882 30200 11888 30252
rect 11940 30240 11946 30252
rect 11977 30243 12035 30249
rect 11977 30240 11989 30243
rect 11940 30212 11989 30240
rect 11940 30200 11946 30212
rect 11977 30209 11989 30212
rect 12023 30240 12035 30243
rect 12023 30212 12112 30240
rect 12023 30209 12035 30212
rect 11977 30203 12035 30209
rect 12084 30184 12112 30212
rect 12802 30200 12808 30252
rect 12860 30200 12866 30252
rect 12986 30200 12992 30252
rect 13044 30240 13050 30252
rect 13446 30240 13452 30252
rect 13044 30212 13452 30240
rect 13044 30200 13050 30212
rect 13446 30200 13452 30212
rect 13504 30200 13510 30252
rect 14277 30243 14335 30249
rect 14277 30209 14289 30243
rect 14323 30240 14335 30243
rect 14458 30240 14464 30252
rect 14323 30212 14464 30240
rect 14323 30209 14335 30212
rect 14277 30203 14335 30209
rect 14458 30200 14464 30212
rect 14516 30200 14522 30252
rect 14844 30249 14872 30280
rect 15562 30268 15568 30280
rect 15620 30308 15626 30320
rect 16040 30308 16068 30339
rect 16390 30336 16396 30348
rect 16448 30336 16454 30388
rect 18230 30336 18236 30388
rect 18288 30376 18294 30388
rect 18288 30348 19564 30376
rect 18288 30336 18294 30348
rect 15620 30280 16068 30308
rect 15620 30268 15626 30280
rect 16114 30268 16120 30320
rect 16172 30308 16178 30320
rect 16172 30280 16712 30308
rect 16172 30268 16178 30280
rect 14829 30243 14887 30249
rect 14829 30209 14841 30243
rect 14875 30209 14887 30243
rect 14829 30203 14887 30209
rect 14921 30243 14979 30249
rect 14921 30209 14933 30243
rect 14967 30209 14979 30243
rect 14921 30203 14979 30209
rect 15289 30243 15347 30249
rect 15289 30209 15301 30243
rect 15335 30240 15347 30243
rect 15657 30243 15715 30249
rect 15657 30240 15669 30243
rect 15335 30212 15669 30240
rect 15335 30209 15347 30212
rect 15289 30203 15347 30209
rect 15657 30209 15669 30212
rect 15703 30240 15715 30243
rect 16206 30240 16212 30252
rect 15703 30212 16212 30240
rect 15703 30209 15715 30212
rect 15657 30203 15715 30209
rect 12066 30132 12072 30184
rect 12124 30132 12130 30184
rect 12820 30104 12848 30200
rect 13998 30132 14004 30184
rect 14056 30172 14062 30184
rect 14369 30175 14427 30181
rect 14369 30172 14381 30175
rect 14056 30144 14381 30172
rect 14056 30132 14062 30144
rect 14369 30141 14381 30144
rect 14415 30141 14427 30175
rect 14369 30135 14427 30141
rect 11808 30076 12848 30104
rect 14645 30107 14703 30113
rect 14645 30073 14657 30107
rect 14691 30104 14703 30107
rect 14734 30104 14740 30116
rect 14691 30076 14740 30104
rect 14691 30073 14703 30076
rect 14645 30067 14703 30073
rect 14734 30064 14740 30076
rect 14792 30064 14798 30116
rect 14936 30104 14964 30203
rect 16206 30200 16212 30212
rect 16264 30200 16270 30252
rect 16684 30249 16712 30280
rect 16669 30243 16727 30249
rect 16669 30209 16681 30243
rect 16715 30209 16727 30243
rect 16669 30203 16727 30209
rect 16850 30200 16856 30252
rect 16908 30200 16914 30252
rect 18248 30249 18276 30336
rect 18782 30308 18788 30320
rect 18340 30280 18788 30308
rect 18233 30243 18291 30249
rect 18233 30209 18245 30243
rect 18279 30209 18291 30243
rect 18233 30203 18291 30209
rect 18340 30184 18368 30280
rect 18782 30268 18788 30280
rect 18840 30268 18846 30320
rect 19426 30308 19432 30320
rect 19168 30280 19432 30308
rect 19168 30249 19196 30280
rect 19426 30268 19432 30280
rect 19484 30268 19490 30320
rect 19536 30308 19564 30348
rect 22094 30336 22100 30388
rect 22152 30376 22158 30388
rect 22830 30376 22836 30388
rect 22152 30348 22836 30376
rect 22152 30336 22158 30348
rect 22830 30336 22836 30348
rect 22888 30336 22894 30388
rect 23014 30336 23020 30388
rect 23072 30376 23078 30388
rect 25038 30376 25044 30388
rect 23072 30348 25044 30376
rect 23072 30336 23078 30348
rect 25038 30336 25044 30348
rect 25096 30376 25102 30388
rect 25314 30376 25320 30388
rect 25096 30348 25320 30376
rect 25096 30336 25102 30348
rect 25314 30336 25320 30348
rect 25372 30336 25378 30388
rect 25498 30336 25504 30388
rect 25556 30376 25562 30388
rect 26053 30379 26111 30385
rect 26053 30376 26065 30379
rect 25556 30348 26065 30376
rect 25556 30336 25562 30348
rect 26053 30345 26065 30348
rect 26099 30345 26111 30379
rect 26053 30339 26111 30345
rect 27982 30336 27988 30388
rect 28040 30376 28046 30388
rect 28810 30376 28816 30388
rect 28040 30348 28816 30376
rect 28040 30336 28046 30348
rect 28810 30336 28816 30348
rect 28868 30376 28874 30388
rect 29822 30376 29828 30388
rect 28868 30348 29828 30376
rect 28868 30336 28874 30348
rect 29822 30336 29828 30348
rect 29880 30336 29886 30388
rect 35894 30336 35900 30388
rect 35952 30336 35958 30388
rect 23293 30311 23351 30317
rect 23293 30308 23305 30311
rect 19536 30280 23305 30308
rect 23293 30277 23305 30280
rect 23339 30277 23351 30311
rect 23661 30311 23719 30317
rect 23293 30271 23351 30277
rect 23401 30280 23612 30308
rect 19153 30243 19211 30249
rect 19153 30209 19165 30243
rect 19199 30209 19211 30243
rect 19153 30203 19211 30209
rect 19334 30200 19340 30252
rect 19392 30200 19398 30252
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30209 19671 30243
rect 19613 30203 19671 30209
rect 18322 30132 18328 30184
rect 18380 30132 18386 30184
rect 18509 30175 18567 30181
rect 18509 30141 18521 30175
rect 18555 30141 18567 30175
rect 18509 30135 18567 30141
rect 18524 30104 18552 30135
rect 18782 30132 18788 30184
rect 18840 30172 18846 30184
rect 19628 30172 19656 30203
rect 19978 30200 19984 30252
rect 20036 30200 20042 30252
rect 20162 30200 20168 30252
rect 20220 30240 20226 30252
rect 21269 30243 21327 30249
rect 21269 30240 21281 30243
rect 20220 30212 21281 30240
rect 20220 30200 20226 30212
rect 21269 30209 21281 30212
rect 21315 30209 21327 30243
rect 21269 30203 21327 30209
rect 21361 30243 21419 30249
rect 21361 30209 21373 30243
rect 21407 30240 21419 30243
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 21407 30212 22017 30240
rect 21407 30209 21419 30212
rect 21361 30203 21419 30209
rect 22005 30209 22017 30212
rect 22051 30240 22063 30243
rect 23017 30243 23075 30249
rect 22051 30212 22692 30240
rect 22051 30209 22063 30212
rect 22005 30203 22063 30209
rect 22664 30184 22692 30212
rect 23017 30209 23029 30243
rect 23063 30209 23075 30243
rect 23017 30203 23075 30209
rect 23201 30243 23259 30249
rect 23201 30209 23213 30243
rect 23247 30240 23259 30243
rect 23401 30240 23429 30280
rect 23584 30252 23612 30280
rect 23661 30277 23673 30311
rect 23707 30308 23719 30311
rect 23707 30280 26188 30308
rect 23707 30277 23719 30280
rect 23661 30271 23719 30277
rect 23247 30212 23429 30240
rect 23247 30209 23259 30212
rect 23201 30203 23259 30209
rect 18840 30144 19656 30172
rect 18840 30132 18846 30144
rect 22278 30132 22284 30184
rect 22336 30132 22342 30184
rect 22646 30132 22652 30184
rect 22704 30132 22710 30184
rect 23032 30172 23060 30203
rect 23474 30200 23480 30252
rect 23532 30200 23538 30252
rect 23566 30200 23572 30252
rect 23624 30200 23630 30252
rect 23676 30172 23704 30271
rect 23753 30243 23811 30249
rect 23753 30209 23765 30243
rect 23799 30240 23811 30243
rect 24394 30240 24400 30252
rect 23799 30212 24400 30240
rect 23799 30209 23811 30212
rect 23753 30203 23811 30209
rect 24394 30200 24400 30212
rect 24452 30200 24458 30252
rect 24688 30184 24716 30280
rect 25038 30200 25044 30252
rect 25096 30240 25102 30252
rect 25608 30249 25636 30280
rect 25133 30243 25191 30249
rect 25133 30240 25145 30243
rect 25096 30212 25145 30240
rect 25096 30200 25102 30212
rect 25133 30209 25145 30212
rect 25179 30209 25191 30243
rect 25133 30203 25191 30209
rect 25317 30243 25375 30249
rect 25317 30209 25329 30243
rect 25363 30240 25375 30243
rect 25593 30243 25651 30249
rect 25363 30212 25544 30240
rect 25363 30209 25375 30212
rect 25317 30203 25375 30209
rect 25516 30184 25544 30212
rect 25593 30209 25605 30243
rect 25639 30209 25651 30243
rect 25593 30203 25651 30209
rect 25869 30243 25927 30249
rect 25869 30209 25881 30243
rect 25915 30240 25927 30243
rect 25958 30240 25964 30252
rect 25915 30212 25964 30240
rect 25915 30209 25927 30212
rect 25869 30203 25927 30209
rect 25958 30200 25964 30212
rect 26016 30240 26022 30252
rect 26160 30249 26188 30280
rect 28166 30268 28172 30320
rect 28224 30308 28230 30320
rect 28626 30308 28632 30320
rect 28224 30280 28632 30308
rect 28224 30268 28230 30280
rect 28626 30268 28632 30280
rect 28684 30268 28690 30320
rect 32398 30268 32404 30320
rect 32456 30268 32462 30320
rect 33796 30280 35388 30308
rect 33796 30252 33824 30280
rect 26053 30243 26111 30249
rect 26053 30240 26065 30243
rect 26016 30212 26065 30240
rect 26016 30200 26022 30212
rect 26053 30209 26065 30212
rect 26099 30209 26111 30243
rect 26053 30203 26111 30209
rect 26145 30243 26203 30249
rect 26145 30209 26157 30243
rect 26191 30209 26203 30243
rect 26145 30203 26203 30209
rect 23032 30144 23704 30172
rect 24670 30132 24676 30184
rect 24728 30132 24734 30184
rect 25498 30132 25504 30184
rect 25556 30132 25562 30184
rect 25685 30175 25743 30181
rect 25685 30141 25697 30175
rect 25731 30141 25743 30175
rect 25685 30135 25743 30141
rect 14936 30076 15976 30104
rect 18524 30076 18920 30104
rect 15948 30048 15976 30076
rect 9033 30039 9091 30045
rect 9033 30005 9045 30039
rect 9079 30036 9091 30039
rect 9214 30036 9220 30048
rect 9079 30008 9220 30036
rect 9079 30005 9091 30008
rect 9033 29999 9091 30005
rect 9214 29996 9220 30008
rect 9272 29996 9278 30048
rect 9766 29996 9772 30048
rect 9824 30036 9830 30048
rect 10134 30036 10140 30048
rect 9824 30008 10140 30036
rect 9824 29996 9830 30008
rect 10134 29996 10140 30008
rect 10192 29996 10198 30048
rect 11054 29996 11060 30048
rect 11112 30036 11118 30048
rect 11882 30036 11888 30048
rect 11112 30008 11888 30036
rect 11112 29996 11118 30008
rect 11882 29996 11888 30008
rect 11940 29996 11946 30048
rect 14461 30039 14519 30045
rect 14461 30005 14473 30039
rect 14507 30036 14519 30039
rect 14826 30036 14832 30048
rect 14507 30008 14832 30036
rect 14507 30005 14519 30008
rect 14461 29999 14519 30005
rect 14826 29996 14832 30008
rect 14884 29996 14890 30048
rect 14918 29996 14924 30048
rect 14976 30036 14982 30048
rect 15289 30039 15347 30045
rect 15289 30036 15301 30039
rect 14976 30008 15301 30036
rect 14976 29996 14982 30008
rect 15289 30005 15301 30008
rect 15335 30005 15347 30039
rect 15289 29999 15347 30005
rect 15378 29996 15384 30048
rect 15436 30036 15442 30048
rect 15473 30039 15531 30045
rect 15473 30036 15485 30039
rect 15436 30008 15485 30036
rect 15436 29996 15442 30008
rect 15473 30005 15485 30008
rect 15519 30005 15531 30039
rect 15473 29999 15531 30005
rect 15930 29996 15936 30048
rect 15988 30036 15994 30048
rect 16025 30039 16083 30045
rect 16025 30036 16037 30039
rect 15988 30008 16037 30036
rect 15988 29996 15994 30008
rect 16025 30005 16037 30008
rect 16071 30005 16083 30039
rect 16025 29999 16083 30005
rect 16206 29996 16212 30048
rect 16264 29996 16270 30048
rect 16850 29996 16856 30048
rect 16908 29996 16914 30048
rect 17034 29996 17040 30048
rect 17092 29996 17098 30048
rect 18230 29996 18236 30048
rect 18288 30036 18294 30048
rect 18325 30039 18383 30045
rect 18325 30036 18337 30039
rect 18288 30008 18337 30036
rect 18288 29996 18294 30008
rect 18325 30005 18337 30008
rect 18371 30005 18383 30039
rect 18325 29999 18383 30005
rect 18414 29996 18420 30048
rect 18472 30036 18478 30048
rect 18785 30039 18843 30045
rect 18785 30036 18797 30039
rect 18472 30008 18797 30036
rect 18472 29996 18478 30008
rect 18785 30005 18797 30008
rect 18831 30005 18843 30039
rect 18892 30036 18920 30076
rect 19150 30064 19156 30116
rect 19208 30104 19214 30116
rect 19794 30104 19800 30116
rect 19208 30076 19800 30104
rect 19208 30064 19214 30076
rect 19794 30064 19800 30076
rect 19852 30064 19858 30116
rect 20254 30064 20260 30116
rect 20312 30064 20318 30116
rect 20714 30064 20720 30116
rect 20772 30104 20778 30116
rect 25700 30104 25728 30135
rect 20772 30076 25728 30104
rect 26068 30104 26096 30203
rect 26602 30200 26608 30252
rect 26660 30240 26666 30252
rect 27798 30240 27804 30252
rect 26660 30212 27804 30240
rect 26660 30200 26666 30212
rect 27798 30200 27804 30212
rect 27856 30200 27862 30252
rect 29641 30243 29699 30249
rect 29641 30209 29653 30243
rect 29687 30240 29699 30243
rect 30282 30240 30288 30252
rect 29687 30212 30288 30240
rect 29687 30209 29699 30212
rect 29641 30203 29699 30209
rect 30282 30200 30288 30212
rect 30340 30200 30346 30252
rect 30742 30200 30748 30252
rect 30800 30200 30806 30252
rect 31205 30243 31263 30249
rect 31205 30209 31217 30243
rect 31251 30209 31263 30243
rect 31205 30203 31263 30209
rect 27154 30132 27160 30184
rect 27212 30172 27218 30184
rect 29914 30172 29920 30184
rect 27212 30144 29920 30172
rect 27212 30132 27218 30144
rect 29914 30132 29920 30144
rect 29972 30132 29978 30184
rect 30098 30132 30104 30184
rect 30156 30172 30162 30184
rect 30377 30175 30435 30181
rect 30377 30172 30389 30175
rect 30156 30144 30389 30172
rect 30156 30132 30162 30144
rect 30377 30141 30389 30144
rect 30423 30141 30435 30175
rect 30377 30135 30435 30141
rect 26510 30104 26516 30116
rect 26068 30076 26516 30104
rect 20772 30064 20778 30076
rect 26510 30064 26516 30076
rect 26568 30064 26574 30116
rect 30760 30104 30788 30200
rect 31220 30172 31248 30203
rect 31570 30200 31576 30252
rect 31628 30200 31634 30252
rect 32674 30200 32680 30252
rect 32732 30200 32738 30252
rect 32861 30243 32919 30249
rect 32861 30209 32873 30243
rect 32907 30240 32919 30243
rect 32950 30240 32956 30252
rect 32907 30212 32956 30240
rect 32907 30209 32919 30212
rect 32861 30203 32919 30209
rect 32950 30200 32956 30212
rect 33008 30200 33014 30252
rect 33137 30243 33195 30249
rect 33137 30209 33149 30243
rect 33183 30240 33195 30243
rect 33226 30240 33232 30252
rect 33183 30212 33232 30240
rect 33183 30209 33195 30212
rect 33137 30203 33195 30209
rect 33226 30200 33232 30212
rect 33284 30200 33290 30252
rect 33413 30243 33471 30249
rect 33413 30209 33425 30243
rect 33459 30240 33471 30243
rect 33502 30240 33508 30252
rect 33459 30212 33508 30240
rect 33459 30209 33471 30212
rect 33413 30203 33471 30209
rect 33502 30200 33508 30212
rect 33560 30200 33566 30252
rect 33594 30200 33600 30252
rect 33652 30200 33658 30252
rect 33778 30200 33784 30252
rect 33836 30200 33842 30252
rect 33965 30243 34023 30249
rect 33965 30209 33977 30243
rect 34011 30209 34023 30243
rect 33965 30203 34023 30209
rect 31294 30172 31300 30184
rect 31220 30144 31300 30172
rect 31294 30132 31300 30144
rect 31352 30172 31358 30184
rect 32125 30175 32183 30181
rect 32125 30172 32137 30175
rect 31352 30144 32137 30172
rect 31352 30132 31358 30144
rect 32125 30141 32137 30144
rect 32171 30172 32183 30175
rect 32214 30172 32220 30184
rect 32171 30144 32220 30172
rect 32171 30141 32183 30144
rect 32125 30135 32183 30141
rect 32214 30132 32220 30144
rect 32272 30132 32278 30184
rect 33612 30172 33640 30200
rect 33980 30172 34008 30203
rect 34146 30200 34152 30252
rect 34204 30240 34210 30252
rect 34425 30243 34483 30249
rect 34425 30240 34437 30243
rect 34204 30212 34437 30240
rect 34204 30200 34210 30212
rect 34425 30209 34437 30212
rect 34471 30209 34483 30243
rect 34425 30203 34483 30209
rect 34514 30200 34520 30252
rect 34572 30240 34578 30252
rect 35360 30249 35388 30280
rect 34793 30243 34851 30249
rect 34793 30240 34805 30243
rect 34572 30212 34805 30240
rect 34572 30200 34578 30212
rect 34793 30209 34805 30212
rect 34839 30209 34851 30243
rect 34793 30203 34851 30209
rect 35345 30243 35403 30249
rect 35345 30209 35357 30243
rect 35391 30209 35403 30243
rect 35345 30203 35403 30209
rect 35713 30243 35771 30249
rect 35713 30209 35725 30243
rect 35759 30209 35771 30243
rect 35713 30203 35771 30209
rect 35250 30172 35256 30184
rect 33612 30144 35256 30172
rect 35250 30132 35256 30144
rect 35308 30132 35314 30184
rect 29932 30076 30788 30104
rect 32324 30076 33732 30104
rect 20732 30036 20760 30064
rect 18892 30008 20760 30036
rect 18785 29999 18843 30005
rect 20806 29996 20812 30048
rect 20864 30036 20870 30048
rect 23017 30039 23075 30045
rect 23017 30036 23029 30039
rect 20864 30008 23029 30036
rect 20864 29996 20870 30008
rect 23017 30005 23029 30008
rect 23063 30005 23075 30039
rect 23017 29999 23075 30005
rect 23474 29996 23480 30048
rect 23532 30036 23538 30048
rect 23750 30036 23756 30048
rect 23532 30008 23756 30036
rect 23532 29996 23538 30008
rect 23750 29996 23756 30008
rect 23808 29996 23814 30048
rect 24026 29996 24032 30048
rect 24084 30036 24090 30048
rect 26602 30036 26608 30048
rect 24084 30008 26608 30036
rect 24084 29996 24090 30008
rect 26602 29996 26608 30008
rect 26660 29996 26666 30048
rect 29932 30045 29960 30076
rect 29917 30039 29975 30045
rect 29917 30005 29929 30039
rect 29963 30005 29975 30039
rect 29917 29999 29975 30005
rect 30098 29996 30104 30048
rect 30156 29996 30162 30048
rect 30190 29996 30196 30048
rect 30248 30036 30254 30048
rect 32324 30036 32352 30076
rect 33704 30045 33732 30076
rect 34606 30064 34612 30116
rect 34664 30104 34670 30116
rect 35728 30104 35756 30203
rect 34664 30076 35756 30104
rect 34664 30064 34670 30076
rect 30248 30008 32352 30036
rect 33689 30039 33747 30045
rect 30248 29996 30254 30008
rect 33689 30005 33701 30039
rect 33735 30005 33747 30039
rect 33689 29999 33747 30005
rect 34790 29996 34796 30048
rect 34848 30036 34854 30048
rect 35526 30036 35532 30048
rect 34848 30008 35532 30036
rect 34848 29996 34854 30008
rect 35526 29996 35532 30008
rect 35584 30036 35590 30048
rect 35621 30039 35679 30045
rect 35621 30036 35633 30039
rect 35584 30008 35633 30036
rect 35584 29996 35590 30008
rect 35621 30005 35633 30008
rect 35667 30005 35679 30039
rect 35621 29999 35679 30005
rect 1104 29946 41400 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 41400 29946
rect 1104 29872 41400 29894
rect 7650 29792 7656 29844
rect 7708 29792 7714 29844
rect 8573 29835 8631 29841
rect 8573 29801 8585 29835
rect 8619 29832 8631 29835
rect 11054 29832 11060 29844
rect 8619 29804 11060 29832
rect 8619 29801 8631 29804
rect 8573 29795 8631 29801
rect 11054 29792 11060 29804
rect 11112 29792 11118 29844
rect 11330 29792 11336 29844
rect 11388 29832 11394 29844
rect 11425 29835 11483 29841
rect 11425 29832 11437 29835
rect 11388 29804 11437 29832
rect 11388 29792 11394 29804
rect 11425 29801 11437 29804
rect 11471 29801 11483 29835
rect 11425 29795 11483 29801
rect 12250 29792 12256 29844
rect 12308 29792 12314 29844
rect 14366 29792 14372 29844
rect 14424 29792 14430 29844
rect 14461 29835 14519 29841
rect 14461 29801 14473 29835
rect 14507 29832 14519 29835
rect 14734 29832 14740 29844
rect 14507 29804 14740 29832
rect 14507 29801 14519 29804
rect 14461 29795 14519 29801
rect 14734 29792 14740 29804
rect 14792 29792 14798 29844
rect 16022 29792 16028 29844
rect 16080 29792 16086 29844
rect 16390 29792 16396 29844
rect 16448 29832 16454 29844
rect 18046 29832 18052 29844
rect 16448 29804 18052 29832
rect 16448 29792 16454 29804
rect 18046 29792 18052 29804
rect 18104 29792 18110 29844
rect 19334 29792 19340 29844
rect 19392 29792 19398 29844
rect 20346 29792 20352 29844
rect 20404 29832 20410 29844
rect 22649 29835 22707 29841
rect 20404 29804 21680 29832
rect 20404 29792 20410 29804
rect 9125 29767 9183 29773
rect 9125 29764 9137 29767
rect 8956 29736 9137 29764
rect 8956 29708 8984 29736
rect 9125 29733 9137 29736
rect 9171 29733 9183 29767
rect 9125 29727 9183 29733
rect 9490 29724 9496 29776
rect 9548 29764 9554 29776
rect 9674 29764 9680 29776
rect 9548 29736 9680 29764
rect 9548 29724 9554 29736
rect 9674 29724 9680 29736
rect 9732 29724 9738 29776
rect 9950 29764 9956 29776
rect 9784 29736 9956 29764
rect 5460 29668 6224 29696
rect 5460 29637 5488 29668
rect 6196 29640 6224 29668
rect 8018 29656 8024 29708
rect 8076 29656 8082 29708
rect 8665 29699 8723 29705
rect 8665 29665 8677 29699
rect 8711 29665 8723 29699
rect 8665 29659 8723 29665
rect 5445 29631 5503 29637
rect 5445 29597 5457 29631
rect 5491 29597 5503 29631
rect 5445 29591 5503 29597
rect 5718 29588 5724 29640
rect 5776 29588 5782 29640
rect 5813 29631 5871 29637
rect 5813 29597 5825 29631
rect 5859 29628 5871 29631
rect 6086 29628 6092 29640
rect 5859 29600 6092 29628
rect 5859 29597 5871 29600
rect 5813 29591 5871 29597
rect 6086 29588 6092 29600
rect 6144 29588 6150 29640
rect 6178 29588 6184 29640
rect 6236 29588 6242 29640
rect 6454 29588 6460 29640
rect 6512 29588 6518 29640
rect 7837 29631 7895 29637
rect 7837 29597 7849 29631
rect 7883 29597 7895 29631
rect 7837 29591 7895 29597
rect 5258 29520 5264 29572
rect 5316 29560 5322 29572
rect 5629 29563 5687 29569
rect 5629 29560 5641 29563
rect 5316 29532 5641 29560
rect 5316 29520 5322 29532
rect 5629 29529 5641 29532
rect 5675 29560 5687 29563
rect 6472 29560 6500 29588
rect 5675 29532 6500 29560
rect 7852 29560 7880 29591
rect 7926 29588 7932 29640
rect 7984 29588 7990 29640
rect 8113 29631 8171 29637
rect 8113 29597 8125 29631
rect 8159 29628 8171 29631
rect 8202 29628 8208 29640
rect 8159 29600 8208 29628
rect 8159 29597 8171 29600
rect 8113 29591 8171 29597
rect 8202 29588 8208 29600
rect 8260 29588 8266 29640
rect 8386 29588 8392 29640
rect 8444 29588 8450 29640
rect 8478 29588 8484 29640
rect 8536 29588 8542 29640
rect 8680 29628 8708 29659
rect 8938 29656 8944 29708
rect 8996 29656 9002 29708
rect 9582 29696 9588 29708
rect 9324 29668 9588 29696
rect 9324 29640 9352 29668
rect 9582 29656 9588 29668
rect 9640 29656 9646 29708
rect 9784 29696 9812 29736
rect 9950 29724 9956 29736
rect 10008 29724 10014 29776
rect 10321 29767 10379 29773
rect 10321 29733 10333 29767
rect 10367 29733 10379 29767
rect 10321 29727 10379 29733
rect 9692 29668 9812 29696
rect 10336 29696 10364 29727
rect 10336 29668 10824 29696
rect 9692 29640 9720 29668
rect 9306 29628 9312 29640
rect 8680 29600 9312 29628
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 9401 29631 9459 29637
rect 9401 29597 9413 29631
rect 9447 29628 9459 29631
rect 9447 29600 9628 29628
rect 9447 29597 9459 29600
rect 9401 29591 9459 29597
rect 8404 29560 8432 29588
rect 9600 29572 9628 29600
rect 9674 29588 9680 29640
rect 9732 29588 9738 29640
rect 9766 29588 9772 29640
rect 9824 29628 9830 29640
rect 9953 29631 10011 29637
rect 9824 29600 9869 29628
rect 9824 29588 9830 29600
rect 9953 29597 9965 29631
rect 9999 29597 10011 29631
rect 9953 29591 10011 29597
rect 7852 29532 8432 29560
rect 5675 29529 5687 29532
rect 5629 29523 5687 29529
rect 8662 29520 8668 29572
rect 8720 29560 8726 29572
rect 8846 29560 8852 29572
rect 8720 29532 8852 29560
rect 8720 29520 8726 29532
rect 8846 29520 8852 29532
rect 8904 29560 8910 29572
rect 9125 29563 9183 29569
rect 9125 29560 9137 29563
rect 8904 29532 9137 29560
rect 8904 29520 8910 29532
rect 9125 29529 9137 29532
rect 9171 29529 9183 29563
rect 9125 29523 9183 29529
rect 9582 29520 9588 29572
rect 9640 29520 9646 29572
rect 9968 29560 9996 29591
rect 10042 29588 10048 29640
rect 10100 29588 10106 29640
rect 10134 29588 10140 29640
rect 10192 29637 10198 29640
rect 10192 29631 10241 29637
rect 10192 29597 10195 29631
rect 10229 29628 10241 29631
rect 10318 29628 10324 29640
rect 10229 29600 10324 29628
rect 10229 29597 10241 29600
rect 10192 29591 10241 29597
rect 10192 29588 10198 29591
rect 10318 29588 10324 29600
rect 10376 29588 10382 29640
rect 10502 29588 10508 29640
rect 10560 29588 10566 29640
rect 10796 29637 10824 29668
rect 11514 29656 11520 29708
rect 11572 29656 11578 29708
rect 12268 29696 12296 29792
rect 14553 29767 14611 29773
rect 14553 29733 14565 29767
rect 14599 29764 14611 29767
rect 15286 29764 15292 29776
rect 14599 29736 15292 29764
rect 14599 29733 14611 29736
rect 14553 29727 14611 29733
rect 15286 29724 15292 29736
rect 15344 29764 15350 29776
rect 16040 29764 16068 29792
rect 15344 29736 16068 29764
rect 15344 29724 15350 29736
rect 16114 29724 16120 29776
rect 16172 29764 16178 29776
rect 16209 29767 16267 29773
rect 16209 29764 16221 29767
rect 16172 29736 16221 29764
rect 16172 29724 16178 29736
rect 16209 29733 16221 29736
rect 16255 29733 16267 29767
rect 16209 29727 16267 29733
rect 17862 29724 17868 29776
rect 17920 29724 17926 29776
rect 18230 29724 18236 29776
rect 18288 29764 18294 29776
rect 19150 29764 19156 29776
rect 18288 29736 19156 29764
rect 18288 29724 18294 29736
rect 19150 29724 19156 29736
rect 19208 29724 19214 29776
rect 19426 29724 19432 29776
rect 19484 29764 19490 29776
rect 21542 29764 21548 29776
rect 19484 29736 21548 29764
rect 19484 29724 19490 29736
rect 21542 29724 21548 29736
rect 21600 29724 21606 29776
rect 21652 29764 21680 29804
rect 22649 29801 22661 29835
rect 22695 29832 22707 29835
rect 22738 29832 22744 29844
rect 22695 29804 22744 29832
rect 22695 29801 22707 29804
rect 22649 29795 22707 29801
rect 22738 29792 22744 29804
rect 22796 29832 22802 29844
rect 23934 29832 23940 29844
rect 22796 29804 23940 29832
rect 22796 29792 22802 29804
rect 23934 29792 23940 29804
rect 23992 29832 23998 29844
rect 23992 29804 26280 29832
rect 23992 29792 23998 29804
rect 26252 29776 26280 29804
rect 27522 29792 27528 29844
rect 27580 29832 27586 29844
rect 30190 29832 30196 29844
rect 27580 29804 30196 29832
rect 27580 29792 27586 29804
rect 30190 29792 30196 29804
rect 30248 29792 30254 29844
rect 35253 29835 35311 29841
rect 35253 29801 35265 29835
rect 35299 29832 35311 29835
rect 35342 29832 35348 29844
rect 35299 29804 35348 29832
rect 35299 29801 35311 29804
rect 35253 29795 35311 29801
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 35434 29792 35440 29844
rect 35492 29792 35498 29844
rect 37550 29792 37556 29844
rect 37608 29792 37614 29844
rect 21652 29736 22140 29764
rect 22112 29708 22140 29736
rect 22278 29724 22284 29776
rect 22336 29764 22342 29776
rect 23017 29767 23075 29773
rect 23017 29764 23029 29767
rect 22336 29736 23029 29764
rect 22336 29724 22342 29736
rect 23017 29733 23029 29736
rect 23063 29733 23075 29767
rect 23017 29727 23075 29733
rect 23566 29724 23572 29776
rect 23624 29764 23630 29776
rect 24578 29764 24584 29776
rect 23624 29736 24584 29764
rect 23624 29724 23630 29736
rect 24578 29724 24584 29736
rect 24636 29724 24642 29776
rect 26234 29724 26240 29776
rect 26292 29724 26298 29776
rect 29822 29764 29828 29776
rect 27586 29736 29828 29764
rect 27586 29708 27614 29736
rect 29822 29724 29828 29736
rect 29880 29724 29886 29776
rect 30558 29724 30564 29776
rect 30616 29724 30622 29776
rect 14918 29696 14924 29708
rect 12268 29668 12848 29696
rect 10781 29631 10839 29637
rect 10781 29597 10793 29631
rect 10827 29597 10839 29631
rect 10781 29591 10839 29597
rect 11333 29631 11391 29637
rect 11333 29597 11345 29631
rect 11379 29628 11391 29631
rect 11532 29628 11560 29656
rect 11379 29600 11560 29628
rect 11379 29597 11391 29600
rect 11333 29591 11391 29597
rect 12434 29588 12440 29640
rect 12492 29628 12498 29640
rect 12820 29637 12848 29668
rect 13740 29668 14924 29696
rect 13740 29640 13768 29668
rect 14918 29656 14924 29668
rect 14976 29656 14982 29708
rect 18690 29696 18696 29708
rect 16132 29668 17632 29696
rect 12713 29631 12771 29637
rect 12713 29628 12725 29631
rect 12492 29600 12725 29628
rect 12492 29588 12498 29600
rect 12713 29597 12725 29600
rect 12759 29597 12771 29631
rect 12713 29591 12771 29597
rect 12805 29631 12863 29637
rect 12805 29597 12817 29631
rect 12851 29597 12863 29631
rect 12805 29591 12863 29597
rect 12894 29588 12900 29640
rect 12952 29588 12958 29640
rect 13081 29631 13139 29637
rect 13081 29597 13093 29631
rect 13127 29628 13139 29631
rect 13170 29628 13176 29640
rect 13127 29600 13176 29628
rect 13127 29597 13139 29600
rect 13081 29591 13139 29597
rect 13170 29588 13176 29600
rect 13228 29588 13234 29640
rect 13722 29588 13728 29640
rect 13780 29588 13786 29640
rect 14366 29588 14372 29640
rect 14424 29628 14430 29640
rect 14829 29631 14887 29637
rect 14829 29628 14841 29631
rect 14424 29600 14841 29628
rect 14424 29588 14430 29600
rect 14829 29597 14841 29600
rect 14875 29597 14887 29631
rect 15105 29631 15163 29637
rect 15105 29628 15117 29631
rect 14829 29591 14887 29597
rect 14936 29600 15117 29628
rect 14936 29572 14964 29600
rect 15105 29597 15117 29600
rect 15151 29597 15163 29631
rect 15105 29591 15163 29597
rect 15378 29588 15384 29640
rect 15436 29588 15442 29640
rect 16132 29637 16160 29668
rect 17604 29640 17632 29668
rect 17972 29668 18696 29696
rect 16025 29631 16083 29637
rect 16025 29628 16037 29631
rect 15580 29600 16037 29628
rect 10689 29563 10747 29569
rect 9968 29532 10088 29560
rect 5994 29452 6000 29504
rect 6052 29452 6058 29504
rect 8294 29452 8300 29504
rect 8352 29492 8358 29504
rect 9030 29492 9036 29504
rect 8352 29464 9036 29492
rect 8352 29452 8358 29464
rect 9030 29452 9036 29464
rect 9088 29452 9094 29504
rect 9398 29452 9404 29504
rect 9456 29492 9462 29504
rect 9950 29492 9956 29504
rect 9456 29464 9956 29492
rect 9456 29452 9462 29464
rect 9950 29452 9956 29464
rect 10008 29492 10014 29504
rect 10060 29492 10088 29532
rect 10689 29529 10701 29563
rect 10735 29529 10747 29563
rect 10689 29523 10747 29529
rect 10008 29464 10088 29492
rect 10704 29492 10732 29523
rect 11054 29520 11060 29572
rect 11112 29560 11118 29572
rect 11241 29563 11299 29569
rect 11241 29560 11253 29563
rect 11112 29532 11253 29560
rect 11112 29520 11118 29532
rect 11241 29529 11253 29532
rect 11287 29529 11299 29563
rect 14093 29563 14151 29569
rect 14093 29560 14105 29563
rect 11241 29523 11299 29529
rect 11348 29532 14105 29560
rect 11348 29492 11376 29532
rect 14093 29529 14105 29532
rect 14139 29529 14151 29563
rect 14093 29523 14151 29529
rect 14918 29520 14924 29572
rect 14976 29520 14982 29572
rect 15289 29563 15347 29569
rect 15289 29529 15301 29563
rect 15335 29529 15347 29563
rect 15289 29523 15347 29529
rect 10704 29464 11376 29492
rect 10008 29452 10014 29464
rect 12434 29452 12440 29504
rect 12492 29452 12498 29504
rect 13906 29452 13912 29504
rect 13964 29492 13970 29504
rect 14737 29495 14795 29501
rect 14737 29492 14749 29495
rect 13964 29464 14749 29492
rect 13964 29452 13970 29464
rect 14737 29461 14749 29464
rect 14783 29492 14795 29495
rect 15304 29492 15332 29523
rect 15580 29504 15608 29600
rect 16025 29597 16037 29600
rect 16071 29597 16083 29631
rect 16025 29591 16083 29597
rect 16117 29631 16175 29637
rect 16117 29597 16129 29631
rect 16163 29597 16175 29631
rect 16117 29591 16175 29597
rect 16298 29588 16304 29640
rect 16356 29588 16362 29640
rect 16390 29588 16396 29640
rect 16448 29628 16454 29640
rect 16485 29631 16543 29637
rect 16485 29628 16497 29631
rect 16448 29600 16497 29628
rect 16448 29588 16454 29600
rect 16485 29597 16497 29600
rect 16531 29597 16543 29631
rect 16485 29591 16543 29597
rect 16574 29588 16580 29640
rect 16632 29588 16638 29640
rect 17034 29588 17040 29640
rect 17092 29588 17098 29640
rect 17126 29588 17132 29640
rect 17184 29628 17190 29640
rect 17497 29631 17555 29637
rect 17497 29628 17509 29631
rect 17184 29600 17509 29628
rect 17184 29588 17190 29600
rect 17497 29597 17509 29600
rect 17543 29597 17555 29631
rect 17497 29591 17555 29597
rect 17586 29588 17592 29640
rect 17644 29588 17650 29640
rect 17865 29631 17923 29637
rect 17865 29597 17877 29631
rect 17911 29597 17923 29631
rect 17865 29591 17923 29597
rect 17880 29560 17908 29591
rect 16040 29532 17908 29560
rect 16040 29504 16068 29532
rect 14783 29464 15332 29492
rect 14783 29461 14795 29464
rect 14737 29455 14795 29461
rect 15562 29452 15568 29504
rect 15620 29452 15626 29504
rect 15838 29452 15844 29504
rect 15896 29452 15902 29504
rect 16022 29452 16028 29504
rect 16080 29452 16086 29504
rect 16114 29452 16120 29504
rect 16172 29492 16178 29504
rect 17310 29492 17316 29504
rect 16172 29464 17316 29492
rect 16172 29452 16178 29464
rect 17310 29452 17316 29464
rect 17368 29492 17374 29504
rect 17972 29492 18000 29668
rect 18690 29656 18696 29668
rect 18748 29656 18754 29708
rect 18892 29668 20392 29696
rect 18230 29588 18236 29640
rect 18288 29588 18294 29640
rect 18892 29637 18920 29668
rect 18877 29631 18935 29637
rect 18877 29597 18889 29631
rect 18923 29597 18935 29631
rect 18877 29591 18935 29597
rect 18966 29588 18972 29640
rect 19024 29628 19030 29640
rect 19245 29631 19303 29637
rect 19245 29628 19257 29631
rect 19024 29600 19257 29628
rect 19024 29588 19030 29600
rect 19245 29597 19257 29600
rect 19291 29597 19303 29631
rect 19245 29591 19303 29597
rect 19334 29588 19340 29640
rect 19392 29628 19398 29640
rect 19521 29631 19579 29637
rect 19521 29628 19533 29631
rect 19392 29600 19533 29628
rect 19392 29588 19398 29600
rect 19521 29597 19533 29600
rect 19567 29597 19579 29631
rect 19521 29591 19579 29597
rect 19886 29588 19892 29640
rect 19944 29588 19950 29640
rect 20364 29637 20392 29668
rect 22094 29656 22100 29708
rect 22152 29656 22158 29708
rect 22462 29656 22468 29708
rect 22520 29656 22526 29708
rect 22830 29696 22836 29708
rect 22572 29668 22836 29696
rect 20073 29631 20131 29637
rect 20073 29597 20085 29631
rect 20119 29628 20131 29631
rect 20349 29631 20407 29637
rect 20119 29600 20300 29628
rect 20119 29597 20131 29600
rect 20073 29591 20131 29597
rect 20272 29560 20300 29600
rect 20349 29597 20361 29631
rect 20395 29628 20407 29631
rect 20714 29628 20720 29640
rect 20395 29600 20720 29628
rect 20395 29597 20407 29600
rect 20349 29591 20407 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 20806 29588 20812 29640
rect 20864 29588 20870 29640
rect 21542 29588 21548 29640
rect 21600 29588 21606 29640
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29597 21787 29631
rect 21729 29591 21787 29597
rect 20824 29560 20852 29588
rect 18156 29532 20236 29560
rect 20272 29532 20852 29560
rect 20993 29563 21051 29569
rect 18156 29504 18184 29532
rect 17368 29464 18000 29492
rect 17368 29452 17374 29464
rect 18138 29452 18144 29504
rect 18196 29452 18202 29504
rect 18230 29452 18236 29504
rect 18288 29492 18294 29504
rect 18690 29492 18696 29504
rect 18288 29464 18696 29492
rect 18288 29452 18294 29464
rect 18690 29452 18696 29464
rect 18748 29452 18754 29504
rect 19061 29495 19119 29501
rect 19061 29461 19073 29495
rect 19107 29492 19119 29495
rect 20070 29492 20076 29504
rect 19107 29464 20076 29492
rect 19107 29461 19119 29464
rect 19061 29455 19119 29461
rect 20070 29452 20076 29464
rect 20128 29452 20134 29504
rect 20208 29492 20236 29532
rect 20993 29529 21005 29563
rect 21039 29560 21051 29563
rect 21082 29560 21088 29572
rect 21039 29532 21088 29560
rect 21039 29529 21051 29532
rect 20993 29523 21051 29529
rect 21082 29520 21088 29532
rect 21140 29520 21146 29572
rect 21744 29560 21772 29591
rect 21910 29588 21916 29640
rect 21968 29628 21974 29640
rect 22005 29631 22063 29637
rect 22005 29628 22017 29631
rect 21968 29600 22017 29628
rect 21968 29588 21974 29600
rect 22005 29597 22017 29600
rect 22051 29628 22063 29631
rect 22572 29628 22600 29668
rect 22830 29656 22836 29668
rect 22888 29656 22894 29708
rect 24026 29696 24032 29708
rect 23400 29668 24032 29696
rect 22051 29600 22600 29628
rect 22051 29597 22063 29600
rect 22005 29591 22063 29597
rect 22646 29588 22652 29640
rect 22704 29588 22710 29640
rect 23017 29631 23075 29637
rect 22278 29560 22284 29572
rect 21744 29532 22284 29560
rect 22278 29520 22284 29532
rect 22336 29520 22342 29572
rect 22373 29563 22431 29569
rect 22373 29529 22385 29563
rect 22419 29560 22431 29563
rect 22830 29560 22836 29606
rect 22419 29554 22836 29560
rect 22888 29554 22894 29606
rect 23017 29597 23029 29631
rect 23063 29628 23075 29631
rect 23198 29628 23204 29640
rect 23063 29600 23204 29628
rect 23063 29597 23075 29600
rect 23017 29591 23075 29597
rect 23198 29588 23204 29600
rect 23256 29588 23262 29640
rect 23290 29588 23296 29640
rect 23348 29588 23354 29640
rect 23400 29560 23428 29668
rect 24026 29656 24032 29668
rect 24084 29656 24090 29708
rect 24302 29656 24308 29708
rect 24360 29696 24366 29708
rect 24946 29696 24952 29708
rect 24360 29668 24952 29696
rect 24360 29656 24366 29668
rect 24872 29637 24900 29668
rect 24946 29656 24952 29668
rect 25004 29656 25010 29708
rect 25590 29656 25596 29708
rect 25648 29696 25654 29708
rect 27433 29699 27491 29705
rect 27433 29696 27445 29699
rect 25648 29668 27445 29696
rect 25648 29656 25654 29668
rect 27433 29665 27445 29668
rect 27479 29665 27491 29699
rect 27433 29659 27491 29665
rect 27522 29656 27528 29708
rect 27580 29668 27614 29708
rect 27709 29699 27767 29705
rect 27580 29656 27586 29668
rect 27709 29665 27721 29699
rect 27755 29696 27767 29699
rect 28994 29696 29000 29708
rect 27755 29668 29000 29696
rect 27755 29665 27767 29668
rect 27709 29659 27767 29665
rect 28994 29656 29000 29668
rect 29052 29656 29058 29708
rect 32033 29699 32091 29705
rect 32033 29696 32045 29699
rect 29656 29668 32045 29696
rect 24857 29631 24915 29637
rect 24857 29597 24869 29631
rect 24903 29597 24915 29631
rect 24857 29591 24915 29597
rect 25035 29631 25093 29637
rect 25035 29597 25047 29631
rect 25081 29628 25176 29631
rect 25958 29628 25964 29640
rect 25081 29603 25964 29628
rect 25081 29597 25093 29603
rect 25148 29600 25964 29603
rect 25035 29591 25093 29597
rect 25958 29588 25964 29600
rect 26016 29628 26022 29640
rect 27614 29628 27620 29640
rect 26016 29600 27620 29628
rect 26016 29588 26022 29600
rect 27614 29588 27620 29600
rect 27672 29588 27678 29640
rect 27798 29588 27804 29640
rect 27856 29628 27862 29640
rect 28077 29631 28135 29637
rect 28077 29628 28089 29631
rect 27856 29600 28089 29628
rect 27856 29588 27862 29600
rect 28077 29597 28089 29600
rect 28123 29628 28135 29631
rect 29656 29628 29684 29668
rect 32033 29665 32045 29668
rect 32079 29665 32091 29699
rect 32033 29659 32091 29665
rect 32214 29656 32220 29708
rect 32272 29696 32278 29708
rect 32272 29668 32996 29696
rect 32272 29656 32278 29668
rect 30098 29628 30104 29640
rect 28123 29600 29684 29628
rect 29748 29600 30104 29628
rect 28123 29597 28135 29600
rect 28077 29591 28135 29597
rect 22419 29532 22876 29554
rect 23216 29532 23428 29560
rect 22419 29529 22431 29532
rect 22373 29523 22431 29529
rect 22462 29492 22468 29504
rect 20208 29464 22468 29492
rect 22462 29452 22468 29464
rect 22520 29452 22526 29504
rect 22830 29452 22836 29504
rect 22888 29452 22894 29504
rect 23216 29501 23244 29532
rect 23566 29520 23572 29572
rect 23624 29560 23630 29572
rect 29748 29560 29776 29600
rect 30098 29588 30104 29600
rect 30156 29588 30162 29640
rect 30282 29588 30288 29640
rect 30340 29588 30346 29640
rect 30374 29588 30380 29640
rect 30432 29628 30438 29640
rect 31294 29628 31300 29640
rect 30432 29600 31300 29628
rect 30432 29588 30438 29600
rect 31294 29588 31300 29600
rect 31352 29588 31358 29640
rect 31478 29588 31484 29640
rect 31536 29628 31542 29640
rect 31685 29634 31825 29638
rect 31685 29628 31840 29634
rect 31536 29610 31794 29628
rect 31536 29600 31713 29610
rect 31536 29588 31542 29600
rect 31782 29594 31794 29610
rect 31828 29594 31840 29628
rect 31782 29588 31840 29594
rect 32585 29631 32643 29637
rect 32585 29597 32597 29631
rect 32631 29628 32643 29631
rect 32674 29628 32680 29640
rect 32631 29600 32680 29628
rect 32631 29597 32643 29600
rect 32585 29591 32643 29597
rect 32674 29588 32680 29600
rect 32732 29588 32738 29640
rect 32968 29637 32996 29668
rect 34072 29668 35296 29696
rect 32953 29631 33011 29637
rect 32953 29597 32965 29631
rect 32999 29628 33011 29631
rect 32999 29600 33088 29628
rect 32999 29597 33011 29600
rect 32953 29591 33011 29597
rect 23624 29532 29776 29560
rect 29825 29563 29883 29569
rect 23624 29520 23630 29532
rect 23201 29495 23259 29501
rect 23201 29461 23213 29495
rect 23247 29461 23259 29495
rect 23201 29455 23259 29461
rect 24762 29452 24768 29504
rect 24820 29492 24826 29504
rect 24949 29495 25007 29501
rect 24949 29492 24961 29495
rect 24820 29464 24961 29492
rect 24820 29452 24826 29464
rect 24949 29461 24961 29464
rect 24995 29461 25007 29495
rect 24949 29455 25007 29461
rect 25038 29452 25044 29504
rect 25096 29492 25102 29504
rect 25590 29492 25596 29504
rect 25096 29464 25596 29492
rect 25096 29452 25102 29464
rect 25590 29452 25596 29464
rect 25648 29452 25654 29504
rect 26234 29452 26240 29504
rect 26292 29492 26298 29504
rect 27522 29492 27528 29504
rect 26292 29464 27528 29492
rect 26292 29452 26298 29464
rect 27522 29452 27528 29464
rect 27580 29452 27586 29504
rect 27816 29501 27844 29532
rect 29825 29529 29837 29563
rect 29871 29560 29883 29563
rect 30742 29560 30748 29572
rect 29871 29532 30748 29560
rect 29871 29529 29883 29532
rect 29825 29523 29883 29529
rect 30742 29520 30748 29532
rect 30800 29560 30806 29572
rect 30837 29563 30895 29569
rect 30837 29560 30849 29563
rect 30800 29532 30849 29560
rect 30800 29520 30806 29532
rect 30837 29529 30849 29532
rect 30883 29529 30895 29563
rect 30837 29523 30895 29529
rect 30926 29520 30932 29572
rect 30984 29520 30990 29572
rect 31389 29563 31447 29569
rect 31389 29529 31401 29563
rect 31435 29560 31447 29563
rect 31570 29560 31576 29572
rect 31435 29532 31576 29560
rect 31435 29529 31447 29532
rect 31389 29523 31447 29529
rect 31570 29520 31576 29532
rect 31628 29520 31634 29572
rect 31797 29560 31825 29588
rect 33060 29560 33088 29600
rect 33226 29588 33232 29640
rect 33284 29588 33290 29640
rect 33594 29588 33600 29640
rect 33652 29588 33658 29640
rect 33778 29588 33784 29640
rect 33836 29628 33842 29640
rect 34072 29637 34100 29668
rect 34057 29631 34115 29637
rect 34057 29628 34069 29631
rect 33836 29600 34069 29628
rect 33836 29588 33842 29600
rect 34057 29597 34069 29600
rect 34103 29597 34115 29631
rect 34057 29591 34115 29597
rect 34333 29631 34391 29637
rect 34333 29597 34345 29631
rect 34379 29628 34391 29631
rect 34514 29628 34520 29640
rect 34379 29600 34520 29628
rect 34379 29597 34391 29600
rect 34333 29591 34391 29597
rect 34348 29560 34376 29591
rect 34514 29588 34520 29600
rect 34572 29588 34578 29640
rect 34790 29588 34796 29640
rect 34848 29588 34854 29640
rect 35268 29637 35296 29668
rect 35802 29656 35808 29708
rect 35860 29696 35866 29708
rect 35860 29668 38148 29696
rect 35860 29656 35866 29668
rect 38120 29640 38148 29668
rect 34885 29631 34943 29637
rect 34885 29597 34897 29631
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 35253 29631 35311 29637
rect 35253 29597 35265 29631
rect 35299 29597 35311 29631
rect 35253 29591 35311 29597
rect 31797 29532 32996 29560
rect 33060 29532 34376 29560
rect 27801 29495 27859 29501
rect 27801 29461 27813 29495
rect 27847 29461 27859 29495
rect 27801 29455 27859 29461
rect 27982 29452 27988 29504
rect 28040 29492 28046 29504
rect 29546 29492 29552 29504
rect 28040 29464 29552 29492
rect 28040 29452 28046 29464
rect 29546 29452 29552 29464
rect 29604 29452 29610 29504
rect 30006 29452 30012 29504
rect 30064 29492 30070 29504
rect 30650 29492 30656 29504
rect 30064 29464 30656 29492
rect 30064 29452 30070 29464
rect 30650 29452 30656 29464
rect 30708 29452 30714 29504
rect 31588 29492 31616 29520
rect 32968 29504 32996 29532
rect 34606 29520 34612 29572
rect 34664 29560 34670 29572
rect 34900 29560 34928 29591
rect 35710 29588 35716 29640
rect 35768 29588 35774 29640
rect 38102 29588 38108 29640
rect 38160 29588 38166 29640
rect 36081 29563 36139 29569
rect 36081 29560 36093 29563
rect 34664 29532 34928 29560
rect 35544 29532 36093 29560
rect 34664 29520 34670 29532
rect 31754 29492 31760 29504
rect 31588 29464 31760 29492
rect 31754 29452 31760 29464
rect 31812 29452 31818 29504
rect 32950 29452 32956 29504
rect 33008 29492 33014 29504
rect 33873 29495 33931 29501
rect 33873 29492 33885 29495
rect 33008 29464 33885 29492
rect 33008 29452 33014 29464
rect 33873 29461 33885 29464
rect 33919 29492 33931 29495
rect 34146 29492 34152 29504
rect 33919 29464 34152 29492
rect 33919 29461 33931 29464
rect 33873 29455 33931 29461
rect 34146 29452 34152 29464
rect 34204 29452 34210 29504
rect 35544 29501 35572 29532
rect 36081 29529 36093 29532
rect 36127 29529 36139 29563
rect 37306 29532 37412 29560
rect 36081 29523 36139 29529
rect 35529 29495 35587 29501
rect 35529 29461 35541 29495
rect 35575 29461 35587 29495
rect 35529 29455 35587 29461
rect 36262 29452 36268 29504
rect 36320 29492 36326 29504
rect 37384 29492 37412 29532
rect 37642 29520 37648 29572
rect 37700 29560 37706 29572
rect 37737 29563 37795 29569
rect 37737 29560 37749 29563
rect 37700 29532 37749 29560
rect 37700 29520 37706 29532
rect 37737 29529 37749 29532
rect 37783 29560 37795 29563
rect 37918 29560 37924 29572
rect 37783 29532 37924 29560
rect 37783 29529 37795 29532
rect 37737 29523 37795 29529
rect 37918 29520 37924 29532
rect 37976 29520 37982 29572
rect 37829 29495 37887 29501
rect 37829 29492 37841 29495
rect 36320 29464 37841 29492
rect 36320 29452 36326 29464
rect 37829 29461 37841 29464
rect 37875 29461 37887 29495
rect 37829 29455 37887 29461
rect 1104 29402 41400 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 41400 29402
rect 1104 29328 41400 29350
rect 7558 29248 7564 29300
rect 7616 29248 7622 29300
rect 7834 29248 7840 29300
rect 7892 29248 7898 29300
rect 8205 29291 8263 29297
rect 8205 29257 8217 29291
rect 8251 29288 8263 29291
rect 8478 29288 8484 29300
rect 8251 29260 8484 29288
rect 8251 29257 8263 29260
rect 8205 29251 8263 29257
rect 8478 29248 8484 29260
rect 8536 29248 8542 29300
rect 8754 29248 8760 29300
rect 8812 29248 8818 29300
rect 9125 29291 9183 29297
rect 9125 29257 9137 29291
rect 9171 29288 9183 29291
rect 9398 29288 9404 29300
rect 9171 29260 9404 29288
rect 9171 29257 9183 29260
rect 9125 29251 9183 29257
rect 9398 29248 9404 29260
rect 9456 29248 9462 29300
rect 10321 29291 10379 29297
rect 10321 29257 10333 29291
rect 10367 29288 10379 29291
rect 10613 29291 10671 29297
rect 10613 29288 10625 29291
rect 10367 29260 10625 29288
rect 10367 29257 10379 29260
rect 10321 29251 10379 29257
rect 10613 29257 10625 29260
rect 10659 29257 10671 29291
rect 10613 29251 10671 29257
rect 11882 29248 11888 29300
rect 11940 29288 11946 29300
rect 12253 29291 12311 29297
rect 12253 29288 12265 29291
rect 11940 29260 12265 29288
rect 11940 29248 11946 29260
rect 12253 29257 12265 29260
rect 12299 29257 12311 29291
rect 12253 29251 12311 29257
rect 12894 29248 12900 29300
rect 12952 29248 12958 29300
rect 13538 29248 13544 29300
rect 13596 29288 13602 29300
rect 13596 29260 14780 29288
rect 13596 29248 13602 29260
rect 5718 29180 5724 29232
rect 5776 29220 5782 29232
rect 6089 29223 6147 29229
rect 6089 29220 6101 29223
rect 5776 29192 6101 29220
rect 5776 29180 5782 29192
rect 6089 29189 6101 29192
rect 6135 29189 6147 29223
rect 7852 29220 7880 29248
rect 7852 29192 8616 29220
rect 6089 29183 6147 29189
rect 5442 29112 5448 29164
rect 5500 29112 5506 29164
rect 7469 29155 7527 29161
rect 7469 29121 7481 29155
rect 7515 29121 7527 29155
rect 7469 29115 7527 29121
rect 3786 29044 3792 29096
rect 3844 29084 3850 29096
rect 4065 29087 4123 29093
rect 4065 29084 4077 29087
rect 3844 29056 4077 29084
rect 3844 29044 3850 29056
rect 4065 29053 4077 29056
rect 4111 29053 4123 29087
rect 4065 29047 4123 29053
rect 5994 28976 6000 29028
rect 6052 28976 6058 29028
rect 7484 29016 7512 29115
rect 7558 29112 7564 29164
rect 7616 29152 7622 29164
rect 7653 29155 7711 29161
rect 7653 29152 7665 29155
rect 7616 29124 7665 29152
rect 7616 29112 7622 29124
rect 7653 29121 7665 29124
rect 7699 29152 7711 29155
rect 8297 29155 8355 29161
rect 8297 29152 8309 29155
rect 7699 29124 8309 29152
rect 7699 29121 7711 29124
rect 7653 29115 7711 29121
rect 8297 29121 8309 29124
rect 8343 29121 8355 29155
rect 8297 29115 8355 29121
rect 7745 29087 7803 29093
rect 7745 29053 7757 29087
rect 7791 29084 7803 29087
rect 7926 29084 7932 29096
rect 7791 29056 7932 29084
rect 7791 29053 7803 29056
rect 7745 29047 7803 29053
rect 7926 29044 7932 29056
rect 7984 29084 7990 29096
rect 8110 29084 8116 29096
rect 7984 29056 8116 29084
rect 7984 29044 7990 29056
rect 8110 29044 8116 29056
rect 8168 29084 8174 29096
rect 8588 29084 8616 29192
rect 8665 29155 8723 29161
rect 8665 29121 8677 29155
rect 8711 29152 8723 29155
rect 8772 29152 8800 29248
rect 9582 29180 9588 29232
rect 9640 29220 9646 29232
rect 9953 29223 10011 29229
rect 9953 29220 9965 29223
rect 9640 29192 9965 29220
rect 9640 29180 9646 29192
rect 9953 29189 9965 29192
rect 9999 29220 10011 29223
rect 10413 29223 10471 29229
rect 9999 29192 10364 29220
rect 9999 29189 10011 29192
rect 9953 29183 10011 29189
rect 8711 29124 8800 29152
rect 8941 29155 8999 29161
rect 8711 29121 8723 29124
rect 8665 29115 8723 29121
rect 8941 29121 8953 29155
rect 8987 29152 8999 29155
rect 9398 29152 9404 29164
rect 8987 29124 9404 29152
rect 8987 29121 8999 29124
rect 8941 29115 8999 29121
rect 8956 29084 8984 29115
rect 9398 29112 9404 29124
rect 9456 29112 9462 29164
rect 9674 29112 9680 29164
rect 9732 29112 9738 29164
rect 9766 29112 9772 29164
rect 9824 29152 9830 29164
rect 10042 29152 10048 29164
rect 9824 29124 9869 29152
rect 9968 29124 10048 29152
rect 9824 29112 9830 29124
rect 9784 29084 9812 29112
rect 8168 29056 8524 29084
rect 8588 29056 8984 29084
rect 9692 29056 9812 29084
rect 8168 29044 8174 29056
rect 8021 29019 8079 29025
rect 8021 29016 8033 29019
rect 7484 28988 8033 29016
rect 8021 28985 8033 28988
rect 8067 29016 8079 29019
rect 8202 29016 8208 29028
rect 8067 28988 8208 29016
rect 8067 28985 8079 28988
rect 8021 28979 8079 28985
rect 8202 28976 8208 28988
rect 8260 28976 8266 29028
rect 8496 29025 8524 29056
rect 9692 29028 9720 29056
rect 8481 29019 8539 29025
rect 8481 28985 8493 29019
rect 8527 29016 8539 29019
rect 8757 29019 8815 29025
rect 8757 29016 8769 29019
rect 8527 28988 8769 29016
rect 8527 28985 8539 28988
rect 8481 28979 8539 28985
rect 8757 28985 8769 28988
rect 8803 29016 8815 29019
rect 9122 29016 9128 29028
rect 8803 28988 9128 29016
rect 8803 28985 8815 28988
rect 8757 28979 8815 28985
rect 9122 28976 9128 28988
rect 9180 28976 9186 29028
rect 9674 28976 9680 29028
rect 9732 28976 9738 29028
rect 9766 28976 9772 29028
rect 9824 29016 9830 29028
rect 9968 29016 9996 29124
rect 10042 29112 10048 29124
rect 10100 29112 10106 29164
rect 10183 29155 10241 29161
rect 10183 29121 10195 29155
rect 10229 29121 10241 29155
rect 10336 29152 10364 29192
rect 10413 29189 10425 29223
rect 10459 29220 10471 29223
rect 10502 29220 10508 29232
rect 10459 29192 10508 29220
rect 10459 29189 10471 29192
rect 10413 29183 10471 29189
rect 10502 29180 10508 29192
rect 10560 29180 10566 29232
rect 14366 29220 14372 29232
rect 12176 29192 14372 29220
rect 12176 29152 12204 29192
rect 14366 29180 14372 29192
rect 14424 29180 14430 29232
rect 14461 29223 14519 29229
rect 14461 29189 14473 29223
rect 14507 29220 14519 29223
rect 14642 29220 14648 29232
rect 14507 29192 14648 29220
rect 14507 29189 14519 29192
rect 14461 29183 14519 29189
rect 14642 29180 14648 29192
rect 14700 29180 14706 29232
rect 14752 29220 14780 29260
rect 14918 29248 14924 29300
rect 14976 29288 14982 29300
rect 15381 29291 15439 29297
rect 15381 29288 15393 29291
rect 14976 29260 15393 29288
rect 14976 29248 14982 29260
rect 15381 29257 15393 29260
rect 15427 29257 15439 29291
rect 16666 29288 16672 29300
rect 15381 29251 15439 29257
rect 15581 29260 16672 29288
rect 15013 29223 15071 29229
rect 15013 29220 15025 29223
rect 14752 29192 15025 29220
rect 15013 29189 15025 29192
rect 15059 29189 15071 29223
rect 15013 29183 15071 29189
rect 15229 29223 15287 29229
rect 15229 29189 15241 29223
rect 15275 29220 15287 29223
rect 15581 29220 15609 29260
rect 16666 29248 16672 29260
rect 16724 29288 16730 29300
rect 17310 29288 17316 29300
rect 16724 29260 17316 29288
rect 16724 29248 16730 29260
rect 17310 29248 17316 29260
rect 17368 29248 17374 29300
rect 18233 29291 18291 29297
rect 18233 29257 18245 29291
rect 18279 29288 18291 29291
rect 18782 29288 18788 29300
rect 18279 29260 18788 29288
rect 18279 29257 18291 29260
rect 18233 29251 18291 29257
rect 18782 29248 18788 29260
rect 18840 29248 18846 29300
rect 19242 29248 19248 29300
rect 19300 29288 19306 29300
rect 23014 29288 23020 29300
rect 19300 29260 20760 29288
rect 19300 29248 19306 29260
rect 15275 29192 15609 29220
rect 15275 29189 15287 29192
rect 15229 29183 15287 29189
rect 15654 29180 15660 29232
rect 15712 29220 15718 29232
rect 15712 29192 16344 29220
rect 15712 29180 15718 29192
rect 16316 29164 16344 29192
rect 16482 29180 16488 29232
rect 16540 29220 16546 29232
rect 19334 29220 19340 29232
rect 16540 29192 19340 29220
rect 16540 29180 16546 29192
rect 19334 29180 19340 29192
rect 19392 29180 19398 29232
rect 20622 29220 20628 29232
rect 19720 29192 20628 29220
rect 13814 29152 13820 29164
rect 10336 29124 12204 29152
rect 12636 29124 13820 29152
rect 10183 29115 10241 29121
rect 10198 29084 10226 29115
rect 11054 29084 11060 29096
rect 10198 29056 11060 29084
rect 11054 29044 11060 29056
rect 11112 29044 11118 29096
rect 12636 29093 12664 29124
rect 13814 29112 13820 29124
rect 13872 29112 13878 29164
rect 13924 29124 14596 29152
rect 12621 29087 12679 29093
rect 12621 29053 12633 29087
rect 12667 29053 12679 29087
rect 12621 29047 12679 29053
rect 12713 29087 12771 29093
rect 12713 29053 12725 29087
rect 12759 29084 12771 29087
rect 12894 29084 12900 29096
rect 12759 29056 12900 29084
rect 12759 29053 12771 29056
rect 12713 29047 12771 29053
rect 12894 29044 12900 29056
rect 12952 29084 12958 29096
rect 13630 29084 13636 29096
rect 12952 29056 13636 29084
rect 12952 29044 12958 29056
rect 13630 29044 13636 29056
rect 13688 29044 13694 29096
rect 13924 29016 13952 29124
rect 9824 28988 9996 29016
rect 10612 28988 13952 29016
rect 14568 29016 14596 29124
rect 14734 29112 14740 29164
rect 14792 29152 14798 29164
rect 14792 29124 15424 29152
rect 14792 29112 14798 29124
rect 14642 29044 14648 29096
rect 14700 29044 14706 29096
rect 14826 29044 14832 29096
rect 14884 29084 14890 29096
rect 15286 29084 15292 29096
rect 14884 29056 15292 29084
rect 14884 29044 14890 29056
rect 15286 29044 15292 29056
rect 15344 29044 15350 29096
rect 15396 29084 15424 29124
rect 15470 29112 15476 29164
rect 15528 29152 15534 29164
rect 15933 29155 15991 29161
rect 15933 29152 15945 29155
rect 15528 29124 15945 29152
rect 15528 29112 15534 29124
rect 15933 29121 15945 29124
rect 15979 29121 15991 29155
rect 15933 29115 15991 29121
rect 16114 29112 16120 29164
rect 16172 29112 16178 29164
rect 16298 29112 16304 29164
rect 16356 29112 16362 29164
rect 16666 29112 16672 29164
rect 16724 29152 16730 29164
rect 16945 29155 17003 29161
rect 16945 29152 16957 29155
rect 16724 29124 16957 29152
rect 16724 29112 16730 29124
rect 16945 29121 16957 29124
rect 16991 29121 17003 29155
rect 16945 29115 17003 29121
rect 17034 29112 17040 29164
rect 17092 29152 17098 29164
rect 17129 29155 17187 29161
rect 17129 29152 17141 29155
rect 17092 29124 17141 29152
rect 17092 29112 17098 29124
rect 17129 29121 17141 29124
rect 17175 29121 17187 29155
rect 17129 29115 17187 29121
rect 17221 29155 17279 29161
rect 17221 29121 17233 29155
rect 17267 29152 17279 29155
rect 17494 29152 17500 29164
rect 17267 29124 17500 29152
rect 17267 29121 17279 29124
rect 17221 29115 17279 29121
rect 17494 29112 17500 29124
rect 17552 29112 17558 29164
rect 18417 29155 18475 29161
rect 18417 29152 18429 29155
rect 17696 29124 18429 29152
rect 15562 29084 15568 29096
rect 15396 29056 15568 29084
rect 15562 29044 15568 29056
rect 15620 29044 15626 29096
rect 15749 29087 15807 29093
rect 15749 29053 15761 29087
rect 15795 29084 15807 29087
rect 16132 29084 16160 29112
rect 15795 29056 16160 29084
rect 15795 29053 15807 29056
rect 15749 29047 15807 29053
rect 14921 29019 14979 29025
rect 14921 29016 14933 29019
rect 14568 28988 14933 29016
rect 9824 28976 9830 28988
rect 4328 28951 4386 28957
rect 4328 28917 4340 28951
rect 4374 28948 4386 28951
rect 6012 28948 6040 28976
rect 10612 28957 10640 28988
rect 14921 28985 14933 28988
rect 14967 28985 14979 29019
rect 14921 28979 14979 28985
rect 16114 28976 16120 29028
rect 16172 28976 16178 29028
rect 16945 29019 17003 29025
rect 16945 28985 16957 29019
rect 16991 29016 17003 29019
rect 17696 29016 17724 29124
rect 18417 29121 18429 29124
rect 18463 29121 18475 29155
rect 18417 29115 18475 29121
rect 18598 29112 18604 29164
rect 18656 29112 18662 29164
rect 18969 29155 19027 29161
rect 18969 29152 18981 29155
rect 18708 29124 18981 29152
rect 18138 29044 18144 29096
rect 18196 29044 18202 29096
rect 18322 29044 18328 29096
rect 18380 29084 18386 29096
rect 18708 29084 18736 29124
rect 18969 29121 18981 29124
rect 19015 29121 19027 29155
rect 18969 29115 19027 29121
rect 19429 29155 19487 29161
rect 19429 29121 19441 29155
rect 19475 29152 19487 29155
rect 19518 29152 19524 29164
rect 19475 29124 19524 29152
rect 19475 29121 19487 29124
rect 19429 29115 19487 29121
rect 19518 29112 19524 29124
rect 19576 29112 19582 29164
rect 19720 29161 19748 29192
rect 20622 29180 20628 29192
rect 20680 29180 20686 29232
rect 20732 29220 20760 29260
rect 21008 29260 23020 29288
rect 21008 29229 21036 29260
rect 23014 29248 23020 29260
rect 23072 29248 23078 29300
rect 23106 29248 23112 29300
rect 23164 29288 23170 29300
rect 23164 29260 24256 29288
rect 23164 29248 23170 29260
rect 20993 29223 21051 29229
rect 20732 29192 20852 29220
rect 19705 29155 19763 29161
rect 19705 29121 19717 29155
rect 19751 29121 19763 29155
rect 19705 29115 19763 29121
rect 19978 29112 19984 29164
rect 20036 29152 20042 29164
rect 20257 29155 20315 29161
rect 20257 29152 20269 29155
rect 20036 29124 20269 29152
rect 20036 29112 20042 29124
rect 20257 29121 20269 29124
rect 20303 29121 20315 29155
rect 20257 29115 20315 29121
rect 18380 29056 18736 29084
rect 18380 29044 18386 29056
rect 18874 29044 18880 29096
rect 18932 29044 18938 29096
rect 20073 29087 20131 29093
rect 20073 29084 20085 29087
rect 18984 29056 20085 29084
rect 16991 28988 17724 29016
rect 16991 28985 17003 28988
rect 16945 28979 17003 28985
rect 17770 28976 17776 29028
rect 17828 29016 17834 29028
rect 18984 29016 19012 29056
rect 20073 29053 20085 29056
rect 20119 29053 20131 29087
rect 20073 29047 20131 29053
rect 19245 29019 19303 29025
rect 19245 29016 19257 29019
rect 17828 28988 19012 29016
rect 19076 28988 19257 29016
rect 17828 28976 17834 28988
rect 4374 28920 6040 28948
rect 10597 28951 10655 28957
rect 4374 28917 4386 28920
rect 4328 28911 4386 28917
rect 10597 28917 10609 28951
rect 10643 28917 10655 28951
rect 10597 28911 10655 28917
rect 10778 28908 10784 28960
rect 10836 28908 10842 28960
rect 13722 28908 13728 28960
rect 13780 28948 13786 28960
rect 14461 28951 14519 28957
rect 14461 28948 14473 28951
rect 13780 28920 14473 28948
rect 13780 28908 13786 28920
rect 14461 28917 14473 28920
rect 14507 28917 14519 28951
rect 14461 28911 14519 28917
rect 15197 28951 15255 28957
rect 15197 28917 15209 28951
rect 15243 28948 15255 28951
rect 15654 28948 15660 28960
rect 15243 28920 15660 28948
rect 15243 28917 15255 28920
rect 15197 28911 15255 28917
rect 15654 28908 15660 28920
rect 15712 28908 15718 28960
rect 16298 28908 16304 28960
rect 16356 28948 16362 28960
rect 17126 28948 17132 28960
rect 16356 28920 17132 28948
rect 16356 28908 16362 28920
rect 17126 28908 17132 28920
rect 17184 28908 17190 28960
rect 17678 28908 17684 28960
rect 17736 28948 17742 28960
rect 19076 28948 19104 28988
rect 19245 28985 19257 28988
rect 19291 28985 19303 29019
rect 19245 28979 19303 28985
rect 19613 29019 19671 29025
rect 19613 28985 19625 29019
rect 19659 29016 19671 29019
rect 20162 29016 20168 29028
rect 19659 28988 20168 29016
rect 19659 28985 19671 28988
rect 19613 28979 19671 28985
rect 20162 28976 20168 28988
rect 20220 28976 20226 29028
rect 20272 29016 20300 29115
rect 20346 29112 20352 29164
rect 20404 29112 20410 29164
rect 20438 29112 20444 29164
rect 20496 29112 20502 29164
rect 20533 29155 20591 29161
rect 20533 29121 20545 29155
rect 20579 29152 20591 29155
rect 20824 29152 20852 29192
rect 20993 29189 21005 29223
rect 21039 29189 21051 29223
rect 20993 29183 21051 29189
rect 21174 29180 21180 29232
rect 21232 29180 21238 29232
rect 21266 29180 21272 29232
rect 21324 29220 21330 29232
rect 23201 29223 23259 29229
rect 23201 29220 23213 29223
rect 21324 29192 23213 29220
rect 21324 29180 21330 29192
rect 22204 29161 22232 29192
rect 23201 29189 23213 29192
rect 23247 29189 23259 29223
rect 23983 29223 24041 29229
rect 23983 29220 23995 29223
rect 23201 29183 23259 29189
rect 23492 29192 23995 29220
rect 21361 29155 21419 29161
rect 21361 29152 21373 29155
rect 20579 29124 20760 29152
rect 20824 29124 21373 29152
rect 20579 29121 20591 29124
rect 20533 29115 20591 29121
rect 20732 29016 20760 29124
rect 21361 29121 21373 29124
rect 21407 29121 21419 29155
rect 21361 29115 21419 29121
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 22462 29112 22468 29164
rect 22520 29112 22526 29164
rect 22649 29155 22707 29161
rect 22649 29121 22661 29155
rect 22695 29121 22707 29155
rect 22649 29115 22707 29121
rect 21634 29044 21640 29096
rect 21692 29084 21698 29096
rect 22373 29087 22431 29093
rect 22373 29084 22385 29087
rect 21692 29056 22385 29084
rect 21692 29044 21698 29056
rect 22373 29053 22385 29056
rect 22419 29053 22431 29087
rect 22664 29084 22692 29115
rect 22738 29112 22744 29164
rect 22796 29112 22802 29164
rect 23109 29155 23167 29161
rect 23109 29121 23121 29155
rect 23155 29152 23167 29155
rect 23492 29152 23520 29192
rect 23983 29189 23995 29192
rect 24029 29220 24041 29223
rect 24029 29192 24164 29220
rect 24029 29189 24041 29192
rect 23983 29183 24041 29189
rect 23155 29124 23520 29152
rect 23569 29155 23627 29161
rect 23155 29121 23167 29124
rect 23109 29115 23167 29121
rect 23569 29121 23581 29155
rect 23615 29152 23627 29155
rect 23615 29124 23980 29152
rect 23615 29121 23627 29124
rect 23569 29115 23627 29121
rect 23952 29096 23980 29124
rect 22373 29047 22431 29053
rect 22480 29056 22692 29084
rect 23017 29087 23075 29093
rect 21358 29016 21364 29028
rect 20272 28988 20622 29016
rect 20732 28988 21364 29016
rect 17736 28920 19104 28948
rect 20594 28948 20622 28988
rect 21358 28976 21364 28988
rect 21416 28976 21422 29028
rect 21910 28976 21916 29028
rect 21968 28976 21974 29028
rect 22002 28976 22008 29028
rect 22060 28976 22066 29028
rect 22278 28976 22284 29028
rect 22336 28976 22342 29028
rect 21928 28948 21956 28976
rect 22480 28960 22508 29056
rect 23017 29053 23029 29087
rect 23063 29053 23075 29087
rect 23017 29047 23075 29053
rect 22554 28976 22560 29028
rect 22612 29016 22618 29028
rect 22612 28988 22692 29016
rect 22612 28976 22618 28988
rect 20594 28920 21956 28948
rect 17736 28908 17742 28920
rect 22462 28908 22468 28960
rect 22520 28908 22526 28960
rect 22664 28948 22692 28988
rect 22738 28976 22744 29028
rect 22796 29016 22802 29028
rect 23032 29016 23060 29047
rect 23198 29044 23204 29096
rect 23256 29084 23262 29096
rect 23256 29056 23704 29084
rect 23256 29044 23262 29056
rect 23676 29016 23704 29056
rect 23934 29044 23940 29096
rect 23992 29044 23998 29096
rect 24136 29084 24164 29192
rect 24228 29161 24256 29260
rect 25590 29248 25596 29300
rect 25648 29288 25654 29300
rect 26053 29291 26111 29297
rect 26053 29288 26065 29291
rect 25648 29260 26065 29288
rect 25648 29248 25654 29260
rect 26053 29257 26065 29260
rect 26099 29257 26111 29291
rect 26053 29251 26111 29257
rect 26510 29248 26516 29300
rect 26568 29288 26574 29300
rect 26694 29288 26700 29300
rect 26568 29260 26700 29288
rect 26568 29248 26574 29260
rect 26694 29248 26700 29260
rect 26752 29248 26758 29300
rect 27249 29291 27307 29297
rect 27249 29257 27261 29291
rect 27295 29288 27307 29291
rect 27338 29288 27344 29300
rect 27295 29260 27344 29288
rect 27295 29257 27307 29260
rect 27249 29251 27307 29257
rect 27338 29248 27344 29260
rect 27396 29248 27402 29300
rect 27890 29248 27896 29300
rect 27948 29288 27954 29300
rect 30469 29291 30527 29297
rect 30469 29288 30481 29291
rect 27948 29260 30481 29288
rect 27948 29248 27954 29260
rect 30469 29257 30481 29260
rect 30515 29257 30527 29291
rect 30469 29251 30527 29257
rect 31665 29291 31723 29297
rect 31665 29257 31677 29291
rect 31711 29288 31723 29291
rect 32214 29288 32220 29300
rect 31711 29260 32220 29288
rect 31711 29257 31723 29260
rect 31665 29251 31723 29257
rect 32214 29248 32220 29260
rect 32272 29248 32278 29300
rect 32674 29248 32680 29300
rect 32732 29288 32738 29300
rect 32732 29260 33916 29288
rect 32732 29248 32738 29260
rect 30098 29220 30104 29232
rect 24412 29192 30104 29220
rect 24213 29155 24271 29161
rect 24213 29121 24225 29155
rect 24259 29121 24271 29155
rect 24213 29115 24271 29121
rect 24302 29112 24308 29164
rect 24360 29112 24366 29164
rect 24412 29084 24440 29192
rect 30098 29180 30104 29192
rect 30156 29180 30162 29232
rect 30282 29180 30288 29232
rect 30340 29229 30346 29232
rect 30340 29223 30368 29229
rect 30356 29220 30368 29223
rect 31573 29223 31631 29229
rect 30356 29192 30604 29220
rect 30356 29189 30368 29192
rect 30340 29183 30368 29189
rect 30340 29180 30346 29183
rect 24486 29112 24492 29164
rect 24544 29112 24550 29164
rect 25133 29158 25191 29161
rect 24964 29155 25191 29158
rect 24964 29130 25145 29155
rect 24136 29056 24440 29084
rect 24578 29044 24584 29096
rect 24636 29084 24642 29096
rect 24857 29087 24915 29093
rect 24857 29084 24869 29087
rect 24636 29056 24869 29084
rect 24636 29044 24642 29056
rect 24857 29053 24869 29056
rect 24903 29053 24915 29087
rect 24964 29084 24992 29130
rect 25133 29121 25145 29130
rect 25179 29121 25191 29155
rect 25133 29115 25191 29121
rect 25222 29112 25228 29164
rect 25280 29152 25286 29164
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 25280 29124 25329 29152
rect 25280 29112 25286 29124
rect 25317 29121 25329 29124
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 25409 29155 25467 29161
rect 25409 29121 25421 29155
rect 25455 29121 25467 29155
rect 25409 29115 25467 29121
rect 25501 29155 25559 29161
rect 25501 29121 25513 29155
rect 25547 29152 25559 29155
rect 25682 29152 25688 29164
rect 25547 29124 25688 29152
rect 25547 29121 25559 29124
rect 25501 29115 25559 29121
rect 25424 29084 25452 29115
rect 25682 29112 25688 29124
rect 25740 29112 25746 29164
rect 25774 29112 25780 29164
rect 25832 29152 25838 29164
rect 25869 29155 25927 29161
rect 25869 29152 25881 29155
rect 25832 29124 25881 29152
rect 25832 29112 25838 29124
rect 25869 29121 25881 29124
rect 25915 29152 25927 29155
rect 25958 29152 25964 29164
rect 25915 29124 25964 29152
rect 25915 29121 25927 29124
rect 25869 29115 25927 29121
rect 25958 29112 25964 29124
rect 26016 29112 26022 29164
rect 26145 29155 26203 29161
rect 26145 29121 26157 29155
rect 26191 29152 26203 29155
rect 26418 29152 26424 29164
rect 26191 29124 26424 29152
rect 26191 29121 26203 29124
rect 26145 29115 26203 29121
rect 26418 29112 26424 29124
rect 26476 29112 26482 29164
rect 26510 29112 26516 29164
rect 26568 29112 26574 29164
rect 26602 29112 26608 29164
rect 26660 29152 26666 29164
rect 27338 29152 27344 29164
rect 26660 29124 27344 29152
rect 26660 29112 26666 29124
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 27433 29155 27491 29161
rect 27433 29121 27445 29155
rect 27479 29121 27491 29155
rect 27433 29115 27491 29121
rect 27617 29155 27675 29161
rect 27617 29121 27629 29155
rect 27663 29152 27675 29155
rect 27982 29152 27988 29164
rect 27663 29124 27988 29152
rect 27663 29121 27675 29124
rect 27617 29115 27675 29121
rect 24964 29056 25084 29084
rect 24857 29047 24915 29053
rect 24765 29019 24823 29025
rect 24765 29016 24777 29019
rect 22796 28988 23520 29016
rect 23676 28988 24777 29016
rect 22796 28976 22802 28988
rect 23385 28951 23443 28957
rect 23385 28948 23397 28951
rect 22664 28920 23397 28948
rect 23385 28917 23397 28920
rect 23431 28917 23443 28951
rect 23492 28948 23520 28988
rect 24765 28985 24777 28988
rect 24811 28985 24823 29019
rect 24765 28979 24823 28985
rect 23937 28951 23995 28957
rect 23937 28948 23949 28951
rect 23492 28920 23949 28948
rect 23385 28911 23443 28917
rect 23937 28917 23949 28920
rect 23983 28948 23995 28951
rect 24946 28948 24952 28960
rect 23983 28920 24952 28948
rect 23983 28917 23995 28920
rect 23937 28911 23995 28917
rect 24946 28908 24952 28920
rect 25004 28948 25010 28960
rect 25056 28948 25084 29056
rect 25332 29056 25452 29084
rect 25332 29028 25360 29056
rect 25590 29044 25596 29096
rect 25648 29084 25654 29096
rect 27448 29084 27476 29115
rect 27982 29112 27988 29124
rect 28040 29112 28046 29164
rect 28166 29112 28172 29164
rect 28224 29112 28230 29164
rect 28442 29112 28448 29164
rect 28500 29152 28506 29164
rect 28537 29155 28595 29161
rect 28537 29152 28549 29155
rect 28500 29124 28549 29152
rect 28500 29112 28506 29124
rect 28537 29121 28549 29124
rect 28583 29121 28595 29155
rect 28537 29115 28595 29121
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29152 29607 29155
rect 30006 29152 30012 29164
rect 29595 29124 30012 29152
rect 29595 29121 29607 29124
rect 29549 29115 29607 29121
rect 30006 29112 30012 29124
rect 30064 29112 30070 29164
rect 30576 29161 30604 29192
rect 31573 29189 31585 29223
rect 31619 29220 31631 29223
rect 32692 29220 32720 29248
rect 31619 29192 32720 29220
rect 31619 29189 31631 29192
rect 31573 29183 31631 29189
rect 30193 29155 30251 29161
rect 30193 29121 30205 29155
rect 30239 29152 30251 29155
rect 30561 29155 30619 29161
rect 30239 29124 30513 29152
rect 30239 29121 30251 29124
rect 30193 29115 30251 29121
rect 27706 29084 27712 29096
rect 25648 29056 25728 29084
rect 25648 29044 25654 29056
rect 25314 28976 25320 29028
rect 25372 28976 25378 29028
rect 25700 29025 25728 29056
rect 25976 29056 27712 29084
rect 25976 29028 26004 29056
rect 27706 29044 27712 29056
rect 27764 29044 27770 29096
rect 28184 29084 28212 29112
rect 28994 29084 29000 29096
rect 28184 29056 29000 29084
rect 28994 29044 29000 29056
rect 29052 29044 29058 29096
rect 29638 29044 29644 29096
rect 29696 29084 29702 29096
rect 29733 29087 29791 29093
rect 29733 29084 29745 29087
rect 29696 29056 29745 29084
rect 29696 29044 29702 29056
rect 29733 29053 29745 29056
rect 29779 29053 29791 29087
rect 29733 29047 29791 29053
rect 29822 29044 29828 29096
rect 29880 29044 29886 29096
rect 30101 29087 30159 29093
rect 30101 29053 30113 29087
rect 30147 29053 30159 29087
rect 30101 29047 30159 29053
rect 25685 29019 25743 29025
rect 25685 28985 25697 29019
rect 25731 28985 25743 29019
rect 25685 28979 25743 28985
rect 25958 28976 25964 29028
rect 26016 28976 26022 29028
rect 26234 28976 26240 29028
rect 26292 29016 26298 29028
rect 27890 29016 27896 29028
rect 26292 28988 27896 29016
rect 26292 28976 26298 28988
rect 27890 28976 27896 28988
rect 27948 28976 27954 29028
rect 28077 29019 28135 29025
rect 28077 28985 28089 29019
rect 28123 29016 28135 29019
rect 28123 28988 28157 29016
rect 28123 28985 28135 28988
rect 28077 28979 28135 28985
rect 25004 28920 25084 28948
rect 25004 28908 25010 28920
rect 25222 28908 25228 28960
rect 25280 28948 25286 28960
rect 25866 28948 25872 28960
rect 25280 28920 25872 28948
rect 25280 28908 25286 28920
rect 25866 28908 25872 28920
rect 25924 28908 25930 28960
rect 27614 28908 27620 28960
rect 27672 28948 27678 28960
rect 28092 28948 28120 28979
rect 29270 28976 29276 29028
rect 29328 29016 29334 29028
rect 30116 29016 30144 29047
rect 30374 29044 30380 29096
rect 30432 29044 30438 29096
rect 30485 29084 30513 29124
rect 30561 29121 30573 29155
rect 30607 29152 30619 29155
rect 31294 29152 31300 29164
rect 30607 29124 31300 29152
rect 30607 29121 30619 29124
rect 30561 29115 30619 29121
rect 31294 29112 31300 29124
rect 31352 29112 31358 29164
rect 30485 29056 30788 29084
rect 30392 29016 30420 29044
rect 30760 29028 30788 29056
rect 29328 28988 30420 29016
rect 29328 28976 29334 28988
rect 30742 28976 30748 29028
rect 30800 29016 30806 29028
rect 30837 29019 30895 29025
rect 30837 29016 30849 29019
rect 30800 28988 30849 29016
rect 30800 28976 30806 28988
rect 30837 28985 30849 28988
rect 30883 29016 30895 29019
rect 31588 29016 31616 29183
rect 31754 29112 31760 29164
rect 31812 29161 31818 29164
rect 31812 29155 31840 29161
rect 31828 29121 31840 29155
rect 31812 29115 31840 29121
rect 31812 29112 31818 29115
rect 32766 29112 32772 29164
rect 32824 29112 32830 29164
rect 33888 29161 33916 29260
rect 35710 29248 35716 29300
rect 35768 29288 35774 29300
rect 35989 29291 36047 29297
rect 35989 29288 36001 29291
rect 35768 29260 36001 29288
rect 35768 29248 35774 29260
rect 35989 29257 36001 29260
rect 36035 29257 36047 29291
rect 35989 29251 36047 29257
rect 36357 29291 36415 29297
rect 36357 29257 36369 29291
rect 36403 29288 36415 29291
rect 37550 29288 37556 29300
rect 36403 29260 37556 29288
rect 36403 29257 36415 29260
rect 36357 29251 36415 29257
rect 37550 29248 37556 29260
rect 37608 29248 37614 29300
rect 40954 29248 40960 29300
rect 41012 29248 41018 29300
rect 33597 29155 33655 29161
rect 33597 29121 33609 29155
rect 33643 29121 33655 29155
rect 33597 29115 33655 29121
rect 33873 29155 33931 29161
rect 33873 29121 33885 29155
rect 33919 29121 33931 29155
rect 33873 29115 33931 29121
rect 33612 29084 33640 29115
rect 34146 29112 34152 29164
rect 34204 29112 34210 29164
rect 34514 29112 34520 29164
rect 34572 29112 34578 29164
rect 40773 29155 40831 29161
rect 40773 29121 40785 29155
rect 40819 29152 40831 29155
rect 40819 29124 41368 29152
rect 40819 29121 40831 29124
rect 40773 29115 40831 29121
rect 34532 29084 34560 29112
rect 33612 29056 34560 29084
rect 36446 29044 36452 29096
rect 36504 29044 36510 29096
rect 36538 29044 36544 29096
rect 36596 29044 36602 29096
rect 41340 29028 41368 29124
rect 31941 29019 31999 29025
rect 31941 29016 31953 29019
rect 30883 28988 31616 29016
rect 31680 28988 31953 29016
rect 30883 28985 30895 28988
rect 30837 28979 30895 28985
rect 27672 28920 28120 28948
rect 27672 28908 27678 28920
rect 30190 28908 30196 28960
rect 30248 28948 30254 28960
rect 31021 28951 31079 28957
rect 31021 28948 31033 28951
rect 30248 28920 31033 28948
rect 30248 28908 30254 28920
rect 31021 28917 31033 28920
rect 31067 28917 31079 28951
rect 31021 28911 31079 28917
rect 31570 28908 31576 28960
rect 31628 28948 31634 28960
rect 31680 28948 31708 28988
rect 31941 28985 31953 28988
rect 31987 28985 31999 29019
rect 31941 28979 31999 28985
rect 41322 28976 41328 29028
rect 41380 28976 41386 29028
rect 31628 28920 31708 28948
rect 31628 28908 31634 28920
rect 32766 28908 32772 28960
rect 32824 28948 32830 28960
rect 33045 28951 33103 28957
rect 33045 28948 33057 28951
rect 32824 28920 33057 28948
rect 32824 28908 32830 28920
rect 33045 28917 33057 28920
rect 33091 28917 33103 28951
rect 33045 28911 33103 28917
rect 1104 28858 41400 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 41400 28858
rect 1104 28784 41400 28806
rect 5258 28704 5264 28756
rect 5316 28704 5322 28756
rect 5537 28747 5595 28753
rect 5537 28713 5549 28747
rect 5583 28744 5595 28747
rect 5886 28747 5944 28753
rect 5886 28744 5898 28747
rect 5583 28716 5898 28744
rect 5583 28713 5595 28716
rect 5537 28707 5595 28713
rect 5886 28713 5898 28716
rect 5932 28713 5944 28747
rect 5886 28707 5944 28713
rect 7377 28747 7435 28753
rect 7377 28713 7389 28747
rect 7423 28744 7435 28747
rect 7558 28744 7564 28756
rect 7423 28716 7564 28744
rect 7423 28713 7435 28716
rect 7377 28707 7435 28713
rect 7558 28704 7564 28716
rect 7616 28704 7622 28756
rect 9217 28747 9275 28753
rect 9217 28713 9229 28747
rect 9263 28744 9275 28747
rect 10226 28744 10232 28756
rect 9263 28716 10232 28744
rect 9263 28713 9275 28716
rect 9217 28707 9275 28713
rect 10226 28704 10232 28716
rect 10284 28704 10290 28756
rect 12250 28704 12256 28756
rect 12308 28744 12314 28756
rect 13998 28744 14004 28756
rect 12308 28716 14004 28744
rect 12308 28704 12314 28716
rect 13998 28704 14004 28716
rect 14056 28704 14062 28756
rect 14090 28704 14096 28756
rect 14148 28744 14154 28756
rect 14369 28747 14427 28753
rect 14369 28744 14381 28747
rect 14148 28716 14381 28744
rect 14148 28704 14154 28716
rect 14369 28713 14381 28716
rect 14415 28713 14427 28747
rect 14369 28707 14427 28713
rect 15654 28704 15660 28756
rect 15712 28704 15718 28756
rect 18598 28704 18604 28756
rect 18656 28744 18662 28756
rect 19426 28744 19432 28756
rect 18656 28716 19432 28744
rect 18656 28704 18662 28716
rect 19426 28704 19432 28716
rect 19484 28704 19490 28756
rect 19521 28747 19579 28753
rect 19521 28713 19533 28747
rect 19567 28744 19579 28747
rect 20622 28744 20628 28756
rect 19567 28716 20628 28744
rect 19567 28713 19579 28716
rect 19521 28707 19579 28713
rect 20622 28704 20628 28716
rect 20680 28704 20686 28756
rect 22738 28704 22744 28756
rect 22796 28744 22802 28756
rect 22833 28747 22891 28753
rect 22833 28744 22845 28747
rect 22796 28716 22845 28744
rect 22796 28704 22802 28716
rect 22833 28713 22845 28716
rect 22879 28744 22891 28747
rect 23198 28744 23204 28756
rect 22879 28716 23204 28744
rect 22879 28713 22891 28716
rect 22833 28707 22891 28713
rect 23198 28704 23204 28716
rect 23256 28704 23262 28756
rect 25038 28704 25044 28756
rect 25096 28744 25102 28756
rect 28902 28744 28908 28756
rect 25096 28716 26004 28744
rect 25096 28704 25102 28716
rect 4985 28543 5043 28549
rect 4985 28509 4997 28543
rect 5031 28509 5043 28543
rect 4985 28503 5043 28509
rect 5169 28543 5227 28549
rect 5169 28509 5181 28543
rect 5215 28540 5227 28543
rect 5276 28540 5304 28704
rect 9122 28636 9128 28688
rect 9180 28676 9186 28688
rect 15672 28676 15700 28704
rect 9180 28648 13216 28676
rect 15672 28648 22908 28676
rect 9180 28636 9186 28648
rect 5994 28608 6000 28620
rect 5368 28580 6000 28608
rect 5368 28549 5396 28580
rect 5994 28568 6000 28580
rect 6052 28568 6058 28620
rect 5215 28512 5304 28540
rect 5353 28543 5411 28549
rect 5215 28509 5227 28512
rect 5169 28503 5227 28509
rect 5353 28509 5365 28543
rect 5399 28509 5411 28543
rect 5353 28503 5411 28509
rect 5000 28404 5028 28503
rect 5534 28500 5540 28552
rect 5592 28540 5598 28552
rect 5629 28543 5687 28549
rect 5629 28540 5641 28543
rect 5592 28512 5641 28540
rect 5592 28500 5598 28512
rect 5629 28509 5641 28512
rect 5675 28509 5687 28543
rect 7282 28540 7288 28552
rect 7038 28512 7288 28540
rect 5629 28503 5687 28509
rect 7282 28500 7288 28512
rect 7340 28500 7346 28552
rect 8754 28500 8760 28552
rect 8812 28540 8818 28552
rect 9140 28549 9168 28636
rect 8941 28543 8999 28549
rect 8941 28540 8953 28543
rect 8812 28512 8953 28540
rect 8812 28500 8818 28512
rect 8941 28509 8953 28512
rect 8987 28509 8999 28543
rect 8941 28503 8999 28509
rect 9125 28543 9183 28549
rect 9125 28509 9137 28543
rect 9171 28509 9183 28543
rect 9125 28503 9183 28509
rect 9398 28500 9404 28552
rect 9456 28506 9462 28552
rect 10336 28549 10364 28648
rect 10410 28568 10416 28620
rect 10468 28608 10474 28620
rect 10468 28580 10916 28608
rect 10468 28568 10474 28580
rect 10321 28543 10379 28549
rect 10321 28509 10333 28543
rect 10367 28509 10379 28543
rect 9456 28500 9536 28506
rect 10321 28503 10379 28509
rect 10778 28500 10784 28552
rect 10836 28500 10842 28552
rect 10888 28540 10916 28580
rect 10962 28568 10968 28620
rect 11020 28608 11026 28620
rect 13081 28611 13139 28617
rect 13081 28608 13093 28611
rect 11020 28580 13093 28608
rect 11020 28568 11026 28580
rect 13081 28577 13093 28580
rect 13127 28577 13139 28611
rect 13081 28571 13139 28577
rect 10888 28512 11836 28540
rect 5261 28475 5319 28481
rect 5261 28441 5273 28475
rect 5307 28472 5319 28475
rect 6178 28472 6184 28484
rect 5307 28444 6184 28472
rect 5307 28441 5319 28444
rect 5261 28435 5319 28441
rect 6178 28432 6184 28444
rect 6236 28432 6242 28484
rect 9416 28478 9536 28500
rect 9508 28472 9536 28478
rect 10505 28475 10563 28481
rect 10505 28472 10517 28475
rect 9508 28444 10517 28472
rect 10505 28441 10517 28444
rect 10551 28441 10563 28475
rect 10505 28435 10563 28441
rect 10612 28444 11376 28472
rect 5902 28404 5908 28416
rect 5000 28376 5908 28404
rect 5902 28364 5908 28376
rect 5960 28404 5966 28416
rect 10612 28404 10640 28444
rect 11348 28416 11376 28444
rect 11514 28432 11520 28484
rect 11572 28432 11578 28484
rect 11808 28472 11836 28512
rect 11882 28500 11888 28552
rect 11940 28500 11946 28552
rect 11977 28543 12035 28549
rect 11977 28509 11989 28543
rect 12023 28509 12035 28543
rect 11977 28503 12035 28509
rect 11992 28472 12020 28503
rect 12158 28500 12164 28552
rect 12216 28500 12222 28552
rect 12253 28543 12311 28549
rect 12253 28509 12265 28543
rect 12299 28509 12311 28543
rect 12253 28503 12311 28509
rect 11808 28444 12020 28472
rect 12066 28432 12072 28484
rect 12124 28472 12130 28484
rect 12268 28472 12296 28503
rect 12526 28500 12532 28552
rect 12584 28540 12590 28552
rect 12713 28543 12771 28549
rect 12713 28540 12725 28543
rect 12584 28512 12725 28540
rect 12584 28500 12590 28512
rect 12713 28509 12725 28512
rect 12759 28509 12771 28543
rect 12713 28503 12771 28509
rect 12124 28444 12296 28472
rect 12728 28472 12756 28503
rect 12894 28500 12900 28552
rect 12952 28500 12958 28552
rect 13188 28540 13216 28648
rect 13354 28568 13360 28620
rect 13412 28608 13418 28620
rect 19334 28608 19340 28620
rect 13412 28580 19340 28608
rect 13412 28568 13418 28580
rect 19334 28568 19340 28580
rect 19392 28568 19398 28620
rect 19429 28611 19487 28617
rect 19429 28577 19441 28611
rect 19475 28608 19487 28611
rect 19475 28580 20208 28608
rect 19475 28577 19487 28580
rect 19429 28571 19487 28577
rect 20180 28552 20208 28580
rect 20824 28580 22094 28608
rect 14277 28543 14335 28549
rect 14277 28540 14289 28543
rect 13188 28512 14289 28540
rect 14277 28509 14289 28512
rect 14323 28540 14335 28543
rect 19521 28543 19579 28549
rect 14323 28512 19380 28540
rect 14323 28509 14335 28512
rect 14277 28503 14335 28509
rect 13538 28472 13544 28484
rect 12728 28444 13544 28472
rect 12124 28432 12130 28444
rect 13538 28432 13544 28444
rect 13596 28432 13602 28484
rect 13722 28432 13728 28484
rect 13780 28472 13786 28484
rect 14093 28475 14151 28481
rect 14093 28472 14105 28475
rect 13780 28444 14105 28472
rect 13780 28432 13786 28444
rect 14093 28441 14105 28444
rect 14139 28472 14151 28475
rect 16758 28472 16764 28484
rect 14139 28444 16764 28472
rect 14139 28441 14151 28444
rect 14093 28435 14151 28441
rect 16758 28432 16764 28444
rect 16816 28432 16822 28484
rect 17218 28432 17224 28484
rect 17276 28472 17282 28484
rect 18230 28472 18236 28484
rect 17276 28444 18236 28472
rect 17276 28432 17282 28444
rect 18230 28432 18236 28444
rect 18288 28432 18294 28484
rect 18966 28432 18972 28484
rect 19024 28472 19030 28484
rect 19242 28472 19248 28484
rect 19024 28444 19248 28472
rect 19024 28432 19030 28444
rect 19242 28432 19248 28444
rect 19300 28432 19306 28484
rect 19352 28472 19380 28512
rect 19521 28509 19533 28543
rect 19567 28540 19579 28543
rect 19978 28540 19984 28552
rect 19567 28512 19984 28540
rect 19567 28509 19579 28512
rect 19521 28503 19579 28509
rect 19978 28500 19984 28512
rect 20036 28500 20042 28552
rect 20162 28500 20168 28552
rect 20220 28500 20226 28552
rect 20349 28543 20407 28549
rect 20349 28509 20361 28543
rect 20395 28540 20407 28543
rect 20438 28540 20444 28552
rect 20395 28512 20444 28540
rect 20395 28509 20407 28512
rect 20349 28503 20407 28509
rect 20438 28500 20444 28512
rect 20496 28500 20502 28552
rect 20533 28543 20591 28549
rect 20533 28509 20545 28543
rect 20579 28540 20591 28543
rect 20622 28540 20628 28552
rect 20579 28512 20628 28540
rect 20579 28509 20591 28512
rect 20533 28503 20591 28509
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 19352 28444 19840 28472
rect 5960 28376 10640 28404
rect 10689 28407 10747 28413
rect 5960 28364 5966 28376
rect 10689 28373 10701 28407
rect 10735 28404 10747 28407
rect 10870 28404 10876 28416
rect 10735 28376 10876 28404
rect 10735 28373 10747 28376
rect 10689 28367 10747 28373
rect 10870 28364 10876 28376
rect 10928 28364 10934 28416
rect 11330 28364 11336 28416
rect 11388 28364 11394 28416
rect 12342 28364 12348 28416
rect 12400 28364 12406 28416
rect 12434 28364 12440 28416
rect 12492 28404 12498 28416
rect 15102 28404 15108 28416
rect 12492 28376 15108 28404
rect 12492 28364 12498 28376
rect 15102 28364 15108 28376
rect 15160 28364 15166 28416
rect 17126 28364 17132 28416
rect 17184 28404 17190 28416
rect 18506 28404 18512 28416
rect 17184 28376 18512 28404
rect 17184 28364 17190 28376
rect 18506 28364 18512 28376
rect 18564 28404 18570 28416
rect 18874 28404 18880 28416
rect 18564 28376 18880 28404
rect 18564 28364 18570 28376
rect 18874 28364 18880 28376
rect 18932 28364 18938 28416
rect 19150 28364 19156 28416
rect 19208 28404 19214 28416
rect 19705 28407 19763 28413
rect 19705 28404 19717 28407
rect 19208 28376 19717 28404
rect 19208 28364 19214 28376
rect 19705 28373 19717 28376
rect 19751 28373 19763 28407
rect 19812 28404 19840 28444
rect 20714 28432 20720 28484
rect 20772 28432 20778 28484
rect 20824 28404 20852 28580
rect 21269 28543 21327 28549
rect 21269 28509 21281 28543
rect 21315 28509 21327 28543
rect 21269 28503 21327 28509
rect 19812 28376 20852 28404
rect 21284 28404 21312 28503
rect 21634 28500 21640 28552
rect 21692 28500 21698 28552
rect 21358 28432 21364 28484
rect 21416 28472 21422 28484
rect 21453 28475 21511 28481
rect 21453 28472 21465 28475
rect 21416 28444 21465 28472
rect 21416 28432 21422 28444
rect 21453 28441 21465 28444
rect 21499 28441 21511 28475
rect 21453 28435 21511 28441
rect 21542 28432 21548 28484
rect 21600 28432 21606 28484
rect 22066 28472 22094 28580
rect 22554 28472 22560 28484
rect 22066 28444 22560 28472
rect 22554 28432 22560 28444
rect 22612 28472 22618 28484
rect 22880 28481 22908 28648
rect 24578 28636 24584 28688
rect 24636 28676 24642 28688
rect 25774 28676 25780 28688
rect 24636 28648 25780 28676
rect 24636 28636 24642 28648
rect 25774 28636 25780 28648
rect 25832 28636 25838 28688
rect 25866 28636 25872 28688
rect 25924 28636 25930 28688
rect 25976 28685 26004 28716
rect 28184 28716 28908 28744
rect 28184 28685 28212 28716
rect 28902 28704 28908 28716
rect 28960 28704 28966 28756
rect 29549 28747 29607 28753
rect 29549 28713 29561 28747
rect 29595 28744 29607 28747
rect 29638 28744 29644 28756
rect 29595 28716 29644 28744
rect 29595 28713 29607 28716
rect 29549 28707 29607 28713
rect 29638 28704 29644 28716
rect 29696 28704 29702 28756
rect 39114 28704 39120 28756
rect 39172 28704 39178 28756
rect 25961 28679 26019 28685
rect 25961 28645 25973 28679
rect 26007 28645 26019 28679
rect 28169 28679 28227 28685
rect 28169 28676 28181 28679
rect 25961 28639 26019 28645
rect 27356 28648 28181 28676
rect 24949 28611 25007 28617
rect 24949 28577 24961 28611
rect 24995 28608 25007 28611
rect 27356 28608 27384 28648
rect 28169 28645 28181 28648
rect 28215 28645 28227 28679
rect 34238 28676 34244 28688
rect 28169 28639 28227 28645
rect 28736 28648 34244 28676
rect 24995 28580 27384 28608
rect 27632 28580 28028 28608
rect 24995 28577 25007 28580
rect 24949 28571 25007 28577
rect 27632 28552 27660 28580
rect 24302 28500 24308 28552
rect 24360 28540 24366 28552
rect 24397 28543 24455 28549
rect 24397 28540 24409 28543
rect 24360 28512 24409 28540
rect 24360 28500 24366 28512
rect 24397 28509 24409 28512
rect 24443 28509 24455 28543
rect 24397 28503 24455 28509
rect 24581 28543 24639 28549
rect 24581 28509 24593 28543
rect 24627 28540 24639 28543
rect 24670 28540 24676 28552
rect 24627 28512 24676 28540
rect 24627 28509 24639 28512
rect 24581 28503 24639 28509
rect 24670 28500 24676 28512
rect 24728 28540 24734 28552
rect 24728 28512 25636 28540
rect 24728 28500 24734 28512
rect 22649 28475 22707 28481
rect 22649 28472 22661 28475
rect 22612 28444 22661 28472
rect 22612 28432 22618 28444
rect 22649 28441 22661 28444
rect 22695 28441 22707 28475
rect 22649 28435 22707 28441
rect 22865 28475 22923 28481
rect 22865 28441 22877 28475
rect 22911 28472 22923 28475
rect 23566 28472 23572 28484
rect 22911 28444 23572 28472
rect 22911 28441 22923 28444
rect 22865 28435 22923 28441
rect 23566 28432 23572 28444
rect 23624 28432 23630 28484
rect 21634 28404 21640 28416
rect 21284 28376 21640 28404
rect 19705 28367 19763 28373
rect 21634 28364 21640 28376
rect 21692 28364 21698 28416
rect 21821 28407 21879 28413
rect 21821 28373 21833 28407
rect 21867 28404 21879 28407
rect 21910 28404 21916 28416
rect 21867 28376 21916 28404
rect 21867 28373 21879 28376
rect 21821 28367 21879 28373
rect 21910 28364 21916 28376
rect 21968 28364 21974 28416
rect 23014 28364 23020 28416
rect 23072 28364 23078 28416
rect 23474 28364 23480 28416
rect 23532 28404 23538 28416
rect 24581 28407 24639 28413
rect 24581 28404 24593 28407
rect 23532 28376 24593 28404
rect 23532 28364 23538 28376
rect 24581 28373 24593 28376
rect 24627 28373 24639 28407
rect 25608 28404 25636 28512
rect 26602 28500 26608 28552
rect 26660 28500 26666 28552
rect 26973 28543 27031 28549
rect 26973 28509 26985 28543
rect 27019 28509 27031 28543
rect 26973 28503 27031 28509
rect 26988 28404 27016 28503
rect 27154 28500 27160 28552
rect 27212 28500 27218 28552
rect 27614 28500 27620 28552
rect 27672 28500 27678 28552
rect 28000 28549 28028 28580
rect 27801 28543 27859 28549
rect 27801 28509 27813 28543
rect 27847 28509 27859 28543
rect 27801 28503 27859 28509
rect 27985 28543 28043 28549
rect 27985 28509 27997 28543
rect 28031 28509 28043 28543
rect 27985 28503 28043 28509
rect 27816 28472 27844 28503
rect 28626 28500 28632 28552
rect 28684 28500 28690 28552
rect 28534 28472 28540 28484
rect 27816 28444 28540 28472
rect 28534 28432 28540 28444
rect 28592 28472 28598 28484
rect 28736 28472 28764 28648
rect 34238 28636 34244 28648
rect 34296 28636 34302 28688
rect 37369 28611 37427 28617
rect 29656 28580 34100 28608
rect 28994 28500 29000 28552
rect 29052 28540 29058 28552
rect 29089 28543 29147 28549
rect 29089 28540 29101 28543
rect 29052 28512 29101 28540
rect 29052 28500 29058 28512
rect 29089 28509 29101 28512
rect 29135 28509 29147 28543
rect 29089 28503 29147 28509
rect 29546 28500 29552 28552
rect 29604 28540 29610 28552
rect 29656 28540 29684 28580
rect 34072 28552 34100 28580
rect 37369 28577 37381 28611
rect 37415 28608 37427 28611
rect 38102 28608 38108 28620
rect 37415 28580 38108 28608
rect 37415 28577 37427 28580
rect 37369 28571 37427 28577
rect 38102 28568 38108 28580
rect 38160 28568 38166 28620
rect 29604 28512 29684 28540
rect 29733 28543 29791 28549
rect 29604 28500 29610 28512
rect 29733 28509 29745 28543
rect 29779 28540 29791 28543
rect 29822 28540 29828 28552
rect 29779 28512 29828 28540
rect 29779 28509 29791 28512
rect 29733 28503 29791 28509
rect 29822 28500 29828 28512
rect 29880 28500 29886 28552
rect 30101 28543 30159 28549
rect 30101 28509 30113 28543
rect 30147 28540 30159 28543
rect 30190 28540 30196 28552
rect 30147 28512 30196 28540
rect 30147 28509 30159 28512
rect 30101 28503 30159 28509
rect 30190 28500 30196 28512
rect 30248 28500 30254 28552
rect 30285 28543 30343 28549
rect 30285 28509 30297 28543
rect 30331 28542 30343 28543
rect 30331 28514 30420 28542
rect 30331 28509 30343 28514
rect 30285 28503 30343 28509
rect 28592 28444 28764 28472
rect 28592 28432 28598 28444
rect 29914 28432 29920 28484
rect 29972 28472 29978 28484
rect 30392 28472 30420 28514
rect 34054 28500 34060 28552
rect 34112 28500 34118 28552
rect 37274 28500 37280 28552
rect 37332 28500 37338 28552
rect 37645 28475 37703 28481
rect 37645 28472 37657 28475
rect 29972 28444 30420 28472
rect 37108 28444 37657 28472
rect 29972 28432 29978 28444
rect 27706 28404 27712 28416
rect 25608 28376 27712 28404
rect 24581 28367 24639 28373
rect 27706 28364 27712 28376
rect 27764 28364 27770 28416
rect 28350 28364 28356 28416
rect 28408 28404 28414 28416
rect 28718 28404 28724 28416
rect 28408 28376 28724 28404
rect 28408 28364 28414 28376
rect 28718 28364 28724 28376
rect 28776 28364 28782 28416
rect 30282 28364 30288 28416
rect 30340 28364 30346 28416
rect 31754 28364 31760 28416
rect 31812 28404 31818 28416
rect 33410 28404 33416 28416
rect 31812 28376 33416 28404
rect 31812 28364 31818 28376
rect 33410 28364 33416 28376
rect 33468 28364 33474 28416
rect 37108 28413 37136 28444
rect 37645 28441 37657 28444
rect 37691 28441 37703 28475
rect 37645 28435 37703 28441
rect 37918 28432 37924 28484
rect 37976 28472 37982 28484
rect 38102 28472 38108 28484
rect 37976 28444 38108 28472
rect 37976 28432 37982 28444
rect 38102 28432 38108 28444
rect 38160 28432 38166 28484
rect 37093 28407 37151 28413
rect 37093 28373 37105 28407
rect 37139 28373 37151 28407
rect 37093 28367 37151 28373
rect 1104 28314 41400 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 41400 28314
rect 1104 28240 41400 28262
rect 8938 28160 8944 28212
rect 8996 28160 9002 28212
rect 10962 28200 10968 28212
rect 10796 28172 10968 28200
rect 8294 28092 8300 28144
rect 8352 28132 8358 28144
rect 8570 28132 8576 28144
rect 8352 28104 8576 28132
rect 8352 28092 8358 28104
rect 8570 28092 8576 28104
rect 8628 28092 8634 28144
rect 9585 28135 9643 28141
rect 9585 28132 9597 28135
rect 8864 28104 9597 28132
rect 1394 28024 1400 28076
rect 1452 28024 1458 28076
rect 4249 28067 4307 28073
rect 4249 28033 4261 28067
rect 4295 28064 4307 28067
rect 4798 28064 4804 28076
rect 4295 28036 4804 28064
rect 4295 28033 4307 28036
rect 4249 28027 4307 28033
rect 4798 28024 4804 28036
rect 4856 28064 4862 28076
rect 5350 28064 5356 28076
rect 4856 28036 5356 28064
rect 4856 28024 4862 28036
rect 5350 28024 5356 28036
rect 5408 28024 5414 28076
rect 8018 28024 8024 28076
rect 8076 28024 8082 28076
rect 8864 28073 8892 28104
rect 9585 28101 9597 28104
rect 9631 28101 9643 28135
rect 9585 28095 9643 28101
rect 8849 28067 8907 28073
rect 8849 28033 8861 28067
rect 8895 28033 8907 28067
rect 8849 28027 8907 28033
rect 9122 28024 9128 28076
rect 9180 28064 9186 28076
rect 9217 28067 9275 28073
rect 9217 28064 9229 28067
rect 9180 28036 9229 28064
rect 9180 28024 9186 28036
rect 9217 28033 9229 28036
rect 9263 28033 9275 28067
rect 9217 28027 9275 28033
rect 9309 28067 9367 28073
rect 9309 28033 9321 28067
rect 9355 28033 9367 28067
rect 9309 28027 9367 28033
rect 9401 28067 9459 28073
rect 9401 28033 9413 28067
rect 9447 28064 9459 28067
rect 10796 28064 10824 28172
rect 10962 28160 10968 28172
rect 11020 28160 11026 28212
rect 11054 28160 11060 28212
rect 11112 28160 11118 28212
rect 11330 28160 11336 28212
rect 11388 28200 11394 28212
rect 18414 28200 18420 28212
rect 11388 28172 12664 28200
rect 11388 28160 11394 28172
rect 9447 28036 10824 28064
rect 9447 28033 9459 28036
rect 9401 28027 9459 28033
rect 3786 27956 3792 28008
rect 3844 27996 3850 28008
rect 4985 27999 5043 28005
rect 4985 27996 4997 27999
rect 3844 27968 4997 27996
rect 3844 27956 3850 27968
rect 4985 27965 4997 27968
rect 5031 27996 5043 27999
rect 5534 27996 5540 28008
rect 5031 27968 5540 27996
rect 5031 27965 5043 27968
rect 4985 27959 5043 27965
rect 5534 27956 5540 27968
rect 5592 27956 5598 28008
rect 8294 27956 8300 28008
rect 8352 27996 8358 28008
rect 9033 27999 9091 28005
rect 9033 27996 9045 27999
rect 8352 27968 9045 27996
rect 8352 27956 8358 27968
rect 9033 27965 9045 27968
rect 9079 27965 9091 27999
rect 9324 27996 9352 28027
rect 9033 27959 9091 27965
rect 9140 27968 9352 27996
rect 934 27888 940 27940
rect 992 27928 998 27940
rect 1581 27931 1639 27937
rect 1581 27928 1593 27931
rect 992 27900 1593 27928
rect 992 27888 998 27900
rect 1581 27897 1593 27900
rect 1627 27897 1639 27931
rect 1581 27891 1639 27897
rect 8938 27888 8944 27940
rect 8996 27928 9002 27940
rect 9140 27928 9168 27968
rect 9490 27956 9496 28008
rect 9548 27996 9554 28008
rect 9585 27999 9643 28005
rect 9585 27996 9597 27999
rect 9548 27968 9597 27996
rect 9548 27956 9554 27968
rect 9585 27965 9597 27968
rect 9631 27965 9643 27999
rect 9585 27959 9643 27965
rect 10594 27956 10600 28008
rect 10652 27956 10658 28008
rect 11072 27996 11100 28160
rect 12526 28092 12532 28144
rect 12584 28092 12590 28144
rect 12434 28073 12440 28076
rect 12253 28067 12311 28073
rect 12253 28033 12265 28067
rect 12299 28033 12311 28067
rect 12253 28027 12311 28033
rect 12401 28067 12440 28073
rect 12401 28033 12413 28067
rect 12401 28027 12440 28033
rect 11146 27996 11152 28008
rect 10796 27968 11008 27996
rect 11072 27968 11152 27996
rect 8996 27900 9168 27928
rect 9217 27931 9275 27937
rect 8996 27888 9002 27900
rect 9217 27897 9229 27931
rect 9263 27928 9275 27931
rect 10796 27928 10824 27968
rect 9263 27900 10824 27928
rect 9263 27897 9275 27900
rect 9217 27891 9275 27897
rect 10870 27888 10876 27940
rect 10928 27888 10934 27940
rect 10980 27928 11008 27968
rect 11146 27956 11152 27968
rect 11204 27956 11210 28008
rect 12268 27996 12296 28027
rect 12434 28024 12440 28027
rect 12492 28024 12498 28076
rect 12636 28073 12664 28172
rect 13648 28172 18420 28200
rect 12621 28067 12679 28073
rect 12621 28033 12633 28067
rect 12667 28033 12679 28067
rect 12621 28027 12679 28033
rect 12759 28067 12817 28073
rect 12759 28033 12771 28067
rect 12805 28064 12817 28067
rect 13648 28064 13676 28172
rect 18414 28160 18420 28172
rect 18472 28160 18478 28212
rect 18785 28203 18843 28209
rect 18785 28169 18797 28203
rect 18831 28169 18843 28203
rect 18785 28163 18843 28169
rect 12805 28036 13676 28064
rect 13740 28104 15148 28132
rect 12805 28033 12817 28036
rect 12759 28027 12817 28033
rect 12526 27996 12532 28008
rect 12268 27968 12532 27996
rect 12526 27956 12532 27968
rect 12584 27956 12590 28008
rect 12636 27996 12664 28027
rect 13630 27996 13636 28008
rect 12636 27968 13636 27996
rect 13630 27956 13636 27968
rect 13688 27956 13694 28008
rect 13740 27928 13768 28104
rect 14826 28024 14832 28076
rect 14884 28024 14890 28076
rect 14918 28024 14924 28076
rect 14976 28024 14982 28076
rect 15120 28073 15148 28104
rect 15654 28092 15660 28144
rect 15712 28132 15718 28144
rect 17957 28135 18015 28141
rect 15712 28104 16344 28132
rect 15712 28092 15718 28104
rect 15105 28067 15163 28073
rect 15105 28033 15117 28067
rect 15151 28033 15163 28067
rect 15105 28027 15163 28033
rect 15194 28024 15200 28076
rect 15252 28024 15258 28076
rect 15470 28024 15476 28076
rect 15528 28064 15534 28076
rect 16316 28073 16344 28104
rect 17957 28101 17969 28135
rect 18003 28132 18015 28135
rect 18003 28104 18276 28132
rect 18003 28101 18015 28104
rect 17957 28095 18015 28101
rect 15749 28067 15807 28073
rect 15749 28064 15761 28067
rect 15528 28036 15761 28064
rect 15528 28024 15534 28036
rect 15749 28033 15761 28036
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28033 15991 28067
rect 15933 28027 15991 28033
rect 16301 28067 16359 28073
rect 16301 28033 16313 28067
rect 16347 28064 16359 28067
rect 17310 28064 17316 28076
rect 16347 28036 17316 28064
rect 16347 28033 16359 28036
rect 16301 28027 16359 28033
rect 15013 27999 15071 28005
rect 15013 27965 15025 27999
rect 15059 27996 15071 27999
rect 15212 27996 15240 28024
rect 15059 27968 15240 27996
rect 15059 27965 15071 27968
rect 15013 27959 15071 27965
rect 10980 27900 13768 27928
rect 13906 27888 13912 27940
rect 13964 27928 13970 27940
rect 14550 27928 14556 27940
rect 13964 27900 14556 27928
rect 13964 27888 13970 27900
rect 14550 27888 14556 27900
rect 14608 27888 14614 27940
rect 14642 27888 14648 27940
rect 14700 27888 14706 27940
rect 14826 27888 14832 27940
rect 14884 27928 14890 27940
rect 15948 27928 15976 28027
rect 17310 28024 17316 28036
rect 17368 28024 17374 28076
rect 18248 28073 18276 28104
rect 17681 28067 17739 28073
rect 17681 28033 17693 28067
rect 17727 28064 17739 28067
rect 18233 28067 18291 28073
rect 17727 28036 18092 28064
rect 17727 28033 17739 28036
rect 17681 28027 17739 28033
rect 16114 27956 16120 28008
rect 16172 27996 16178 28008
rect 17954 27996 17960 28008
rect 16172 27968 17960 27996
rect 16172 27956 16178 27968
rect 17954 27956 17960 27968
rect 18012 27956 18018 28008
rect 17586 27928 17592 27940
rect 14884 27900 17592 27928
rect 14884 27888 14890 27900
rect 17586 27888 17592 27900
rect 17644 27888 17650 27940
rect 18064 27928 18092 28036
rect 18233 28033 18245 28067
rect 18279 28033 18291 28067
rect 18233 28027 18291 28033
rect 18601 28067 18659 28073
rect 18601 28033 18613 28067
rect 18647 28033 18659 28067
rect 18601 28027 18659 28033
rect 18138 27956 18144 28008
rect 18196 27956 18202 28008
rect 18616 27996 18644 28027
rect 18544 27968 18644 27996
rect 18800 27996 18828 28163
rect 18874 28160 18880 28212
rect 18932 28160 18938 28212
rect 19058 28160 19064 28212
rect 19116 28200 19122 28212
rect 19518 28200 19524 28212
rect 19116 28172 19524 28200
rect 19116 28160 19122 28172
rect 19518 28160 19524 28172
rect 19576 28160 19582 28212
rect 20346 28160 20352 28212
rect 20404 28200 20410 28212
rect 27154 28200 27160 28212
rect 20404 28172 27160 28200
rect 20404 28160 20410 28172
rect 27154 28160 27160 28172
rect 27212 28160 27218 28212
rect 27338 28160 27344 28212
rect 27396 28200 27402 28212
rect 27798 28200 27804 28212
rect 27396 28172 27804 28200
rect 27396 28160 27402 28172
rect 27798 28160 27804 28172
rect 27856 28160 27862 28212
rect 31938 28200 31944 28212
rect 30668 28172 31944 28200
rect 18892 28132 18920 28160
rect 18892 28104 19012 28132
rect 18874 28024 18880 28076
rect 18932 28024 18938 28076
rect 18984 28073 19012 28104
rect 19242 28092 19248 28144
rect 19300 28092 19306 28144
rect 22738 28092 22744 28144
rect 22796 28132 22802 28144
rect 26602 28132 26608 28144
rect 22796 28104 26608 28132
rect 22796 28092 22802 28104
rect 26602 28092 26608 28104
rect 26660 28092 26666 28144
rect 27816 28132 27844 28160
rect 27632 28104 27844 28132
rect 18970 28067 19028 28073
rect 18970 28033 18982 28067
rect 19016 28033 19028 28067
rect 18970 28027 19028 28033
rect 19150 28024 19156 28076
rect 19208 28024 19214 28076
rect 19342 28067 19400 28073
rect 19342 28033 19354 28067
rect 19388 28033 19400 28067
rect 19342 28027 19400 28033
rect 19352 27996 19380 28027
rect 20438 28024 20444 28076
rect 20496 28024 20502 28076
rect 20714 28024 20720 28076
rect 20772 28064 20778 28076
rect 25038 28064 25044 28076
rect 20772 28036 25044 28064
rect 20772 28024 20778 28036
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 25314 28024 25320 28076
rect 25372 28064 25378 28076
rect 26142 28064 26148 28076
rect 25372 28036 26148 28064
rect 25372 28024 25378 28036
rect 26142 28024 26148 28036
rect 26200 28024 26206 28076
rect 26510 28024 26516 28076
rect 26568 28064 26574 28076
rect 27341 28067 27399 28073
rect 27341 28064 27353 28067
rect 26568 28036 27353 28064
rect 26568 28024 26574 28036
rect 27341 28033 27353 28036
rect 27387 28064 27399 28067
rect 27430 28064 27436 28076
rect 27387 28036 27436 28064
rect 27387 28033 27399 28036
rect 27341 28027 27399 28033
rect 27430 28024 27436 28036
rect 27488 28024 27494 28076
rect 27525 28067 27583 28073
rect 27525 28033 27537 28067
rect 27571 28064 27583 28067
rect 27632 28064 27660 28104
rect 27982 28092 27988 28144
rect 28040 28132 28046 28144
rect 30668 28141 30696 28172
rect 31938 28160 31944 28172
rect 31996 28160 32002 28212
rect 32674 28160 32680 28212
rect 32732 28160 32738 28212
rect 32858 28160 32864 28212
rect 32916 28160 32922 28212
rect 33410 28160 33416 28212
rect 33468 28160 33474 28212
rect 33597 28203 33655 28209
rect 33597 28169 33609 28203
rect 33643 28200 33655 28203
rect 34054 28200 34060 28212
rect 33643 28172 34060 28200
rect 33643 28169 33655 28172
rect 33597 28163 33655 28169
rect 34054 28160 34060 28172
rect 34112 28160 34118 28212
rect 34238 28160 34244 28212
rect 34296 28160 34302 28212
rect 34517 28203 34575 28209
rect 34517 28169 34529 28203
rect 34563 28200 34575 28203
rect 34885 28203 34943 28209
rect 34885 28200 34897 28203
rect 34563 28172 34897 28200
rect 34563 28169 34575 28172
rect 34517 28163 34575 28169
rect 34885 28169 34897 28172
rect 34931 28169 34943 28203
rect 34885 28163 34943 28169
rect 37274 28160 37280 28212
rect 37332 28200 37338 28212
rect 37369 28203 37427 28209
rect 37369 28200 37381 28203
rect 37332 28172 37381 28200
rect 37332 28160 37338 28172
rect 37369 28169 37381 28172
rect 37415 28169 37427 28203
rect 37369 28163 37427 28169
rect 37737 28203 37795 28209
rect 37737 28169 37749 28203
rect 37783 28200 37795 28203
rect 39117 28203 39175 28209
rect 39117 28200 39129 28203
rect 37783 28172 39129 28200
rect 37783 28169 37795 28172
rect 37737 28163 37795 28169
rect 39117 28169 39129 28172
rect 39163 28169 39175 28203
rect 39117 28163 39175 28169
rect 30653 28135 30711 28141
rect 28040 28104 30144 28132
rect 28040 28092 28046 28104
rect 27571 28036 27660 28064
rect 27571 28033 27583 28036
rect 27525 28027 27583 28033
rect 27706 28024 27712 28076
rect 27764 28064 27770 28076
rect 29825 28067 29883 28073
rect 29825 28064 29837 28067
rect 27764 28036 29837 28064
rect 27764 28024 27770 28036
rect 29825 28033 29837 28036
rect 29871 28064 29883 28067
rect 30116 28064 30144 28104
rect 30653 28101 30665 28135
rect 30699 28101 30711 28135
rect 30653 28095 30711 28101
rect 30834 28092 30840 28144
rect 30892 28092 30898 28144
rect 31018 28092 31024 28144
rect 31076 28092 31082 28144
rect 33045 28135 33103 28141
rect 33045 28132 33057 28135
rect 31680 28104 33057 28132
rect 31110 28064 31116 28076
rect 29871 28036 30052 28064
rect 30116 28036 31116 28064
rect 29871 28033 29883 28036
rect 29825 28027 29883 28033
rect 18800 27968 19380 27996
rect 18414 27928 18420 27940
rect 18064 27900 18420 27928
rect 18414 27888 18420 27900
rect 18472 27888 18478 27940
rect 18544 27928 18572 27968
rect 20456 27928 20484 28024
rect 20622 27956 20628 28008
rect 20680 27996 20686 28008
rect 20898 27996 20904 28008
rect 20680 27968 20904 27996
rect 20680 27956 20686 27968
rect 20898 27956 20904 27968
rect 20956 27956 20962 28008
rect 21450 27956 21456 28008
rect 21508 27996 21514 28008
rect 27614 27996 27620 28008
rect 21508 27968 27620 27996
rect 21508 27956 21514 27968
rect 27614 27956 27620 27968
rect 27672 27956 27678 28008
rect 29362 27956 29368 28008
rect 29420 27996 29426 28008
rect 29917 27999 29975 28005
rect 29917 27996 29929 27999
rect 29420 27968 29929 27996
rect 29420 27956 29426 27968
rect 29917 27965 29929 27968
rect 29963 27965 29975 27999
rect 30024 27996 30052 28036
rect 31110 28024 31116 28036
rect 31168 28024 31174 28076
rect 31680 28073 31708 28104
rect 33045 28101 33057 28104
rect 33091 28101 33103 28135
rect 33045 28095 33103 28101
rect 31665 28067 31723 28073
rect 31665 28033 31677 28067
rect 31711 28033 31723 28067
rect 31665 28027 31723 28033
rect 31849 28067 31907 28073
rect 31849 28033 31861 28067
rect 31895 28064 31907 28067
rect 32309 28067 32367 28073
rect 32309 28064 32321 28067
rect 31895 28036 32321 28064
rect 31895 28033 31907 28036
rect 31849 28027 31907 28033
rect 32309 28033 32321 28036
rect 32355 28033 32367 28067
rect 32309 28027 32367 28033
rect 32398 28024 32404 28076
rect 32456 28064 32462 28076
rect 32493 28067 32551 28073
rect 32493 28064 32505 28067
rect 32456 28036 32505 28064
rect 32456 28024 32462 28036
rect 32493 28033 32505 28036
rect 32539 28033 32551 28067
rect 32493 28027 32551 28033
rect 32585 28067 32643 28073
rect 32585 28033 32597 28067
rect 32631 28064 32643 28067
rect 32766 28064 32772 28076
rect 32631 28036 32772 28064
rect 32631 28033 32643 28036
rect 32585 28027 32643 28033
rect 30024 27968 31754 27996
rect 29917 27959 29975 27965
rect 18544 27900 20484 27928
rect 22646 27888 22652 27940
rect 22704 27928 22710 27940
rect 26510 27928 26516 27940
rect 22704 27900 26516 27928
rect 22704 27888 22710 27900
rect 26510 27888 26516 27900
rect 26568 27888 26574 27940
rect 26602 27888 26608 27940
rect 26660 27928 26666 27940
rect 28626 27928 28632 27940
rect 26660 27900 28632 27928
rect 26660 27888 26666 27900
rect 28626 27888 28632 27900
rect 28684 27928 28690 27940
rect 29546 27928 29552 27940
rect 28684 27900 29552 27928
rect 28684 27888 28690 27900
rect 29546 27888 29552 27900
rect 29604 27888 29610 27940
rect 29822 27888 29828 27940
rect 29880 27928 29886 27940
rect 30834 27928 30840 27940
rect 29880 27900 30840 27928
rect 29880 27888 29886 27900
rect 5166 27820 5172 27872
rect 5224 27860 5230 27872
rect 11514 27860 11520 27872
rect 5224 27832 11520 27860
rect 5224 27820 5230 27832
rect 11514 27820 11520 27832
rect 11572 27820 11578 27872
rect 12894 27820 12900 27872
rect 12952 27820 12958 27872
rect 13814 27820 13820 27872
rect 13872 27860 13878 27872
rect 15746 27860 15752 27872
rect 13872 27832 15752 27860
rect 13872 27820 13878 27832
rect 15746 27820 15752 27832
rect 15804 27820 15810 27872
rect 15930 27820 15936 27872
rect 15988 27860 15994 27872
rect 16209 27863 16267 27869
rect 16209 27860 16221 27863
rect 15988 27832 16221 27860
rect 15988 27820 15994 27832
rect 16209 27829 16221 27832
rect 16255 27829 16267 27863
rect 16209 27823 16267 27829
rect 17770 27820 17776 27872
rect 17828 27820 17834 27872
rect 18230 27820 18236 27872
rect 18288 27860 18294 27872
rect 18509 27863 18567 27869
rect 18509 27860 18521 27863
rect 18288 27832 18521 27860
rect 18288 27820 18294 27832
rect 18509 27829 18521 27832
rect 18555 27829 18567 27863
rect 18509 27823 18567 27829
rect 19288 27820 19294 27872
rect 19346 27860 19352 27872
rect 19521 27863 19579 27869
rect 19521 27860 19533 27863
rect 19346 27832 19533 27860
rect 19346 27820 19352 27832
rect 19521 27829 19533 27832
rect 19567 27829 19579 27863
rect 19521 27823 19579 27829
rect 21634 27820 21640 27872
rect 21692 27860 21698 27872
rect 29270 27860 29276 27872
rect 21692 27832 29276 27860
rect 21692 27820 21698 27832
rect 29270 27820 29276 27832
rect 29328 27820 29334 27872
rect 29932 27869 29960 27900
rect 30834 27888 30840 27900
rect 30892 27888 30898 27940
rect 31726 27928 31754 27968
rect 31938 27956 31944 28008
rect 31996 27956 32002 28008
rect 32030 27956 32036 28008
rect 32088 27956 32094 28008
rect 32508 27996 32536 28027
rect 32766 28024 32772 28036
rect 32824 28024 32830 28076
rect 33229 28067 33287 28073
rect 33229 28064 33241 28067
rect 32876 28036 33241 28064
rect 32876 27996 32904 28036
rect 33229 28033 33241 28036
rect 33275 28033 33287 28067
rect 33229 28027 33287 28033
rect 33321 28067 33379 28073
rect 33321 28033 33333 28067
rect 33367 28064 33379 28067
rect 33870 28064 33876 28076
rect 33367 28036 33876 28064
rect 33367 28033 33379 28036
rect 33321 28027 33379 28033
rect 32508 27968 32904 27996
rect 32953 27999 33011 28005
rect 32953 27965 32965 27999
rect 32999 27965 33011 27999
rect 32953 27959 33011 27965
rect 32048 27928 32076 27956
rect 32968 27928 32996 27959
rect 31726 27900 31984 27928
rect 32048 27900 32996 27928
rect 29917 27863 29975 27869
rect 29917 27829 29929 27863
rect 29963 27829 29975 27863
rect 29917 27823 29975 27829
rect 30190 27820 30196 27872
rect 30248 27820 30254 27872
rect 30374 27820 30380 27872
rect 30432 27860 30438 27872
rect 31754 27860 31760 27872
rect 30432 27832 31760 27860
rect 30432 27820 30438 27832
rect 31754 27820 31760 27832
rect 31812 27820 31818 27872
rect 31956 27860 31984 27900
rect 33336 27860 33364 28027
rect 33870 28024 33876 28036
rect 33928 28024 33934 28076
rect 33962 28024 33968 28076
rect 34020 28024 34026 28076
rect 34256 28064 34284 28160
rect 34422 28092 34428 28144
rect 34480 28132 34486 28144
rect 37829 28135 37887 28141
rect 37829 28132 37841 28135
rect 34480 28104 37841 28132
rect 34480 28092 34486 28104
rect 37829 28101 37841 28104
rect 37875 28101 37887 28135
rect 37829 28095 37887 28101
rect 34072 28036 34284 28064
rect 33594 27956 33600 28008
rect 33652 27956 33658 28008
rect 33689 27999 33747 28005
rect 33689 27965 33701 27999
rect 33735 27996 33747 27999
rect 34072 27996 34100 28036
rect 35158 28024 35164 28076
rect 35216 28064 35222 28076
rect 35710 28064 35716 28076
rect 35216 28036 35716 28064
rect 35216 28024 35222 28036
rect 35710 28024 35716 28036
rect 35768 28064 35774 28076
rect 38565 28067 38623 28073
rect 35768 28036 37964 28064
rect 35768 28024 35774 28036
rect 33735 27968 34100 27996
rect 34241 27999 34299 28005
rect 33735 27965 33747 27968
rect 33689 27959 33747 27965
rect 34241 27965 34253 27999
rect 34287 27996 34299 27999
rect 35253 27999 35311 28005
rect 35253 27996 35265 27999
rect 34287 27968 35265 27996
rect 34287 27965 34299 27968
rect 34241 27959 34299 27965
rect 35253 27965 35265 27968
rect 35299 27965 35311 27999
rect 35253 27959 35311 27965
rect 35345 27999 35403 28005
rect 35345 27965 35357 27999
rect 35391 27996 35403 27999
rect 35434 27996 35440 28008
rect 35391 27968 35440 27996
rect 35391 27965 35403 27968
rect 35345 27959 35403 27965
rect 33612 27928 33640 27956
rect 34256 27928 34284 27959
rect 33612 27900 34284 27928
rect 35268 27928 35296 27959
rect 35434 27956 35440 27968
rect 35492 27956 35498 28008
rect 37936 28005 37964 28036
rect 38565 28033 38577 28067
rect 38611 28064 38623 28067
rect 39114 28064 39120 28076
rect 38611 28036 39120 28064
rect 38611 28033 38623 28036
rect 38565 28027 38623 28033
rect 39114 28024 39120 28036
rect 39172 28024 39178 28076
rect 37921 27999 37979 28005
rect 37921 27965 37933 27999
rect 37967 27965 37979 27999
rect 37921 27959 37979 27965
rect 36814 27928 36820 27940
rect 35268 27900 36820 27928
rect 36814 27888 36820 27900
rect 36872 27888 36878 27940
rect 31956 27832 33364 27860
rect 34330 27820 34336 27872
rect 34388 27820 34394 27872
rect 35526 27820 35532 27872
rect 35584 27820 35590 27872
rect 1104 27770 41400 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 41400 27770
rect 1104 27696 41400 27718
rect 5537 27659 5595 27665
rect 5537 27625 5549 27659
rect 5583 27656 5595 27659
rect 5626 27656 5632 27668
rect 5583 27628 5632 27656
rect 5583 27625 5595 27628
rect 5537 27619 5595 27625
rect 5626 27616 5632 27628
rect 5684 27616 5690 27668
rect 9030 27616 9036 27668
rect 9088 27656 9094 27668
rect 10226 27656 10232 27668
rect 9088 27628 10232 27656
rect 9088 27616 9094 27628
rect 10226 27616 10232 27628
rect 10284 27656 10290 27668
rect 11882 27656 11888 27668
rect 10284 27628 11888 27656
rect 10284 27616 10290 27628
rect 11882 27616 11888 27628
rect 11940 27616 11946 27668
rect 12250 27616 12256 27668
rect 12308 27616 12314 27668
rect 12526 27616 12532 27668
rect 12584 27616 12590 27668
rect 12897 27659 12955 27665
rect 12897 27625 12909 27659
rect 12943 27625 12955 27659
rect 12897 27619 12955 27625
rect 5644 27529 5672 27616
rect 6086 27548 6092 27600
rect 6144 27588 6150 27600
rect 6730 27588 6736 27600
rect 6144 27560 6736 27588
rect 6144 27548 6150 27560
rect 6730 27548 6736 27560
rect 6788 27548 6794 27600
rect 8938 27548 8944 27600
rect 8996 27588 9002 27600
rect 8996 27548 9030 27588
rect 9214 27548 9220 27600
rect 9272 27588 9278 27600
rect 12434 27588 12440 27600
rect 9272 27560 12440 27588
rect 9272 27548 9278 27560
rect 12434 27548 12440 27560
rect 12492 27548 12498 27600
rect 12544 27588 12572 27616
rect 12621 27591 12679 27597
rect 12621 27588 12633 27591
rect 12544 27560 12633 27588
rect 12621 27557 12633 27560
rect 12667 27557 12679 27591
rect 12912 27588 12940 27619
rect 13170 27616 13176 27668
rect 13228 27656 13234 27668
rect 13449 27659 13507 27665
rect 13449 27656 13461 27659
rect 13228 27628 13461 27656
rect 13228 27616 13234 27628
rect 13449 27625 13461 27628
rect 13495 27656 13507 27659
rect 14093 27659 14151 27665
rect 13495 27628 14044 27656
rect 13495 27625 13507 27628
rect 13449 27619 13507 27625
rect 13262 27588 13268 27600
rect 12912 27560 13268 27588
rect 12621 27551 12679 27557
rect 13262 27548 13268 27560
rect 13320 27548 13326 27600
rect 14016 27588 14044 27628
rect 14093 27625 14105 27659
rect 14139 27656 14151 27659
rect 14918 27656 14924 27668
rect 14139 27628 14924 27656
rect 14139 27625 14151 27628
rect 14093 27619 14151 27625
rect 14918 27616 14924 27628
rect 14976 27616 14982 27668
rect 15102 27616 15108 27668
rect 15160 27656 15166 27668
rect 17126 27656 17132 27668
rect 15160 27628 15700 27656
rect 15160 27616 15166 27628
rect 14642 27588 14648 27600
rect 14016 27560 14648 27588
rect 14642 27548 14648 27560
rect 14700 27548 14706 27600
rect 15013 27591 15071 27597
rect 15013 27557 15025 27591
rect 15059 27588 15071 27591
rect 15378 27588 15384 27600
rect 15059 27560 15384 27588
rect 15059 27557 15071 27560
rect 15013 27551 15071 27557
rect 15378 27548 15384 27560
rect 15436 27548 15442 27600
rect 5629 27523 5687 27529
rect 5629 27489 5641 27523
rect 5675 27489 5687 27523
rect 5629 27483 5687 27489
rect 6178 27480 6184 27532
rect 6236 27520 6242 27532
rect 8478 27520 8484 27532
rect 6236 27492 8484 27520
rect 6236 27480 6242 27492
rect 3786 27412 3792 27464
rect 3844 27412 3850 27464
rect 5442 27452 5448 27464
rect 5198 27424 5448 27452
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 6270 27412 6276 27464
rect 6328 27412 6334 27464
rect 6380 27461 6408 27492
rect 8478 27480 8484 27492
rect 8536 27480 8542 27532
rect 9002 27520 9030 27548
rect 9398 27520 9404 27532
rect 9002 27492 9404 27520
rect 6365 27455 6423 27461
rect 6365 27421 6377 27455
rect 6411 27421 6423 27455
rect 6365 27415 6423 27421
rect 6454 27412 6460 27464
rect 6512 27452 6518 27464
rect 6549 27455 6607 27461
rect 6549 27452 6561 27455
rect 6512 27424 6561 27452
rect 6512 27412 6518 27424
rect 6549 27421 6561 27424
rect 6595 27421 6607 27455
rect 6549 27415 6607 27421
rect 6730 27412 6736 27464
rect 6788 27412 6794 27464
rect 8846 27412 8852 27464
rect 8904 27452 8910 27464
rect 9232 27461 9260 27492
rect 9398 27480 9404 27492
rect 9456 27480 9462 27532
rect 9490 27480 9496 27532
rect 9548 27520 9554 27532
rect 9548 27492 9905 27520
rect 9548 27480 9554 27492
rect 8941 27455 8999 27461
rect 8941 27452 8953 27455
rect 8904 27424 8953 27452
rect 8904 27412 8910 27424
rect 8941 27421 8953 27424
rect 8987 27421 8999 27455
rect 8941 27415 8999 27421
rect 9217 27455 9275 27461
rect 9217 27421 9229 27455
rect 9263 27421 9275 27455
rect 9217 27415 9275 27421
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27446 9367 27455
rect 9508 27446 9536 27480
rect 9355 27421 9536 27446
rect 9309 27418 9536 27421
rect 9309 27415 9367 27418
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 9766 27452 9772 27464
rect 9640 27424 9772 27452
rect 9640 27412 9646 27424
rect 9766 27412 9772 27424
rect 9824 27412 9830 27464
rect 4062 27344 4068 27396
rect 4120 27344 4126 27396
rect 6288 27384 6316 27412
rect 6641 27387 6699 27393
rect 6641 27384 6653 27387
rect 6288 27356 6653 27384
rect 6641 27353 6653 27356
rect 6687 27384 6699 27387
rect 6822 27384 6828 27396
rect 6687 27356 6828 27384
rect 6687 27353 6699 27356
rect 6641 27347 6699 27353
rect 6822 27344 6828 27356
rect 6880 27344 6886 27396
rect 9125 27387 9183 27393
rect 9125 27353 9137 27387
rect 9171 27384 9183 27387
rect 9877 27384 9905 27492
rect 12268 27492 13860 27520
rect 10042 27412 10048 27464
rect 10100 27452 10106 27464
rect 12268 27461 12296 27492
rect 12253 27455 12311 27461
rect 10100 27424 12112 27452
rect 10100 27412 10106 27424
rect 10778 27384 10784 27396
rect 9171 27356 9674 27384
rect 9877 27356 10784 27384
rect 9171 27353 9183 27356
rect 9125 27347 9183 27353
rect 6270 27276 6276 27328
rect 6328 27276 6334 27328
rect 6914 27276 6920 27328
rect 6972 27276 6978 27328
rect 9490 27276 9496 27328
rect 9548 27276 9554 27328
rect 9646 27316 9674 27356
rect 10778 27344 10784 27356
rect 10836 27344 10842 27396
rect 10594 27316 10600 27328
rect 9646 27288 10600 27316
rect 10594 27276 10600 27288
rect 10652 27276 10658 27328
rect 12084 27316 12112 27424
rect 12253 27421 12265 27455
rect 12299 27421 12311 27455
rect 12253 27415 12311 27421
rect 12345 27455 12403 27461
rect 12345 27421 12357 27455
rect 12391 27421 12403 27455
rect 12345 27415 12403 27421
rect 12820 27424 13492 27452
rect 12158 27344 12164 27396
rect 12216 27384 12222 27396
rect 12360 27384 12388 27415
rect 12216 27356 12388 27384
rect 12216 27344 12222 27356
rect 12526 27344 12532 27396
rect 12584 27384 12590 27396
rect 12722 27387 12780 27393
rect 12722 27384 12734 27387
rect 12584 27356 12734 27384
rect 12584 27344 12590 27356
rect 12722 27353 12734 27356
rect 12768 27353 12780 27387
rect 12722 27347 12780 27353
rect 12820 27316 12848 27424
rect 13464 27396 13492 27424
rect 12897 27387 12955 27393
rect 12897 27353 12909 27387
rect 12943 27384 12955 27387
rect 13170 27384 13176 27396
rect 12943 27356 13176 27384
rect 12943 27353 12955 27356
rect 12897 27347 12955 27353
rect 13170 27344 13176 27356
rect 13228 27344 13234 27396
rect 13262 27344 13268 27396
rect 13320 27344 13326 27396
rect 13446 27344 13452 27396
rect 13504 27344 13510 27396
rect 13722 27384 13728 27396
rect 13556 27356 13728 27384
rect 12084 27288 12848 27316
rect 13081 27319 13139 27325
rect 13081 27285 13093 27319
rect 13127 27316 13139 27319
rect 13556 27316 13584 27356
rect 13722 27344 13728 27356
rect 13780 27344 13786 27396
rect 13127 27288 13584 27316
rect 13633 27319 13691 27325
rect 13127 27285 13139 27288
rect 13081 27279 13139 27285
rect 13633 27285 13645 27319
rect 13679 27316 13691 27319
rect 13832 27316 13860 27492
rect 14090 27480 14096 27532
rect 14148 27520 14154 27532
rect 14369 27523 14427 27529
rect 14369 27520 14381 27523
rect 14148 27492 14381 27520
rect 14148 27480 14154 27492
rect 14369 27489 14381 27492
rect 14415 27520 14427 27523
rect 15672 27520 15700 27628
rect 15764 27628 17132 27656
rect 15764 27600 15792 27628
rect 17126 27616 17132 27628
rect 17184 27616 17190 27668
rect 17586 27616 17592 27668
rect 17644 27656 17650 27668
rect 18506 27656 18512 27668
rect 17644 27628 18512 27656
rect 17644 27616 17650 27628
rect 18506 27616 18512 27628
rect 18564 27616 18570 27668
rect 18966 27616 18972 27668
rect 19024 27656 19030 27668
rect 19061 27659 19119 27665
rect 19061 27656 19073 27659
rect 19024 27628 19073 27656
rect 19024 27616 19030 27628
rect 19061 27625 19073 27628
rect 19107 27625 19119 27659
rect 19061 27619 19119 27625
rect 20901 27659 20959 27665
rect 20901 27625 20913 27659
rect 20947 27625 20959 27659
rect 22833 27659 22891 27665
rect 22833 27656 22845 27659
rect 20901 27619 20959 27625
rect 21284 27628 22845 27656
rect 15746 27548 15752 27600
rect 15804 27548 15810 27600
rect 14415 27492 15608 27520
rect 15672 27492 16620 27520
rect 14415 27489 14427 27492
rect 14369 27483 14427 27489
rect 14277 27455 14335 27461
rect 14277 27421 14289 27455
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14292 27384 14320 27415
rect 14458 27412 14464 27464
rect 14516 27412 14522 27464
rect 14550 27412 14556 27464
rect 14608 27452 14614 27464
rect 14826 27452 14832 27464
rect 14608 27424 14832 27452
rect 14608 27412 14614 27424
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 15194 27412 15200 27464
rect 15252 27412 15258 27464
rect 15580 27461 15608 27492
rect 15289 27455 15347 27461
rect 15289 27421 15301 27455
rect 15335 27452 15347 27455
rect 15565 27455 15623 27461
rect 15335 27424 15516 27452
rect 15335 27421 15347 27424
rect 15289 27415 15347 27421
rect 15381 27387 15439 27393
rect 14292 27356 14596 27384
rect 14568 27328 14596 27356
rect 15381 27353 15393 27387
rect 15427 27353 15439 27387
rect 15488 27384 15516 27424
rect 15565 27421 15577 27455
rect 15611 27421 15623 27455
rect 15565 27415 15623 27421
rect 15657 27455 15715 27461
rect 15657 27421 15669 27455
rect 15703 27452 15715 27455
rect 16117 27455 16175 27461
rect 15703 27424 16068 27452
rect 15703 27421 15715 27424
rect 15657 27415 15715 27421
rect 16040 27396 16068 27424
rect 16117 27421 16129 27455
rect 16163 27452 16175 27455
rect 16592 27452 16620 27492
rect 16666 27480 16672 27532
rect 16724 27520 16730 27532
rect 17144 27529 17172 27616
rect 20622 27548 20628 27600
rect 20680 27588 20686 27600
rect 20916 27588 20944 27619
rect 20680 27560 20944 27588
rect 20680 27548 20686 27560
rect 17132 27523 17190 27529
rect 16724 27492 17080 27520
rect 16724 27480 16730 27492
rect 16853 27455 16911 27461
rect 16853 27452 16865 27455
rect 16163 27424 16528 27452
rect 16592 27424 16865 27452
rect 16163 27421 16175 27424
rect 16117 27415 16175 27421
rect 15488 27356 15884 27384
rect 15381 27347 15439 27353
rect 13906 27316 13912 27328
rect 13679 27288 13912 27316
rect 13679 27285 13691 27288
rect 13633 27279 13691 27285
rect 13906 27276 13912 27288
rect 13964 27276 13970 27328
rect 14550 27276 14556 27328
rect 14608 27276 14614 27328
rect 15396 27316 15424 27347
rect 15856 27328 15884 27356
rect 16022 27344 16028 27396
rect 16080 27344 16086 27396
rect 16500 27328 16528 27424
rect 16853 27421 16865 27424
rect 16899 27421 16911 27455
rect 16853 27415 16911 27421
rect 16942 27412 16948 27464
rect 17000 27412 17006 27464
rect 17052 27452 17080 27492
rect 17132 27489 17144 27523
rect 17178 27489 17190 27523
rect 17132 27483 17190 27489
rect 17972 27492 18828 27520
rect 17972 27464 18000 27492
rect 17221 27455 17279 27461
rect 17221 27452 17233 27455
rect 17052 27424 17233 27452
rect 17221 27421 17233 27424
rect 17267 27421 17279 27455
rect 17221 27415 17279 27421
rect 17310 27412 17316 27464
rect 17368 27452 17374 27464
rect 17405 27455 17463 27461
rect 17405 27452 17417 27455
rect 17368 27424 17417 27452
rect 17368 27412 17374 27424
rect 17405 27421 17417 27424
rect 17451 27421 17463 27455
rect 17405 27415 17463 27421
rect 17954 27412 17960 27464
rect 18012 27412 18018 27464
rect 18506 27412 18512 27464
rect 18564 27412 18570 27464
rect 18800 27461 18828 27492
rect 20806 27480 20812 27532
rect 20864 27520 20870 27532
rect 20990 27520 20996 27532
rect 20864 27492 20996 27520
rect 20864 27480 20870 27492
rect 20990 27480 20996 27492
rect 21048 27480 21054 27532
rect 21284 27520 21312 27628
rect 22833 27625 22845 27628
rect 22879 27625 22891 27659
rect 22833 27619 22891 27625
rect 23109 27659 23167 27665
rect 23109 27625 23121 27659
rect 23155 27656 23167 27659
rect 23198 27656 23204 27668
rect 23155 27628 23204 27656
rect 23155 27625 23167 27628
rect 23109 27619 23167 27625
rect 23198 27616 23204 27628
rect 23256 27616 23262 27668
rect 25406 27656 25412 27668
rect 23676 27628 25412 27656
rect 21358 27548 21364 27600
rect 21416 27588 21422 27600
rect 22097 27591 22155 27597
rect 21416 27560 21496 27588
rect 21416 27548 21422 27560
rect 21284 27492 21404 27520
rect 21376 27464 21404 27492
rect 18693 27455 18751 27461
rect 18693 27421 18705 27455
rect 18739 27421 18751 27455
rect 18693 27415 18751 27421
rect 18785 27455 18843 27461
rect 18785 27421 18797 27455
rect 18831 27421 18843 27455
rect 18785 27415 18843 27421
rect 18877 27455 18935 27461
rect 18877 27421 18889 27455
rect 18923 27454 18935 27455
rect 18923 27452 19196 27454
rect 21082 27452 21088 27464
rect 18923 27426 21088 27452
rect 18923 27421 18935 27426
rect 19168 27424 21088 27426
rect 18877 27415 18935 27421
rect 16758 27344 16764 27396
rect 16816 27384 16822 27396
rect 18230 27384 18236 27396
rect 16816 27356 18236 27384
rect 16816 27344 16822 27356
rect 18230 27344 18236 27356
rect 18288 27344 18294 27396
rect 18708 27384 18736 27415
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 21177 27455 21235 27461
rect 21177 27421 21189 27455
rect 21223 27452 21235 27455
rect 21266 27452 21272 27464
rect 21223 27424 21272 27452
rect 21223 27421 21235 27424
rect 21177 27415 21235 27421
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 21358 27412 21364 27464
rect 21416 27412 21422 27464
rect 21468 27461 21496 27560
rect 22097 27557 22109 27591
rect 22143 27588 22155 27591
rect 22922 27588 22928 27600
rect 22143 27560 22928 27588
rect 22143 27557 22155 27560
rect 22097 27551 22155 27557
rect 22922 27548 22928 27560
rect 22980 27548 22986 27600
rect 23293 27591 23351 27597
rect 23293 27557 23305 27591
rect 23339 27557 23351 27591
rect 23293 27551 23351 27557
rect 23308 27464 23336 27551
rect 23676 27520 23704 27628
rect 25406 27616 25412 27628
rect 25464 27656 25470 27668
rect 25464 27628 27850 27656
rect 25464 27616 25470 27628
rect 23750 27548 23756 27600
rect 23808 27588 23814 27600
rect 27706 27588 27712 27600
rect 23808 27560 27712 27588
rect 23808 27548 23814 27560
rect 23676 27492 23888 27520
rect 21453 27455 21511 27461
rect 21453 27421 21465 27455
rect 21499 27421 21511 27455
rect 21453 27415 21511 27421
rect 22020 27424 22508 27452
rect 18966 27384 18972 27396
rect 18708 27356 18972 27384
rect 18966 27344 18972 27356
rect 19024 27384 19030 27396
rect 19426 27384 19432 27396
rect 19024 27356 19432 27384
rect 19024 27344 19030 27356
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 20622 27344 20628 27396
rect 20680 27384 20686 27396
rect 22020 27384 22048 27424
rect 20680 27356 22048 27384
rect 22097 27387 22155 27393
rect 20680 27344 20686 27356
rect 22097 27353 22109 27387
rect 22143 27384 22155 27387
rect 22370 27384 22376 27396
rect 22143 27356 22376 27384
rect 22143 27353 22155 27356
rect 22097 27347 22155 27353
rect 22370 27344 22376 27356
rect 22428 27344 22434 27396
rect 22480 27384 22508 27424
rect 22554 27412 22560 27464
rect 22612 27452 22618 27464
rect 22612 27424 22968 27452
rect 22612 27412 22618 27424
rect 22940 27393 22968 27424
rect 23290 27412 23296 27464
rect 23348 27412 23354 27464
rect 23566 27412 23572 27464
rect 23624 27452 23630 27464
rect 23860 27461 23888 27492
rect 24228 27461 24256 27560
rect 27706 27548 27712 27560
rect 27764 27548 27770 27600
rect 27822 27588 27850 27628
rect 27890 27616 27896 27668
rect 27948 27656 27954 27668
rect 28445 27659 28503 27665
rect 28445 27656 28457 27659
rect 27948 27628 28457 27656
rect 27948 27616 27954 27628
rect 28445 27625 28457 27628
rect 28491 27625 28503 27659
rect 28445 27619 28503 27625
rect 28994 27616 29000 27668
rect 29052 27656 29058 27668
rect 30285 27659 30343 27665
rect 29052 27628 30236 27656
rect 29052 27616 29058 27628
rect 27982 27588 27988 27600
rect 27822 27560 27988 27588
rect 27982 27548 27988 27560
rect 28040 27548 28046 27600
rect 28629 27591 28687 27597
rect 28629 27557 28641 27591
rect 28675 27588 28687 27591
rect 29089 27591 29147 27597
rect 29089 27588 29101 27591
rect 28675 27560 29101 27588
rect 28675 27557 28687 27560
rect 28629 27551 28687 27557
rect 29089 27557 29101 27560
rect 29135 27557 29147 27591
rect 29089 27551 29147 27557
rect 24688 27492 26740 27520
rect 24688 27464 24716 27492
rect 23661 27455 23719 27461
rect 23661 27452 23673 27455
rect 23624 27424 23673 27452
rect 23624 27412 23630 27424
rect 23661 27421 23673 27424
rect 23707 27421 23719 27455
rect 23661 27415 23719 27421
rect 23845 27455 23903 27461
rect 23845 27421 23857 27455
rect 23891 27421 23903 27455
rect 23845 27415 23903 27421
rect 24213 27455 24271 27461
rect 24213 27421 24225 27455
rect 24259 27421 24271 27455
rect 24213 27415 24271 27421
rect 24670 27412 24676 27464
rect 24728 27412 24734 27464
rect 25041 27455 25099 27461
rect 25041 27421 25053 27455
rect 25087 27421 25099 27455
rect 25041 27415 25099 27421
rect 25225 27455 25283 27461
rect 25225 27421 25237 27455
rect 25271 27452 25283 27455
rect 25406 27452 25412 27464
rect 25271 27424 25412 27452
rect 25271 27421 25283 27424
rect 25225 27415 25283 27421
rect 22925 27387 22983 27393
rect 22480 27356 22784 27384
rect 15746 27316 15752 27328
rect 15396 27288 15752 27316
rect 15746 27276 15752 27288
rect 15804 27276 15810 27328
rect 15838 27276 15844 27328
rect 15896 27276 15902 27328
rect 16298 27276 16304 27328
rect 16356 27276 16362 27328
rect 16482 27276 16488 27328
rect 16540 27276 16546 27328
rect 17126 27276 17132 27328
rect 17184 27276 17190 27328
rect 17405 27319 17463 27325
rect 17405 27285 17417 27319
rect 17451 27316 17463 27319
rect 18138 27316 18144 27328
rect 17451 27288 18144 27316
rect 17451 27285 17463 27288
rect 17405 27279 17463 27285
rect 18138 27276 18144 27288
rect 18196 27276 18202 27328
rect 18248 27316 18276 27344
rect 22278 27316 22284 27328
rect 18248 27288 22284 27316
rect 22278 27276 22284 27288
rect 22336 27276 22342 27328
rect 22646 27276 22652 27328
rect 22704 27276 22710 27328
rect 22756 27316 22784 27356
rect 22925 27353 22937 27387
rect 22971 27353 22983 27387
rect 22925 27347 22983 27353
rect 23382 27344 23388 27396
rect 23440 27384 23446 27396
rect 25056 27384 25084 27415
rect 25406 27412 25412 27424
rect 25464 27412 25470 27464
rect 25498 27412 25504 27464
rect 25556 27412 25562 27464
rect 25608 27461 25636 27492
rect 25593 27455 25651 27461
rect 25593 27421 25605 27455
rect 25639 27421 25651 27455
rect 25593 27415 25651 27421
rect 25958 27412 25964 27464
rect 26016 27412 26022 27464
rect 26418 27412 26424 27464
rect 26476 27452 26482 27464
rect 26513 27455 26571 27461
rect 26513 27452 26525 27455
rect 26476 27424 26525 27452
rect 26476 27412 26482 27424
rect 26513 27421 26525 27424
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 26602 27412 26608 27464
rect 26660 27412 26666 27464
rect 26712 27461 26740 27492
rect 26878 27480 26884 27532
rect 26936 27520 26942 27532
rect 27065 27523 27123 27529
rect 27065 27520 27077 27523
rect 26936 27492 27077 27520
rect 26936 27480 26942 27492
rect 27065 27489 27077 27492
rect 27111 27489 27123 27523
rect 27065 27483 27123 27489
rect 27249 27523 27307 27529
rect 27249 27489 27261 27523
rect 27295 27520 27307 27523
rect 28721 27523 28779 27529
rect 28721 27520 28733 27523
rect 27295 27492 28733 27520
rect 27295 27489 27307 27492
rect 27249 27483 27307 27489
rect 28721 27489 28733 27492
rect 28767 27489 28779 27523
rect 28721 27483 28779 27489
rect 29270 27480 29276 27532
rect 29328 27520 29334 27532
rect 29546 27520 29552 27532
rect 29328 27492 29552 27520
rect 29328 27480 29334 27492
rect 29546 27480 29552 27492
rect 29604 27520 29610 27532
rect 30208 27529 30236 27628
rect 30285 27625 30297 27659
rect 30331 27656 30343 27659
rect 30374 27656 30380 27668
rect 30331 27628 30380 27656
rect 30331 27625 30343 27628
rect 30285 27619 30343 27625
rect 30374 27616 30380 27628
rect 30432 27616 30438 27668
rect 30834 27616 30840 27668
rect 30892 27616 30898 27668
rect 31110 27616 31116 27668
rect 31168 27656 31174 27668
rect 32674 27656 32680 27668
rect 31168 27628 32680 27656
rect 31168 27616 31174 27628
rect 32674 27616 32680 27628
rect 32732 27616 32738 27668
rect 35056 27659 35114 27665
rect 35056 27625 35068 27659
rect 35102 27656 35114 27659
rect 35526 27656 35532 27668
rect 35102 27628 35532 27656
rect 35102 27625 35114 27628
rect 35056 27619 35114 27625
rect 35526 27616 35532 27628
rect 35584 27616 35590 27668
rect 30852 27588 30880 27616
rect 30852 27560 31432 27588
rect 30193 27523 30251 27529
rect 29604 27492 30052 27520
rect 29604 27480 29610 27492
rect 26697 27455 26755 27461
rect 26697 27421 26709 27455
rect 26743 27452 26755 27455
rect 26789 27455 26847 27461
rect 26789 27452 26801 27455
rect 26743 27424 26801 27452
rect 26743 27421 26755 27424
rect 26697 27415 26755 27421
rect 26789 27421 26801 27424
rect 26835 27421 26847 27455
rect 26789 27415 26847 27421
rect 26973 27455 27031 27461
rect 26973 27421 26985 27455
rect 27019 27452 27031 27455
rect 27338 27452 27344 27464
rect 27019 27424 27344 27452
rect 27019 27421 27031 27424
rect 26973 27415 27031 27421
rect 27338 27412 27344 27424
rect 27396 27412 27402 27464
rect 27522 27412 27528 27464
rect 27580 27412 27586 27464
rect 28534 27452 28540 27464
rect 27632 27424 28540 27452
rect 27632 27384 27660 27424
rect 28534 27412 28540 27424
rect 28592 27412 28598 27464
rect 28810 27412 28816 27464
rect 28868 27452 28874 27464
rect 28905 27455 28963 27461
rect 28905 27452 28917 27455
rect 28868 27424 28917 27452
rect 28868 27412 28874 27424
rect 28905 27421 28917 27424
rect 28951 27421 28963 27455
rect 28905 27415 28963 27421
rect 28994 27412 29000 27464
rect 29052 27412 29058 27464
rect 29181 27455 29239 27461
rect 29181 27421 29193 27455
rect 29227 27421 29239 27455
rect 29181 27415 29239 27421
rect 29365 27455 29423 27461
rect 29365 27421 29377 27455
rect 29411 27452 29423 27455
rect 29638 27452 29644 27464
rect 29411 27424 29644 27452
rect 29411 27421 29423 27424
rect 29365 27415 29423 27421
rect 23440 27356 24348 27384
rect 25056 27356 27660 27384
rect 23440 27344 23446 27356
rect 23125 27319 23183 27325
rect 23125 27316 23137 27319
rect 22756 27288 23137 27316
rect 23125 27285 23137 27288
rect 23171 27316 23183 27319
rect 24026 27316 24032 27328
rect 23171 27288 24032 27316
rect 23171 27285 23183 27288
rect 23125 27279 23183 27285
rect 24026 27276 24032 27288
rect 24084 27276 24090 27328
rect 24121 27319 24179 27325
rect 24121 27285 24133 27319
rect 24167 27316 24179 27319
rect 24210 27316 24216 27328
rect 24167 27288 24216 27316
rect 24167 27285 24179 27288
rect 24121 27279 24179 27285
rect 24210 27276 24216 27288
rect 24268 27276 24274 27328
rect 24320 27316 24348 27356
rect 27890 27344 27896 27396
rect 27948 27384 27954 27396
rect 28261 27387 28319 27393
rect 28261 27384 28273 27387
rect 27948 27356 28273 27384
rect 27948 27344 27954 27356
rect 28261 27353 28273 27356
rect 28307 27384 28319 27387
rect 28350 27384 28356 27396
rect 28307 27356 28356 27384
rect 28307 27353 28319 27356
rect 28261 27347 28319 27353
rect 28350 27344 28356 27356
rect 28408 27344 28414 27396
rect 29196 27384 29224 27415
rect 29638 27412 29644 27424
rect 29696 27412 29702 27464
rect 30024 27452 30052 27492
rect 30193 27489 30205 27523
rect 30239 27520 30251 27523
rect 30929 27523 30987 27529
rect 30929 27520 30941 27523
rect 30239 27492 30941 27520
rect 30239 27489 30251 27492
rect 30193 27483 30251 27489
rect 30929 27489 30941 27492
rect 30975 27489 30987 27523
rect 30929 27483 30987 27489
rect 31404 27461 31432 27560
rect 31665 27523 31723 27529
rect 31665 27489 31677 27523
rect 31711 27520 31723 27523
rect 31754 27520 31760 27532
rect 31711 27492 31760 27520
rect 31711 27489 31723 27492
rect 31665 27483 31723 27489
rect 31754 27480 31760 27492
rect 31812 27520 31818 27532
rect 32398 27520 32404 27532
rect 31812 27492 32404 27520
rect 31812 27480 31818 27492
rect 32398 27480 32404 27492
rect 32456 27480 32462 27532
rect 34790 27480 34796 27532
rect 34848 27520 34854 27532
rect 35802 27520 35808 27532
rect 34848 27492 35808 27520
rect 34848 27480 34854 27492
rect 35802 27480 35808 27492
rect 35860 27480 35866 27532
rect 36814 27480 36820 27532
rect 36872 27480 36878 27532
rect 30377 27455 30435 27461
rect 30377 27452 30389 27455
rect 30024 27424 30389 27452
rect 30377 27421 30389 27424
rect 30423 27452 30435 27455
rect 31113 27455 31171 27461
rect 31113 27452 31125 27455
rect 30423 27424 31125 27452
rect 30423 27421 30435 27424
rect 30377 27415 30435 27421
rect 31113 27421 31125 27424
rect 31159 27421 31171 27455
rect 31113 27415 31171 27421
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27421 31447 27455
rect 31389 27415 31447 27421
rect 33505 27455 33563 27461
rect 33505 27421 33517 27455
rect 33551 27452 33563 27455
rect 34330 27452 34336 27464
rect 33551 27424 34336 27452
rect 33551 27421 33563 27424
rect 33505 27415 33563 27421
rect 34330 27412 34336 27424
rect 34388 27412 34394 27464
rect 29917 27387 29975 27393
rect 29917 27384 29929 27387
rect 29196 27356 29408 27384
rect 29380 27328 29408 27356
rect 29564 27356 29929 27384
rect 29564 27328 29592 27356
rect 29917 27353 29929 27356
rect 29963 27353 29975 27387
rect 29917 27347 29975 27353
rect 30098 27344 30104 27396
rect 30156 27384 30162 27396
rect 30653 27387 30711 27393
rect 30653 27384 30665 27387
rect 30156 27356 30665 27384
rect 30156 27344 30162 27356
rect 30653 27353 30665 27356
rect 30699 27353 30711 27387
rect 30653 27347 30711 27353
rect 35452 27356 35558 27384
rect 35452 27328 35480 27356
rect 25774 27316 25780 27328
rect 24320 27288 25780 27316
rect 25774 27276 25780 27288
rect 25832 27316 25838 27328
rect 25961 27319 26019 27325
rect 25961 27316 25973 27319
rect 25832 27288 25973 27316
rect 25832 27276 25838 27288
rect 25961 27285 25973 27288
rect 26007 27285 26019 27319
rect 25961 27279 26019 27285
rect 26142 27276 26148 27328
rect 26200 27316 26206 27328
rect 28461 27319 28519 27325
rect 28461 27316 28473 27319
rect 26200 27288 28473 27316
rect 26200 27276 26206 27288
rect 28461 27285 28473 27288
rect 28507 27316 28519 27319
rect 28718 27316 28724 27328
rect 28507 27288 28724 27316
rect 28507 27285 28519 27288
rect 28461 27279 28519 27285
rect 28718 27276 28724 27288
rect 28776 27276 28782 27328
rect 29362 27276 29368 27328
rect 29420 27276 29426 27328
rect 29546 27276 29552 27328
rect 29604 27276 29610 27328
rect 30558 27276 30564 27328
rect 30616 27276 30622 27328
rect 31294 27276 31300 27328
rect 31352 27276 31358 27328
rect 33502 27276 33508 27328
rect 33560 27316 33566 27328
rect 34057 27319 34115 27325
rect 34057 27316 34069 27319
rect 33560 27288 34069 27316
rect 33560 27276 33566 27288
rect 34057 27285 34069 27288
rect 34103 27285 34115 27319
rect 34057 27279 34115 27285
rect 35434 27276 35440 27328
rect 35492 27316 35498 27328
rect 38102 27316 38108 27328
rect 35492 27288 38108 27316
rect 35492 27276 35498 27288
rect 38102 27276 38108 27288
rect 38160 27276 38166 27328
rect 1104 27226 41400 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 41400 27226
rect 1104 27152 41400 27174
rect 3973 27115 4031 27121
rect 3973 27081 3985 27115
rect 4019 27112 4031 27115
rect 4062 27112 4068 27124
rect 4019 27084 4068 27112
rect 4019 27081 4031 27084
rect 3973 27075 4031 27081
rect 4062 27072 4068 27084
rect 4120 27072 4126 27124
rect 4893 27115 4951 27121
rect 4893 27081 4905 27115
rect 4939 27112 4951 27115
rect 6270 27112 6276 27124
rect 4939 27084 6276 27112
rect 4939 27081 4951 27084
rect 4893 27075 4951 27081
rect 6270 27072 6276 27084
rect 6328 27072 6334 27124
rect 6914 27112 6920 27124
rect 6656 27084 6920 27112
rect 6656 27053 6684 27084
rect 6914 27072 6920 27084
rect 6972 27072 6978 27124
rect 11606 27112 11612 27124
rect 8404 27084 11612 27112
rect 6641 27047 6699 27053
rect 6641 27013 6653 27047
rect 6687 27013 6699 27047
rect 6641 27007 6699 27013
rect 7282 27004 7288 27056
rect 7340 27004 7346 27056
rect 8202 27004 8208 27056
rect 8260 27044 8266 27056
rect 8404 27053 8432 27084
rect 11606 27072 11612 27084
rect 11664 27072 11670 27124
rect 11698 27072 11704 27124
rect 11756 27072 11762 27124
rect 11882 27072 11888 27124
rect 11940 27112 11946 27124
rect 11940 27084 12296 27112
rect 11940 27072 11946 27084
rect 8389 27047 8447 27053
rect 8389 27044 8401 27047
rect 8260 27016 8401 27044
rect 8260 27004 8266 27016
rect 8389 27013 8401 27016
rect 8435 27013 8447 27047
rect 8846 27044 8852 27056
rect 8389 27007 8447 27013
rect 8588 27016 8852 27044
rect 4157 26979 4215 26985
rect 4157 26945 4169 26979
rect 4203 26976 4215 26979
rect 4203 26948 4568 26976
rect 4203 26945 4215 26948
rect 4157 26939 4215 26945
rect 4540 26849 4568 26948
rect 5534 26936 5540 26988
rect 5592 26976 5598 26988
rect 8588 26985 8616 27016
rect 8846 27004 8852 27016
rect 8904 27004 8910 27056
rect 9398 27044 9404 27056
rect 8956 27016 9404 27044
rect 6365 26979 6423 26985
rect 6365 26976 6377 26979
rect 5592 26948 6377 26976
rect 5592 26936 5598 26948
rect 6365 26945 6377 26948
rect 6411 26945 6423 26979
rect 6365 26939 6423 26945
rect 8573 26979 8631 26985
rect 8573 26945 8585 26979
rect 8619 26945 8631 26979
rect 8573 26939 8631 26945
rect 8757 26979 8815 26985
rect 8757 26945 8769 26979
rect 8803 26976 8815 26979
rect 8956 26976 8984 27016
rect 9398 27004 9404 27016
rect 9456 27004 9462 27056
rect 9490 27004 9496 27056
rect 9548 27004 9554 27056
rect 10134 27044 10140 27056
rect 9692 27016 10140 27044
rect 8803 26948 8984 26976
rect 8803 26945 8815 26948
rect 8757 26939 8815 26945
rect 9030 26936 9036 26988
rect 9088 26936 9094 26988
rect 9309 26979 9367 26985
rect 9309 26945 9321 26979
rect 9355 26976 9367 26979
rect 9508 26976 9536 27004
rect 9692 26985 9720 27016
rect 10134 27004 10140 27016
rect 10192 27044 10198 27056
rect 10870 27044 10876 27056
rect 10192 27016 10876 27044
rect 10192 27004 10198 27016
rect 10870 27004 10876 27016
rect 10928 27004 10934 27056
rect 11716 27044 11744 27072
rect 11716 27016 12204 27044
rect 9355 26948 9536 26976
rect 9677 26979 9735 26985
rect 9355 26945 9367 26948
rect 9309 26939 9367 26945
rect 9677 26945 9689 26979
rect 9723 26945 9735 26979
rect 9677 26939 9735 26945
rect 9766 26936 9772 26988
rect 9824 26936 9830 26988
rect 9858 26936 9864 26988
rect 9916 26976 9922 26988
rect 9953 26979 10011 26985
rect 9953 26976 9965 26979
rect 9916 26948 9965 26976
rect 9916 26936 9922 26948
rect 9953 26945 9965 26948
rect 9999 26945 10011 26979
rect 9953 26939 10011 26945
rect 10045 26979 10103 26985
rect 10045 26945 10057 26979
rect 10091 26976 10103 26979
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 10091 26948 10272 26976
rect 10091 26945 10103 26948
rect 10045 26939 10103 26945
rect 10244 26920 10272 26948
rect 10704 26948 11713 26976
rect 4982 26868 4988 26920
rect 5040 26868 5046 26920
rect 5166 26868 5172 26920
rect 5224 26868 5230 26920
rect 9125 26911 9183 26917
rect 9125 26877 9137 26911
rect 9171 26877 9183 26911
rect 9125 26871 9183 26877
rect 9217 26911 9275 26917
rect 9217 26877 9229 26911
rect 9263 26908 9275 26911
rect 10134 26908 10140 26920
rect 9263 26880 10140 26908
rect 9263 26877 9275 26880
rect 9217 26871 9275 26877
rect 4525 26843 4583 26849
rect 4525 26809 4537 26843
rect 4571 26809 4583 26843
rect 9140 26840 9168 26871
rect 10134 26868 10140 26880
rect 10192 26868 10198 26920
rect 10226 26868 10232 26920
rect 10284 26868 10290 26920
rect 9950 26840 9956 26852
rect 9140 26812 9956 26840
rect 4525 26803 4583 26809
rect 9950 26800 9956 26812
rect 10008 26800 10014 26852
rect 8294 26732 8300 26784
rect 8352 26772 8358 26784
rect 8665 26775 8723 26781
rect 8665 26772 8677 26775
rect 8352 26744 8677 26772
rect 8352 26732 8358 26744
rect 8665 26741 8677 26744
rect 8711 26741 8723 26775
rect 8665 26735 8723 26741
rect 8846 26732 8852 26784
rect 8904 26732 8910 26784
rect 9493 26775 9551 26781
rect 9493 26741 9505 26775
rect 9539 26772 9551 26775
rect 9674 26772 9680 26784
rect 9539 26744 9680 26772
rect 9539 26741 9551 26744
rect 9493 26735 9551 26741
rect 9674 26732 9680 26744
rect 9732 26732 9738 26784
rect 9766 26732 9772 26784
rect 9824 26772 9830 26784
rect 10704 26772 10732 26948
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 12066 26936 12072 26988
rect 12124 26936 12130 26988
rect 12176 26985 12204 27016
rect 12161 26979 12219 26985
rect 12161 26945 12173 26979
rect 12207 26945 12219 26979
rect 12268 26976 12296 27084
rect 12434 27072 12440 27124
rect 12492 27112 12498 27124
rect 12492 27084 12848 27112
rect 12492 27072 12498 27084
rect 12710 27004 12716 27056
rect 12768 27004 12774 27056
rect 12820 27044 12848 27084
rect 12894 27072 12900 27124
rect 12952 27121 12958 27124
rect 12952 27115 12971 27121
rect 12959 27081 12971 27115
rect 12952 27075 12971 27081
rect 12952 27072 12958 27075
rect 14366 27072 14372 27124
rect 14424 27112 14430 27124
rect 14461 27115 14519 27121
rect 14461 27112 14473 27115
rect 14424 27084 14473 27112
rect 14424 27072 14430 27084
rect 14461 27081 14473 27084
rect 14507 27081 14519 27115
rect 14461 27075 14519 27081
rect 15473 27115 15531 27121
rect 15473 27081 15485 27115
rect 15519 27112 15531 27115
rect 16390 27112 16396 27124
rect 15519 27084 16396 27112
rect 15519 27081 15531 27084
rect 15473 27075 15531 27081
rect 16390 27072 16396 27084
rect 16448 27072 16454 27124
rect 17144 27084 18184 27112
rect 13078 27044 13084 27056
rect 12820 27016 13084 27044
rect 13078 27004 13084 27016
rect 13136 27044 13142 27056
rect 13136 27016 15056 27044
rect 13136 27004 13142 27016
rect 14093 26979 14151 26985
rect 14093 26976 14105 26979
rect 12268 26948 14105 26976
rect 12161 26939 12219 26945
rect 14093 26945 14105 26948
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 14921 26979 14979 26985
rect 14921 26945 14933 26979
rect 14967 26945 14979 26979
rect 15028 26976 15056 27016
rect 15102 27004 15108 27056
rect 15160 27044 15166 27056
rect 15289 27047 15347 27053
rect 15289 27044 15301 27047
rect 15160 27016 15301 27044
rect 15160 27004 15166 27016
rect 15289 27013 15301 27016
rect 15335 27013 15347 27047
rect 17034 27044 17040 27056
rect 15289 27007 15347 27013
rect 15672 27016 17040 27044
rect 15473 26979 15531 26985
rect 15473 26976 15485 26979
rect 15028 26948 15485 26976
rect 14921 26939 14979 26945
rect 15473 26945 15485 26948
rect 15519 26976 15531 26979
rect 15672 26976 15700 27016
rect 17034 27004 17040 27016
rect 17092 27004 17098 27056
rect 17144 27053 17172 27084
rect 18156 27056 18184 27084
rect 18598 27072 18604 27124
rect 18656 27112 18662 27124
rect 18719 27115 18777 27121
rect 18719 27112 18731 27115
rect 18656 27084 18731 27112
rect 18656 27072 18662 27084
rect 18719 27081 18731 27084
rect 18765 27112 18777 27115
rect 20622 27112 20628 27124
rect 18765 27084 20628 27112
rect 18765 27081 18777 27084
rect 18719 27075 18777 27081
rect 20622 27072 20628 27084
rect 20680 27072 20686 27124
rect 21266 27072 21272 27124
rect 21324 27112 21330 27124
rect 25130 27112 25136 27124
rect 21324 27084 21496 27112
rect 21324 27072 21330 27084
rect 17129 27047 17187 27053
rect 17129 27013 17141 27047
rect 17175 27013 17187 27047
rect 17129 27007 17187 27013
rect 17359 27013 17417 27019
rect 17359 27010 17371 27013
rect 15519 26948 15700 26976
rect 15519 26945 15531 26948
rect 15473 26939 15531 26945
rect 10778 26868 10784 26920
rect 10836 26908 10842 26920
rect 11517 26911 11575 26917
rect 11517 26908 11529 26911
rect 10836 26880 11529 26908
rect 10836 26868 10842 26880
rect 11517 26877 11529 26880
rect 11563 26877 11575 26911
rect 11517 26871 11575 26877
rect 13446 26868 13452 26920
rect 13504 26908 13510 26920
rect 13998 26908 14004 26920
rect 13504 26880 14004 26908
rect 13504 26868 13510 26880
rect 13998 26868 14004 26880
rect 14056 26868 14062 26920
rect 14185 26911 14243 26917
rect 14185 26877 14197 26911
rect 14231 26908 14243 26911
rect 14642 26908 14648 26920
rect 14231 26880 14648 26908
rect 14231 26877 14243 26880
rect 14185 26871 14243 26877
rect 14642 26868 14648 26880
rect 14700 26908 14706 26920
rect 14737 26911 14795 26917
rect 14737 26908 14749 26911
rect 14700 26880 14749 26908
rect 14700 26868 14706 26880
rect 14737 26877 14749 26880
rect 14783 26877 14795 26911
rect 14936 26908 14964 26939
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 15933 26979 15991 26985
rect 15933 26976 15945 26979
rect 15896 26948 15945 26976
rect 15896 26936 15902 26948
rect 15933 26945 15945 26948
rect 15979 26945 15991 26979
rect 15933 26939 15991 26945
rect 16298 26936 16304 26988
rect 16356 26936 16362 26988
rect 16669 26979 16727 26985
rect 16669 26945 16681 26979
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 17344 26979 17371 27010
rect 17405 26979 17417 27013
rect 18138 27004 18144 27056
rect 18196 27004 18202 27056
rect 18230 27004 18236 27056
rect 18288 27044 18294 27056
rect 18509 27047 18567 27053
rect 18509 27044 18521 27047
rect 18288 27016 18521 27044
rect 18288 27004 18294 27016
rect 18509 27013 18521 27016
rect 18555 27013 18567 27047
rect 18509 27007 18567 27013
rect 19978 27004 19984 27056
rect 20036 27044 20042 27056
rect 20036 27016 20668 27044
rect 20036 27004 20042 27016
rect 17344 26973 17417 26979
rect 15010 26908 15016 26920
rect 14737 26871 14795 26877
rect 14844 26880 15016 26908
rect 12158 26840 12164 26852
rect 11256 26812 12164 26840
rect 11256 26784 11284 26812
rect 12158 26800 12164 26812
rect 12216 26840 12222 26852
rect 12216 26812 12296 26840
rect 12216 26800 12222 26812
rect 9824 26744 10732 26772
rect 9824 26732 9830 26744
rect 11238 26732 11244 26784
rect 11296 26732 11302 26784
rect 11974 26732 11980 26784
rect 12032 26732 12038 26784
rect 12268 26781 12296 26812
rect 12526 26800 12532 26852
rect 12584 26840 12590 26852
rect 14844 26840 14872 26880
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 15197 26911 15255 26917
rect 15197 26877 15209 26911
rect 15243 26908 15255 26911
rect 16684 26908 16712 26939
rect 17344 26908 17372 26973
rect 18782 26936 18788 26988
rect 18840 26936 18846 26988
rect 19153 26979 19211 26985
rect 19153 26945 19165 26979
rect 19199 26976 19211 26979
rect 19334 26976 19340 26988
rect 19199 26948 19340 26976
rect 19199 26945 19211 26948
rect 19153 26939 19211 26945
rect 19334 26936 19340 26948
rect 19392 26936 19398 26988
rect 20530 26976 20536 26988
rect 19904 26948 20536 26976
rect 18800 26908 18828 26936
rect 15243 26880 16712 26908
rect 16776 26880 17372 26908
rect 18524 26880 18828 26908
rect 19245 26911 19303 26917
rect 15243 26877 15255 26880
rect 15197 26871 15255 26877
rect 12584 26812 14872 26840
rect 12584 26800 12590 26812
rect 12253 26775 12311 26781
rect 12253 26741 12265 26775
rect 12299 26741 12311 26775
rect 12253 26735 12311 26741
rect 12621 26775 12679 26781
rect 12621 26741 12633 26775
rect 12667 26772 12679 26775
rect 12897 26775 12955 26781
rect 12897 26772 12909 26775
rect 12667 26744 12909 26772
rect 12667 26741 12679 26744
rect 12621 26735 12679 26741
rect 12897 26741 12909 26744
rect 12943 26741 12955 26775
rect 12897 26735 12955 26741
rect 13078 26732 13084 26784
rect 13136 26732 13142 26784
rect 13262 26732 13268 26784
rect 13320 26772 13326 26784
rect 14093 26775 14151 26781
rect 14093 26772 14105 26775
rect 13320 26744 14105 26772
rect 13320 26732 13326 26744
rect 14093 26741 14105 26744
rect 14139 26772 14151 26775
rect 14274 26772 14280 26784
rect 14139 26744 14280 26772
rect 14139 26741 14151 26744
rect 14093 26735 14151 26741
rect 14274 26732 14280 26744
rect 14332 26732 14338 26784
rect 14734 26732 14740 26784
rect 14792 26772 14798 26784
rect 15212 26772 15240 26871
rect 15930 26800 15936 26852
rect 15988 26840 15994 26852
rect 16776 26840 16804 26880
rect 15988 26812 16804 26840
rect 15988 26800 15994 26812
rect 17126 26800 17132 26852
rect 17184 26840 17190 26852
rect 17184 26812 17356 26840
rect 17184 26800 17190 26812
rect 14792 26744 15240 26772
rect 14792 26732 14798 26744
rect 16758 26732 16764 26784
rect 16816 26732 16822 26784
rect 17328 26781 17356 26812
rect 17313 26775 17371 26781
rect 17313 26741 17325 26775
rect 17359 26741 17371 26775
rect 17313 26735 17371 26741
rect 17494 26732 17500 26784
rect 17552 26732 17558 26784
rect 18524 26772 18552 26880
rect 19245 26877 19257 26911
rect 19291 26908 19303 26911
rect 19904 26908 19932 26948
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 20640 26985 20668 27016
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26945 20683 26979
rect 20625 26939 20683 26945
rect 20714 26936 20720 26988
rect 20772 26976 20778 26988
rect 20809 26979 20867 26985
rect 20809 26976 20821 26979
rect 20772 26948 20821 26976
rect 20772 26936 20778 26948
rect 20809 26945 20821 26948
rect 20855 26945 20867 26979
rect 20809 26939 20867 26945
rect 21177 26979 21235 26985
rect 21177 26945 21189 26979
rect 21223 26976 21235 26979
rect 21266 26976 21272 26988
rect 21223 26948 21272 26976
rect 21223 26945 21235 26948
rect 21177 26939 21235 26945
rect 21266 26936 21272 26948
rect 21324 26936 21330 26988
rect 21468 26985 21496 27084
rect 24596 27084 25136 27112
rect 24596 27044 24624 27084
rect 25130 27072 25136 27084
rect 25188 27072 25194 27124
rect 25498 27112 25504 27124
rect 25332 27084 25504 27112
rect 23584 27016 24624 27044
rect 21453 26979 21511 26985
rect 21453 26945 21465 26979
rect 21499 26976 21511 26979
rect 21542 26976 21548 26988
rect 21499 26948 21548 26976
rect 21499 26945 21511 26948
rect 21453 26939 21511 26945
rect 21542 26936 21548 26948
rect 21600 26936 21606 26988
rect 21637 26979 21695 26985
rect 21637 26945 21649 26979
rect 21683 26976 21695 26979
rect 22738 26976 22744 26988
rect 21683 26948 22744 26976
rect 21683 26945 21695 26948
rect 21637 26939 21695 26945
rect 22738 26936 22744 26948
rect 22796 26936 22802 26988
rect 22833 26979 22891 26985
rect 22833 26945 22845 26979
rect 22879 26976 22891 26979
rect 22922 26976 22928 26988
rect 22879 26948 22928 26976
rect 22879 26945 22891 26948
rect 22833 26939 22891 26945
rect 22922 26936 22928 26948
rect 22980 26936 22986 26988
rect 23198 26936 23204 26988
rect 23256 26936 23262 26988
rect 23584 26985 23612 27016
rect 23569 26979 23627 26985
rect 23569 26945 23581 26979
rect 23615 26945 23627 26979
rect 23569 26939 23627 26945
rect 24394 26936 24400 26988
rect 24452 26936 24458 26988
rect 24596 26985 24624 27016
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26945 24639 26979
rect 24581 26939 24639 26945
rect 24946 26936 24952 26988
rect 25004 26936 25010 26988
rect 25130 26936 25136 26988
rect 25188 26936 25194 26988
rect 25332 26985 25360 27084
rect 25498 27072 25504 27084
rect 25556 27112 25562 27124
rect 25556 27084 25636 27112
rect 25556 27072 25562 27084
rect 25608 27044 25636 27084
rect 25682 27072 25688 27124
rect 25740 27112 25746 27124
rect 25740 27084 26464 27112
rect 25740 27072 25746 27084
rect 26436 27044 26464 27084
rect 26510 27072 26516 27124
rect 26568 27112 26574 27124
rect 27157 27115 27215 27121
rect 27157 27112 27169 27115
rect 26568 27084 27169 27112
rect 26568 27072 26574 27084
rect 27157 27081 27169 27084
rect 27203 27081 27215 27115
rect 27157 27075 27215 27081
rect 27893 27115 27951 27121
rect 27893 27081 27905 27115
rect 27939 27112 27951 27115
rect 28258 27112 28264 27124
rect 27939 27084 28264 27112
rect 27939 27081 27951 27084
rect 27893 27075 27951 27081
rect 28258 27072 28264 27084
rect 28316 27072 28322 27124
rect 28537 27115 28595 27121
rect 28537 27081 28549 27115
rect 28583 27112 28595 27115
rect 28810 27112 28816 27124
rect 28583 27084 28816 27112
rect 28583 27081 28595 27084
rect 28537 27075 28595 27081
rect 28810 27072 28816 27084
rect 28868 27072 28874 27124
rect 28905 27115 28963 27121
rect 28905 27081 28917 27115
rect 28951 27112 28963 27115
rect 28994 27112 29000 27124
rect 28951 27084 29000 27112
rect 28951 27081 28963 27084
rect 28905 27075 28963 27081
rect 28994 27072 29000 27084
rect 29052 27072 29058 27124
rect 30190 27072 30196 27124
rect 30248 27112 30254 27124
rect 30285 27115 30343 27121
rect 30285 27112 30297 27115
rect 30248 27084 30297 27112
rect 30248 27072 30254 27084
rect 30285 27081 30297 27084
rect 30331 27081 30343 27115
rect 33502 27112 33508 27124
rect 30285 27075 30343 27081
rect 33060 27084 33508 27112
rect 32858 27044 32864 27056
rect 25608 27016 26096 27044
rect 26436 27016 28120 27044
rect 25317 26979 25375 26985
rect 25317 26945 25329 26979
rect 25363 26945 25375 26979
rect 25317 26939 25375 26945
rect 25682 26936 25688 26988
rect 25740 26936 25746 26988
rect 26068 26976 26096 27016
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26068 26948 27169 26976
rect 27157 26945 27169 26948
rect 27203 26976 27215 26979
rect 27246 26976 27252 26988
rect 27203 26948 27252 26976
rect 27203 26945 27215 26948
rect 27157 26939 27215 26945
rect 27246 26936 27252 26948
rect 27304 26936 27310 26988
rect 27338 26936 27344 26988
rect 27396 26976 27402 26988
rect 27396 26948 27660 26976
rect 27396 26936 27402 26948
rect 19291 26880 19932 26908
rect 20441 26911 20499 26917
rect 19291 26877 19303 26880
rect 19245 26871 19303 26877
rect 20441 26877 20453 26911
rect 20487 26908 20499 26911
rect 20487 26880 23704 26908
rect 20487 26877 20499 26880
rect 20441 26871 20499 26877
rect 18598 26800 18604 26852
rect 18656 26840 18662 26852
rect 20073 26843 20131 26849
rect 20073 26840 20085 26843
rect 18656 26812 20085 26840
rect 18656 26800 18662 26812
rect 18693 26775 18751 26781
rect 18693 26772 18705 26775
rect 18524 26744 18705 26772
rect 18693 26741 18705 26744
rect 18739 26741 18751 26775
rect 18693 26735 18751 26741
rect 18782 26732 18788 26784
rect 18840 26772 18846 26784
rect 18877 26775 18935 26781
rect 18877 26772 18889 26775
rect 18840 26744 18889 26772
rect 18840 26732 18846 26744
rect 18877 26741 18889 26744
rect 18923 26772 18935 26775
rect 19058 26772 19064 26784
rect 18923 26744 19064 26772
rect 18923 26741 18935 26744
rect 18877 26735 18935 26741
rect 19058 26732 19064 26744
rect 19116 26732 19122 26784
rect 19352 26781 19380 26812
rect 20073 26809 20085 26812
rect 20119 26809 20131 26843
rect 20073 26803 20131 26809
rect 20533 26843 20591 26849
rect 20533 26809 20545 26843
rect 20579 26840 20591 26843
rect 23382 26840 23388 26852
rect 20579 26812 23388 26840
rect 20579 26809 20591 26812
rect 20533 26803 20591 26809
rect 23382 26800 23388 26812
rect 23440 26800 23446 26852
rect 23676 26840 23704 26880
rect 23750 26868 23756 26920
rect 23808 26868 23814 26920
rect 23952 26880 24808 26908
rect 23952 26840 23980 26880
rect 23676 26812 23980 26840
rect 24029 26843 24087 26849
rect 24029 26809 24041 26843
rect 24075 26840 24087 26843
rect 24118 26840 24124 26852
rect 24075 26812 24124 26840
rect 24075 26809 24087 26812
rect 24029 26803 24087 26809
rect 24118 26800 24124 26812
rect 24176 26800 24182 26852
rect 24578 26800 24584 26852
rect 24636 26800 24642 26852
rect 24670 26800 24676 26852
rect 24728 26800 24734 26852
rect 24780 26840 24808 26880
rect 24854 26868 24860 26920
rect 24912 26908 24918 26920
rect 25958 26908 25964 26920
rect 24912 26880 25964 26908
rect 24912 26868 24918 26880
rect 25958 26868 25964 26880
rect 26016 26868 26022 26920
rect 26970 26868 26976 26920
rect 27028 26868 27034 26920
rect 27430 26868 27436 26920
rect 27488 26908 27494 26920
rect 27525 26911 27583 26917
rect 27525 26908 27537 26911
rect 27488 26880 27537 26908
rect 27488 26868 27494 26880
rect 27525 26877 27537 26880
rect 27571 26877 27583 26911
rect 27632 26908 27660 26948
rect 27706 26936 27712 26988
rect 27764 26936 27770 26988
rect 28092 26985 28120 27016
rect 28920 27016 32864 27044
rect 27801 26979 27859 26985
rect 27801 26945 27813 26979
rect 27847 26945 27859 26979
rect 27801 26939 27859 26945
rect 28077 26979 28135 26985
rect 28077 26945 28089 26979
rect 28123 26976 28135 26979
rect 28166 26976 28172 26988
rect 28123 26948 28172 26976
rect 28123 26945 28135 26948
rect 28077 26939 28135 26945
rect 27816 26908 27844 26939
rect 28166 26936 28172 26948
rect 28224 26936 28230 26988
rect 28261 26979 28319 26985
rect 28261 26945 28273 26979
rect 28307 26945 28319 26979
rect 28261 26939 28319 26945
rect 28276 26908 28304 26939
rect 28350 26936 28356 26988
rect 28408 26936 28414 26988
rect 28534 26936 28540 26988
rect 28592 26936 28598 26988
rect 28718 26936 28724 26988
rect 28776 26976 28782 26988
rect 28920 26985 28948 27016
rect 32858 27004 32864 27016
rect 32916 27004 32922 27056
rect 28905 26979 28963 26985
rect 28905 26976 28917 26979
rect 28776 26948 28917 26976
rect 28776 26936 28782 26948
rect 28905 26945 28917 26948
rect 28951 26945 28963 26979
rect 28905 26939 28963 26945
rect 28997 26979 29055 26985
rect 28997 26945 29009 26979
rect 29043 26976 29055 26979
rect 29822 26976 29828 26988
rect 29043 26948 29828 26976
rect 29043 26945 29055 26948
rect 28997 26939 29055 26945
rect 27632 26880 27844 26908
rect 28184 26880 28304 26908
rect 28368 26908 28396 26936
rect 28813 26911 28871 26917
rect 28813 26908 28825 26911
rect 28368 26880 28825 26908
rect 27525 26871 27583 26877
rect 25866 26840 25872 26852
rect 24780 26812 25872 26840
rect 25866 26800 25872 26812
rect 25924 26800 25930 26852
rect 26234 26800 26240 26852
rect 26292 26800 26298 26852
rect 26988 26840 27016 26868
rect 28184 26840 28212 26880
rect 28813 26877 28825 26880
rect 28859 26877 28871 26911
rect 28813 26871 28871 26877
rect 29012 26852 29040 26939
rect 29822 26936 29828 26948
rect 29880 26936 29886 26988
rect 30193 26979 30251 26985
rect 30193 26945 30205 26979
rect 30239 26976 30251 26979
rect 30558 26976 30564 26988
rect 30239 26948 30564 26976
rect 30239 26945 30251 26948
rect 30193 26939 30251 26945
rect 30558 26936 30564 26948
rect 30616 26936 30622 26988
rect 31294 26936 31300 26988
rect 31352 26936 31358 26988
rect 33060 26985 33088 27084
rect 33502 27072 33508 27084
rect 33560 27072 33566 27124
rect 34790 27112 34796 27124
rect 33704 27084 34796 27112
rect 33318 27004 33324 27056
rect 33376 27044 33382 27056
rect 33594 27044 33600 27056
rect 33376 27016 33600 27044
rect 33376 27004 33382 27016
rect 33594 27004 33600 27016
rect 33652 27004 33658 27056
rect 33045 26979 33103 26985
rect 33045 26945 33057 26979
rect 33091 26945 33103 26979
rect 33045 26939 33103 26945
rect 33134 26936 33140 26988
rect 33192 26976 33198 26988
rect 33229 26979 33287 26985
rect 33229 26976 33241 26979
rect 33192 26948 33241 26976
rect 33192 26936 33198 26948
rect 33229 26945 33241 26948
rect 33275 26945 33287 26979
rect 33229 26939 33287 26945
rect 33413 26979 33471 26985
rect 33413 26945 33425 26979
rect 33459 26976 33471 26979
rect 33502 26976 33508 26988
rect 33459 26948 33508 26976
rect 33459 26945 33471 26948
rect 33413 26939 33471 26945
rect 33502 26936 33508 26948
rect 33560 26936 33566 26988
rect 33704 26985 33732 27084
rect 34790 27072 34796 27084
rect 34848 27072 34854 27124
rect 35434 27044 35440 27056
rect 35190 27016 35440 27044
rect 35434 27004 35440 27016
rect 35492 27004 35498 27056
rect 33689 26979 33747 26985
rect 33689 26945 33701 26979
rect 33735 26945 33747 26979
rect 33689 26939 33747 26945
rect 29181 26911 29239 26917
rect 29181 26877 29193 26911
rect 29227 26908 29239 26911
rect 29546 26908 29552 26920
rect 29227 26880 29552 26908
rect 29227 26877 29239 26880
rect 29181 26871 29239 26877
rect 26988 26812 28212 26840
rect 28350 26800 28356 26852
rect 28408 26800 28414 26852
rect 28629 26843 28687 26849
rect 28629 26809 28641 26843
rect 28675 26840 28687 26843
rect 28994 26840 29000 26852
rect 28675 26812 29000 26840
rect 28675 26809 28687 26812
rect 28629 26803 28687 26809
rect 28994 26800 29000 26812
rect 29052 26800 29058 26852
rect 19337 26775 19395 26781
rect 19337 26741 19349 26775
rect 19383 26741 19395 26775
rect 19337 26735 19395 26741
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 19521 26775 19579 26781
rect 19521 26772 19533 26775
rect 19484 26744 19533 26772
rect 19484 26732 19490 26744
rect 19521 26741 19533 26744
rect 19567 26741 19579 26775
rect 19521 26735 19579 26741
rect 20162 26732 20168 26784
rect 20220 26772 20226 26784
rect 20349 26775 20407 26781
rect 20349 26772 20361 26775
rect 20220 26744 20361 26772
rect 20220 26732 20226 26744
rect 20349 26741 20361 26744
rect 20395 26741 20407 26775
rect 20349 26735 20407 26741
rect 20622 26732 20628 26784
rect 20680 26772 20686 26784
rect 20901 26775 20959 26781
rect 20901 26772 20913 26775
rect 20680 26744 20913 26772
rect 20680 26732 20686 26744
rect 20901 26741 20913 26744
rect 20947 26741 20959 26775
rect 20901 26735 20959 26741
rect 20990 26732 20996 26784
rect 21048 26772 21054 26784
rect 21266 26772 21272 26784
rect 21048 26744 21272 26772
rect 21048 26732 21054 26744
rect 21266 26732 21272 26744
rect 21324 26732 21330 26784
rect 21361 26775 21419 26781
rect 21361 26741 21373 26775
rect 21407 26772 21419 26775
rect 22002 26772 22008 26784
rect 21407 26744 22008 26772
rect 21407 26741 21419 26744
rect 21361 26735 21419 26741
rect 22002 26732 22008 26744
rect 22060 26732 22066 26784
rect 23198 26732 23204 26784
rect 23256 26772 23262 26784
rect 24946 26772 24952 26784
rect 23256 26744 24952 26772
rect 23256 26732 23262 26744
rect 24946 26732 24952 26744
rect 25004 26732 25010 26784
rect 25774 26732 25780 26784
rect 25832 26772 25838 26784
rect 26142 26772 26148 26784
rect 25832 26744 26148 26772
rect 25832 26732 25838 26744
rect 26142 26732 26148 26744
rect 26200 26732 26206 26784
rect 26252 26772 26280 26800
rect 28368 26772 28396 26800
rect 26252 26744 28396 26772
rect 28534 26732 28540 26784
rect 28592 26772 28598 26784
rect 29196 26772 29224 26871
rect 29546 26868 29552 26880
rect 29604 26868 29610 26920
rect 30469 26911 30527 26917
rect 30469 26877 30481 26911
rect 30515 26908 30527 26911
rect 31312 26908 31340 26936
rect 33965 26911 34023 26917
rect 33965 26908 33977 26911
rect 30515 26880 31340 26908
rect 33612 26880 33977 26908
rect 30515 26877 30527 26880
rect 30469 26871 30527 26877
rect 30098 26840 30104 26852
rect 29656 26812 30104 26840
rect 29656 26784 29684 26812
rect 30098 26800 30104 26812
rect 30156 26840 30162 26852
rect 30561 26843 30619 26849
rect 30156 26812 30420 26840
rect 30156 26800 30162 26812
rect 28592 26744 29224 26772
rect 28592 26732 28598 26744
rect 29638 26732 29644 26784
rect 29696 26732 29702 26784
rect 30006 26732 30012 26784
rect 30064 26732 30070 26784
rect 30392 26772 30420 26812
rect 30561 26809 30573 26843
rect 30607 26840 30619 26843
rect 31018 26840 31024 26852
rect 30607 26812 31024 26840
rect 30607 26809 30619 26812
rect 30561 26803 30619 26809
rect 31018 26800 31024 26812
rect 31076 26800 31082 26852
rect 33612 26849 33640 26880
rect 33965 26877 33977 26880
rect 34011 26877 34023 26911
rect 33965 26871 34023 26877
rect 34330 26868 34336 26920
rect 34388 26908 34394 26920
rect 35437 26911 35495 26917
rect 35437 26908 35449 26911
rect 34388 26880 35449 26908
rect 34388 26868 34394 26880
rect 35437 26877 35449 26880
rect 35483 26877 35495 26911
rect 35437 26871 35495 26877
rect 33597 26843 33655 26849
rect 33597 26809 33609 26843
rect 33643 26809 33655 26843
rect 33597 26803 33655 26809
rect 30753 26775 30811 26781
rect 30753 26772 30765 26775
rect 30392 26744 30765 26772
rect 30753 26741 30765 26744
rect 30799 26741 30811 26775
rect 30753 26735 30811 26741
rect 32582 26732 32588 26784
rect 32640 26772 32646 26784
rect 34422 26772 34428 26784
rect 32640 26744 34428 26772
rect 32640 26732 32646 26744
rect 34422 26732 34428 26744
rect 34480 26732 34486 26784
rect 1104 26682 41400 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 41400 26682
rect 1104 26608 41400 26630
rect 6822 26528 6828 26580
rect 6880 26568 6886 26580
rect 7929 26571 7987 26577
rect 7929 26568 7941 26571
rect 6880 26540 7941 26568
rect 6880 26528 6886 26540
rect 7929 26537 7941 26540
rect 7975 26568 7987 26571
rect 13262 26568 13268 26580
rect 7975 26540 13268 26568
rect 7975 26537 7987 26540
rect 7929 26531 7987 26537
rect 13262 26528 13268 26540
rect 13320 26528 13326 26580
rect 14090 26528 14096 26580
rect 14148 26568 14154 26580
rect 16298 26568 16304 26580
rect 14148 26540 16304 26568
rect 14148 26528 14154 26540
rect 16298 26528 16304 26540
rect 16356 26528 16362 26580
rect 16758 26528 16764 26580
rect 16816 26568 16822 26580
rect 19705 26571 19763 26577
rect 16816 26540 19656 26568
rect 16816 26528 16822 26540
rect 5353 26503 5411 26509
rect 5353 26469 5365 26503
rect 5399 26469 5411 26503
rect 5353 26463 5411 26469
rect 1670 26324 1676 26376
rect 1728 26324 1734 26376
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26364 5319 26367
rect 5368 26364 5396 26463
rect 9490 26460 9496 26512
rect 9548 26460 9554 26512
rect 10505 26503 10563 26509
rect 10505 26469 10517 26503
rect 10551 26500 10563 26503
rect 11054 26500 11060 26512
rect 10551 26472 11060 26500
rect 10551 26469 10563 26472
rect 10505 26463 10563 26469
rect 11054 26460 11060 26472
rect 11112 26460 11118 26512
rect 11425 26503 11483 26509
rect 11425 26469 11437 26503
rect 11471 26500 11483 26503
rect 11471 26472 18920 26500
rect 11471 26469 11483 26472
rect 11425 26463 11483 26469
rect 5997 26435 6055 26441
rect 5997 26401 6009 26435
rect 6043 26432 6055 26435
rect 6730 26432 6736 26444
rect 6043 26404 6736 26432
rect 6043 26401 6055 26404
rect 5997 26395 6055 26401
rect 6730 26392 6736 26404
rect 6788 26432 6794 26444
rect 8386 26432 8392 26444
rect 6788 26404 8392 26432
rect 6788 26392 6794 26404
rect 8386 26392 8392 26404
rect 8444 26392 8450 26444
rect 9508 26432 9536 26460
rect 9140 26404 9536 26432
rect 9585 26435 9643 26441
rect 5307 26336 5396 26364
rect 7653 26367 7711 26373
rect 5307 26333 5319 26336
rect 5261 26327 5319 26333
rect 7653 26333 7665 26367
rect 7699 26364 7711 26367
rect 8202 26364 8208 26376
rect 7699 26336 8208 26364
rect 7699 26333 7711 26336
rect 7653 26327 7711 26333
rect 8202 26324 8208 26336
rect 8260 26324 8266 26376
rect 9140 26373 9168 26404
rect 9585 26401 9597 26435
rect 9631 26432 9643 26435
rect 9766 26432 9772 26444
rect 9631 26404 9772 26432
rect 9631 26401 9643 26404
rect 9585 26395 9643 26401
rect 9766 26392 9772 26404
rect 9824 26392 9830 26444
rect 10594 26432 10600 26444
rect 9876 26404 10600 26432
rect 9125 26367 9183 26373
rect 9125 26333 9137 26367
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 9214 26324 9220 26376
rect 9272 26324 9278 26376
rect 9398 26364 9404 26376
rect 9456 26373 9462 26376
rect 9456 26367 9485 26373
rect 9385 26336 9404 26364
rect 9398 26324 9404 26336
rect 9473 26364 9485 26367
rect 9876 26364 9904 26404
rect 10594 26392 10600 26404
rect 10652 26432 10658 26444
rect 11072 26432 11100 26460
rect 10652 26404 10824 26432
rect 11072 26404 11560 26432
rect 10652 26392 10658 26404
rect 9473 26336 9904 26364
rect 9473 26333 9485 26336
rect 9456 26327 9485 26333
rect 9456 26324 9462 26327
rect 9950 26324 9956 26376
rect 10008 26364 10014 26376
rect 10686 26364 10692 26376
rect 10008 26336 10692 26364
rect 10008 26324 10014 26336
rect 10686 26324 10692 26336
rect 10744 26324 10750 26376
rect 10796 26373 10824 26404
rect 11532 26373 11560 26404
rect 11698 26392 11704 26444
rect 11756 26392 11762 26444
rect 15105 26435 15163 26441
rect 15105 26401 15117 26435
rect 15151 26432 15163 26435
rect 15194 26432 15200 26444
rect 15151 26404 15200 26432
rect 15151 26401 15163 26404
rect 15105 26395 15163 26401
rect 15194 26392 15200 26404
rect 15252 26392 15258 26444
rect 15378 26392 15384 26444
rect 15436 26392 15442 26444
rect 15749 26435 15807 26441
rect 15749 26401 15761 26435
rect 15795 26432 15807 26435
rect 15838 26432 15844 26444
rect 15795 26404 15844 26432
rect 15795 26401 15807 26404
rect 15749 26395 15807 26401
rect 15838 26392 15844 26404
rect 15896 26392 15902 26444
rect 16022 26392 16028 26444
rect 16080 26432 16086 26444
rect 16080 26404 16620 26432
rect 16080 26392 16086 26404
rect 10781 26367 10839 26373
rect 10781 26333 10793 26367
rect 10827 26333 10839 26367
rect 10781 26327 10839 26333
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26333 11391 26367
rect 11333 26327 11391 26333
rect 11517 26367 11575 26373
rect 11517 26333 11529 26367
rect 11563 26333 11575 26367
rect 11517 26327 11575 26333
rect 1688 26296 1716 26324
rect 5721 26299 5779 26305
rect 5721 26296 5733 26299
rect 1688 26268 5733 26296
rect 5721 26265 5733 26268
rect 5767 26296 5779 26299
rect 6914 26296 6920 26308
rect 5767 26268 6920 26296
rect 5767 26265 5779 26268
rect 5721 26259 5779 26265
rect 6914 26256 6920 26268
rect 6972 26256 6978 26308
rect 8662 26256 8668 26308
rect 8720 26296 8726 26308
rect 8941 26299 8999 26305
rect 8941 26296 8953 26299
rect 8720 26268 8953 26296
rect 8720 26256 8726 26268
rect 8941 26265 8953 26268
rect 8987 26265 8999 26299
rect 8941 26259 8999 26265
rect 9309 26299 9367 26305
rect 9309 26265 9321 26299
rect 9355 26265 9367 26299
rect 9309 26259 9367 26265
rect 5074 26188 5080 26240
rect 5132 26188 5138 26240
rect 5813 26231 5871 26237
rect 5813 26197 5825 26231
rect 5859 26228 5871 26231
rect 6546 26228 6552 26240
rect 5859 26200 6552 26228
rect 5859 26197 5871 26200
rect 5813 26191 5871 26197
rect 6546 26188 6552 26200
rect 6604 26188 6610 26240
rect 8478 26188 8484 26240
rect 8536 26228 8542 26240
rect 9324 26228 9352 26259
rect 10226 26256 10232 26308
rect 10284 26296 10290 26308
rect 10502 26296 10508 26308
rect 10284 26268 10508 26296
rect 10284 26256 10290 26268
rect 10502 26256 10508 26268
rect 10560 26296 10566 26308
rect 10962 26296 10968 26308
rect 10560 26268 10968 26296
rect 10560 26256 10566 26268
rect 10962 26256 10968 26268
rect 11020 26256 11026 26308
rect 11348 26296 11376 26327
rect 11716 26296 11744 26392
rect 14918 26324 14924 26376
rect 14976 26324 14982 26376
rect 15286 26324 15292 26376
rect 15344 26324 15350 26376
rect 15473 26367 15531 26373
rect 15473 26364 15485 26367
rect 15397 26336 15485 26364
rect 11348 26268 11744 26296
rect 12158 26256 12164 26308
rect 12216 26256 12222 26308
rect 14274 26256 14280 26308
rect 14332 26256 14338 26308
rect 14936 26296 14964 26324
rect 15397 26296 15425 26336
rect 15473 26333 15485 26336
rect 15519 26333 15531 26367
rect 15473 26327 15531 26333
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26333 15623 26367
rect 15565 26327 15623 26333
rect 15933 26367 15991 26373
rect 15933 26333 15945 26367
rect 15979 26364 15991 26367
rect 16482 26364 16488 26376
rect 15979 26336 16488 26364
rect 15979 26333 15991 26336
rect 15933 26327 15991 26333
rect 15580 26296 15608 26327
rect 16482 26324 16488 26336
rect 16540 26324 16546 26376
rect 14936 26268 15425 26296
rect 15488 26268 15608 26296
rect 16592 26296 16620 26404
rect 16942 26392 16948 26444
rect 17000 26432 17006 26444
rect 18233 26435 18291 26441
rect 18233 26432 18245 26435
rect 17000 26404 18245 26432
rect 17000 26392 17006 26404
rect 18233 26401 18245 26404
rect 18279 26401 18291 26435
rect 18233 26395 18291 26401
rect 18598 26392 18604 26444
rect 18656 26392 18662 26444
rect 17126 26324 17132 26376
rect 17184 26364 17190 26376
rect 17402 26364 17408 26376
rect 17184 26336 17408 26364
rect 17184 26324 17190 26336
rect 17402 26324 17408 26336
rect 17460 26324 17466 26376
rect 17954 26324 17960 26376
rect 18012 26324 18018 26376
rect 18616 26364 18644 26392
rect 18892 26373 18920 26472
rect 19058 26460 19064 26512
rect 19116 26460 19122 26512
rect 19628 26500 19656 26540
rect 19705 26537 19717 26571
rect 19751 26568 19763 26571
rect 22646 26568 22652 26580
rect 19751 26540 22652 26568
rect 19751 26537 19763 26540
rect 19705 26531 19763 26537
rect 22646 26528 22652 26540
rect 22704 26568 22710 26580
rect 23290 26568 23296 26580
rect 22704 26540 23296 26568
rect 22704 26528 22710 26540
rect 23290 26528 23296 26540
rect 23348 26528 23354 26580
rect 25682 26568 25688 26580
rect 25424 26540 25688 26568
rect 19628 26472 20944 26500
rect 19076 26432 19104 26460
rect 19613 26435 19671 26441
rect 19613 26432 19625 26435
rect 19076 26404 19625 26432
rect 19613 26401 19625 26404
rect 19659 26401 19671 26435
rect 19613 26395 19671 26401
rect 19797 26435 19855 26441
rect 19797 26401 19809 26435
rect 19843 26432 19855 26435
rect 20806 26432 20812 26444
rect 19843 26404 20392 26432
rect 19843 26401 19855 26404
rect 19797 26395 19855 26401
rect 18693 26367 18751 26373
rect 18693 26364 18705 26367
rect 18616 26336 18705 26364
rect 18693 26333 18705 26336
rect 18739 26333 18751 26367
rect 18693 26327 18751 26333
rect 18785 26367 18843 26373
rect 18785 26333 18797 26367
rect 18831 26333 18843 26367
rect 18785 26327 18843 26333
rect 18877 26367 18935 26373
rect 18877 26333 18889 26367
rect 18923 26333 18935 26367
rect 18877 26327 18935 26333
rect 19061 26367 19119 26373
rect 19061 26333 19073 26367
rect 19107 26364 19119 26367
rect 19107 26336 19278 26364
rect 19107 26333 19119 26336
rect 19061 26327 19119 26333
rect 17862 26296 17868 26308
rect 16592 26268 17868 26296
rect 12176 26228 12204 26256
rect 8536 26200 12204 26228
rect 14292 26228 14320 26256
rect 15488 26240 15516 26268
rect 17862 26256 17868 26268
rect 17920 26256 17926 26308
rect 18230 26256 18236 26308
rect 18288 26296 18294 26308
rect 18417 26299 18475 26305
rect 18417 26296 18429 26299
rect 18288 26268 18429 26296
rect 18288 26256 18294 26268
rect 18417 26265 18429 26268
rect 18463 26265 18475 26299
rect 18800 26296 18828 26327
rect 19150 26296 19156 26308
rect 18800 26268 19156 26296
rect 18417 26259 18475 26265
rect 19150 26256 19156 26268
rect 19208 26256 19214 26308
rect 15286 26228 15292 26240
rect 14292 26200 15292 26228
rect 8536 26188 8542 26200
rect 15286 26188 15292 26200
rect 15344 26188 15350 26240
rect 15470 26188 15476 26240
rect 15528 26188 15534 26240
rect 15838 26188 15844 26240
rect 15896 26228 15902 26240
rect 16117 26231 16175 26237
rect 16117 26228 16129 26231
rect 15896 26200 16129 26228
rect 15896 26188 15902 26200
rect 16117 26197 16129 26200
rect 16163 26197 16175 26231
rect 16117 26191 16175 26197
rect 17034 26188 17040 26240
rect 17092 26228 17098 26240
rect 18046 26228 18052 26240
rect 17092 26200 18052 26228
rect 17092 26188 17098 26200
rect 18046 26188 18052 26200
rect 18104 26228 18110 26240
rect 19058 26228 19064 26240
rect 18104 26200 19064 26228
rect 18104 26188 18110 26200
rect 19058 26188 19064 26200
rect 19116 26228 19122 26240
rect 19250 26228 19278 26336
rect 19518 26324 19524 26376
rect 19576 26324 19582 26376
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 19978 26364 19984 26376
rect 19935 26336 19984 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 20073 26367 20131 26373
rect 20073 26333 20085 26367
rect 20119 26333 20131 26367
rect 20073 26327 20131 26333
rect 19536 26296 19564 26324
rect 20088 26296 20116 26327
rect 20364 26308 20392 26404
rect 20640 26404 20812 26432
rect 20640 26373 20668 26404
rect 20806 26392 20812 26404
rect 20864 26392 20870 26444
rect 20916 26373 20944 26472
rect 21358 26460 21364 26512
rect 21416 26460 21422 26512
rect 22189 26503 22247 26509
rect 22189 26469 22201 26503
rect 22235 26469 22247 26503
rect 22189 26463 22247 26469
rect 21376 26432 21404 26460
rect 21008 26404 21404 26432
rect 22204 26432 22232 26463
rect 22738 26460 22744 26512
rect 22796 26500 22802 26512
rect 22833 26503 22891 26509
rect 22833 26500 22845 26503
rect 22796 26472 22845 26500
rect 22796 26460 22802 26472
rect 22833 26469 22845 26472
rect 22879 26469 22891 26503
rect 22833 26463 22891 26469
rect 22922 26460 22928 26512
rect 22980 26500 22986 26512
rect 23842 26500 23848 26512
rect 22980 26472 23152 26500
rect 22980 26460 22986 26472
rect 23124 26441 23152 26472
rect 23492 26472 23848 26500
rect 23109 26435 23167 26441
rect 23109 26432 23121 26435
rect 22204 26404 23121 26432
rect 21008 26373 21036 26404
rect 23109 26401 23121 26404
rect 23155 26401 23167 26435
rect 23109 26395 23167 26401
rect 20625 26367 20683 26373
rect 20625 26333 20637 26367
rect 20671 26333 20683 26367
rect 20625 26327 20683 26333
rect 20717 26367 20775 26373
rect 20717 26333 20729 26367
rect 20763 26333 20775 26367
rect 20717 26327 20775 26333
rect 20901 26367 20959 26373
rect 20901 26333 20913 26367
rect 20947 26333 20959 26367
rect 20901 26327 20959 26333
rect 20993 26367 21051 26373
rect 20993 26333 21005 26367
rect 21039 26333 21051 26367
rect 20993 26327 21051 26333
rect 19536 26268 20116 26296
rect 20346 26256 20352 26308
rect 20404 26256 20410 26308
rect 20732 26296 20760 26327
rect 21174 26324 21180 26376
rect 21232 26324 21238 26376
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26364 22155 26367
rect 22278 26364 22284 26376
rect 22143 26336 22284 26364
rect 22143 26333 22155 26336
rect 22097 26327 22155 26333
rect 22278 26324 22284 26336
rect 22336 26324 22342 26376
rect 22833 26367 22891 26373
rect 22833 26333 22845 26367
rect 22879 26333 22891 26367
rect 22833 26327 22891 26333
rect 22925 26367 22983 26373
rect 22925 26333 22937 26367
rect 22971 26364 22983 26367
rect 23492 26364 23520 26472
rect 23842 26460 23848 26472
rect 23900 26500 23906 26512
rect 24670 26500 24676 26512
rect 23900 26472 24676 26500
rect 23900 26460 23906 26472
rect 24670 26460 24676 26472
rect 24728 26460 24734 26512
rect 23566 26392 23572 26444
rect 23624 26432 23630 26444
rect 25424 26432 25452 26540
rect 25682 26528 25688 26540
rect 25740 26528 25746 26580
rect 25866 26528 25872 26580
rect 25924 26528 25930 26580
rect 27338 26528 27344 26580
rect 27396 26528 27402 26580
rect 27430 26528 27436 26580
rect 27488 26568 27494 26580
rect 28994 26568 29000 26580
rect 27488 26540 29000 26568
rect 27488 26528 27494 26540
rect 28994 26528 29000 26540
rect 29052 26528 29058 26580
rect 32122 26528 32128 26580
rect 32180 26528 32186 26580
rect 33134 26528 33140 26580
rect 33192 26528 33198 26580
rect 35529 26571 35587 26577
rect 35529 26568 35541 26571
rect 34716 26540 35541 26568
rect 23624 26404 24348 26432
rect 23624 26392 23630 26404
rect 22971 26336 23520 26364
rect 22971 26333 22983 26336
rect 22925 26327 22983 26333
rect 21192 26296 21220 26324
rect 20732 26268 21220 26296
rect 19116 26200 19278 26228
rect 19116 26188 19122 26200
rect 19334 26188 19340 26240
rect 19392 26228 19398 26240
rect 19978 26228 19984 26240
rect 19392 26200 19984 26228
rect 19392 26188 19398 26200
rect 19978 26188 19984 26200
rect 20036 26188 20042 26240
rect 20438 26188 20444 26240
rect 20496 26188 20502 26240
rect 22848 26228 22876 26327
rect 24320 26296 24348 26404
rect 24596 26404 25452 26432
rect 24596 26373 24624 26404
rect 25498 26392 25504 26444
rect 25556 26432 25562 26444
rect 25593 26435 25651 26441
rect 25593 26432 25605 26435
rect 25556 26404 25605 26432
rect 25556 26392 25562 26404
rect 25593 26401 25605 26404
rect 25639 26401 25651 26435
rect 25884 26432 25912 26528
rect 25958 26460 25964 26512
rect 26016 26500 26022 26512
rect 26016 26472 26464 26500
rect 26016 26460 26022 26472
rect 26436 26432 26464 26472
rect 26510 26460 26516 26512
rect 26568 26460 26574 26512
rect 25884 26404 26081 26432
rect 25593 26395 25651 26401
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 24946 26324 24952 26376
rect 25004 26324 25010 26376
rect 25409 26367 25467 26373
rect 25409 26333 25421 26367
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 25424 26296 25452 26327
rect 25774 26324 25780 26376
rect 25832 26324 25838 26376
rect 25866 26324 25872 26376
rect 25924 26324 25930 26376
rect 26053 26373 26081 26404
rect 26436 26404 27108 26432
rect 26038 26367 26096 26373
rect 26038 26333 26050 26367
rect 26084 26333 26096 26367
rect 26038 26327 26096 26333
rect 26142 26324 26148 26376
rect 26200 26324 26206 26376
rect 26436 26373 26464 26404
rect 27080 26376 27108 26404
rect 26421 26367 26479 26373
rect 26421 26333 26433 26367
rect 26467 26333 26479 26367
rect 26421 26327 26479 26333
rect 26510 26324 26516 26376
rect 26568 26364 26574 26376
rect 26605 26367 26663 26373
rect 26605 26364 26617 26367
rect 26568 26336 26617 26364
rect 26568 26324 26574 26336
rect 26605 26333 26617 26336
rect 26651 26333 26663 26367
rect 26605 26327 26663 26333
rect 26697 26367 26755 26373
rect 26697 26333 26709 26367
rect 26743 26364 26755 26367
rect 26970 26364 26976 26376
rect 26743 26336 26976 26364
rect 26743 26333 26755 26336
rect 26697 26327 26755 26333
rect 26970 26324 26976 26336
rect 27028 26324 27034 26376
rect 27062 26324 27068 26376
rect 27120 26324 27126 26376
rect 27356 26296 27384 26528
rect 28166 26460 28172 26512
rect 28224 26500 28230 26512
rect 31754 26500 31760 26512
rect 28224 26472 31760 26500
rect 28224 26460 28230 26472
rect 31754 26460 31760 26472
rect 31812 26460 31818 26512
rect 30466 26392 30472 26444
rect 30524 26392 30530 26444
rect 32140 26432 32168 26528
rect 32490 26460 32496 26512
rect 32548 26460 32554 26512
rect 33226 26460 33232 26512
rect 33284 26460 33290 26512
rect 32508 26432 32536 26460
rect 32140 26404 32444 26432
rect 32508 26404 33548 26432
rect 30484 26296 30512 26392
rect 32125 26367 32183 26373
rect 32125 26364 32137 26367
rect 24320 26268 27384 26296
rect 27448 26268 30512 26296
rect 31726 26336 32137 26364
rect 24302 26228 24308 26240
rect 22848 26200 24308 26228
rect 24302 26188 24308 26200
rect 24360 26188 24366 26240
rect 24486 26188 24492 26240
rect 24544 26188 24550 26240
rect 26237 26231 26295 26237
rect 26237 26197 26249 26231
rect 26283 26228 26295 26231
rect 26418 26228 26424 26240
rect 26283 26200 26424 26228
rect 26283 26197 26295 26200
rect 26237 26191 26295 26197
rect 26418 26188 26424 26200
rect 26476 26188 26482 26240
rect 26602 26188 26608 26240
rect 26660 26228 26666 26240
rect 27448 26228 27476 26268
rect 26660 26200 27476 26228
rect 26660 26188 26666 26200
rect 28350 26188 28356 26240
rect 28408 26228 28414 26240
rect 31726 26228 31754 26336
rect 32125 26333 32137 26336
rect 32171 26364 32183 26367
rect 32214 26364 32220 26376
rect 32171 26336 32220 26364
rect 32171 26333 32183 26336
rect 32125 26327 32183 26333
rect 32214 26324 32220 26336
rect 32272 26324 32278 26376
rect 32416 26364 32444 26404
rect 33520 26373 33548 26404
rect 32493 26367 32551 26373
rect 32493 26364 32505 26367
rect 32416 26336 32505 26364
rect 32493 26333 32505 26336
rect 32539 26364 32551 26367
rect 33413 26367 33471 26373
rect 33413 26364 33425 26367
rect 32539 26336 33425 26364
rect 32539 26333 32551 26336
rect 32493 26327 32551 26333
rect 33413 26333 33425 26336
rect 33459 26333 33471 26367
rect 33413 26327 33471 26333
rect 33505 26367 33563 26373
rect 33505 26333 33517 26367
rect 33551 26333 33563 26367
rect 33505 26327 33563 26333
rect 34606 26324 34612 26376
rect 34664 26364 34670 26376
rect 34716 26373 34744 26540
rect 35529 26537 35541 26540
rect 35575 26537 35587 26571
rect 35529 26531 35587 26537
rect 39666 26432 39672 26444
rect 35452 26404 39672 26432
rect 35452 26373 35480 26404
rect 39666 26392 39672 26404
rect 39724 26392 39730 26444
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 34664 26336 34713 26364
rect 34664 26324 34670 26336
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 34701 26327 34759 26333
rect 35437 26367 35495 26373
rect 35437 26333 35449 26367
rect 35483 26333 35495 26367
rect 35437 26327 35495 26333
rect 35802 26324 35808 26376
rect 35860 26324 35866 26376
rect 35897 26367 35955 26373
rect 35897 26333 35909 26367
rect 35943 26333 35955 26367
rect 35897 26327 35955 26333
rect 31938 26256 31944 26308
rect 31996 26296 32002 26308
rect 32309 26299 32367 26305
rect 32309 26296 32321 26299
rect 31996 26268 32321 26296
rect 31996 26256 32002 26268
rect 32309 26265 32321 26268
rect 32355 26265 32367 26299
rect 32309 26259 32367 26265
rect 28408 26200 31754 26228
rect 32324 26228 32352 26259
rect 32398 26256 32404 26308
rect 32456 26256 32462 26308
rect 32769 26299 32827 26305
rect 32769 26296 32781 26299
rect 32508 26268 32781 26296
rect 32508 26228 32536 26268
rect 32769 26265 32781 26268
rect 32815 26265 32827 26299
rect 32769 26259 32827 26265
rect 32961 26299 33019 26305
rect 32961 26265 32973 26299
rect 33007 26296 33019 26299
rect 33229 26299 33287 26305
rect 33007 26268 33088 26296
rect 33007 26265 33019 26268
rect 32961 26259 33019 26265
rect 32324 26200 32536 26228
rect 28408 26188 28414 26200
rect 32674 26188 32680 26240
rect 32732 26188 32738 26240
rect 33060 26228 33088 26268
rect 33229 26265 33241 26299
rect 33275 26296 33287 26299
rect 35345 26299 35403 26305
rect 35345 26296 35357 26299
rect 33275 26268 35357 26296
rect 33275 26265 33287 26268
rect 33229 26259 33287 26265
rect 35345 26265 35357 26268
rect 35391 26265 35403 26299
rect 35345 26259 35403 26265
rect 33318 26228 33324 26240
rect 33060 26200 33324 26228
rect 33318 26188 33324 26200
rect 33376 26188 33382 26240
rect 34330 26188 34336 26240
rect 34388 26228 34394 26240
rect 35912 26228 35940 26327
rect 34388 26200 35940 26228
rect 34388 26188 34394 26200
rect 36078 26188 36084 26240
rect 36136 26188 36142 26240
rect 1104 26138 41400 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 41400 26138
rect 1104 26064 41400 26086
rect 5074 26024 5080 26036
rect 4724 25996 5080 26024
rect 4724 25965 4752 25996
rect 5074 25984 5080 25996
rect 5132 25984 5138 26036
rect 6914 25984 6920 26036
rect 6972 25984 6978 26036
rect 8389 26027 8447 26033
rect 8389 25993 8401 26027
rect 8435 26024 8447 26027
rect 8478 26024 8484 26036
rect 8435 25996 8484 26024
rect 8435 25993 8447 25996
rect 8389 25987 8447 25993
rect 8478 25984 8484 25996
rect 8536 25984 8542 26036
rect 8754 25984 8760 26036
rect 8812 25984 8818 26036
rect 9416 25996 10318 26024
rect 4709 25959 4767 25965
rect 4709 25925 4721 25959
rect 4755 25925 4767 25959
rect 4709 25919 4767 25925
rect 5442 25916 5448 25968
rect 5500 25916 5506 25968
rect 6932 25888 6960 25984
rect 8018 25916 8024 25968
rect 8076 25956 8082 25968
rect 8772 25956 8800 25984
rect 8076 25928 9076 25956
rect 8076 25916 8082 25928
rect 7193 25891 7251 25897
rect 7193 25888 7205 25891
rect 6932 25860 7205 25888
rect 7193 25857 7205 25860
rect 7239 25857 7251 25891
rect 7193 25851 7251 25857
rect 8113 25891 8171 25897
rect 8113 25857 8125 25891
rect 8159 25888 8171 25891
rect 8570 25888 8576 25900
rect 8159 25860 8576 25888
rect 8159 25857 8171 25860
rect 8113 25851 8171 25857
rect 8570 25848 8576 25860
rect 8628 25848 8634 25900
rect 8754 25848 8760 25900
rect 8812 25848 8818 25900
rect 8846 25848 8852 25900
rect 8904 25848 8910 25900
rect 3786 25780 3792 25832
rect 3844 25820 3850 25832
rect 4433 25823 4491 25829
rect 4433 25820 4445 25823
rect 3844 25792 4445 25820
rect 3844 25780 3850 25792
rect 4433 25789 4445 25792
rect 4479 25789 4491 25823
rect 4433 25783 4491 25789
rect 6181 25823 6239 25829
rect 6181 25789 6193 25823
rect 6227 25820 6239 25823
rect 6457 25823 6515 25829
rect 6457 25820 6469 25823
rect 6227 25792 6469 25820
rect 6227 25789 6239 25792
rect 6181 25783 6239 25789
rect 6457 25789 6469 25792
rect 6503 25789 6515 25823
rect 6457 25783 6515 25789
rect 6546 25780 6552 25832
rect 6604 25820 6610 25832
rect 9048 25829 9076 25928
rect 9416 25900 9444 25996
rect 9674 25916 9680 25968
rect 9732 25956 9738 25968
rect 9732 25928 9812 25956
rect 9732 25916 9738 25928
rect 9398 25848 9404 25900
rect 9456 25848 9462 25900
rect 9784 25897 9812 25928
rect 10042 25916 10048 25968
rect 10100 25916 10106 25968
rect 9950 25897 9956 25900
rect 9769 25891 9827 25897
rect 9769 25857 9781 25891
rect 9815 25857 9827 25891
rect 9917 25891 9956 25897
rect 9917 25888 9929 25891
rect 9863 25860 9929 25888
rect 9769 25851 9827 25857
rect 9917 25857 9929 25860
rect 9917 25851 9956 25857
rect 9950 25848 9956 25851
rect 10008 25848 10014 25900
rect 10290 25897 10318 25996
rect 11054 25984 11060 26036
rect 11112 25984 11118 26036
rect 11149 26027 11207 26033
rect 11149 25993 11161 26027
rect 11195 26024 11207 26027
rect 11422 26024 11428 26036
rect 11195 25996 11428 26024
rect 11195 25993 11207 25996
rect 11149 25987 11207 25993
rect 11422 25984 11428 25996
rect 11480 26024 11486 26036
rect 13170 26024 13176 26036
rect 11480 25996 13176 26024
rect 11480 25984 11486 25996
rect 13170 25984 13176 25996
rect 13228 25984 13234 26036
rect 14277 26027 14335 26033
rect 14277 25993 14289 26027
rect 14323 26024 14335 26027
rect 14458 26024 14464 26036
rect 14323 25996 14464 26024
rect 14323 25993 14335 25996
rect 14277 25987 14335 25993
rect 14458 25984 14464 25996
rect 14516 25984 14522 26036
rect 14568 25996 19104 26024
rect 11072 25897 11100 25984
rect 11793 25959 11851 25965
rect 11793 25925 11805 25959
rect 11839 25956 11851 25959
rect 13078 25956 13084 25968
rect 11839 25928 13084 25956
rect 11839 25925 11851 25928
rect 11793 25919 11851 25925
rect 13078 25916 13084 25928
rect 13136 25916 13142 25968
rect 14090 25916 14096 25968
rect 14148 25956 14154 25968
rect 14568 25956 14596 25996
rect 16114 25956 16120 25968
rect 14148 25928 14596 25956
rect 15580 25928 16120 25956
rect 14148 25916 14154 25928
rect 15580 25900 15608 25928
rect 16114 25916 16120 25928
rect 16172 25916 16178 25968
rect 16868 25928 17264 25956
rect 16868 25900 16896 25928
rect 10137 25891 10195 25897
rect 10137 25857 10149 25891
rect 10183 25857 10195 25891
rect 10137 25851 10195 25857
rect 10275 25891 10333 25897
rect 10275 25857 10287 25891
rect 10321 25857 10333 25891
rect 10275 25851 10333 25857
rect 11057 25891 11115 25897
rect 11057 25857 11069 25891
rect 11103 25857 11115 25891
rect 11057 25851 11115 25857
rect 7101 25823 7159 25829
rect 7101 25820 7113 25823
rect 6604 25792 7113 25820
rect 6604 25780 6610 25792
rect 7101 25789 7113 25792
rect 7147 25789 7159 25823
rect 7101 25783 7159 25789
rect 9033 25823 9091 25829
rect 9033 25789 9045 25823
rect 9079 25820 9091 25823
rect 9582 25820 9588 25832
rect 9079 25792 9588 25820
rect 9079 25789 9091 25792
rect 9033 25783 9091 25789
rect 9582 25780 9588 25792
rect 9640 25780 9646 25832
rect 9677 25823 9735 25829
rect 9677 25789 9689 25823
rect 9723 25820 9735 25823
rect 9968 25820 9996 25848
rect 9723 25792 9996 25820
rect 9723 25789 9735 25792
rect 9677 25783 9735 25789
rect 9950 25752 9956 25764
rect 8956 25724 9956 25752
rect 7282 25644 7288 25696
rect 7340 25644 7346 25696
rect 8956 25693 8984 25724
rect 9950 25712 9956 25724
rect 10008 25712 10014 25764
rect 8941 25687 8999 25693
rect 8941 25653 8953 25687
rect 8987 25653 8999 25687
rect 8941 25647 8999 25653
rect 9214 25644 9220 25696
rect 9272 25644 9278 25696
rect 9306 25644 9312 25696
rect 9364 25684 9370 25696
rect 9582 25684 9588 25696
rect 9364 25656 9588 25684
rect 9364 25644 9370 25656
rect 9582 25644 9588 25656
rect 9640 25684 9646 25696
rect 10152 25684 10180 25851
rect 10290 25820 10318 25851
rect 11146 25848 11152 25900
rect 11204 25848 11210 25900
rect 12805 25891 12863 25897
rect 12805 25857 12817 25891
rect 12851 25888 12863 25891
rect 12986 25888 12992 25900
rect 12851 25860 12992 25888
rect 12851 25857 12863 25860
rect 12805 25851 12863 25857
rect 12986 25848 12992 25860
rect 13044 25848 13050 25900
rect 13538 25848 13544 25900
rect 13596 25888 13602 25900
rect 14461 25891 14519 25897
rect 14461 25888 14473 25891
rect 13596 25860 14473 25888
rect 13596 25848 13602 25860
rect 14461 25857 14473 25860
rect 14507 25888 14519 25891
rect 14918 25888 14924 25900
rect 14507 25860 14924 25888
rect 14507 25857 14519 25860
rect 14461 25851 14519 25857
rect 14918 25848 14924 25860
rect 14976 25888 14982 25900
rect 15562 25888 15568 25900
rect 14976 25860 15568 25888
rect 14976 25848 14982 25860
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 15654 25848 15660 25900
rect 15712 25888 15718 25900
rect 15712 25860 16574 25888
rect 15712 25848 15718 25860
rect 11164 25820 11192 25848
rect 10290 25792 11192 25820
rect 11238 25780 11244 25832
rect 11296 25820 11302 25832
rect 12621 25823 12679 25829
rect 12621 25820 12633 25823
rect 11296 25792 12633 25820
rect 11296 25780 11302 25792
rect 12621 25789 12633 25792
rect 12667 25820 12679 25823
rect 12710 25820 12716 25832
rect 12667 25792 12716 25820
rect 12667 25789 12679 25792
rect 12621 25783 12679 25789
rect 12710 25780 12716 25792
rect 12768 25780 12774 25832
rect 12894 25780 12900 25832
rect 12952 25820 12958 25832
rect 13081 25823 13139 25829
rect 13081 25820 13093 25823
rect 12952 25792 13093 25820
rect 12952 25780 12958 25792
rect 13081 25789 13093 25792
rect 13127 25820 13139 25823
rect 13262 25820 13268 25832
rect 13127 25792 13268 25820
rect 13127 25789 13139 25792
rect 13081 25783 13139 25789
rect 13262 25780 13268 25792
rect 13320 25820 13326 25832
rect 14550 25820 14556 25832
rect 13320 25792 14556 25820
rect 13320 25780 13326 25792
rect 14550 25780 14556 25792
rect 14608 25780 14614 25832
rect 14737 25823 14795 25829
rect 14737 25789 14749 25823
rect 14783 25820 14795 25823
rect 15102 25820 15108 25832
rect 14783 25792 15108 25820
rect 14783 25789 14795 25792
rect 14737 25783 14795 25789
rect 15102 25780 15108 25792
rect 15160 25820 15166 25832
rect 15838 25820 15844 25832
rect 15160 25792 15844 25820
rect 15160 25780 15166 25792
rect 15838 25780 15844 25792
rect 15896 25780 15902 25832
rect 16546 25820 16574 25860
rect 16850 25848 16856 25900
rect 16908 25848 16914 25900
rect 17034 25848 17040 25900
rect 17092 25848 17098 25900
rect 17236 25897 17264 25928
rect 17310 25916 17316 25968
rect 17368 25916 17374 25968
rect 18874 25956 18880 25968
rect 17880 25928 18880 25956
rect 17314 25913 17372 25916
rect 17221 25891 17279 25897
rect 17221 25857 17233 25891
rect 17267 25857 17279 25891
rect 17314 25879 17326 25913
rect 17360 25879 17372 25913
rect 17314 25873 17372 25879
rect 17439 25891 17497 25897
rect 17221 25851 17279 25857
rect 17439 25857 17451 25891
rect 17485 25888 17497 25891
rect 17880 25888 17908 25928
rect 18874 25916 18880 25928
rect 18932 25916 18938 25968
rect 19076 25965 19104 25996
rect 19886 25984 19892 26036
rect 19944 26024 19950 26036
rect 21542 26024 21548 26036
rect 19944 25996 21548 26024
rect 19944 25984 19950 25996
rect 21542 25984 21548 25996
rect 21600 25984 21606 26036
rect 27338 26024 27344 26036
rect 24688 25996 27344 26024
rect 19061 25959 19119 25965
rect 19061 25925 19073 25959
rect 19107 25925 19119 25959
rect 20438 25956 20444 25968
rect 19061 25919 19119 25925
rect 19812 25928 20444 25956
rect 17485 25860 17908 25888
rect 17485 25857 17497 25860
rect 17439 25851 17497 25857
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18322 25888 18328 25900
rect 18012 25860 18328 25888
rect 18012 25848 18018 25860
rect 18322 25848 18328 25860
rect 18380 25848 18386 25900
rect 19812 25897 19840 25928
rect 20438 25916 20444 25928
rect 20496 25916 20502 25968
rect 20530 25916 20536 25968
rect 20588 25916 20594 25968
rect 24688 25956 24716 25996
rect 20732 25928 24716 25956
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25888 18567 25891
rect 19797 25891 19855 25897
rect 18555 25860 19748 25888
rect 18555 25857 18567 25860
rect 18509 25851 18567 25857
rect 17586 25820 17592 25832
rect 16546 25792 17592 25820
rect 17586 25780 17592 25792
rect 17644 25780 17650 25832
rect 17862 25780 17868 25832
rect 17920 25820 17926 25832
rect 18233 25823 18291 25829
rect 18233 25820 18245 25823
rect 17920 25792 18245 25820
rect 17920 25780 17926 25792
rect 18233 25789 18245 25792
rect 18279 25789 18291 25823
rect 18233 25783 18291 25789
rect 18417 25823 18475 25829
rect 18417 25789 18429 25823
rect 18463 25789 18475 25823
rect 18417 25783 18475 25789
rect 12158 25712 12164 25764
rect 12216 25752 12222 25764
rect 17034 25752 17040 25764
rect 12216 25724 17040 25752
rect 12216 25712 12222 25724
rect 17034 25712 17040 25724
rect 17092 25712 17098 25764
rect 17310 25712 17316 25764
rect 17368 25752 17374 25764
rect 17681 25755 17739 25761
rect 17681 25752 17693 25755
rect 17368 25724 17693 25752
rect 17368 25712 17374 25724
rect 17681 25721 17693 25724
rect 17727 25721 17739 25755
rect 18432 25752 18460 25783
rect 19334 25780 19340 25832
rect 19392 25820 19398 25832
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 19392 25792 19625 25820
rect 19392 25780 19398 25792
rect 19613 25789 19625 25792
rect 19659 25789 19671 25823
rect 19720 25820 19748 25860
rect 19797 25857 19809 25891
rect 19843 25857 19855 25891
rect 19797 25851 19855 25857
rect 19978 25848 19984 25900
rect 20036 25848 20042 25900
rect 20073 25891 20131 25897
rect 20073 25857 20085 25891
rect 20119 25888 20131 25891
rect 20548 25888 20576 25916
rect 20732 25900 20760 25928
rect 25038 25916 25044 25968
rect 25096 25956 25102 25968
rect 25133 25959 25191 25965
rect 25133 25956 25145 25959
rect 25096 25928 25145 25956
rect 25096 25916 25102 25928
rect 25133 25925 25145 25928
rect 25179 25925 25191 25959
rect 25133 25919 25191 25925
rect 20119 25860 20576 25888
rect 20119 25857 20131 25860
rect 20073 25851 20131 25857
rect 20622 25848 20628 25900
rect 20680 25848 20686 25900
rect 20714 25848 20720 25900
rect 20772 25848 20778 25900
rect 20898 25848 20904 25900
rect 20956 25888 20962 25900
rect 21726 25888 21732 25900
rect 20956 25860 21732 25888
rect 20956 25848 20962 25860
rect 21726 25848 21732 25860
rect 21784 25848 21790 25900
rect 24578 25848 24584 25900
rect 24636 25888 24642 25900
rect 25240 25897 25268 25996
rect 27338 25984 27344 25996
rect 27396 25984 27402 26036
rect 27985 26027 28043 26033
rect 27985 26024 27997 26027
rect 27448 25996 27997 26024
rect 26050 25956 26056 25968
rect 25884 25928 26056 25956
rect 25884 25900 25912 25928
rect 26050 25916 26056 25928
rect 26108 25956 26114 25968
rect 26970 25956 26976 25968
rect 26108 25928 26976 25956
rect 26108 25916 26114 25928
rect 26970 25916 26976 25928
rect 27028 25916 27034 25968
rect 24857 25891 24915 25897
rect 24857 25888 24869 25891
rect 24636 25860 24869 25888
rect 24636 25848 24642 25860
rect 24857 25857 24869 25860
rect 24903 25857 24915 25891
rect 24857 25851 24915 25857
rect 24950 25891 25008 25897
rect 24950 25857 24962 25891
rect 24996 25857 25008 25891
rect 24950 25851 25008 25857
rect 25225 25891 25283 25897
rect 25225 25857 25237 25891
rect 25271 25857 25283 25891
rect 25225 25851 25283 25857
rect 20640 25820 20668 25848
rect 19720 25792 20668 25820
rect 19613 25783 19671 25789
rect 21358 25780 21364 25832
rect 21416 25820 21422 25832
rect 24596 25820 24624 25848
rect 21416 25792 24624 25820
rect 24964 25820 24992 25851
rect 25314 25848 25320 25900
rect 25372 25897 25378 25900
rect 25372 25888 25380 25897
rect 25866 25888 25872 25900
rect 25372 25860 25417 25888
rect 25608 25860 25872 25888
rect 25372 25851 25380 25860
rect 25372 25848 25378 25851
rect 25608 25820 25636 25860
rect 25866 25848 25872 25860
rect 25924 25848 25930 25900
rect 26326 25848 26332 25900
rect 26384 25848 26390 25900
rect 26418 25848 26424 25900
rect 26476 25848 26482 25900
rect 26605 25891 26663 25897
rect 26605 25857 26617 25891
rect 26651 25857 26663 25891
rect 26605 25851 26663 25857
rect 24964 25792 25636 25820
rect 21416 25780 21422 25792
rect 17681 25715 17739 25721
rect 17972 25724 20392 25752
rect 9640 25656 10180 25684
rect 9640 25644 9646 25656
rect 10410 25644 10416 25696
rect 10468 25644 10474 25696
rect 10870 25644 10876 25696
rect 10928 25684 10934 25696
rect 12434 25684 12440 25696
rect 10928 25656 12440 25684
rect 10928 25644 10934 25656
rect 12434 25644 12440 25656
rect 12492 25644 12498 25696
rect 12894 25644 12900 25696
rect 12952 25644 12958 25696
rect 12986 25644 12992 25696
rect 13044 25644 13050 25696
rect 14366 25644 14372 25696
rect 14424 25684 14430 25696
rect 14645 25687 14703 25693
rect 14645 25684 14657 25687
rect 14424 25656 14657 25684
rect 14424 25644 14430 25656
rect 14645 25653 14657 25656
rect 14691 25653 14703 25687
rect 14645 25647 14703 25653
rect 14918 25644 14924 25696
rect 14976 25684 14982 25696
rect 17972 25684 18000 25724
rect 14976 25656 18000 25684
rect 14976 25644 14982 25656
rect 18046 25644 18052 25696
rect 18104 25644 18110 25696
rect 20364 25684 20392 25724
rect 20438 25712 20444 25764
rect 20496 25752 20502 25764
rect 22738 25752 22744 25764
rect 20496 25724 22744 25752
rect 20496 25712 20502 25724
rect 22738 25712 22744 25724
rect 22796 25712 22802 25764
rect 24964 25752 24992 25792
rect 25682 25780 25688 25832
rect 25740 25780 25746 25832
rect 26142 25780 26148 25832
rect 26200 25780 26206 25832
rect 24596 25724 24992 25752
rect 24596 25696 24624 25724
rect 25498 25712 25504 25764
rect 25556 25752 25562 25764
rect 26620 25752 26648 25851
rect 26694 25848 26700 25900
rect 26752 25848 26758 25900
rect 27448 25897 27476 25996
rect 27985 25993 27997 25996
rect 28031 26024 28043 26027
rect 28553 26027 28611 26033
rect 28553 26024 28565 26027
rect 28031 25996 28565 26024
rect 28031 25993 28043 25996
rect 27985 25987 28043 25993
rect 28553 25993 28565 25996
rect 28599 25993 28611 26027
rect 28553 25987 28611 25993
rect 31297 26027 31355 26033
rect 31297 25993 31309 26027
rect 31343 26024 31355 26027
rect 31662 26024 31668 26036
rect 31343 25996 31668 26024
rect 31343 25993 31355 25996
rect 31297 25987 31355 25993
rect 27614 25916 27620 25968
rect 27672 25956 27678 25968
rect 28353 25959 28411 25965
rect 28353 25956 28365 25959
rect 27672 25928 28365 25956
rect 27672 25916 27678 25928
rect 28353 25925 28365 25928
rect 28399 25925 28411 25959
rect 30745 25959 30803 25965
rect 30745 25956 30757 25959
rect 28353 25919 28411 25925
rect 30392 25928 30757 25956
rect 30392 25900 30420 25928
rect 30745 25925 30757 25928
rect 30791 25925 30803 25959
rect 30745 25919 30803 25925
rect 27433 25891 27491 25897
rect 27433 25888 27445 25891
rect 26988 25860 27445 25888
rect 25556 25724 26648 25752
rect 26712 25752 26740 25848
rect 26988 25832 27016 25860
rect 27433 25857 27445 25860
rect 27479 25857 27491 25891
rect 27433 25851 27491 25857
rect 27522 25848 27528 25900
rect 27580 25848 27586 25900
rect 27893 25891 27951 25897
rect 27893 25857 27905 25891
rect 27939 25857 27951 25891
rect 27893 25851 27951 25857
rect 26970 25780 26976 25832
rect 27028 25780 27034 25832
rect 27338 25780 27344 25832
rect 27396 25780 27402 25832
rect 27617 25823 27675 25829
rect 27617 25789 27629 25823
rect 27663 25820 27675 25823
rect 27798 25820 27804 25832
rect 27663 25792 27804 25820
rect 27663 25789 27675 25792
rect 27617 25783 27675 25789
rect 27798 25780 27804 25792
rect 27856 25780 27862 25832
rect 27908 25752 27936 25851
rect 30374 25848 30380 25900
rect 30432 25848 30438 25900
rect 30558 25848 30564 25900
rect 30616 25848 30622 25900
rect 30926 25848 30932 25900
rect 30984 25848 30990 25900
rect 31496 25888 31524 25996
rect 31662 25984 31668 25996
rect 31720 25984 31726 26036
rect 31938 25984 31944 26036
rect 31996 25984 32002 26036
rect 32490 25984 32496 26036
rect 32548 26024 32554 26036
rect 32953 26027 33011 26033
rect 32953 26024 32965 26027
rect 32548 25996 32965 26024
rect 32548 25984 32554 25996
rect 32953 25993 32965 25996
rect 32999 25993 33011 26027
rect 34882 26024 34888 26036
rect 32953 25987 33011 25993
rect 33336 25996 34888 26024
rect 33336 25956 33364 25996
rect 34882 25984 34888 25996
rect 34940 25984 34946 26036
rect 35437 26027 35495 26033
rect 35437 25993 35449 26027
rect 35483 26024 35495 26027
rect 36078 26024 36084 26036
rect 35483 25996 36084 26024
rect 35483 25993 35495 25996
rect 35437 25987 35495 25993
rect 36078 25984 36084 25996
rect 36136 25984 36142 26036
rect 32508 25928 33364 25956
rect 33413 25959 33471 25965
rect 32508 25897 32536 25928
rect 33413 25925 33425 25959
rect 33459 25956 33471 25959
rect 33873 25959 33931 25965
rect 33873 25956 33885 25959
rect 33459 25928 33885 25956
rect 33459 25925 33471 25928
rect 33413 25919 33471 25925
rect 33873 25925 33885 25928
rect 33919 25925 33931 25959
rect 36262 25956 36268 25968
rect 35098 25928 36268 25956
rect 33873 25919 33931 25925
rect 36262 25916 36268 25928
rect 36320 25916 36326 25968
rect 31573 25891 31631 25897
rect 31573 25888 31585 25891
rect 31496 25860 31585 25888
rect 31573 25857 31585 25860
rect 31619 25857 31631 25891
rect 32493 25891 32551 25897
rect 32493 25888 32505 25891
rect 31573 25851 31631 25857
rect 31772 25860 32505 25888
rect 31772 25832 31800 25860
rect 32493 25857 32505 25860
rect 32539 25857 32551 25891
rect 32493 25851 32551 25857
rect 32769 25891 32827 25897
rect 32769 25857 32781 25891
rect 32815 25888 32827 25891
rect 32815 25860 32904 25888
rect 32815 25857 32827 25860
rect 32769 25851 32827 25857
rect 29546 25780 29552 25832
rect 29604 25820 29610 25832
rect 31665 25823 31723 25829
rect 31665 25820 31677 25823
rect 29604 25792 31677 25820
rect 29604 25780 29610 25792
rect 31665 25789 31677 25792
rect 31711 25789 31723 25823
rect 31665 25783 31723 25789
rect 31754 25780 31760 25832
rect 31812 25780 31818 25832
rect 31938 25780 31944 25832
rect 31996 25820 32002 25832
rect 32876 25820 32904 25860
rect 33226 25848 33232 25900
rect 33284 25888 33290 25900
rect 33321 25891 33379 25897
rect 33321 25888 33333 25891
rect 33284 25860 33333 25888
rect 33284 25848 33290 25860
rect 33321 25857 33333 25860
rect 33367 25857 33379 25891
rect 33321 25851 33379 25857
rect 33502 25848 33508 25900
rect 33560 25848 33566 25900
rect 35526 25848 35532 25900
rect 35584 25848 35590 25900
rect 35805 25891 35863 25897
rect 35805 25857 35817 25891
rect 35851 25888 35863 25891
rect 36817 25891 36875 25897
rect 36817 25888 36829 25891
rect 35851 25860 36829 25888
rect 35851 25857 35863 25860
rect 35805 25851 35863 25857
rect 36817 25857 36829 25860
rect 36863 25857 36875 25891
rect 36817 25851 36875 25857
rect 31996 25792 32904 25820
rect 31996 25780 32002 25792
rect 26712 25724 27936 25752
rect 28552 25724 30052 25752
rect 25556 25712 25562 25724
rect 20898 25684 20904 25696
rect 20364 25656 20904 25684
rect 20898 25644 20904 25656
rect 20956 25644 20962 25696
rect 24578 25644 24584 25696
rect 24636 25644 24642 25696
rect 27154 25644 27160 25696
rect 27212 25644 27218 25696
rect 28166 25644 28172 25696
rect 28224 25684 28230 25696
rect 28552 25693 28580 25724
rect 28537 25687 28595 25693
rect 28537 25684 28549 25687
rect 28224 25656 28549 25684
rect 28224 25644 28230 25656
rect 28537 25653 28549 25656
rect 28583 25653 28595 25687
rect 28537 25647 28595 25653
rect 28718 25644 28724 25696
rect 28776 25644 28782 25696
rect 30024 25684 30052 25724
rect 32398 25712 32404 25764
rect 32456 25752 32462 25764
rect 32585 25755 32643 25761
rect 32585 25752 32597 25755
rect 32456 25724 32597 25752
rect 32456 25712 32462 25724
rect 32585 25721 32597 25724
rect 32631 25721 32643 25755
rect 32876 25752 32904 25792
rect 33597 25823 33655 25829
rect 33597 25789 33609 25823
rect 33643 25820 33655 25823
rect 34422 25820 34428 25832
rect 33643 25792 34428 25820
rect 33643 25789 33655 25792
rect 33597 25783 33655 25789
rect 34422 25780 34428 25792
rect 34480 25780 34486 25832
rect 35544 25820 35572 25848
rect 35897 25823 35955 25829
rect 35897 25820 35909 25823
rect 35544 25792 35909 25820
rect 35897 25789 35909 25792
rect 35943 25789 35955 25823
rect 35897 25783 35955 25789
rect 36173 25823 36231 25829
rect 36173 25789 36185 25823
rect 36219 25789 36231 25823
rect 36173 25783 36231 25789
rect 33318 25752 33324 25764
rect 32876 25724 33324 25752
rect 32585 25715 32643 25721
rect 33318 25712 33324 25724
rect 33376 25712 33382 25764
rect 34882 25712 34888 25764
rect 34940 25752 34946 25764
rect 35802 25752 35808 25764
rect 34940 25724 35808 25752
rect 34940 25712 34946 25724
rect 35802 25712 35808 25724
rect 35860 25752 35866 25764
rect 36188 25752 36216 25783
rect 36814 25752 36820 25764
rect 35860 25724 36820 25752
rect 35860 25712 35866 25724
rect 36814 25712 36820 25724
rect 36872 25712 36878 25764
rect 31573 25687 31631 25693
rect 31573 25684 31585 25687
rect 30024 25656 31585 25684
rect 31573 25653 31585 25656
rect 31619 25684 31631 25687
rect 34606 25684 34612 25696
rect 31619 25656 34612 25684
rect 31619 25653 31631 25656
rect 31573 25647 31631 25653
rect 34606 25644 34612 25656
rect 34664 25684 34670 25696
rect 35345 25687 35403 25693
rect 35345 25684 35357 25687
rect 34664 25656 35357 25684
rect 34664 25644 34670 25656
rect 35345 25653 35357 25656
rect 35391 25653 35403 25687
rect 35345 25647 35403 25653
rect 36078 25644 36084 25696
rect 36136 25644 36142 25696
rect 1104 25594 41400 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 41400 25594
rect 1104 25520 41400 25542
rect 4706 25440 4712 25492
rect 4764 25480 4770 25492
rect 5537 25483 5595 25489
rect 5537 25480 5549 25483
rect 4764 25452 5549 25480
rect 4764 25440 4770 25452
rect 5537 25449 5549 25452
rect 5583 25449 5595 25483
rect 5537 25443 5595 25449
rect 6546 25440 6552 25492
rect 6604 25440 6610 25492
rect 7282 25440 7288 25492
rect 7340 25440 7346 25492
rect 7760 25452 8708 25480
rect 3786 25304 3792 25356
rect 3844 25304 3850 25356
rect 6564 25344 6592 25440
rect 6641 25347 6699 25353
rect 6641 25344 6653 25347
rect 6564 25316 6653 25344
rect 6641 25313 6653 25316
rect 6687 25313 6699 25347
rect 6641 25307 6699 25313
rect 6733 25347 6791 25353
rect 6733 25313 6745 25347
rect 6779 25344 6791 25347
rect 7300 25344 7328 25440
rect 6779 25316 7328 25344
rect 6779 25313 6791 25316
rect 6733 25307 6791 25313
rect 5442 25276 5448 25288
rect 5198 25248 5448 25276
rect 5442 25236 5448 25248
rect 5500 25236 5506 25288
rect 6549 25279 6607 25285
rect 6549 25245 6561 25279
rect 6595 25245 6607 25279
rect 6549 25239 6607 25245
rect 4062 25168 4068 25220
rect 4120 25168 4126 25220
rect 6564 25208 6592 25239
rect 6822 25236 6828 25288
rect 6880 25236 6886 25288
rect 7760 25208 7788 25452
rect 7837 25415 7895 25421
rect 7837 25381 7849 25415
rect 7883 25381 7895 25415
rect 8680 25412 8708 25452
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 9125 25483 9183 25489
rect 9125 25480 9137 25483
rect 8812 25452 9137 25480
rect 8812 25440 8818 25452
rect 9125 25449 9137 25452
rect 9171 25449 9183 25483
rect 9125 25443 9183 25449
rect 9677 25483 9735 25489
rect 9677 25449 9689 25483
rect 9723 25480 9735 25483
rect 9766 25480 9772 25492
rect 9723 25452 9772 25480
rect 9723 25449 9735 25452
rect 9677 25443 9735 25449
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 14918 25480 14924 25492
rect 14568 25452 14924 25480
rect 9030 25412 9036 25424
rect 8680 25384 9036 25412
rect 7837 25375 7895 25381
rect 7852 25344 7880 25375
rect 9030 25372 9036 25384
rect 9088 25372 9094 25424
rect 9493 25415 9551 25421
rect 9493 25381 9505 25415
rect 9539 25412 9551 25415
rect 9582 25412 9588 25424
rect 9539 25384 9588 25412
rect 9539 25381 9551 25384
rect 9493 25375 9551 25381
rect 9582 25372 9588 25384
rect 9640 25412 9646 25424
rect 9640 25384 11376 25412
rect 9640 25372 9646 25384
rect 8202 25344 8208 25356
rect 7852 25316 8208 25344
rect 8202 25304 8208 25316
rect 8260 25304 8266 25356
rect 9122 25344 9128 25356
rect 8312 25316 9128 25344
rect 7837 25279 7895 25285
rect 7837 25245 7849 25279
rect 7883 25276 7895 25279
rect 8018 25276 8024 25288
rect 7883 25248 8024 25276
rect 7883 25245 7895 25248
rect 7837 25239 7895 25245
rect 8018 25236 8024 25248
rect 8076 25236 8082 25288
rect 8110 25236 8116 25288
rect 8168 25236 8174 25288
rect 8312 25217 8340 25316
rect 8496 25288 8524 25316
rect 9122 25304 9128 25316
rect 9180 25304 9186 25356
rect 9214 25304 9220 25356
rect 9272 25344 9278 25356
rect 9272 25316 9904 25344
rect 9272 25304 9278 25316
rect 8478 25236 8484 25288
rect 8536 25236 8542 25288
rect 8665 25279 8723 25285
rect 8665 25245 8677 25279
rect 8711 25276 8723 25279
rect 9309 25279 9367 25285
rect 8711 25248 9168 25276
rect 8711 25245 8723 25248
rect 8665 25239 8723 25245
rect 6564 25180 7788 25208
rect 8297 25211 8355 25217
rect 8297 25177 8309 25211
rect 8343 25177 8355 25211
rect 8297 25171 8355 25177
rect 8386 25168 8392 25220
rect 8444 25208 8450 25220
rect 8680 25208 8708 25239
rect 8444 25180 8708 25208
rect 8444 25168 8450 25180
rect 9030 25168 9036 25220
rect 9088 25168 9094 25220
rect 6362 25100 6368 25152
rect 6420 25100 6426 25152
rect 8021 25143 8079 25149
rect 8021 25109 8033 25143
rect 8067 25140 8079 25143
rect 9048 25140 9076 25168
rect 8067 25112 9076 25140
rect 9140 25140 9168 25248
rect 9309 25245 9321 25279
rect 9355 25276 9367 25279
rect 9398 25276 9404 25288
rect 9355 25248 9404 25276
rect 9355 25245 9367 25248
rect 9309 25239 9367 25245
rect 9398 25236 9404 25248
rect 9456 25236 9462 25288
rect 9490 25236 9496 25288
rect 9548 25276 9554 25288
rect 9585 25279 9643 25285
rect 9585 25276 9597 25279
rect 9548 25248 9597 25276
rect 9548 25236 9554 25248
rect 9585 25245 9597 25248
rect 9631 25245 9643 25279
rect 9585 25239 9643 25245
rect 9674 25236 9680 25288
rect 9732 25236 9738 25288
rect 9876 25285 9904 25316
rect 9861 25279 9919 25285
rect 9861 25245 9873 25279
rect 9907 25245 9919 25279
rect 9861 25239 9919 25245
rect 11146 25236 11152 25288
rect 11204 25236 11210 25288
rect 11348 25285 11376 25384
rect 14568 25353 14596 25452
rect 14918 25440 14924 25452
rect 14976 25440 14982 25492
rect 15194 25440 15200 25492
rect 15252 25480 15258 25492
rect 15381 25483 15439 25489
rect 15381 25480 15393 25483
rect 15252 25452 15393 25480
rect 15252 25440 15258 25452
rect 15381 25449 15393 25452
rect 15427 25449 15439 25483
rect 15381 25443 15439 25449
rect 15562 25440 15568 25492
rect 15620 25440 15626 25492
rect 15746 25440 15752 25492
rect 15804 25480 15810 25492
rect 16574 25480 16580 25492
rect 15804 25452 16580 25480
rect 15804 25440 15810 25452
rect 16574 25440 16580 25452
rect 16632 25440 16638 25492
rect 16669 25483 16727 25489
rect 16669 25449 16681 25483
rect 16715 25480 16727 25483
rect 16850 25480 16856 25492
rect 16715 25452 16856 25480
rect 16715 25449 16727 25452
rect 16669 25443 16727 25449
rect 16850 25440 16856 25452
rect 16908 25440 16914 25492
rect 20714 25480 20720 25492
rect 17926 25452 20720 25480
rect 14660 25384 15608 25412
rect 14553 25347 14611 25353
rect 14553 25344 14565 25347
rect 11532 25316 14565 25344
rect 11532 25288 11560 25316
rect 14553 25313 14565 25316
rect 14599 25313 14611 25347
rect 14553 25307 14611 25313
rect 11333 25279 11391 25285
rect 11333 25245 11345 25279
rect 11379 25245 11391 25279
rect 11333 25239 11391 25245
rect 11514 25236 11520 25288
rect 11572 25236 11578 25288
rect 11698 25236 11704 25288
rect 11756 25276 11762 25288
rect 13354 25276 13360 25288
rect 11756 25248 13360 25276
rect 11756 25236 11762 25248
rect 13354 25236 13360 25248
rect 13412 25236 13418 25288
rect 14660 25276 14688 25384
rect 14921 25347 14979 25353
rect 14921 25313 14933 25347
rect 14967 25344 14979 25347
rect 15378 25344 15384 25356
rect 14967 25316 15384 25344
rect 14967 25313 14979 25316
rect 14921 25307 14979 25313
rect 15378 25304 15384 25316
rect 15436 25304 15442 25356
rect 15580 25344 15608 25384
rect 16758 25372 16764 25424
rect 16816 25412 16822 25424
rect 17926 25412 17954 25452
rect 20714 25440 20720 25452
rect 20772 25440 20778 25492
rect 21174 25440 21180 25492
rect 21232 25480 21238 25492
rect 21232 25452 25176 25480
rect 21232 25440 21238 25452
rect 16816 25384 16896 25412
rect 16816 25372 16822 25384
rect 15654 25344 15660 25356
rect 15580 25316 15660 25344
rect 15654 25304 15660 25316
rect 15712 25304 15718 25356
rect 16022 25304 16028 25356
rect 16080 25304 16086 25356
rect 16298 25304 16304 25356
rect 16356 25304 16362 25356
rect 16868 25353 16896 25384
rect 17144 25384 17954 25412
rect 18233 25415 18291 25421
rect 16853 25347 16911 25353
rect 16853 25313 16865 25347
rect 16899 25313 16911 25347
rect 16853 25307 16911 25313
rect 17034 25304 17040 25356
rect 17092 25344 17098 25356
rect 17144 25344 17172 25384
rect 18233 25381 18245 25415
rect 18279 25412 18291 25415
rect 19242 25412 19248 25424
rect 18279 25384 19248 25412
rect 18279 25381 18291 25384
rect 18233 25375 18291 25381
rect 19242 25372 19248 25384
rect 19300 25372 19306 25424
rect 20622 25372 20628 25424
rect 20680 25412 20686 25424
rect 20680 25384 22968 25412
rect 20680 25372 20686 25384
rect 17092 25316 17172 25344
rect 17092 25304 17098 25316
rect 17954 25304 17960 25356
rect 18012 25304 18018 25356
rect 18046 25304 18052 25356
rect 18104 25304 18110 25356
rect 18325 25347 18383 25353
rect 18325 25313 18337 25347
rect 18371 25344 18383 25347
rect 19426 25344 19432 25356
rect 18371 25316 19432 25344
rect 18371 25313 18383 25316
rect 18325 25307 18383 25313
rect 19426 25304 19432 25316
rect 19484 25304 19490 25356
rect 21450 25344 21456 25356
rect 20916 25316 21456 25344
rect 14292 25248 14688 25276
rect 14737 25279 14795 25285
rect 11882 25168 11888 25220
rect 11940 25208 11946 25220
rect 14292 25208 14320 25248
rect 14737 25245 14749 25279
rect 14783 25245 14795 25279
rect 14737 25239 14795 25245
rect 11940 25180 14320 25208
rect 11940 25168 11946 25180
rect 14366 25168 14372 25220
rect 14424 25208 14430 25220
rect 14752 25208 14780 25239
rect 14826 25236 14832 25288
rect 14884 25276 14890 25288
rect 15197 25279 15255 25285
rect 15197 25276 15209 25279
rect 14884 25248 15209 25276
rect 14884 25236 14890 25248
rect 15197 25245 15209 25248
rect 15243 25245 15255 25279
rect 15197 25239 15255 25245
rect 14424 25180 14780 25208
rect 15212 25208 15240 25239
rect 15286 25236 15292 25288
rect 15344 25276 15350 25288
rect 15473 25279 15531 25285
rect 15473 25276 15485 25279
rect 15344 25248 15485 25276
rect 15344 25236 15350 25248
rect 15473 25245 15485 25248
rect 15519 25276 15531 25279
rect 15565 25279 15623 25285
rect 15565 25276 15577 25279
rect 15519 25248 15577 25276
rect 15519 25245 15531 25248
rect 15473 25239 15531 25245
rect 15565 25245 15577 25248
rect 15611 25276 15623 25279
rect 15838 25276 15844 25288
rect 15611 25248 15844 25276
rect 15611 25245 15623 25248
rect 15565 25239 15623 25245
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 15930 25236 15936 25288
rect 15988 25276 15994 25288
rect 16209 25279 16267 25285
rect 16209 25276 16221 25279
rect 15988 25248 16221 25276
rect 15988 25236 15994 25248
rect 16209 25245 16221 25248
rect 16255 25245 16267 25279
rect 16316 25276 16344 25304
rect 16758 25276 16764 25288
rect 16316 25248 16764 25276
rect 16209 25239 16267 25245
rect 16758 25236 16764 25248
rect 16816 25276 16822 25288
rect 16816 25248 16896 25276
rect 16816 25236 16822 25248
rect 16022 25208 16028 25220
rect 15212 25180 16028 25208
rect 14424 25168 14430 25180
rect 16022 25168 16028 25180
rect 16080 25168 16086 25220
rect 16482 25168 16488 25220
rect 16540 25168 16546 25220
rect 16577 25211 16635 25217
rect 16577 25177 16589 25211
rect 16623 25177 16635 25211
rect 16868 25208 16896 25248
rect 16942 25236 16948 25288
rect 17000 25236 17006 25288
rect 17129 25279 17187 25285
rect 17129 25245 17141 25279
rect 17175 25245 17187 25279
rect 17129 25239 17187 25245
rect 17144 25208 17172 25239
rect 17402 25236 17408 25288
rect 17460 25236 17466 25288
rect 18064 25276 18092 25304
rect 20916 25288 20944 25316
rect 18141 25279 18199 25285
rect 18141 25276 18153 25279
rect 18064 25248 18153 25276
rect 18141 25245 18153 25248
rect 18187 25245 18199 25279
rect 18141 25239 18199 25245
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25276 18475 25279
rect 18506 25276 18512 25288
rect 18463 25248 18512 25276
rect 18463 25245 18475 25248
rect 18417 25239 18475 25245
rect 18506 25236 18512 25248
rect 18564 25236 18570 25288
rect 18601 25279 18659 25285
rect 18601 25245 18613 25279
rect 18647 25245 18659 25279
rect 18601 25239 18659 25245
rect 16868 25180 17172 25208
rect 17420 25208 17448 25236
rect 18616 25208 18644 25239
rect 20898 25236 20904 25288
rect 20956 25236 20962 25288
rect 21284 25285 21312 25316
rect 21450 25304 21456 25316
rect 21508 25344 21514 25356
rect 22940 25344 22968 25384
rect 25148 25344 25176 25452
rect 25498 25440 25504 25492
rect 25556 25440 25562 25492
rect 25774 25440 25780 25492
rect 25832 25480 25838 25492
rect 26510 25480 26516 25492
rect 25832 25452 26516 25480
rect 25832 25440 25838 25452
rect 26510 25440 26516 25452
rect 26568 25440 26574 25492
rect 27338 25440 27344 25492
rect 27396 25480 27402 25492
rect 28077 25483 28135 25489
rect 28077 25480 28089 25483
rect 27396 25452 28089 25480
rect 27396 25440 27402 25452
rect 28077 25449 28089 25452
rect 28123 25449 28135 25483
rect 28077 25443 28135 25449
rect 30650 25440 30656 25492
rect 30708 25480 30714 25492
rect 31021 25483 31079 25489
rect 31021 25480 31033 25483
rect 30708 25452 31033 25480
rect 30708 25440 30714 25452
rect 31021 25449 31033 25452
rect 31067 25449 31079 25483
rect 31021 25443 31079 25449
rect 32214 25440 32220 25492
rect 32272 25480 32278 25492
rect 32272 25452 34376 25480
rect 32272 25440 32278 25452
rect 25516 25344 25544 25440
rect 28166 25372 28172 25424
rect 28224 25372 28230 25424
rect 28644 25384 31340 25412
rect 21508 25316 22784 25344
rect 21508 25304 21514 25316
rect 20993 25279 21051 25285
rect 20993 25245 21005 25279
rect 21039 25245 21051 25279
rect 20993 25239 21051 25245
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 17420 25180 18644 25208
rect 16577 25171 16635 25177
rect 9398 25140 9404 25152
rect 9140 25112 9404 25140
rect 8067 25109 8079 25112
rect 8021 25103 8079 25109
rect 9398 25100 9404 25112
rect 9456 25100 9462 25152
rect 11333 25143 11391 25149
rect 11333 25109 11345 25143
rect 11379 25140 11391 25143
rect 12250 25140 12256 25152
rect 11379 25112 12256 25140
rect 11379 25109 11391 25112
rect 11333 25103 11391 25109
rect 12250 25100 12256 25112
rect 12308 25100 12314 25152
rect 12526 25100 12532 25152
rect 12584 25140 12590 25152
rect 13446 25140 13452 25152
rect 12584 25112 13452 25140
rect 12584 25100 12590 25112
rect 13446 25100 13452 25112
rect 13504 25100 13510 25152
rect 13630 25100 13636 25152
rect 13688 25140 13694 25152
rect 14274 25140 14280 25152
rect 13688 25112 14280 25140
rect 13688 25100 13694 25112
rect 14274 25100 14280 25112
rect 14332 25100 14338 25152
rect 14918 25100 14924 25152
rect 14976 25140 14982 25152
rect 15013 25143 15071 25149
rect 15013 25140 15025 25143
rect 14976 25112 15025 25140
rect 14976 25100 14982 25112
rect 15013 25109 15025 25112
rect 15059 25109 15071 25143
rect 15013 25103 15071 25109
rect 15562 25100 15568 25152
rect 15620 25140 15626 25152
rect 15930 25140 15936 25152
rect 15620 25112 15936 25140
rect 15620 25100 15626 25112
rect 15930 25100 15936 25112
rect 15988 25100 15994 25152
rect 16040 25140 16068 25168
rect 16592 25140 16620 25171
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 19886 25208 19892 25220
rect 19484 25180 19892 25208
rect 19484 25168 19490 25180
rect 19886 25168 19892 25180
rect 19944 25208 19950 25220
rect 21008 25208 21036 25239
rect 21358 25236 21364 25288
rect 21416 25236 21422 25288
rect 22186 25276 22192 25288
rect 22066 25248 22192 25276
rect 19944 25180 21036 25208
rect 21177 25211 21235 25217
rect 19944 25168 19950 25180
rect 21177 25177 21189 25211
rect 21223 25177 21235 25211
rect 22066 25208 22094 25248
rect 22186 25236 22192 25248
rect 22244 25236 22250 25288
rect 22756 25285 22784 25316
rect 22940 25316 24164 25344
rect 25148 25316 25268 25344
rect 22940 25285 22968 25316
rect 24136 25288 24164 25316
rect 22649 25279 22707 25285
rect 22649 25245 22661 25279
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 22741 25279 22799 25285
rect 22741 25245 22753 25279
rect 22787 25245 22799 25279
rect 22741 25239 22799 25245
rect 22925 25279 22983 25285
rect 22925 25245 22937 25279
rect 22971 25245 22983 25279
rect 22925 25239 22983 25245
rect 21177 25171 21235 25177
rect 21468 25180 22094 25208
rect 22664 25208 22692 25239
rect 23014 25236 23020 25288
rect 23072 25236 23078 25288
rect 23658 25276 23664 25288
rect 23124 25248 23664 25276
rect 23124 25208 23152 25248
rect 23658 25236 23664 25248
rect 23716 25236 23722 25288
rect 24118 25236 24124 25288
rect 24176 25236 24182 25288
rect 25130 25236 25136 25288
rect 25188 25236 25194 25288
rect 25240 25285 25268 25316
rect 25424 25316 25544 25344
rect 25424 25285 25452 25316
rect 26326 25304 26332 25356
rect 26384 25344 26390 25356
rect 28258 25344 28264 25356
rect 26384 25316 28264 25344
rect 26384 25304 26390 25316
rect 28258 25304 28264 25316
rect 28316 25304 28322 25356
rect 28350 25304 28356 25356
rect 28408 25304 28414 25356
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25245 25283 25279
rect 25225 25239 25283 25245
rect 25409 25279 25467 25285
rect 25409 25245 25421 25279
rect 25455 25245 25467 25279
rect 25409 25239 25467 25245
rect 25501 25279 25559 25285
rect 25501 25245 25513 25279
rect 25547 25276 25559 25279
rect 25590 25276 25596 25288
rect 25547 25248 25596 25276
rect 25547 25245 25559 25248
rect 25501 25239 25559 25245
rect 22664 25180 23152 25208
rect 25240 25208 25268 25239
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 28077 25279 28135 25285
rect 28077 25276 28089 25279
rect 27586 25248 28089 25276
rect 26970 25208 26976 25220
rect 25240 25180 26976 25208
rect 16942 25140 16948 25152
rect 16040 25112 16948 25140
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 17586 25100 17592 25152
rect 17644 25140 17650 25152
rect 18874 25140 18880 25152
rect 17644 25112 18880 25140
rect 17644 25100 17650 25112
rect 18874 25100 18880 25112
rect 18932 25100 18938 25152
rect 21192 25140 21220 25171
rect 21468 25140 21496 25180
rect 26970 25168 26976 25180
rect 27028 25168 27034 25220
rect 21192 25112 21496 25140
rect 21542 25100 21548 25152
rect 21600 25100 21606 25152
rect 22186 25100 22192 25152
rect 22244 25140 22250 25152
rect 22465 25143 22523 25149
rect 22465 25140 22477 25143
rect 22244 25112 22477 25140
rect 22244 25100 22250 25112
rect 22465 25109 22477 25112
rect 22511 25109 22523 25143
rect 22465 25103 22523 25109
rect 24949 25143 25007 25149
rect 24949 25109 24961 25143
rect 24995 25140 25007 25143
rect 25314 25140 25320 25152
rect 24995 25112 25320 25140
rect 24995 25109 25007 25112
rect 24949 25103 25007 25109
rect 25314 25100 25320 25112
rect 25372 25100 25378 25152
rect 25958 25100 25964 25152
rect 26016 25140 26022 25152
rect 27586 25140 27614 25248
rect 28077 25245 28089 25248
rect 28123 25276 28135 25279
rect 28644 25276 28672 25384
rect 29641 25347 29699 25353
rect 29641 25313 29653 25347
rect 29687 25344 29699 25347
rect 30558 25344 30564 25356
rect 29687 25316 30564 25344
rect 29687 25313 29699 25316
rect 29641 25307 29699 25313
rect 28123 25248 28672 25276
rect 28123 25245 28135 25248
rect 28077 25239 28135 25245
rect 28718 25236 28724 25288
rect 28776 25236 28782 25288
rect 28997 25279 29055 25285
rect 28997 25245 29009 25279
rect 29043 25276 29055 25279
rect 29086 25276 29092 25288
rect 29043 25248 29092 25276
rect 29043 25245 29055 25248
rect 28997 25239 29055 25245
rect 29086 25236 29092 25248
rect 29144 25236 29150 25288
rect 29549 25279 29607 25285
rect 29257 25273 29315 25279
rect 29549 25276 29561 25279
rect 29257 25270 29269 25273
rect 29196 25242 29269 25270
rect 28736 25208 28764 25236
rect 29196 25208 29224 25242
rect 29257 25239 29269 25242
rect 29303 25270 29315 25273
rect 29303 25254 29316 25270
rect 29472 25254 29561 25276
rect 29303 25248 29561 25254
rect 29303 25239 29500 25248
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 29257 25233 29500 25239
rect 29730 25236 29736 25288
rect 29788 25236 29794 25288
rect 30300 25285 30328 25316
rect 30558 25304 30564 25316
rect 30616 25304 30622 25356
rect 31312 25353 31340 25384
rect 31297 25347 31355 25353
rect 31297 25313 31309 25347
rect 31343 25344 31355 25347
rect 31938 25344 31944 25356
rect 31343 25316 31944 25344
rect 31343 25313 31355 25316
rect 31297 25307 31355 25313
rect 31938 25304 31944 25316
rect 31996 25304 32002 25356
rect 32214 25304 32220 25356
rect 32272 25344 32278 25356
rect 32493 25347 32551 25353
rect 32493 25344 32505 25347
rect 32272 25316 32505 25344
rect 32272 25304 32278 25316
rect 32493 25313 32505 25316
rect 32539 25344 32551 25347
rect 34348 25344 34376 25452
rect 36078 25440 36084 25492
rect 36136 25440 36142 25492
rect 34517 25347 34575 25353
rect 34517 25344 34529 25347
rect 32539 25316 34284 25344
rect 34348 25316 34529 25344
rect 32539 25313 32551 25316
rect 32493 25307 32551 25313
rect 30285 25279 30343 25285
rect 30285 25245 30297 25279
rect 30331 25245 30343 25279
rect 30285 25239 30343 25245
rect 30374 25236 30380 25288
rect 30432 25276 30438 25288
rect 30469 25279 30527 25285
rect 30469 25276 30481 25279
rect 30432 25248 30481 25276
rect 30432 25236 30438 25248
rect 30469 25245 30481 25248
rect 30515 25245 30527 25279
rect 30469 25239 30527 25245
rect 31021 25279 31079 25285
rect 31021 25245 31033 25279
rect 31067 25245 31079 25279
rect 31021 25239 31079 25245
rect 29288 25226 29500 25233
rect 28736 25180 29224 25208
rect 31036 25208 31064 25239
rect 31110 25236 31116 25288
rect 31168 25236 31174 25288
rect 34256 25276 34284 25316
rect 34517 25313 34529 25316
rect 34563 25313 34575 25347
rect 34517 25307 34575 25313
rect 35069 25347 35127 25353
rect 35069 25313 35081 25347
rect 35115 25344 35127 25347
rect 36096 25344 36124 25440
rect 35115 25316 36124 25344
rect 35115 25313 35127 25316
rect 35069 25307 35127 25313
rect 36262 25304 36268 25356
rect 36320 25304 36326 25356
rect 34422 25276 34428 25288
rect 34256 25248 34428 25276
rect 34422 25236 34428 25248
rect 34480 25276 34486 25288
rect 34790 25276 34796 25288
rect 34480 25248 34796 25276
rect 34480 25236 34486 25248
rect 34790 25236 34796 25248
rect 34848 25236 34854 25288
rect 36280 25276 36308 25304
rect 36202 25262 36308 25276
rect 36188 25248 36308 25262
rect 31662 25208 31668 25220
rect 31036 25180 31668 25208
rect 31662 25168 31668 25180
rect 31720 25168 31726 25220
rect 32674 25168 32680 25220
rect 32732 25208 32738 25220
rect 32769 25211 32827 25217
rect 32769 25208 32781 25211
rect 32732 25180 32781 25208
rect 32732 25168 32738 25180
rect 32769 25177 32781 25180
rect 32815 25177 32827 25211
rect 34054 25208 34060 25220
rect 33994 25180 34060 25208
rect 32769 25171 32827 25177
rect 34054 25168 34060 25180
rect 34112 25208 34118 25220
rect 34112 25180 34836 25208
rect 34112 25168 34118 25180
rect 26016 25112 27614 25140
rect 26016 25100 26022 25112
rect 28810 25100 28816 25152
rect 28868 25100 28874 25152
rect 28994 25100 29000 25152
rect 29052 25140 29058 25152
rect 29181 25143 29239 25149
rect 29181 25140 29193 25143
rect 29052 25112 29193 25140
rect 29052 25100 29058 25112
rect 29181 25109 29193 25112
rect 29227 25109 29239 25143
rect 29181 25103 29239 25109
rect 29730 25100 29736 25152
rect 29788 25140 29794 25152
rect 30377 25143 30435 25149
rect 30377 25140 30389 25143
rect 29788 25112 30389 25140
rect 29788 25100 29794 25112
rect 30377 25109 30389 25112
rect 30423 25140 30435 25143
rect 33502 25140 33508 25152
rect 30423 25112 33508 25140
rect 30423 25109 30435 25112
rect 30377 25103 30435 25109
rect 33502 25100 33508 25112
rect 33560 25100 33566 25152
rect 34808 25140 34836 25180
rect 35802 25140 35808 25152
rect 34808 25112 35808 25140
rect 35802 25100 35808 25112
rect 35860 25140 35866 25152
rect 36188 25140 36216 25248
rect 36814 25236 36820 25288
rect 36872 25236 36878 25288
rect 35860 25112 36216 25140
rect 35860 25100 35866 25112
rect 1104 25050 41400 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 41400 25050
rect 1104 24976 41400 24998
rect 3697 24939 3755 24945
rect 3697 24905 3709 24939
rect 3743 24936 3755 24939
rect 4062 24936 4068 24948
rect 3743 24908 4068 24936
rect 3743 24905 3755 24908
rect 3697 24899 3755 24905
rect 4062 24896 4068 24908
rect 4120 24896 4126 24948
rect 4617 24939 4675 24945
rect 4617 24905 4629 24939
rect 4663 24936 4675 24939
rect 4706 24936 4712 24948
rect 4663 24908 4712 24936
rect 4663 24905 4675 24908
rect 4617 24899 4675 24905
rect 4706 24896 4712 24908
rect 4764 24896 4770 24948
rect 8294 24936 8300 24948
rect 8220 24908 8300 24936
rect 3881 24803 3939 24809
rect 3881 24769 3893 24803
rect 3927 24800 3939 24803
rect 8021 24803 8079 24809
rect 3927 24772 4292 24800
rect 3927 24769 3939 24772
rect 3881 24763 3939 24769
rect 4264 24673 4292 24772
rect 8021 24769 8033 24803
rect 8067 24769 8079 24803
rect 8021 24763 8079 24769
rect 8113 24803 8171 24809
rect 8113 24769 8125 24803
rect 8159 24800 8171 24803
rect 8220 24800 8248 24908
rect 8294 24896 8300 24908
rect 8352 24896 8358 24948
rect 8478 24936 8484 24948
rect 8404 24908 8484 24936
rect 8404 24868 8432 24908
rect 8478 24896 8484 24908
rect 8536 24896 8542 24948
rect 8570 24896 8576 24948
rect 8628 24936 8634 24948
rect 11514 24936 11520 24948
rect 8628 24908 11520 24936
rect 8628 24896 8634 24908
rect 11514 24896 11520 24908
rect 11572 24896 11578 24948
rect 12158 24896 12164 24948
rect 12216 24936 12222 24948
rect 12216 24908 12848 24936
rect 12216 24896 12222 24908
rect 8312 24840 8432 24868
rect 8312 24809 8340 24840
rect 10042 24828 10048 24880
rect 10100 24868 10106 24880
rect 12253 24871 12311 24877
rect 12253 24868 12265 24871
rect 10100 24840 12265 24868
rect 10100 24828 10106 24840
rect 12253 24837 12265 24840
rect 12299 24837 12311 24871
rect 12253 24831 12311 24837
rect 12345 24871 12403 24877
rect 12345 24837 12357 24871
rect 12391 24868 12403 24871
rect 12526 24868 12532 24880
rect 12391 24840 12532 24868
rect 12391 24837 12403 24840
rect 12345 24831 12403 24837
rect 12526 24828 12532 24840
rect 12584 24828 12590 24880
rect 8159 24772 8248 24800
rect 8297 24803 8355 24809
rect 8159 24769 8171 24772
rect 8113 24763 8171 24769
rect 8297 24769 8309 24803
rect 8343 24769 8355 24803
rect 8297 24763 8355 24769
rect 4706 24692 4712 24744
rect 4764 24692 4770 24744
rect 4890 24692 4896 24744
rect 4948 24692 4954 24744
rect 8036 24732 8064 24763
rect 8386 24760 8392 24812
rect 8444 24760 8450 24812
rect 8662 24809 8668 24812
rect 8481 24803 8539 24809
rect 8481 24769 8493 24803
rect 8527 24769 8539 24803
rect 8481 24763 8539 24769
rect 8629 24803 8668 24809
rect 8629 24769 8641 24803
rect 8629 24763 8668 24769
rect 8202 24732 8208 24744
rect 8036 24704 8208 24732
rect 8202 24692 8208 24704
rect 8260 24692 8266 24744
rect 8496 24732 8524 24763
rect 8662 24760 8668 24763
rect 8720 24760 8726 24812
rect 8754 24760 8760 24812
rect 8812 24760 8818 24812
rect 8846 24760 8852 24812
rect 8904 24760 8910 24812
rect 8987 24804 9045 24809
rect 9122 24804 9128 24812
rect 8987 24803 9128 24804
rect 8987 24769 8999 24803
rect 9033 24776 9128 24803
rect 9033 24769 9045 24776
rect 8987 24763 9045 24769
rect 9122 24760 9128 24776
rect 9180 24760 9186 24812
rect 11422 24800 11428 24812
rect 9232 24772 11428 24800
rect 9232 24732 9260 24772
rect 11422 24760 11428 24772
rect 11480 24760 11486 24812
rect 11977 24803 12035 24809
rect 11977 24769 11989 24803
rect 12023 24769 12035 24803
rect 11977 24763 12035 24769
rect 12125 24803 12183 24809
rect 12125 24769 12137 24803
rect 12171 24800 12183 24803
rect 12171 24772 12296 24800
rect 12171 24769 12183 24772
rect 12125 24763 12183 24769
rect 8496 24704 9260 24732
rect 9306 24692 9312 24744
rect 9364 24732 9370 24744
rect 11054 24732 11060 24744
rect 9364 24704 11060 24732
rect 9364 24692 9370 24704
rect 11054 24692 11060 24704
rect 11112 24692 11118 24744
rect 4249 24667 4307 24673
rect 4249 24633 4261 24667
rect 4295 24633 4307 24667
rect 4249 24627 4307 24633
rect 9950 24624 9956 24676
rect 10008 24664 10014 24676
rect 11606 24664 11612 24676
rect 10008 24636 11612 24664
rect 10008 24624 10014 24636
rect 11606 24624 11612 24636
rect 11664 24624 11670 24676
rect 11992 24608 12020 24763
rect 12268 24664 12296 24772
rect 12434 24760 12440 24812
rect 12492 24809 12498 24812
rect 12820 24809 12848 24908
rect 13446 24896 13452 24948
rect 13504 24936 13510 24948
rect 14826 24936 14832 24948
rect 13504 24908 14832 24936
rect 13504 24896 13510 24908
rect 13630 24828 13636 24880
rect 13688 24828 13694 24880
rect 13740 24877 13768 24908
rect 14826 24896 14832 24908
rect 14884 24896 14890 24948
rect 15120 24908 15516 24936
rect 13725 24871 13783 24877
rect 13725 24837 13737 24871
rect 13771 24837 13783 24871
rect 15120 24868 15148 24908
rect 13725 24831 13783 24837
rect 14016 24840 15148 24868
rect 15212 24840 15425 24868
rect 14016 24812 14044 24840
rect 12492 24763 12500 24809
rect 12713 24803 12771 24809
rect 12713 24800 12725 24803
rect 12709 24769 12725 24800
rect 12759 24769 12771 24803
rect 12709 24763 12771 24769
rect 12806 24803 12864 24809
rect 12806 24769 12818 24803
rect 12852 24769 12864 24803
rect 12806 24763 12864 24769
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 12492 24760 12498 24763
rect 12526 24692 12532 24744
rect 12584 24732 12590 24744
rect 12709 24732 12737 24763
rect 12584 24704 12737 24732
rect 13004 24732 13032 24763
rect 13078 24760 13084 24812
rect 13136 24760 13142 24812
rect 13170 24760 13176 24812
rect 13228 24809 13234 24812
rect 13228 24800 13236 24809
rect 13449 24803 13507 24809
rect 13228 24772 13273 24800
rect 13228 24763 13236 24772
rect 13449 24769 13461 24803
rect 13495 24800 13507 24803
rect 13817 24806 13875 24809
rect 13998 24806 14004 24812
rect 13817 24803 14004 24806
rect 13495 24772 13768 24800
rect 13495 24769 13507 24772
rect 13449 24763 13507 24769
rect 13228 24760 13234 24763
rect 13004 24704 13124 24732
rect 12584 24692 12590 24704
rect 13096 24664 13124 24704
rect 13464 24664 13492 24763
rect 13740 24732 13768 24772
rect 13817 24769 13829 24803
rect 13863 24778 14004 24803
rect 13863 24769 13875 24778
rect 13817 24763 13875 24769
rect 13998 24760 14004 24778
rect 14056 24760 14062 24812
rect 14182 24760 14188 24812
rect 14240 24760 14246 24812
rect 14274 24760 14280 24812
rect 14332 24760 14338 24812
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24769 14427 24803
rect 14369 24763 14427 24769
rect 14553 24803 14611 24809
rect 14553 24769 14565 24803
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 14645 24803 14703 24809
rect 14645 24769 14657 24803
rect 14691 24769 14703 24803
rect 14645 24763 14703 24769
rect 14200 24732 14228 24760
rect 14384 24732 14412 24763
rect 13740 24704 14412 24732
rect 12268 24636 13492 24664
rect 14568 24664 14596 24763
rect 14660 24732 14688 24763
rect 15010 24760 15016 24812
rect 15068 24800 15074 24812
rect 15212 24800 15240 24840
rect 15068 24772 15240 24800
rect 15068 24760 15074 24772
rect 15286 24760 15292 24812
rect 15344 24760 15350 24812
rect 15397 24809 15425 24840
rect 15382 24803 15440 24809
rect 15382 24769 15394 24803
rect 15428 24769 15440 24803
rect 15488 24800 15516 24908
rect 18322 24896 18328 24948
rect 18380 24896 18386 24948
rect 18414 24896 18420 24948
rect 18472 24936 18478 24948
rect 18472 24908 19012 24936
rect 18472 24896 18478 24908
rect 15562 24828 15568 24880
rect 15620 24828 15626 24880
rect 15654 24828 15660 24880
rect 15712 24868 15718 24880
rect 17126 24868 17132 24880
rect 15712 24840 17132 24868
rect 15712 24828 15718 24840
rect 17126 24828 17132 24840
rect 17184 24828 17190 24880
rect 18340 24868 18368 24896
rect 18984 24868 19012 24908
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19392 24908 21128 24936
rect 19392 24896 19398 24908
rect 18340 24840 18920 24868
rect 18984 24840 20293 24868
rect 15754 24803 15812 24809
rect 15754 24800 15766 24803
rect 15488 24772 15766 24800
rect 15382 24763 15440 24769
rect 15754 24769 15766 24772
rect 15800 24769 15812 24803
rect 15754 24763 15812 24769
rect 16574 24760 16580 24812
rect 16632 24760 16638 24812
rect 17313 24803 17371 24809
rect 17313 24769 17325 24803
rect 17359 24800 17371 24803
rect 18230 24800 18236 24812
rect 17359 24772 18236 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 18892 24800 18920 24840
rect 19153 24803 19211 24809
rect 19153 24800 19165 24803
rect 18892 24772 19165 24800
rect 19153 24769 19165 24772
rect 19199 24769 19211 24803
rect 19153 24763 19211 24769
rect 19334 24760 19340 24812
rect 19392 24760 19398 24812
rect 19794 24760 19800 24812
rect 19852 24800 19858 24812
rect 19981 24803 20039 24809
rect 19981 24800 19993 24803
rect 19852 24772 19993 24800
rect 19852 24760 19858 24772
rect 19981 24769 19993 24772
rect 20027 24800 20039 24803
rect 20070 24800 20076 24812
rect 20027 24772 20076 24800
rect 20027 24769 20039 24772
rect 19981 24763 20039 24769
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20162 24760 20168 24812
rect 20220 24760 20226 24812
rect 14826 24732 14832 24744
rect 14660 24704 14832 24732
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 15194 24692 15200 24744
rect 15252 24692 15258 24744
rect 15838 24692 15844 24744
rect 15896 24692 15902 24744
rect 16592 24732 16620 24760
rect 17589 24735 17647 24741
rect 17589 24732 17601 24735
rect 16592 24704 17601 24732
rect 17589 24701 17601 24704
rect 17635 24732 17647 24735
rect 19518 24732 19524 24744
rect 17635 24704 19524 24732
rect 17635 24701 17647 24704
rect 17589 24695 17647 24701
rect 19518 24692 19524 24704
rect 19576 24692 19582 24744
rect 19702 24692 19708 24744
rect 19760 24732 19766 24744
rect 20180 24732 20208 24760
rect 19760 24704 20208 24732
rect 19760 24692 19766 24704
rect 15212 24664 15240 24692
rect 14568 24636 15240 24664
rect 15856 24664 15884 24692
rect 17497 24667 17555 24673
rect 17497 24664 17509 24667
rect 15856 24636 17509 24664
rect 17497 24633 17509 24636
rect 17543 24633 17555 24667
rect 17497 24627 17555 24633
rect 19613 24667 19671 24673
rect 19613 24633 19625 24667
rect 19659 24664 19671 24667
rect 20070 24664 20076 24676
rect 19659 24636 20076 24664
rect 19659 24633 19671 24636
rect 19613 24627 19671 24633
rect 20070 24624 20076 24636
rect 20128 24624 20134 24676
rect 20265 24664 20293 24840
rect 20349 24803 20407 24809
rect 20349 24769 20361 24803
rect 20395 24800 20407 24803
rect 20438 24800 20444 24812
rect 20395 24772 20444 24800
rect 20395 24769 20407 24772
rect 20349 24763 20407 24769
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 20714 24760 20720 24812
rect 20772 24760 20778 24812
rect 21100 24809 21128 24908
rect 21634 24896 21640 24948
rect 21692 24936 21698 24948
rect 25130 24936 25136 24948
rect 21692 24908 25136 24936
rect 21692 24896 21698 24908
rect 25130 24896 25136 24908
rect 25188 24896 25194 24948
rect 27522 24896 27528 24948
rect 27580 24896 27586 24948
rect 29270 24936 29276 24948
rect 28966 24908 29276 24936
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24800 21143 24803
rect 21266 24800 21272 24812
rect 21131 24772 21272 24800
rect 21131 24769 21143 24772
rect 21085 24763 21143 24769
rect 21266 24760 21272 24772
rect 21324 24760 21330 24812
rect 21652 24809 21680 24896
rect 21637 24803 21695 24809
rect 21637 24769 21649 24803
rect 21683 24769 21695 24803
rect 21637 24763 21695 24769
rect 21913 24803 21971 24809
rect 21913 24769 21925 24803
rect 21959 24800 21971 24803
rect 22186 24800 22192 24812
rect 21959 24772 22192 24800
rect 21959 24769 21971 24772
rect 21913 24763 21971 24769
rect 22186 24760 22192 24772
rect 22244 24760 22250 24812
rect 22373 24803 22431 24809
rect 22373 24769 22385 24803
rect 22419 24800 22431 24803
rect 22830 24800 22836 24812
rect 22419 24772 22836 24800
rect 22419 24769 22431 24772
rect 22373 24763 22431 24769
rect 22830 24760 22836 24772
rect 22888 24760 22894 24812
rect 23658 24760 23664 24812
rect 23716 24760 23722 24812
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24769 23995 24803
rect 23937 24763 23995 24769
rect 20809 24735 20867 24741
rect 20809 24701 20821 24735
rect 20855 24732 20867 24735
rect 20898 24732 20904 24744
rect 20855 24704 20904 24732
rect 20855 24701 20867 24704
rect 20809 24695 20867 24701
rect 20898 24692 20904 24704
rect 20956 24692 20962 24744
rect 22094 24692 22100 24744
rect 22152 24692 22158 24744
rect 22278 24692 22284 24744
rect 22336 24692 22342 24744
rect 22649 24735 22707 24741
rect 22649 24701 22661 24735
rect 22695 24732 22707 24735
rect 22738 24732 22744 24744
rect 22695 24704 22744 24732
rect 22695 24701 22707 24704
rect 22649 24695 22707 24701
rect 22738 24692 22744 24704
rect 22796 24692 22802 24744
rect 22189 24667 22247 24673
rect 20265 24636 22048 24664
rect 7834 24556 7840 24608
rect 7892 24556 7898 24608
rect 9122 24556 9128 24608
rect 9180 24556 9186 24608
rect 11974 24556 11980 24608
rect 12032 24556 12038 24608
rect 12621 24599 12679 24605
rect 12621 24565 12633 24599
rect 12667 24596 12679 24599
rect 13262 24596 13268 24608
rect 12667 24568 13268 24596
rect 12667 24565 12679 24568
rect 12621 24559 12679 24565
rect 13262 24556 13268 24568
rect 13320 24556 13326 24608
rect 13354 24556 13360 24608
rect 13412 24556 13418 24608
rect 13998 24556 14004 24608
rect 14056 24556 14062 24608
rect 14093 24599 14151 24605
rect 14093 24565 14105 24599
rect 14139 24596 14151 24599
rect 14918 24596 14924 24608
rect 14139 24568 14924 24596
rect 14139 24565 14151 24568
rect 14093 24559 14151 24565
rect 14918 24556 14924 24568
rect 14976 24556 14982 24608
rect 15930 24556 15936 24608
rect 15988 24556 15994 24608
rect 16942 24556 16948 24608
rect 17000 24596 17006 24608
rect 17129 24599 17187 24605
rect 17129 24596 17141 24599
rect 17000 24568 17141 24596
rect 17000 24556 17006 24568
rect 17129 24565 17141 24568
rect 17175 24565 17187 24599
rect 17129 24559 17187 24565
rect 17586 24556 17592 24608
rect 17644 24596 17650 24608
rect 17862 24596 17868 24608
rect 17644 24568 17868 24596
rect 17644 24556 17650 24568
rect 17862 24556 17868 24568
rect 17920 24556 17926 24608
rect 18506 24556 18512 24608
rect 18564 24596 18570 24608
rect 20346 24596 20352 24608
rect 18564 24568 20352 24596
rect 18564 24556 18570 24568
rect 20346 24556 20352 24568
rect 20404 24556 20410 24608
rect 21634 24556 21640 24608
rect 21692 24596 21698 24608
rect 21913 24599 21971 24605
rect 21913 24596 21925 24599
rect 21692 24568 21925 24596
rect 21692 24556 21698 24568
rect 21913 24565 21925 24568
rect 21959 24565 21971 24599
rect 22020 24596 22048 24636
rect 22189 24633 22201 24667
rect 22235 24664 22247 24667
rect 22925 24667 22983 24673
rect 22925 24664 22937 24667
rect 22235 24636 22937 24664
rect 22235 24633 22247 24636
rect 22189 24627 22247 24633
rect 22925 24633 22937 24636
rect 22971 24633 22983 24667
rect 22925 24627 22983 24633
rect 23474 24624 23480 24676
rect 23532 24664 23538 24676
rect 23676 24664 23704 24760
rect 23952 24732 23980 24763
rect 24026 24760 24032 24812
rect 24084 24800 24090 24812
rect 24213 24803 24271 24809
rect 24213 24800 24225 24803
rect 24084 24772 24225 24800
rect 24084 24760 24090 24772
rect 24213 24769 24225 24772
rect 24259 24769 24271 24803
rect 24213 24763 24271 24769
rect 26878 24760 26884 24812
rect 26936 24760 26942 24812
rect 27062 24760 27068 24812
rect 27120 24760 27126 24812
rect 27249 24803 27307 24809
rect 27249 24769 27261 24803
rect 27295 24800 27307 24803
rect 27540 24800 27568 24896
rect 28353 24871 28411 24877
rect 28353 24837 28365 24871
rect 28399 24868 28411 24871
rect 28718 24868 28724 24880
rect 28399 24840 28724 24868
rect 28399 24837 28411 24840
rect 28353 24831 28411 24837
rect 28718 24828 28724 24840
rect 28776 24828 28782 24880
rect 27295 24772 27568 24800
rect 27295 24769 27307 24772
rect 27249 24763 27307 24769
rect 28074 24760 28080 24812
rect 28132 24760 28138 24812
rect 28537 24803 28595 24809
rect 28537 24769 28549 24803
rect 28583 24769 28595 24803
rect 28537 24763 28595 24769
rect 28629 24803 28687 24809
rect 28629 24769 28641 24803
rect 28675 24800 28687 24803
rect 28966 24800 28994 24908
rect 29270 24896 29276 24908
rect 29328 24896 29334 24948
rect 28675 24772 28994 24800
rect 28675 24769 28687 24772
rect 28629 24763 28687 24769
rect 24762 24732 24768 24744
rect 23952 24704 24768 24732
rect 24762 24692 24768 24704
rect 24820 24692 24826 24744
rect 26896 24732 26924 24760
rect 27433 24735 27491 24741
rect 27433 24732 27445 24735
rect 26896 24704 27445 24732
rect 24029 24667 24087 24673
rect 24029 24664 24041 24667
rect 23532 24636 24041 24664
rect 23532 24624 23538 24636
rect 24029 24633 24041 24636
rect 24075 24633 24087 24667
rect 24029 24627 24087 24633
rect 24121 24667 24179 24673
rect 24121 24633 24133 24667
rect 24167 24664 24179 24667
rect 26896 24664 26924 24704
rect 27433 24701 27445 24704
rect 27479 24701 27491 24735
rect 27433 24695 27491 24701
rect 27525 24735 27583 24741
rect 27525 24701 27537 24735
rect 27571 24732 27583 24735
rect 28092 24732 28120 24760
rect 27571 24704 28120 24732
rect 27571 24701 27583 24704
rect 27525 24695 27583 24701
rect 24167 24636 26924 24664
rect 24167 24633 24179 24636
rect 24121 24627 24179 24633
rect 26970 24624 26976 24676
rect 27028 24664 27034 24676
rect 28552 24664 28580 24763
rect 30374 24760 30380 24812
rect 30432 24800 30438 24812
rect 31297 24803 31355 24809
rect 31297 24800 31309 24803
rect 30432 24772 31309 24800
rect 30432 24760 30438 24772
rect 31297 24769 31309 24772
rect 31343 24769 31355 24803
rect 31297 24763 31355 24769
rect 40865 24803 40923 24809
rect 40865 24769 40877 24803
rect 40911 24800 40923 24803
rect 40911 24772 41368 24800
rect 40911 24769 40923 24772
rect 40865 24763 40923 24769
rect 30742 24692 30748 24744
rect 30800 24732 30806 24744
rect 31110 24732 31116 24744
rect 30800 24704 31116 24732
rect 30800 24692 30806 24704
rect 31110 24692 31116 24704
rect 31168 24732 31174 24744
rect 31168 24704 32444 24732
rect 31168 24692 31174 24704
rect 31846 24664 31852 24676
rect 27028 24636 28580 24664
rect 29196 24636 31852 24664
rect 27028 24624 27034 24636
rect 29196 24608 29224 24636
rect 31846 24624 31852 24636
rect 31904 24624 31910 24676
rect 32416 24608 32444 24704
rect 41340 24676 41368 24772
rect 41322 24624 41328 24676
rect 41380 24624 41386 24676
rect 22465 24599 22523 24605
rect 22465 24596 22477 24599
rect 22020 24568 22477 24596
rect 21913 24559 21971 24565
rect 22465 24565 22477 24568
rect 22511 24565 22523 24599
rect 22465 24559 22523 24565
rect 23750 24556 23756 24608
rect 23808 24556 23814 24608
rect 24302 24556 24308 24608
rect 24360 24596 24366 24608
rect 24486 24596 24492 24608
rect 24360 24568 24492 24596
rect 24360 24556 24366 24568
rect 24486 24556 24492 24568
rect 24544 24556 24550 24608
rect 24854 24556 24860 24608
rect 24912 24596 24918 24608
rect 26786 24596 26792 24608
rect 24912 24568 26792 24596
rect 24912 24556 24918 24568
rect 26786 24556 26792 24568
rect 26844 24556 26850 24608
rect 28353 24599 28411 24605
rect 28353 24565 28365 24599
rect 28399 24596 28411 24599
rect 28810 24596 28816 24608
rect 28399 24568 28816 24596
rect 28399 24565 28411 24568
rect 28353 24559 28411 24565
rect 28810 24556 28816 24568
rect 28868 24556 28874 24608
rect 29178 24556 29184 24608
rect 29236 24556 29242 24608
rect 31478 24556 31484 24608
rect 31536 24556 31542 24608
rect 32398 24556 32404 24608
rect 32456 24556 32462 24608
rect 41046 24556 41052 24608
rect 41104 24556 41110 24608
rect 1104 24506 41400 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 41400 24506
rect 1104 24432 41400 24454
rect 4890 24352 4896 24404
rect 4948 24392 4954 24404
rect 11238 24392 11244 24404
rect 4948 24364 11244 24392
rect 4948 24352 4954 24364
rect 11238 24352 11244 24364
rect 11296 24352 11302 24404
rect 11698 24352 11704 24404
rect 11756 24352 11762 24404
rect 13170 24392 13176 24404
rect 12457 24364 13176 24392
rect 7374 24284 7380 24336
rect 7432 24324 7438 24336
rect 11514 24324 11520 24336
rect 7432 24296 9444 24324
rect 7432 24284 7438 24296
rect 8202 24216 8208 24268
rect 8260 24256 8266 24268
rect 9416 24265 9444 24296
rect 10796 24296 11520 24324
rect 10796 24265 10824 24296
rect 11514 24284 11520 24296
rect 11572 24324 11578 24336
rect 11716 24324 11744 24352
rect 11572 24296 11744 24324
rect 11885 24327 11943 24333
rect 11572 24284 11578 24296
rect 11885 24293 11897 24327
rect 11931 24293 11943 24327
rect 11885 24287 11943 24293
rect 8941 24259 8999 24265
rect 8941 24256 8953 24259
rect 8260 24228 8953 24256
rect 8260 24216 8266 24228
rect 8941 24225 8953 24228
rect 8987 24225 8999 24259
rect 8941 24219 8999 24225
rect 9401 24259 9459 24265
rect 9401 24225 9413 24259
rect 9447 24225 9459 24259
rect 9401 24219 9459 24225
rect 10781 24259 10839 24265
rect 10781 24225 10793 24259
rect 10827 24225 10839 24259
rect 10781 24219 10839 24225
rect 11333 24259 11391 24265
rect 11333 24225 11345 24259
rect 11379 24256 11391 24259
rect 11900 24256 11928 24287
rect 11379 24228 11928 24256
rect 11379 24225 11391 24228
rect 11333 24219 11391 24225
rect 1489 24191 1547 24197
rect 1489 24157 1501 24191
rect 1535 24188 1547 24191
rect 6086 24188 6092 24200
rect 1535 24160 6092 24188
rect 1535 24157 1547 24160
rect 1489 24151 1547 24157
rect 6086 24148 6092 24160
rect 6144 24188 6150 24200
rect 6181 24191 6239 24197
rect 6181 24188 6193 24191
rect 6144 24160 6193 24188
rect 6144 24148 6150 24160
rect 6181 24157 6193 24160
rect 6227 24157 6239 24191
rect 6181 24151 6239 24157
rect 7098 24148 7104 24200
rect 7156 24148 7162 24200
rect 8846 24148 8852 24200
rect 8904 24188 8910 24200
rect 9306 24188 9312 24200
rect 8904 24160 9312 24188
rect 8904 24148 8910 24160
rect 9306 24148 9312 24160
rect 9364 24148 9370 24200
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 10321 24191 10379 24197
rect 10321 24188 10333 24191
rect 10192 24160 10333 24188
rect 10192 24148 10198 24160
rect 10321 24157 10333 24160
rect 10367 24157 10379 24191
rect 10321 24151 10379 24157
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24188 10655 24191
rect 10962 24188 10968 24200
rect 10643 24160 10968 24188
rect 10643 24157 10655 24160
rect 10597 24151 10655 24157
rect 4706 24080 4712 24132
rect 4764 24120 4770 24132
rect 9490 24120 9496 24132
rect 4764 24092 9496 24120
rect 4764 24080 4770 24092
rect 9490 24080 9496 24092
rect 9548 24080 9554 24132
rect 10336 24120 10364 24151
rect 10962 24148 10968 24160
rect 11020 24148 11026 24200
rect 11238 24148 11244 24200
rect 11296 24148 11302 24200
rect 11422 24148 11428 24200
rect 11480 24148 11486 24200
rect 11517 24191 11575 24197
rect 11517 24157 11529 24191
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 11256 24120 11284 24148
rect 10336 24092 11284 24120
rect 11532 24120 11560 24151
rect 11606 24148 11612 24200
rect 11664 24148 11670 24200
rect 11790 24148 11796 24200
rect 11848 24148 11854 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 11974 24188 11980 24200
rect 11931 24160 11980 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 11808 24120 11836 24148
rect 11532 24092 11836 24120
rect 11900 24120 11928 24151
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 12069 24191 12127 24197
rect 12069 24157 12081 24191
rect 12115 24188 12127 24191
rect 12345 24191 12403 24197
rect 12345 24188 12357 24191
rect 12115 24160 12357 24188
rect 12115 24157 12127 24160
rect 12069 24151 12127 24157
rect 12345 24157 12357 24160
rect 12391 24157 12403 24191
rect 12457 24188 12485 24364
rect 13170 24352 13176 24364
rect 13228 24352 13234 24404
rect 13357 24395 13415 24401
rect 13357 24361 13369 24395
rect 13403 24392 13415 24395
rect 13538 24392 13544 24404
rect 13403 24364 13544 24392
rect 13403 24361 13415 24364
rect 13357 24355 13415 24361
rect 13538 24352 13544 24364
rect 13596 24392 13602 24404
rect 15194 24392 15200 24404
rect 13596 24364 15200 24392
rect 13596 24352 13602 24364
rect 15194 24352 15200 24364
rect 15252 24352 15258 24404
rect 15286 24352 15292 24404
rect 15344 24352 15350 24404
rect 15930 24352 15936 24404
rect 15988 24352 15994 24404
rect 16592 24364 17448 24392
rect 12526 24284 12532 24336
rect 12584 24284 12590 24336
rect 13722 24324 13728 24336
rect 12820 24296 13728 24324
rect 12544 24256 12572 24284
rect 12544 24228 12664 24256
rect 12636 24197 12664 24228
rect 12820 24197 12848 24296
rect 13722 24284 13728 24296
rect 13780 24324 13786 24336
rect 14826 24324 14832 24336
rect 13780 24296 14832 24324
rect 13780 24284 13786 24296
rect 14826 24284 14832 24296
rect 14884 24284 14890 24336
rect 15304 24324 15332 24352
rect 16592 24324 16620 24364
rect 17034 24324 17040 24336
rect 15304 24296 16620 24324
rect 16960 24296 17040 24324
rect 13998 24256 14004 24268
rect 12912 24228 14004 24256
rect 12912 24197 12940 24228
rect 13998 24216 14004 24228
rect 14056 24216 14062 24268
rect 16025 24259 16083 24265
rect 16025 24256 16037 24259
rect 14108 24228 16037 24256
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12457 24160 12541 24188
rect 12345 24151 12403 24157
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 12621 24191 12679 24197
rect 12621 24157 12633 24191
rect 12667 24157 12679 24191
rect 12621 24151 12679 24157
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24157 12863 24191
rect 12805 24151 12863 24157
rect 12897 24191 12955 24197
rect 12897 24157 12909 24191
rect 12943 24157 12955 24191
rect 12897 24151 12955 24157
rect 12986 24148 12992 24200
rect 13044 24148 13050 24200
rect 13262 24148 13268 24200
rect 13320 24148 13326 24200
rect 14108 24120 14136 24228
rect 16025 24225 16037 24228
rect 16071 24256 16083 24259
rect 16577 24259 16635 24265
rect 16577 24256 16589 24259
rect 16071 24228 16589 24256
rect 16071 24225 16083 24228
rect 16025 24219 16083 24225
rect 16577 24225 16589 24228
rect 16623 24225 16635 24259
rect 16577 24219 16635 24225
rect 15838 24148 15844 24200
rect 15896 24148 15902 24200
rect 16114 24148 16120 24200
rect 16172 24148 16178 24200
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24157 16359 24191
rect 16301 24151 16359 24157
rect 11900 24092 14136 24120
rect 14182 24080 14188 24132
rect 14240 24080 14246 24132
rect 16316 24120 16344 24151
rect 16758 24148 16764 24200
rect 16816 24148 16822 24200
rect 16960 24188 16988 24296
rect 17034 24284 17040 24296
rect 17092 24284 17098 24336
rect 17218 24324 17224 24336
rect 17147 24296 17224 24324
rect 17147 24222 17175 24296
rect 17218 24284 17224 24296
rect 17276 24284 17282 24336
rect 17420 24324 17448 24364
rect 17862 24352 17868 24404
rect 17920 24392 17926 24404
rect 18141 24395 18199 24401
rect 18141 24392 18153 24395
rect 17920 24364 18153 24392
rect 17920 24352 17926 24364
rect 18141 24361 18153 24364
rect 18187 24361 18199 24395
rect 18141 24355 18199 24361
rect 19613 24395 19671 24401
rect 19613 24361 19625 24395
rect 19659 24392 19671 24395
rect 20346 24392 20352 24404
rect 19659 24364 20352 24392
rect 19659 24361 19671 24364
rect 19613 24355 19671 24361
rect 20346 24352 20352 24364
rect 20404 24352 20410 24404
rect 20530 24352 20536 24404
rect 20588 24392 20594 24404
rect 23014 24392 23020 24404
rect 20588 24364 21864 24392
rect 20588 24352 20594 24364
rect 17773 24327 17831 24333
rect 17773 24324 17785 24327
rect 17420 24296 17785 24324
rect 17773 24293 17785 24296
rect 17819 24293 17831 24327
rect 17773 24287 17831 24293
rect 18322 24284 18328 24336
rect 18380 24324 18386 24336
rect 19334 24324 19340 24336
rect 18380 24296 19340 24324
rect 18380 24284 18386 24296
rect 19334 24284 19340 24296
rect 19392 24284 19398 24336
rect 19797 24327 19855 24333
rect 19797 24293 19809 24327
rect 19843 24293 19855 24327
rect 21174 24324 21180 24336
rect 19797 24287 19855 24293
rect 19904 24296 21180 24324
rect 17144 24197 17175 24222
rect 17402 24216 17408 24268
rect 17460 24256 17466 24268
rect 17460 24228 17954 24256
rect 17460 24216 17466 24228
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 16960 24160 17049 24188
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 17129 24191 17187 24197
rect 17129 24157 17141 24191
rect 17175 24157 17187 24191
rect 17129 24151 17187 24157
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24178 17371 24191
rect 17926 24188 17954 24228
rect 18598 24216 18604 24268
rect 18656 24256 18662 24268
rect 18877 24259 18935 24265
rect 18877 24256 18889 24259
rect 18656 24228 18889 24256
rect 18656 24216 18662 24228
rect 18877 24225 18889 24228
rect 18923 24256 18935 24259
rect 19812 24256 19840 24287
rect 18923 24228 19840 24256
rect 18923 24225 18935 24228
rect 18877 24219 18935 24225
rect 17987 24191 18045 24197
rect 17987 24188 17999 24191
rect 17359 24157 17448 24178
rect 17926 24160 17999 24188
rect 17313 24151 17448 24157
rect 17987 24157 17999 24160
rect 18033 24157 18045 24191
rect 17987 24151 18045 24157
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24188 18291 24191
rect 18690 24188 18696 24200
rect 18279 24160 18696 24188
rect 18279 24157 18291 24160
rect 18233 24151 18291 24157
rect 17329 24150 17448 24151
rect 16316 24092 17080 24120
rect 934 24012 940 24064
rect 992 24052 998 24064
rect 1581 24055 1639 24061
rect 1581 24052 1593 24055
rect 992 24024 1593 24052
rect 992 24012 998 24024
rect 1581 24021 1593 24024
rect 1627 24021 1639 24055
rect 1581 24015 1639 24021
rect 6822 24012 6828 24064
rect 6880 24012 6886 24064
rect 6917 24055 6975 24061
rect 6917 24021 6929 24055
rect 6963 24052 6975 24055
rect 7006 24052 7012 24064
rect 6963 24024 7012 24052
rect 6963 24021 6975 24024
rect 6917 24015 6975 24021
rect 7006 24012 7012 24024
rect 7064 24012 7070 24064
rect 9585 24055 9643 24061
rect 9585 24021 9597 24055
rect 9631 24052 9643 24055
rect 10042 24052 10048 24064
rect 9631 24024 10048 24052
rect 9631 24021 9643 24024
rect 9585 24015 9643 24021
rect 10042 24012 10048 24024
rect 10100 24012 10106 24064
rect 10686 24012 10692 24064
rect 10744 24052 10750 24064
rect 11149 24055 11207 24061
rect 11149 24052 11161 24055
rect 10744 24024 11161 24052
rect 10744 24012 10750 24024
rect 11149 24021 11161 24024
rect 11195 24021 11207 24055
rect 11149 24015 11207 24021
rect 11974 24012 11980 24064
rect 12032 24052 12038 24064
rect 13541 24055 13599 24061
rect 13541 24052 13553 24055
rect 12032 24024 13553 24052
rect 12032 24012 12038 24024
rect 13541 24021 13553 24024
rect 13587 24021 13599 24055
rect 13541 24015 13599 24021
rect 14461 24055 14519 24061
rect 14461 24021 14473 24055
rect 14507 24052 14519 24055
rect 14550 24052 14556 24064
rect 14507 24024 14556 24052
rect 14507 24021 14519 24024
rect 14461 24015 14519 24021
rect 14550 24012 14556 24024
rect 14608 24012 14614 24064
rect 14826 24012 14832 24064
rect 14884 24052 14890 24064
rect 15565 24055 15623 24061
rect 15565 24052 15577 24055
rect 14884 24024 15577 24052
rect 14884 24012 14890 24024
rect 15565 24021 15577 24024
rect 15611 24021 15623 24055
rect 15565 24015 15623 24021
rect 16666 24012 16672 24064
rect 16724 24052 16730 24064
rect 16945 24055 17003 24061
rect 16945 24052 16957 24055
rect 16724 24024 16957 24052
rect 16724 24012 16730 24024
rect 16945 24021 16957 24024
rect 16991 24021 17003 24055
rect 17052 24052 17080 24092
rect 17218 24080 17224 24132
rect 17276 24080 17282 24132
rect 17420 24120 17448 24150
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 19084 24182 19385 24188
rect 19084 24160 19472 24182
rect 17770 24120 17776 24132
rect 17420 24092 17776 24120
rect 17770 24080 17776 24092
rect 17828 24120 17834 24132
rect 18509 24123 18567 24129
rect 18509 24120 18521 24123
rect 17828 24092 18521 24120
rect 17828 24080 17834 24092
rect 18509 24089 18521 24092
rect 18555 24120 18567 24123
rect 19084 24120 19112 24160
rect 19357 24154 19472 24160
rect 18555 24092 19112 24120
rect 19444 24120 19472 24154
rect 19518 24148 19524 24200
rect 19576 24148 19582 24200
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24190 19763 24191
rect 19794 24190 19800 24200
rect 19751 24162 19800 24190
rect 19751 24157 19763 24162
rect 19705 24151 19763 24157
rect 19794 24148 19800 24162
rect 19852 24148 19858 24200
rect 19904 24120 19932 24296
rect 21174 24284 21180 24296
rect 21232 24284 21238 24336
rect 21361 24327 21419 24333
rect 21361 24293 21373 24327
rect 21407 24324 21419 24327
rect 21726 24324 21732 24336
rect 21407 24296 21732 24324
rect 21407 24293 21419 24296
rect 21361 24287 21419 24293
rect 21726 24284 21732 24296
rect 21784 24284 21790 24336
rect 20990 24256 20996 24268
rect 19996 24228 20996 24256
rect 19996 24197 20024 24228
rect 20990 24216 20996 24228
rect 21048 24216 21054 24268
rect 21100 24228 21404 24256
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20070 24148 20076 24200
rect 20128 24188 20134 24200
rect 20533 24191 20591 24197
rect 20533 24188 20545 24191
rect 20128 24160 20545 24188
rect 20128 24148 20134 24160
rect 20533 24157 20545 24160
rect 20579 24157 20591 24191
rect 20533 24151 20591 24157
rect 20757 24191 20815 24197
rect 20757 24157 20769 24191
rect 20803 24188 20815 24191
rect 21100 24188 21128 24228
rect 20803 24160 21128 24188
rect 21177 24191 21235 24197
rect 20803 24157 20815 24160
rect 20757 24151 20815 24157
rect 21177 24157 21189 24191
rect 21223 24188 21235 24191
rect 21266 24188 21272 24200
rect 21223 24160 21272 24188
rect 21223 24157 21235 24160
rect 21177 24151 21235 24157
rect 21266 24148 21272 24160
rect 21324 24148 21330 24200
rect 21376 24188 21404 24228
rect 21450 24216 21456 24268
rect 21508 24216 21514 24268
rect 21836 24256 21864 24364
rect 22296 24364 23020 24392
rect 22186 24284 22192 24336
rect 22244 24324 22250 24336
rect 22296 24333 22324 24364
rect 23014 24352 23020 24364
rect 23072 24352 23078 24404
rect 23201 24395 23259 24401
rect 23201 24361 23213 24395
rect 23247 24392 23259 24395
rect 23290 24392 23296 24404
rect 23247 24364 23296 24392
rect 23247 24361 23259 24364
rect 23201 24355 23259 24361
rect 23290 24352 23296 24364
rect 23348 24352 23354 24404
rect 24302 24352 24308 24404
rect 24360 24352 24366 24404
rect 24596 24364 25084 24392
rect 22281 24327 22339 24333
rect 22281 24324 22293 24327
rect 22244 24296 22293 24324
rect 22244 24284 22250 24296
rect 22281 24293 22293 24296
rect 22327 24293 22339 24327
rect 23385 24327 23443 24333
rect 23385 24324 23397 24327
rect 22281 24287 22339 24293
rect 22388 24296 23397 24324
rect 22388 24265 22416 24296
rect 23385 24293 23397 24296
rect 23431 24293 23443 24327
rect 23385 24287 23443 24293
rect 23658 24284 23664 24336
rect 23716 24324 23722 24336
rect 23753 24327 23811 24333
rect 23753 24324 23765 24327
rect 23716 24296 23765 24324
rect 23716 24284 23722 24296
rect 23753 24293 23765 24296
rect 23799 24293 23811 24327
rect 23753 24287 23811 24293
rect 23845 24327 23903 24333
rect 23845 24293 23857 24327
rect 23891 24324 23903 24327
rect 24320 24324 24348 24352
rect 23891 24296 24348 24324
rect 23891 24293 23903 24296
rect 23845 24287 23903 24293
rect 22373 24259 22431 24265
rect 21836 24228 22324 24256
rect 21634 24188 21640 24200
rect 21376 24160 21640 24188
rect 21634 24148 21640 24160
rect 21692 24148 21698 24200
rect 22094 24148 22100 24200
rect 22152 24148 22158 24200
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24157 22247 24191
rect 22296 24188 22324 24228
rect 22373 24225 22385 24259
rect 22419 24225 22431 24259
rect 24596 24256 24624 24364
rect 24670 24284 24676 24336
rect 24728 24324 24734 24336
rect 24765 24327 24823 24333
rect 24765 24324 24777 24327
rect 24728 24296 24777 24324
rect 24728 24284 24734 24296
rect 24765 24293 24777 24296
rect 24811 24293 24823 24327
rect 24765 24287 24823 24293
rect 24854 24284 24860 24336
rect 24912 24284 24918 24336
rect 24872 24256 24900 24284
rect 22373 24219 22431 24225
rect 22480 24228 24624 24256
rect 24688 24228 24900 24256
rect 22480 24197 22508 24228
rect 22465 24191 22523 24197
rect 22465 24188 22477 24191
rect 22296 24160 22477 24188
rect 22189 24151 22247 24157
rect 22465 24157 22477 24160
rect 22511 24157 22523 24191
rect 22465 24151 22523 24157
rect 19444 24092 19932 24120
rect 20349 24123 20407 24129
rect 18555 24089 18567 24092
rect 18509 24083 18567 24089
rect 20349 24089 20361 24123
rect 20395 24120 20407 24123
rect 20395 24092 20852 24120
rect 20395 24089 20407 24092
rect 20349 24083 20407 24089
rect 18966 24052 18972 24064
rect 17052 24024 18972 24052
rect 16945 24015 17003 24021
rect 18966 24012 18972 24024
rect 19024 24012 19030 24064
rect 19242 24012 19248 24064
rect 19300 24012 19306 24064
rect 19334 24012 19340 24064
rect 19392 24052 19398 24064
rect 19702 24052 19708 24064
rect 19392 24024 19708 24052
rect 19392 24012 19398 24024
rect 19702 24012 19708 24024
rect 19760 24012 19766 24064
rect 20438 24012 20444 24064
rect 20496 24052 20502 24064
rect 20625 24055 20683 24061
rect 20625 24052 20637 24055
rect 20496 24024 20637 24052
rect 20496 24012 20502 24024
rect 20625 24021 20637 24024
rect 20671 24021 20683 24055
rect 20824 24052 20852 24092
rect 20898 24080 20904 24132
rect 20956 24080 20962 24132
rect 20993 24123 21051 24129
rect 20993 24089 21005 24123
rect 21039 24120 21051 24123
rect 21450 24120 21456 24132
rect 21039 24092 21456 24120
rect 21039 24089 21051 24092
rect 20993 24083 21051 24089
rect 21450 24080 21456 24092
rect 21508 24080 21514 24132
rect 21726 24052 21732 24064
rect 20824 24024 21732 24052
rect 20625 24015 20683 24021
rect 21726 24012 21732 24024
rect 21784 24012 21790 24064
rect 22002 24012 22008 24064
rect 22060 24012 22066 24064
rect 22112 24052 22140 24148
rect 22204 24120 22232 24151
rect 22646 24148 22652 24200
rect 22704 24148 22710 24200
rect 22738 24148 22744 24200
rect 22796 24148 22802 24200
rect 23106 24148 23112 24200
rect 23164 24148 23170 24200
rect 23201 24191 23259 24197
rect 23201 24157 23213 24191
rect 23247 24188 23259 24191
rect 23474 24188 23480 24200
rect 23247 24160 23480 24188
rect 23247 24157 23259 24160
rect 23201 24151 23259 24157
rect 23474 24148 23480 24160
rect 23532 24148 23538 24200
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 23937 24191 23995 24197
rect 23937 24157 23949 24191
rect 23983 24188 23995 24191
rect 24026 24188 24032 24200
rect 23983 24160 24032 24188
rect 23983 24157 23995 24160
rect 23937 24151 23995 24157
rect 22370 24120 22376 24132
rect 22204 24092 22376 24120
rect 22370 24080 22376 24092
rect 22428 24080 22434 24132
rect 23676 24120 23704 24151
rect 24026 24148 24032 24160
rect 24084 24148 24090 24200
rect 24302 24148 24308 24200
rect 24360 24188 24366 24200
rect 24688 24197 24716 24228
rect 25056 24197 25084 24364
rect 26050 24352 26056 24404
rect 26108 24352 26114 24404
rect 26620 24364 28580 24392
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 24360 24160 24409 24188
rect 24360 24148 24366 24160
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 24397 24151 24455 24157
rect 24581 24191 24639 24197
rect 24581 24157 24593 24191
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 24673 24191 24731 24197
rect 24673 24157 24685 24191
rect 24719 24157 24731 24191
rect 24673 24151 24731 24157
rect 24857 24191 24915 24197
rect 24857 24157 24869 24191
rect 24903 24188 24915 24191
rect 25041 24191 25099 24197
rect 24903 24157 24926 24188
rect 24857 24151 24926 24157
rect 25041 24157 25053 24191
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 24596 24120 24624 24151
rect 23676 24092 24624 24120
rect 24898 24120 24926 24151
rect 26620 24120 26648 24364
rect 28552 24336 28580 24364
rect 38010 24352 38016 24404
rect 38068 24352 38074 24404
rect 26878 24284 26884 24336
rect 26936 24284 26942 24336
rect 27246 24284 27252 24336
rect 27304 24284 27310 24336
rect 27430 24284 27436 24336
rect 27488 24324 27494 24336
rect 27525 24327 27583 24333
rect 27525 24324 27537 24327
rect 27488 24296 27537 24324
rect 27488 24284 27494 24296
rect 27525 24293 27537 24296
rect 27571 24293 27583 24327
rect 27525 24287 27583 24293
rect 28534 24284 28540 24336
rect 28592 24284 28598 24336
rect 30190 24284 30196 24336
rect 30248 24284 30254 24336
rect 30926 24284 30932 24336
rect 30984 24284 30990 24336
rect 26697 24259 26755 24265
rect 26697 24225 26709 24259
rect 26743 24256 26755 24259
rect 26786 24256 26792 24268
rect 26743 24228 26792 24256
rect 26743 24225 26755 24228
rect 26697 24219 26755 24225
rect 26786 24216 26792 24228
rect 26844 24216 26850 24268
rect 26881 24191 26939 24197
rect 26881 24157 26893 24191
rect 26927 24188 26939 24191
rect 27062 24188 27068 24200
rect 26927 24160 27068 24188
rect 26927 24157 26939 24160
rect 26881 24151 26939 24157
rect 27062 24148 27068 24160
rect 27120 24148 27126 24200
rect 27157 24191 27215 24197
rect 27157 24157 27169 24191
rect 27203 24188 27215 24191
rect 27264 24188 27292 24284
rect 27617 24259 27675 24265
rect 27617 24225 27629 24259
rect 27663 24256 27675 24259
rect 29273 24259 29331 24265
rect 29273 24256 29285 24259
rect 27663 24228 29285 24256
rect 27663 24225 27675 24228
rect 27617 24219 27675 24225
rect 29273 24225 29285 24228
rect 29319 24256 29331 24259
rect 29319 24228 30236 24256
rect 29319 24225 29331 24228
rect 29273 24219 29331 24225
rect 27203 24160 27292 24188
rect 27203 24157 27215 24160
rect 27157 24151 27215 24157
rect 27430 24148 27436 24200
rect 27488 24148 27494 24200
rect 30208 24197 30236 24228
rect 30282 24216 30288 24268
rect 30340 24216 30346 24268
rect 30944 24228 32352 24256
rect 30944 24200 30972 24228
rect 32324 24200 32352 24228
rect 34790 24216 34796 24268
rect 34848 24256 34854 24268
rect 36265 24259 36323 24265
rect 36265 24256 36277 24259
rect 34848 24228 36277 24256
rect 34848 24216 34854 24228
rect 36265 24225 36277 24228
rect 36311 24256 36323 24259
rect 36311 24228 38332 24256
rect 36311 24225 36323 24228
rect 36265 24219 36323 24225
rect 38304 24200 38332 24228
rect 27709 24191 27767 24197
rect 27709 24157 27721 24191
rect 27755 24157 27767 24191
rect 29181 24191 29239 24197
rect 27709 24151 27767 24157
rect 27890 24169 27948 24175
rect 27249 24123 27307 24129
rect 27249 24120 27261 24123
rect 24898 24092 26648 24120
rect 26988 24092 27261 24120
rect 23477 24055 23535 24061
rect 23477 24052 23489 24055
rect 22112 24024 23489 24052
rect 23477 24021 23489 24024
rect 23523 24021 23535 24055
rect 24596 24052 24624 24092
rect 25866 24052 25872 24064
rect 24596 24024 25872 24052
rect 23477 24015 23535 24021
rect 25866 24012 25872 24024
rect 25924 24012 25930 24064
rect 26418 24012 26424 24064
rect 26476 24012 26482 24064
rect 26513 24055 26571 24061
rect 26513 24021 26525 24055
rect 26559 24052 26571 24055
rect 26988 24052 27016 24092
rect 27249 24089 27261 24092
rect 27295 24089 27307 24123
rect 27249 24083 27307 24089
rect 27614 24080 27620 24132
rect 27672 24120 27678 24132
rect 27724 24120 27752 24151
rect 27672 24092 27752 24120
rect 27890 24135 27902 24169
rect 27936 24135 27948 24169
rect 29181 24157 29193 24191
rect 29227 24188 29239 24191
rect 30193 24191 30251 24197
rect 29227 24160 29316 24188
rect 29227 24157 29239 24160
rect 29181 24151 29239 24157
rect 27890 24132 27948 24135
rect 29288 24132 29316 24160
rect 30193 24157 30205 24191
rect 30239 24157 30251 24191
rect 30193 24151 30251 24157
rect 30742 24148 30748 24200
rect 30800 24148 30806 24200
rect 30926 24148 30932 24200
rect 30984 24148 30990 24200
rect 31478 24148 31484 24200
rect 31536 24188 31542 24200
rect 31941 24191 31999 24197
rect 31941 24188 31953 24191
rect 31536 24160 31953 24188
rect 31536 24148 31542 24160
rect 31941 24157 31953 24160
rect 31987 24157 31999 24191
rect 31941 24151 31999 24157
rect 32306 24148 32312 24200
rect 32364 24148 32370 24200
rect 38286 24148 38292 24200
rect 38344 24148 38350 24200
rect 27672 24080 27678 24092
rect 27890 24080 27896 24132
rect 27948 24080 27954 24132
rect 29270 24080 29276 24132
rect 29328 24080 29334 24132
rect 30561 24123 30619 24129
rect 30561 24089 30573 24123
rect 30607 24120 30619 24123
rect 31570 24120 31576 24132
rect 30607 24092 31576 24120
rect 30607 24089 30619 24092
rect 30561 24083 30619 24089
rect 31570 24080 31576 24092
rect 31628 24080 31634 24132
rect 36538 24080 36544 24132
rect 36596 24080 36602 24132
rect 36998 24120 37004 24132
rect 36648 24092 37004 24120
rect 26559 24024 27016 24052
rect 26559 24021 26571 24024
rect 26513 24015 26571 24021
rect 27062 24012 27068 24064
rect 27120 24012 27126 24064
rect 27522 24012 27528 24064
rect 27580 24052 27586 24064
rect 28902 24052 28908 24064
rect 27580 24024 28908 24052
rect 27580 24012 27586 24024
rect 28902 24012 28908 24024
rect 28960 24012 28966 24064
rect 31754 24012 31760 24064
rect 31812 24012 31818 24064
rect 35802 24012 35808 24064
rect 35860 24052 35866 24064
rect 36648 24052 36676 24092
rect 36998 24080 37004 24092
rect 37056 24080 37062 24132
rect 35860 24024 36676 24052
rect 35860 24012 35866 24024
rect 1104 23962 41400 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 41400 23962
rect 1104 23888 41400 23910
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 5592 23820 5764 23848
rect 5592 23808 5598 23820
rect 4614 23740 4620 23792
rect 4672 23740 4678 23792
rect 5736 23712 5764 23820
rect 6086 23808 6092 23860
rect 6144 23808 6150 23860
rect 8754 23808 8760 23860
rect 8812 23808 8818 23860
rect 10060 23820 10364 23848
rect 6196 23752 7130 23780
rect 6196 23712 6224 23752
rect 8297 23715 8355 23721
rect 8297 23712 8309 23715
rect 5736 23698 6224 23712
rect 5750 23684 6224 23698
rect 8128 23684 8309 23712
rect 4062 23604 4068 23656
rect 4120 23644 4126 23656
rect 4341 23647 4399 23653
rect 4341 23644 4353 23647
rect 4120 23616 4353 23644
rect 4120 23604 4126 23616
rect 4341 23613 4353 23616
rect 4387 23644 4399 23647
rect 6365 23647 6423 23653
rect 6365 23644 6377 23647
rect 4387 23616 6377 23644
rect 4387 23613 4399 23616
rect 4341 23607 4399 23613
rect 6365 23613 6377 23616
rect 6411 23613 6423 23647
rect 6365 23607 6423 23613
rect 6641 23647 6699 23653
rect 6641 23613 6653 23647
rect 6687 23644 6699 23647
rect 7006 23644 7012 23656
rect 6687 23616 7012 23644
rect 6687 23613 6699 23616
rect 6641 23607 6699 23613
rect 7006 23604 7012 23616
rect 7064 23604 7070 23656
rect 8128 23653 8156 23684
rect 8297 23681 8309 23684
rect 8343 23712 8355 23715
rect 8772 23712 8800 23808
rect 10060 23789 10088 23820
rect 10045 23783 10103 23789
rect 10045 23749 10057 23783
rect 10091 23749 10103 23783
rect 10245 23783 10303 23789
rect 10245 23780 10257 23783
rect 10045 23743 10103 23749
rect 10244 23749 10257 23780
rect 10291 23749 10303 23783
rect 10244 23743 10303 23749
rect 8343 23684 8800 23712
rect 8343 23681 8355 23684
rect 8297 23675 8355 23681
rect 8113 23647 8171 23653
rect 8113 23613 8125 23647
rect 8159 23613 8171 23647
rect 8113 23607 8171 23613
rect 10244 23576 10272 23743
rect 10336 23644 10364 23820
rect 10410 23808 10416 23860
rect 10468 23808 10474 23860
rect 12161 23851 12219 23857
rect 12161 23817 12173 23851
rect 12207 23817 12219 23851
rect 13722 23848 13728 23860
rect 12161 23811 12219 23817
rect 12820 23820 13728 23848
rect 10428 23712 10456 23808
rect 12176 23780 12204 23811
rect 10796 23752 12204 23780
rect 10689 23715 10747 23721
rect 10689 23712 10701 23715
rect 10428 23684 10701 23712
rect 10689 23681 10701 23684
rect 10735 23681 10747 23715
rect 10689 23675 10747 23681
rect 10505 23647 10563 23653
rect 10505 23644 10517 23647
rect 10336 23616 10517 23644
rect 10505 23613 10517 23616
rect 10551 23644 10563 23647
rect 10594 23644 10600 23656
rect 10551 23616 10600 23644
rect 10551 23613 10563 23616
rect 10505 23607 10563 23613
rect 10594 23604 10600 23616
rect 10652 23604 10658 23656
rect 10796 23576 10824 23752
rect 11609 23715 11667 23721
rect 11609 23681 11621 23715
rect 11655 23712 11667 23715
rect 11790 23712 11796 23724
rect 11655 23684 11796 23712
rect 11655 23681 11667 23684
rect 11609 23675 11667 23681
rect 11790 23672 11796 23684
rect 11848 23672 11854 23724
rect 11974 23672 11980 23724
rect 12032 23672 12038 23724
rect 12618 23672 12624 23724
rect 12676 23712 12682 23724
rect 12820 23721 12848 23820
rect 13722 23808 13728 23820
rect 13780 23848 13786 23860
rect 14182 23848 14188 23860
rect 13780 23820 14188 23848
rect 13780 23808 13786 23820
rect 14182 23808 14188 23820
rect 14240 23848 14246 23860
rect 15289 23851 15347 23857
rect 15289 23848 15301 23851
rect 14240 23820 15301 23848
rect 14240 23808 14246 23820
rect 15289 23817 15301 23820
rect 15335 23817 15347 23851
rect 15289 23811 15347 23817
rect 15838 23808 15844 23860
rect 15896 23848 15902 23860
rect 16209 23851 16267 23857
rect 16209 23848 16221 23851
rect 15896 23820 16221 23848
rect 15896 23808 15902 23820
rect 16209 23817 16221 23820
rect 16255 23817 16267 23851
rect 16209 23811 16267 23817
rect 16776 23820 17402 23848
rect 16776 23792 16804 23820
rect 13354 23740 13360 23792
rect 13412 23740 13418 23792
rect 16758 23780 16764 23792
rect 14660 23752 16344 23780
rect 12713 23715 12771 23721
rect 12713 23712 12725 23715
rect 12676 23684 12725 23712
rect 12676 23672 12682 23684
rect 12713 23681 12725 23684
rect 12759 23681 12771 23715
rect 12713 23675 12771 23681
rect 12805 23715 12863 23721
rect 12805 23681 12817 23715
rect 12851 23681 12863 23715
rect 12805 23675 12863 23681
rect 12986 23672 12992 23724
rect 13044 23672 13050 23724
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23712 13139 23715
rect 13372 23712 13400 23740
rect 14660 23712 14688 23752
rect 13127 23684 13400 23712
rect 13464 23684 14688 23712
rect 14921 23715 14979 23721
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 10873 23647 10931 23653
rect 10873 23613 10885 23647
rect 10919 23644 10931 23647
rect 13262 23644 13268 23656
rect 10919 23616 13268 23644
rect 10919 23613 10931 23616
rect 10873 23607 10931 23613
rect 13262 23604 13268 23616
rect 13320 23604 13326 23656
rect 10244 23548 10824 23576
rect 11238 23536 11244 23588
rect 11296 23576 11302 23588
rect 13464 23576 13492 23684
rect 14921 23681 14933 23715
rect 14967 23712 14979 23715
rect 15102 23712 15108 23724
rect 14967 23684 15108 23712
rect 14967 23681 14979 23684
rect 14921 23675 14979 23681
rect 15102 23672 15108 23684
rect 15160 23672 15166 23724
rect 15930 23672 15936 23724
rect 15988 23712 15994 23724
rect 16316 23721 16344 23752
rect 16408 23752 16764 23780
rect 16117 23715 16175 23721
rect 16117 23712 16129 23715
rect 15988 23684 16129 23712
rect 15988 23672 15994 23684
rect 16117 23681 16129 23684
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23681 16359 23715
rect 16301 23675 16359 23681
rect 13630 23604 13636 23656
rect 13688 23644 13694 23656
rect 16408 23644 16436 23752
rect 16758 23740 16764 23752
rect 16816 23740 16822 23792
rect 17034 23740 17040 23792
rect 17092 23789 17098 23792
rect 17092 23780 17102 23789
rect 17092 23752 17137 23780
rect 17092 23743 17102 23752
rect 17092 23740 17098 23743
rect 17374 23721 17402 23820
rect 17678 23808 17684 23860
rect 17736 23848 17742 23860
rect 17862 23848 17868 23860
rect 17736 23820 17868 23848
rect 17736 23808 17742 23820
rect 17862 23808 17868 23820
rect 17920 23808 17926 23860
rect 18598 23808 18604 23860
rect 18656 23808 18662 23860
rect 18892 23820 19104 23848
rect 18616 23721 18644 23808
rect 18892 23780 18920 23820
rect 18800 23752 18920 23780
rect 19076 23780 19104 23820
rect 19242 23808 19248 23860
rect 19300 23848 19306 23860
rect 24670 23848 24676 23860
rect 19300 23820 24676 23848
rect 19300 23808 19306 23820
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 26234 23848 26240 23860
rect 24780 23820 26240 23848
rect 19076 23752 20668 23780
rect 18800 23721 18828 23752
rect 17353 23715 17411 23721
rect 17353 23681 17365 23715
rect 17399 23681 17411 23715
rect 17353 23675 17411 23681
rect 18601 23715 18659 23721
rect 18601 23681 18613 23715
rect 18647 23681 18659 23715
rect 18601 23675 18659 23681
rect 18785 23715 18843 23721
rect 18785 23681 18797 23715
rect 18831 23681 18843 23715
rect 18785 23675 18843 23681
rect 13688 23616 16436 23644
rect 13688 23604 13694 23616
rect 17126 23604 17132 23656
rect 17184 23604 17190 23656
rect 17221 23647 17279 23653
rect 17221 23613 17233 23647
rect 17267 23644 17279 23647
rect 17267 23616 17356 23644
rect 17267 23613 17279 23616
rect 17221 23607 17279 23613
rect 15838 23576 15844 23588
rect 11296 23548 13492 23576
rect 15304 23548 15844 23576
rect 11296 23536 11302 23548
rect 8846 23468 8852 23520
rect 8904 23468 8910 23520
rect 9122 23468 9128 23520
rect 9180 23508 9186 23520
rect 10229 23511 10287 23517
rect 10229 23508 10241 23511
rect 9180 23480 10241 23508
rect 9180 23468 9186 23480
rect 10229 23477 10241 23480
rect 10275 23477 10287 23511
rect 10229 23471 10287 23477
rect 10410 23468 10416 23520
rect 10468 23468 10474 23520
rect 11330 23468 11336 23520
rect 11388 23508 11394 23520
rect 11701 23511 11759 23517
rect 11701 23508 11713 23511
rect 11388 23480 11713 23508
rect 11388 23468 11394 23480
rect 11701 23477 11713 23480
rect 11747 23477 11759 23511
rect 11701 23471 11759 23477
rect 12526 23468 12532 23520
rect 12584 23468 12590 23520
rect 15304 23517 15332 23548
rect 15838 23536 15844 23548
rect 15896 23576 15902 23588
rect 17147 23576 17175 23604
rect 15896 23548 16896 23576
rect 15896 23536 15902 23548
rect 16868 23520 16896 23548
rect 17052 23548 17175 23576
rect 17328 23576 17356 23616
rect 17678 23604 17684 23656
rect 17736 23644 17742 23656
rect 18800 23644 18828 23675
rect 18874 23672 18880 23724
rect 18932 23672 18938 23724
rect 20162 23672 20168 23724
rect 20220 23712 20226 23724
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 20220 23684 20269 23712
rect 20220 23672 20226 23684
rect 20257 23681 20269 23684
rect 20303 23712 20315 23715
rect 20438 23712 20444 23724
rect 20303 23684 20444 23712
rect 20303 23681 20315 23684
rect 20257 23675 20315 23681
rect 20438 23672 20444 23684
rect 20496 23672 20502 23724
rect 17736 23616 18828 23644
rect 18892 23644 18920 23672
rect 19058 23644 19064 23656
rect 18892 23616 19064 23644
rect 17736 23604 17742 23616
rect 19058 23604 19064 23616
rect 19116 23644 19122 23656
rect 20533 23647 20591 23653
rect 20533 23644 20545 23647
rect 19116 23616 20545 23644
rect 19116 23604 19122 23616
rect 20272 23588 20300 23616
rect 20533 23613 20545 23616
rect 20579 23613 20591 23647
rect 20640 23644 20668 23752
rect 20806 23740 20812 23792
rect 20864 23740 20870 23792
rect 20990 23672 20996 23724
rect 21048 23672 21054 23724
rect 21266 23672 21272 23724
rect 21324 23672 21330 23724
rect 24210 23672 24216 23724
rect 24268 23672 24274 23724
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23712 24455 23715
rect 24780 23712 24808 23820
rect 26234 23808 26240 23820
rect 26292 23808 26298 23860
rect 26878 23808 26884 23860
rect 26936 23848 26942 23860
rect 26973 23851 27031 23857
rect 26973 23848 26985 23851
rect 26936 23820 26985 23848
rect 26936 23808 26942 23820
rect 26973 23817 26985 23820
rect 27019 23848 27031 23851
rect 27019 23820 27200 23848
rect 27019 23817 27031 23820
rect 26973 23811 27031 23817
rect 27172 23780 27200 23820
rect 27246 23808 27252 23860
rect 27304 23848 27310 23860
rect 29825 23851 29883 23857
rect 27304 23820 27936 23848
rect 27304 23808 27310 23820
rect 27709 23783 27767 23789
rect 27709 23780 27721 23783
rect 25516 23752 25820 23780
rect 27172 23752 27721 23780
rect 24443 23684 24808 23712
rect 24443 23681 24455 23684
rect 24397 23675 24455 23681
rect 24854 23672 24860 23724
rect 24912 23712 24918 23724
rect 25133 23715 25191 23721
rect 25516 23718 25544 23752
rect 25133 23712 25145 23715
rect 24912 23684 25145 23712
rect 24912 23672 24918 23684
rect 25133 23681 25145 23684
rect 25179 23712 25191 23715
rect 25332 23712 25544 23718
rect 25179 23690 25544 23712
rect 25179 23684 25360 23690
rect 25179 23681 25191 23684
rect 25133 23675 25191 23681
rect 25590 23672 25596 23724
rect 25648 23712 25654 23724
rect 25685 23715 25743 23721
rect 25685 23712 25697 23715
rect 25648 23684 25697 23712
rect 25648 23672 25654 23684
rect 25685 23681 25697 23684
rect 25731 23681 25743 23715
rect 25792 23712 25820 23752
rect 27709 23749 27721 23752
rect 27755 23749 27767 23783
rect 27709 23743 27767 23749
rect 27908 23780 27936 23820
rect 29825 23817 29837 23851
rect 29871 23848 29883 23851
rect 30926 23848 30932 23860
rect 29871 23820 30932 23848
rect 29871 23817 29883 23820
rect 29825 23811 29883 23817
rect 30926 23808 30932 23820
rect 30984 23808 30990 23860
rect 32233 23820 32812 23848
rect 28258 23780 28264 23792
rect 27908 23752 28264 23780
rect 25961 23715 26019 23721
rect 25961 23712 25973 23715
rect 25792 23684 25973 23712
rect 25685 23675 25743 23681
rect 25961 23681 25973 23684
rect 26007 23712 26019 23715
rect 26142 23712 26148 23724
rect 26007 23684 26148 23712
rect 26007 23681 26019 23684
rect 25961 23675 26019 23681
rect 26142 23672 26148 23684
rect 26200 23672 26206 23724
rect 26326 23672 26332 23724
rect 26384 23712 26390 23724
rect 27908 23721 27936 23752
rect 28258 23740 28264 23752
rect 28316 23740 28322 23792
rect 32233 23780 32261 23820
rect 31510 23752 32261 23780
rect 32784 23780 32812 23820
rect 33042 23808 33048 23860
rect 33100 23848 33106 23860
rect 34698 23848 34704 23860
rect 33100 23820 34704 23848
rect 33100 23808 33106 23820
rect 34698 23808 34704 23820
rect 34756 23848 34762 23860
rect 35989 23851 36047 23857
rect 35989 23848 36001 23851
rect 34756 23820 36001 23848
rect 34756 23808 34762 23820
rect 35989 23817 36001 23820
rect 36035 23817 36047 23851
rect 35989 23811 36047 23817
rect 36538 23808 36544 23860
rect 36596 23848 36602 23860
rect 37277 23851 37335 23857
rect 37277 23848 37289 23851
rect 36596 23820 37289 23848
rect 36596 23808 36602 23820
rect 37277 23817 37289 23820
rect 37323 23817 37335 23851
rect 38010 23848 38016 23860
rect 37277 23811 37335 23817
rect 37568 23820 38016 23848
rect 34054 23780 34060 23792
rect 32784 23752 32890 23780
rect 33534 23752 34060 23780
rect 34054 23740 34060 23752
rect 34112 23740 34118 23792
rect 34790 23780 34796 23792
rect 34256 23752 34796 23780
rect 26513 23715 26571 23721
rect 26513 23712 26525 23715
rect 26384 23684 26525 23712
rect 26384 23672 26390 23684
rect 26513 23681 26525 23684
rect 26559 23712 26571 23715
rect 27893 23715 27951 23721
rect 26559 23684 27016 23712
rect 26559 23681 26571 23684
rect 26513 23675 26571 23681
rect 20640 23616 21036 23644
rect 20533 23607 20591 23613
rect 18506 23576 18512 23588
rect 17328 23548 18512 23576
rect 15289 23511 15347 23517
rect 15289 23477 15301 23511
rect 15335 23477 15347 23511
rect 15289 23471 15347 23477
rect 15378 23468 15384 23520
rect 15436 23508 15442 23520
rect 15473 23511 15531 23517
rect 15473 23508 15485 23511
rect 15436 23480 15485 23508
rect 15436 23468 15442 23480
rect 15473 23477 15485 23480
rect 15519 23477 15531 23511
rect 15473 23471 15531 23477
rect 15562 23468 15568 23520
rect 15620 23508 15626 23520
rect 16758 23508 16764 23520
rect 15620 23480 16764 23508
rect 15620 23468 15626 23480
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 16850 23468 16856 23520
rect 16908 23468 16914 23520
rect 17052 23517 17080 23548
rect 18506 23536 18512 23548
rect 18564 23536 18570 23588
rect 18693 23579 18751 23585
rect 18693 23545 18705 23579
rect 18739 23576 18751 23579
rect 18966 23576 18972 23588
rect 18739 23548 18972 23576
rect 18739 23545 18751 23548
rect 18693 23539 18751 23545
rect 18966 23536 18972 23548
rect 19024 23576 19030 23588
rect 19886 23576 19892 23588
rect 19024 23548 19892 23576
rect 19024 23536 19030 23548
rect 19886 23536 19892 23548
rect 19944 23536 19950 23588
rect 20254 23536 20260 23588
rect 20312 23536 20318 23588
rect 20349 23579 20407 23585
rect 20349 23545 20361 23579
rect 20395 23576 20407 23579
rect 21008 23576 21036 23616
rect 21082 23604 21088 23656
rect 21140 23604 21146 23656
rect 21174 23604 21180 23656
rect 21232 23604 21238 23656
rect 23290 23604 23296 23656
rect 23348 23644 23354 23656
rect 24486 23644 24492 23656
rect 23348 23616 24492 23644
rect 23348 23604 23354 23616
rect 24486 23604 24492 23616
rect 24544 23604 24550 23656
rect 25409 23647 25467 23653
rect 25409 23644 25421 23647
rect 25332 23616 25421 23644
rect 24581 23579 24639 23585
rect 24581 23576 24593 23579
rect 20395 23548 20944 23576
rect 21008 23548 24593 23576
rect 20395 23545 20407 23548
rect 20349 23539 20407 23545
rect 17037 23511 17095 23517
rect 17037 23477 17049 23511
rect 17083 23477 17095 23511
rect 17037 23471 17095 23477
rect 17126 23468 17132 23520
rect 17184 23508 17190 23520
rect 17497 23511 17555 23517
rect 17497 23508 17509 23511
rect 17184 23480 17509 23508
rect 17184 23468 17190 23480
rect 17497 23477 17509 23480
rect 17543 23477 17555 23511
rect 17497 23471 17555 23477
rect 18414 23468 18420 23520
rect 18472 23468 18478 23520
rect 18524 23508 18552 23536
rect 18874 23508 18880 23520
rect 18524 23480 18880 23508
rect 18874 23468 18880 23480
rect 18932 23468 18938 23520
rect 20438 23468 20444 23520
rect 20496 23468 20502 23520
rect 20916 23508 20944 23548
rect 24581 23545 24593 23548
rect 24627 23545 24639 23579
rect 24581 23539 24639 23545
rect 24670 23536 24676 23588
rect 24728 23576 24734 23588
rect 25332 23576 25360 23616
rect 25409 23613 25421 23616
rect 25455 23613 25467 23647
rect 25409 23607 25467 23613
rect 25501 23647 25559 23653
rect 25501 23613 25513 23647
rect 25547 23644 25559 23647
rect 26694 23644 26700 23656
rect 25547 23616 26700 23644
rect 25547 23613 25559 23616
rect 25501 23607 25559 23613
rect 26694 23604 26700 23616
rect 26752 23604 26758 23656
rect 26789 23647 26847 23653
rect 26789 23613 26801 23647
rect 26835 23644 26847 23647
rect 26878 23644 26884 23656
rect 26835 23616 26884 23644
rect 26835 23613 26847 23616
rect 26789 23607 26847 23613
rect 26878 23604 26884 23616
rect 26936 23604 26942 23656
rect 26988 23644 27016 23684
rect 27893 23681 27905 23715
rect 27939 23681 27951 23715
rect 27893 23675 27951 23681
rect 27982 23672 27988 23724
rect 28040 23712 28046 23724
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 28040 23684 29745 23712
rect 28040 23672 28046 23684
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 31754 23672 31760 23724
rect 31812 23672 31818 23724
rect 34256 23721 34284 23752
rect 34790 23740 34796 23752
rect 34848 23740 34854 23792
rect 35802 23780 35808 23792
rect 35742 23752 35808 23780
rect 35802 23740 35808 23752
rect 35860 23740 35866 23792
rect 37568 23780 37596 23820
rect 38010 23808 38016 23820
rect 38068 23808 38074 23860
rect 36556 23752 37596 23780
rect 36556 23721 36584 23752
rect 37734 23740 37740 23792
rect 37792 23740 37798 23792
rect 32125 23715 32183 23721
rect 32125 23681 32137 23715
rect 32171 23712 32183 23715
rect 34241 23715 34299 23721
rect 32171 23684 32628 23712
rect 32171 23681 32183 23684
rect 32125 23675 32183 23681
rect 27341 23647 27399 23653
rect 27341 23644 27353 23647
rect 26988 23616 27353 23644
rect 27341 23613 27353 23616
rect 27387 23613 27399 23647
rect 27341 23607 27399 23613
rect 27433 23647 27491 23653
rect 27433 23613 27445 23647
rect 27479 23644 27491 23647
rect 27522 23644 27528 23656
rect 27479 23616 27528 23644
rect 27479 23613 27491 23616
rect 27433 23607 27491 23613
rect 27522 23604 27528 23616
rect 27580 23644 27586 23656
rect 29178 23644 29184 23656
rect 27580 23616 29184 23644
rect 27580 23604 27586 23616
rect 29178 23604 29184 23616
rect 29236 23604 29242 23656
rect 30006 23604 30012 23656
rect 30064 23604 30070 23656
rect 30285 23647 30343 23653
rect 30285 23613 30297 23647
rect 30331 23644 30343 23647
rect 30650 23644 30656 23656
rect 30331 23616 30656 23644
rect 30331 23613 30343 23616
rect 30285 23607 30343 23613
rect 30650 23604 30656 23616
rect 30708 23604 30714 23656
rect 31772 23644 31800 23672
rect 32493 23647 32551 23653
rect 32493 23644 32505 23647
rect 31772 23616 32505 23644
rect 32493 23613 32505 23616
rect 32539 23613 32551 23647
rect 32600 23644 32628 23684
rect 34241 23681 34253 23715
rect 34287 23681 34299 23715
rect 34241 23675 34299 23681
rect 36541 23715 36599 23721
rect 36541 23681 36553 23715
rect 36587 23681 36599 23715
rect 36541 23675 36599 23681
rect 37461 23715 37519 23721
rect 37461 23681 37473 23715
rect 37507 23681 37519 23715
rect 37461 23675 37519 23681
rect 32674 23644 32680 23656
rect 32600 23616 32680 23644
rect 32493 23607 32551 23613
rect 32674 23604 32680 23616
rect 32732 23604 32738 23656
rect 34514 23604 34520 23656
rect 34572 23604 34578 23656
rect 36630 23604 36636 23656
rect 36688 23604 36694 23656
rect 36722 23604 36728 23656
rect 36780 23604 36786 23656
rect 25590 23576 25596 23588
rect 24728 23548 25360 23576
rect 25516 23548 25596 23576
rect 24728 23536 24734 23548
rect 23106 23508 23112 23520
rect 20916 23480 23112 23508
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 23658 23468 23664 23520
rect 23716 23508 23722 23520
rect 24213 23511 24271 23517
rect 24213 23508 24225 23511
rect 23716 23480 24225 23508
rect 23716 23468 23722 23480
rect 24213 23477 24225 23480
rect 24259 23477 24271 23511
rect 24213 23471 24271 23477
rect 24762 23468 24768 23520
rect 24820 23508 24826 23520
rect 24949 23511 25007 23517
rect 24949 23508 24961 23511
rect 24820 23480 24961 23508
rect 24820 23468 24826 23480
rect 24949 23477 24961 23480
rect 24995 23477 25007 23511
rect 24949 23471 25007 23477
rect 25317 23511 25375 23517
rect 25317 23477 25329 23511
rect 25363 23508 25375 23511
rect 25516 23508 25544 23548
rect 25590 23536 25596 23548
rect 25648 23576 25654 23588
rect 25777 23579 25835 23585
rect 25777 23576 25789 23579
rect 25648 23548 25789 23576
rect 25648 23536 25654 23548
rect 25777 23545 25789 23548
rect 25823 23545 25835 23579
rect 25777 23539 25835 23545
rect 25869 23579 25927 23585
rect 25869 23545 25881 23579
rect 25915 23576 25927 23579
rect 27617 23579 27675 23585
rect 27617 23576 27629 23579
rect 25915 23548 27629 23576
rect 25915 23545 25927 23548
rect 25869 23539 25927 23545
rect 27617 23545 27629 23548
rect 27663 23545 27675 23579
rect 27617 23539 27675 23545
rect 31757 23579 31815 23585
rect 31757 23545 31769 23579
rect 31803 23576 31815 23579
rect 31846 23576 31852 23588
rect 31803 23548 31852 23576
rect 31803 23545 31815 23548
rect 31757 23539 31815 23545
rect 31846 23536 31852 23548
rect 31904 23536 31910 23588
rect 36173 23579 36231 23585
rect 36173 23545 36185 23579
rect 36219 23576 36231 23579
rect 37476 23576 37504 23675
rect 38286 23604 38292 23656
rect 38344 23644 38350 23656
rect 38473 23647 38531 23653
rect 38473 23644 38485 23647
rect 38344 23616 38485 23644
rect 38344 23604 38350 23616
rect 38473 23613 38485 23616
rect 38519 23613 38531 23647
rect 38473 23607 38531 23613
rect 36219 23548 37504 23576
rect 36219 23545 36231 23548
rect 36173 23539 36231 23545
rect 25363 23480 25544 23508
rect 25363 23477 25375 23480
rect 25317 23471 25375 23477
rect 26326 23468 26332 23520
rect 26384 23468 26390 23520
rect 26418 23468 26424 23520
rect 26476 23508 26482 23520
rect 26697 23511 26755 23517
rect 26697 23508 26709 23511
rect 26476 23480 26709 23508
rect 26476 23468 26482 23480
rect 26697 23477 26709 23480
rect 26743 23477 26755 23511
rect 26697 23471 26755 23477
rect 26786 23468 26792 23520
rect 26844 23508 26850 23520
rect 28077 23511 28135 23517
rect 28077 23508 28089 23511
rect 26844 23480 28089 23508
rect 26844 23468 26850 23480
rect 28077 23477 28089 23480
rect 28123 23477 28135 23511
rect 28077 23471 28135 23477
rect 32398 23468 32404 23520
rect 32456 23508 32462 23520
rect 33873 23511 33931 23517
rect 33873 23508 33885 23511
rect 32456 23480 33885 23508
rect 32456 23468 32462 23480
rect 33873 23477 33885 23480
rect 33919 23477 33931 23511
rect 33873 23471 33931 23477
rect 1104 23418 41400 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 41400 23418
rect 1104 23344 41400 23366
rect 1394 23264 1400 23316
rect 1452 23304 1458 23316
rect 2041 23307 2099 23313
rect 2041 23304 2053 23307
rect 1452 23276 2053 23304
rect 1452 23264 1458 23276
rect 2041 23273 2053 23276
rect 2087 23273 2099 23307
rect 2041 23267 2099 23273
rect 4614 23264 4620 23316
rect 4672 23304 4678 23316
rect 5077 23307 5135 23313
rect 5077 23304 5089 23307
rect 4672 23276 5089 23304
rect 4672 23264 4678 23276
rect 5077 23273 5089 23276
rect 5123 23273 5135 23307
rect 5077 23267 5135 23273
rect 7098 23264 7104 23316
rect 7156 23264 7162 23316
rect 11422 23264 11428 23316
rect 11480 23304 11486 23316
rect 11698 23304 11704 23316
rect 11480 23276 11704 23304
rect 11480 23264 11486 23276
rect 11698 23264 11704 23276
rect 11756 23264 11762 23316
rect 12894 23264 12900 23316
rect 12952 23264 12958 23316
rect 14829 23307 14887 23313
rect 14829 23273 14841 23307
rect 14875 23304 14887 23307
rect 17126 23304 17132 23316
rect 14875 23276 17132 23304
rect 14875 23273 14887 23276
rect 14829 23267 14887 23273
rect 17126 23264 17132 23276
rect 17184 23264 17190 23316
rect 20717 23307 20775 23313
rect 17236 23276 20392 23304
rect 9214 23236 9220 23248
rect 6380 23208 9220 23236
rect 6380 23177 6408 23208
rect 9214 23196 9220 23208
rect 9272 23196 9278 23248
rect 10413 23239 10471 23245
rect 10413 23205 10425 23239
rect 10459 23236 10471 23239
rect 10594 23236 10600 23248
rect 10459 23208 10600 23236
rect 10459 23205 10471 23208
rect 10413 23199 10471 23205
rect 10594 23196 10600 23208
rect 10652 23196 10658 23248
rect 12912 23236 12940 23264
rect 15562 23236 15568 23248
rect 12912 23208 15568 23236
rect 6365 23171 6423 23177
rect 6365 23137 6377 23171
rect 6411 23137 6423 23171
rect 6365 23131 6423 23137
rect 7745 23171 7803 23177
rect 7745 23137 7757 23171
rect 7791 23168 7803 23171
rect 7834 23168 7840 23180
rect 7791 23140 7840 23168
rect 7791 23137 7803 23140
rect 7745 23131 7803 23137
rect 7834 23128 7840 23140
rect 7892 23128 7898 23180
rect 8846 23128 8852 23180
rect 8904 23128 8910 23180
rect 12434 23168 12440 23180
rect 9048 23140 12440 23168
rect 1854 23060 1860 23112
rect 1912 23060 1918 23112
rect 5261 23103 5319 23109
rect 5261 23069 5273 23103
rect 5307 23100 5319 23103
rect 6089 23103 6147 23109
rect 5307 23072 5764 23100
rect 5307 23069 5319 23072
rect 5261 23063 5319 23069
rect 5736 22973 5764 23072
rect 6089 23069 6101 23103
rect 6135 23100 6147 23103
rect 6822 23100 6828 23112
rect 6135 23072 6828 23100
rect 6135 23069 6147 23072
rect 6089 23063 6147 23069
rect 6822 23060 6828 23072
rect 6880 23060 6886 23112
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23100 7619 23103
rect 8864 23100 8892 23128
rect 9048 23109 9076 23140
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 13078 23128 13084 23180
rect 13136 23168 13142 23180
rect 13136 23140 15424 23168
rect 13136 23128 13142 23140
rect 7607 23072 8892 23100
rect 9033 23103 9091 23109
rect 7607 23069 7619 23072
rect 7561 23063 7619 23069
rect 9033 23069 9045 23103
rect 9079 23069 9091 23103
rect 9033 23063 9091 23069
rect 10042 23060 10048 23112
rect 10100 23100 10106 23112
rect 10597 23103 10655 23109
rect 10597 23100 10609 23103
rect 10100 23072 10609 23100
rect 10100 23060 10106 23072
rect 10597 23069 10609 23072
rect 10643 23069 10655 23103
rect 10597 23063 10655 23069
rect 10686 23060 10692 23112
rect 10744 23060 10750 23112
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23100 10839 23103
rect 13906 23100 13912 23112
rect 10827 23072 13912 23100
rect 10827 23069 10839 23072
rect 10781 23063 10839 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 14737 23103 14795 23109
rect 14737 23069 14749 23103
rect 14783 23069 14795 23103
rect 14737 23063 14795 23069
rect 14921 23103 14979 23109
rect 14921 23069 14933 23103
rect 14967 23069 14979 23103
rect 14921 23063 14979 23069
rect 8018 23032 8024 23044
rect 6196 23004 8024 23032
rect 6196 22973 6224 23004
rect 8018 22992 8024 23004
rect 8076 22992 8082 23044
rect 9306 23032 9312 23044
rect 9232 23004 9312 23032
rect 5721 22967 5779 22973
rect 5721 22933 5733 22967
rect 5767 22933 5779 22967
rect 5721 22927 5779 22933
rect 6181 22967 6239 22973
rect 6181 22933 6193 22967
rect 6227 22933 6239 22967
rect 6181 22927 6239 22933
rect 7469 22967 7527 22973
rect 7469 22933 7481 22967
rect 7515 22964 7527 22967
rect 8110 22964 8116 22976
rect 7515 22936 8116 22964
rect 7515 22933 7527 22936
rect 7469 22927 7527 22933
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 9232 22973 9260 23004
rect 9306 22992 9312 23004
rect 9364 23032 9370 23044
rect 11149 23035 11207 23041
rect 11149 23032 11161 23035
rect 9364 23004 11161 23032
rect 9364 22992 9370 23004
rect 11149 23001 11161 23004
rect 11195 23032 11207 23035
rect 13078 23032 13084 23044
rect 11195 23004 13084 23032
rect 11195 23001 11207 23004
rect 11149 22995 11207 23001
rect 13078 22992 13084 23004
rect 13136 22992 13142 23044
rect 13262 22992 13268 23044
rect 13320 23032 13326 23044
rect 14752 23032 14780 23063
rect 13320 23004 14780 23032
rect 14936 23032 14964 23063
rect 15010 23060 15016 23112
rect 15068 23060 15074 23112
rect 15197 23103 15255 23109
rect 15197 23069 15209 23103
rect 15243 23100 15255 23103
rect 15286 23100 15292 23112
rect 15243 23072 15292 23100
rect 15243 23069 15255 23072
rect 15197 23063 15255 23069
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 15396 23032 15424 23140
rect 15488 23109 15516 23208
rect 15562 23196 15568 23208
rect 15620 23196 15626 23248
rect 16022 23236 16028 23248
rect 15672 23208 16028 23236
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23069 15531 23103
rect 15473 23063 15531 23069
rect 15565 23103 15623 23109
rect 15565 23069 15577 23103
rect 15611 23100 15623 23103
rect 15672 23100 15700 23208
rect 16022 23196 16028 23208
rect 16080 23196 16086 23248
rect 16758 23196 16764 23248
rect 16816 23236 16822 23248
rect 17236 23236 17264 23276
rect 20364 23248 20392 23276
rect 20717 23273 20729 23307
rect 20763 23304 20775 23307
rect 27982 23304 27988 23316
rect 20763 23276 27988 23304
rect 20763 23273 20775 23276
rect 20717 23267 20775 23273
rect 27982 23264 27988 23276
rect 28040 23264 28046 23316
rect 30006 23264 30012 23316
rect 30064 23304 30070 23316
rect 32674 23304 32680 23316
rect 30064 23276 32680 23304
rect 30064 23264 30070 23276
rect 32674 23264 32680 23276
rect 32732 23264 32738 23316
rect 16816 23208 17264 23236
rect 16816 23196 16822 23208
rect 17402 23196 17408 23248
rect 17460 23236 17466 23248
rect 20073 23239 20131 23245
rect 20073 23236 20085 23239
rect 17460 23208 20085 23236
rect 17460 23196 17466 23208
rect 20073 23205 20085 23208
rect 20119 23205 20131 23239
rect 20073 23199 20131 23205
rect 20346 23196 20352 23248
rect 20404 23236 20410 23248
rect 20441 23239 20499 23245
rect 20441 23236 20453 23239
rect 20404 23208 20453 23236
rect 20404 23196 20410 23208
rect 20441 23205 20453 23208
rect 20487 23236 20499 23239
rect 21174 23236 21180 23248
rect 20487 23208 21180 23236
rect 20487 23205 20499 23208
rect 20441 23199 20499 23205
rect 21174 23196 21180 23208
rect 21232 23196 21238 23248
rect 24026 23236 24032 23248
rect 23400 23208 24032 23236
rect 16301 23171 16359 23177
rect 16301 23168 16313 23171
rect 15764 23140 16313 23168
rect 15764 23109 15792 23140
rect 16301 23137 16313 23140
rect 16347 23137 16359 23171
rect 17678 23168 17684 23180
rect 16301 23131 16359 23137
rect 16868 23140 17684 23168
rect 15611 23072 15700 23100
rect 15749 23103 15807 23109
rect 15611 23069 15623 23072
rect 15565 23063 15623 23069
rect 15749 23069 15761 23103
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 15841 23103 15899 23109
rect 15841 23069 15853 23103
rect 15887 23069 15899 23103
rect 15841 23063 15899 23069
rect 15580 23032 15608 23063
rect 14936 23004 15332 23032
rect 15396 23004 15608 23032
rect 15856 23032 15884 23063
rect 16022 23060 16028 23112
rect 16080 23060 16086 23112
rect 16117 23103 16175 23109
rect 16117 23069 16129 23103
rect 16163 23100 16175 23103
rect 16868 23100 16896 23140
rect 17678 23128 17684 23140
rect 17736 23128 17742 23180
rect 17972 23140 22508 23168
rect 16163 23072 16896 23100
rect 16163 23069 16175 23072
rect 16117 23063 16175 23069
rect 16942 23060 16948 23112
rect 17000 23100 17006 23112
rect 17972 23109 18000 23140
rect 22480 23112 22508 23140
rect 22738 23128 22744 23180
rect 22796 23168 22802 23180
rect 23400 23168 23428 23208
rect 24026 23196 24032 23208
rect 24084 23196 24090 23248
rect 25038 23196 25044 23248
rect 25096 23196 25102 23248
rect 25222 23196 25228 23248
rect 25280 23196 25286 23248
rect 27522 23236 27528 23248
rect 26206 23208 27528 23236
rect 23842 23168 23848 23180
rect 22796 23140 23428 23168
rect 22796 23128 22802 23140
rect 17773 23103 17831 23109
rect 17773 23100 17785 23103
rect 17000 23072 17785 23100
rect 17000 23060 17006 23072
rect 17773 23069 17785 23072
rect 17819 23069 17831 23103
rect 17773 23063 17831 23069
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 18598 23060 18604 23112
rect 18656 23100 18662 23112
rect 19058 23100 19064 23112
rect 18656 23072 19064 23100
rect 18656 23060 18662 23072
rect 19058 23060 19064 23072
rect 19116 23060 19122 23112
rect 20070 23060 20076 23112
rect 20128 23100 20134 23112
rect 20257 23103 20315 23109
rect 20257 23100 20269 23103
rect 20128 23072 20269 23100
rect 20128 23060 20134 23072
rect 20257 23069 20269 23072
rect 20303 23069 20315 23103
rect 20257 23063 20315 23069
rect 20349 23103 20407 23109
rect 20349 23069 20361 23103
rect 20395 23100 20407 23103
rect 20533 23103 20591 23109
rect 20395 23072 20484 23100
rect 20395 23069 20407 23072
rect 20349 23063 20407 23069
rect 20162 23032 20168 23044
rect 15856 23004 20168 23032
rect 13320 22992 13326 23004
rect 9217 22967 9275 22973
rect 9217 22933 9229 22967
rect 9263 22933 9275 22967
rect 9217 22927 9275 22933
rect 10965 22967 11023 22973
rect 10965 22933 10977 22967
rect 11011 22964 11023 22967
rect 11054 22964 11060 22976
rect 11011 22936 11060 22964
rect 11011 22933 11023 22936
rect 10965 22927 11023 22933
rect 11054 22924 11060 22936
rect 11112 22924 11118 22976
rect 11882 22924 11888 22976
rect 11940 22964 11946 22976
rect 14274 22964 14280 22976
rect 11940 22936 14280 22964
rect 11940 22924 11946 22936
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 14458 22924 14464 22976
rect 14516 22924 14522 22976
rect 15304 22973 15332 23004
rect 15289 22967 15347 22973
rect 15289 22933 15301 22967
rect 15335 22964 15347 22967
rect 15470 22964 15476 22976
rect 15335 22936 15476 22964
rect 15335 22933 15347 22936
rect 15289 22927 15347 22933
rect 15470 22924 15476 22936
rect 15528 22924 15534 22976
rect 15562 22924 15568 22976
rect 15620 22964 15626 22976
rect 15856 22964 15884 23004
rect 20162 22992 20168 23004
rect 20220 22992 20226 23044
rect 15620 22936 15884 22964
rect 15620 22924 15626 22936
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 17770 22964 17776 22976
rect 16724 22936 17776 22964
rect 16724 22924 16730 22936
rect 17770 22924 17776 22936
rect 17828 22924 17834 22976
rect 18138 22924 18144 22976
rect 18196 22924 18202 22976
rect 18782 22924 18788 22976
rect 18840 22964 18846 22976
rect 19058 22964 19064 22976
rect 18840 22936 19064 22964
rect 18840 22924 18846 22936
rect 19058 22924 19064 22936
rect 19116 22964 19122 22976
rect 20346 22964 20352 22976
rect 19116 22936 20352 22964
rect 19116 22924 19122 22936
rect 20346 22924 20352 22936
rect 20404 22924 20410 22976
rect 20456 22964 20484 23072
rect 20533 23069 20545 23103
rect 20579 23100 20591 23103
rect 20622 23100 20628 23112
rect 20579 23072 20628 23100
rect 20579 23069 20591 23072
rect 20533 23063 20591 23069
rect 20622 23060 20628 23072
rect 20680 23060 20686 23112
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 20901 23103 20959 23109
rect 20901 23100 20913 23103
rect 20864 23072 20913 23100
rect 20864 23060 20870 23072
rect 20901 23069 20913 23072
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 20990 23060 20996 23112
rect 21048 23060 21054 23112
rect 21082 23060 21088 23112
rect 21140 23060 21146 23112
rect 21174 23060 21180 23112
rect 21232 23060 21238 23112
rect 22462 23060 22468 23112
rect 22520 23100 22526 23112
rect 23400 23109 23428 23140
rect 23492 23140 23848 23168
rect 23492 23109 23520 23140
rect 23842 23128 23848 23140
rect 23900 23128 23906 23180
rect 23201 23103 23259 23109
rect 23201 23100 23213 23103
rect 22520 23072 23213 23100
rect 22520 23060 22526 23072
rect 23201 23069 23213 23072
rect 23247 23069 23259 23103
rect 23201 23063 23259 23069
rect 23385 23103 23443 23109
rect 23385 23069 23397 23103
rect 23431 23069 23443 23103
rect 23385 23063 23443 23069
rect 23477 23103 23535 23109
rect 23477 23069 23489 23103
rect 23523 23069 23535 23103
rect 24044 23100 24072 23196
rect 24949 23103 25007 23109
rect 24949 23100 24961 23103
rect 24044 23072 24961 23100
rect 23477 23063 23535 23069
rect 24949 23069 24961 23072
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 25133 23103 25191 23109
rect 25133 23069 25145 23103
rect 25179 23069 25191 23103
rect 25133 23063 25191 23069
rect 20640 23032 20668 23060
rect 21358 23032 21364 23044
rect 20640 23004 21364 23032
rect 21358 22992 21364 23004
rect 21416 22992 21422 23044
rect 23017 23035 23075 23041
rect 23017 23001 23029 23035
rect 23063 23032 23075 23035
rect 23658 23032 23664 23044
rect 23063 23004 23664 23032
rect 23063 23001 23075 23004
rect 23017 22995 23075 23001
rect 23658 22992 23664 23004
rect 23716 22992 23722 23044
rect 24578 22992 24584 23044
rect 24636 23032 24642 23044
rect 25148 23032 25176 23063
rect 25222 23060 25228 23112
rect 25280 23100 25286 23112
rect 25409 23103 25467 23109
rect 25409 23100 25421 23103
rect 25280 23072 25421 23100
rect 25280 23060 25286 23072
rect 25409 23069 25421 23072
rect 25455 23100 25467 23103
rect 26206 23100 26234 23208
rect 27522 23196 27528 23208
rect 27580 23196 27586 23248
rect 27706 23196 27712 23248
rect 27764 23196 27770 23248
rect 27893 23239 27951 23245
rect 27893 23205 27905 23239
rect 27939 23236 27951 23239
rect 29825 23239 29883 23245
rect 27939 23208 29040 23236
rect 27939 23205 27951 23208
rect 27893 23199 27951 23205
rect 26344 23140 27292 23168
rect 26344 23112 26372 23140
rect 25455 23072 26234 23100
rect 25455 23069 25467 23072
rect 25409 23063 25467 23069
rect 26326 23060 26332 23112
rect 26384 23060 26390 23112
rect 27264 23109 27292 23140
rect 27430 23128 27436 23180
rect 27488 23128 27494 23180
rect 27724 23109 27752 23196
rect 29012 23180 29040 23208
rect 29825 23205 29837 23239
rect 29871 23205 29883 23239
rect 29825 23199 29883 23205
rect 28994 23128 29000 23180
rect 29052 23128 29058 23180
rect 26973 23103 27031 23109
rect 26973 23069 26985 23103
rect 27019 23069 27031 23103
rect 26973 23063 27031 23069
rect 27249 23103 27307 23109
rect 27249 23069 27261 23103
rect 27295 23069 27307 23103
rect 27249 23063 27307 23069
rect 27525 23103 27583 23109
rect 27525 23069 27537 23103
rect 27571 23069 27583 23103
rect 27525 23063 27583 23069
rect 27709 23103 27767 23109
rect 27709 23069 27721 23103
rect 27755 23069 27767 23103
rect 27709 23063 27767 23069
rect 27985 23103 28043 23109
rect 27985 23069 27997 23103
rect 28031 23069 28043 23103
rect 28169 23103 28227 23109
rect 28169 23100 28181 23103
rect 27985 23063 28043 23069
rect 28092 23072 28181 23100
rect 25774 23032 25780 23044
rect 24636 23004 25780 23032
rect 24636 22992 24642 23004
rect 25774 22992 25780 23004
rect 25832 22992 25838 23044
rect 26418 22992 26424 23044
rect 26476 22992 26482 23044
rect 26988 23032 27016 23063
rect 27540 23032 27568 23063
rect 26988 23004 27568 23032
rect 27724 23032 27752 23063
rect 28000 23032 28028 23063
rect 27724 23004 28028 23032
rect 23290 22964 23296 22976
rect 20456 22936 23296 22964
rect 23290 22924 23296 22936
rect 23348 22924 23354 22976
rect 23566 22924 23572 22976
rect 23624 22964 23630 22976
rect 24673 22967 24731 22973
rect 24673 22964 24685 22967
rect 23624 22936 24685 22964
rect 23624 22924 23630 22936
rect 24673 22933 24685 22936
rect 24719 22933 24731 22967
rect 24673 22927 24731 22933
rect 24854 22924 24860 22976
rect 24912 22964 24918 22976
rect 26988 22964 27016 23004
rect 24912 22936 27016 22964
rect 27540 22964 27568 23004
rect 28092 22964 28120 23072
rect 28169 23069 28181 23072
rect 28215 23069 28227 23103
rect 28169 23063 28227 23069
rect 28258 23060 28264 23112
rect 28316 23100 28322 23112
rect 28721 23103 28779 23109
rect 28721 23100 28733 23103
rect 28316 23072 28733 23100
rect 28316 23060 28322 23072
rect 28721 23069 28733 23072
rect 28767 23069 28779 23103
rect 28721 23063 28779 23069
rect 28810 23060 28816 23112
rect 28868 23060 28874 23112
rect 28905 23103 28963 23109
rect 28905 23069 28917 23103
rect 28951 23069 28963 23103
rect 28905 23063 28963 23069
rect 28920 23032 28948 23063
rect 29086 23060 29092 23112
rect 29144 23100 29150 23112
rect 29546 23100 29552 23112
rect 29144 23072 29552 23100
rect 29144 23060 29150 23072
rect 29546 23060 29552 23072
rect 29604 23060 29610 23112
rect 29840 23100 29868 23199
rect 29914 23196 29920 23248
rect 29972 23236 29978 23248
rect 29972 23208 30328 23236
rect 29972 23196 29978 23208
rect 30300 23177 30328 23208
rect 30650 23196 30656 23248
rect 30708 23196 30714 23248
rect 31570 23196 31576 23248
rect 31628 23196 31634 23248
rect 30285 23171 30343 23177
rect 30285 23137 30297 23171
rect 30331 23137 30343 23171
rect 30285 23131 30343 23137
rect 30374 23128 30380 23180
rect 30432 23128 30438 23180
rect 30466 23128 30472 23180
rect 30524 23168 30530 23180
rect 32953 23171 33011 23177
rect 32953 23168 32965 23171
rect 30524 23140 32965 23168
rect 30524 23128 30530 23140
rect 32953 23137 32965 23140
rect 32999 23137 33011 23171
rect 32953 23131 33011 23137
rect 35345 23171 35403 23177
rect 35345 23137 35357 23171
rect 35391 23168 35403 23171
rect 35710 23168 35716 23180
rect 35391 23140 35716 23168
rect 35391 23137 35403 23140
rect 35345 23131 35403 23137
rect 35710 23128 35716 23140
rect 35768 23128 35774 23180
rect 30837 23103 30895 23109
rect 30837 23100 30849 23103
rect 29840 23072 30849 23100
rect 30837 23069 30849 23072
rect 30883 23069 30895 23103
rect 30837 23063 30895 23069
rect 31662 23060 31668 23112
rect 31720 23060 31726 23112
rect 31849 23103 31907 23109
rect 31849 23069 31861 23103
rect 31895 23100 31907 23103
rect 31938 23100 31944 23112
rect 31895 23072 31944 23100
rect 31895 23069 31907 23072
rect 31849 23063 31907 23069
rect 31938 23060 31944 23072
rect 31996 23060 32002 23112
rect 32125 23103 32183 23109
rect 32125 23069 32137 23103
rect 32171 23100 32183 23103
rect 32306 23100 32312 23112
rect 32171 23072 32312 23100
rect 32171 23069 32183 23072
rect 32125 23063 32183 23069
rect 32306 23060 32312 23072
rect 32364 23060 32370 23112
rect 32398 23060 32404 23112
rect 32456 23060 32462 23112
rect 32674 23060 32680 23112
rect 32732 23060 32738 23112
rect 34054 23060 34060 23112
rect 34112 23060 34118 23112
rect 34698 23060 34704 23112
rect 34756 23100 34762 23112
rect 35069 23103 35127 23109
rect 35069 23100 35081 23103
rect 34756 23072 35081 23100
rect 34756 23060 34762 23072
rect 35069 23069 35081 23072
rect 35115 23069 35127 23103
rect 35069 23063 35127 23069
rect 28184 23004 28948 23032
rect 29564 23032 29592 23060
rect 29564 23004 32904 23032
rect 28184 22976 28212 23004
rect 27540 22936 28120 22964
rect 24912 22924 24918 22936
rect 28166 22924 28172 22976
rect 28224 22924 28230 22976
rect 28442 22924 28448 22976
rect 28500 22924 28506 22976
rect 30193 22967 30251 22973
rect 30193 22933 30205 22967
rect 30239 22964 30251 22967
rect 30558 22964 30564 22976
rect 30239 22936 30564 22964
rect 30239 22933 30251 22936
rect 30193 22927 30251 22933
rect 30558 22924 30564 22936
rect 30616 22924 30622 22976
rect 32876 22964 32904 23004
rect 34330 22964 34336 22976
rect 32876 22936 34336 22964
rect 34330 22924 34336 22936
rect 34388 22964 34394 22976
rect 34425 22967 34483 22973
rect 34425 22964 34437 22967
rect 34388 22936 34437 22964
rect 34388 22924 34394 22936
rect 34425 22933 34437 22936
rect 34471 22933 34483 22967
rect 34425 22927 34483 22933
rect 34698 22924 34704 22976
rect 34756 22924 34762 22976
rect 35161 22967 35219 22973
rect 35161 22933 35173 22967
rect 35207 22964 35219 22967
rect 37366 22964 37372 22976
rect 35207 22936 37372 22964
rect 35207 22933 35219 22936
rect 35161 22927 35219 22933
rect 37366 22924 37372 22936
rect 37424 22924 37430 22976
rect 1104 22874 41400 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 41400 22874
rect 1104 22800 41400 22822
rect 9214 22760 9220 22772
rect 8128 22732 9220 22760
rect 8128 22692 8156 22732
rect 9214 22720 9220 22732
rect 9272 22720 9278 22772
rect 11790 22720 11796 22772
rect 11848 22720 11854 22772
rect 11882 22720 11888 22772
rect 11940 22760 11946 22772
rect 12345 22763 12403 22769
rect 11940 22732 12112 22760
rect 11940 22720 11946 22732
rect 7116 22664 8234 22692
rect 11716 22664 12020 22692
rect 7116 22636 7144 22664
rect 5261 22627 5319 22633
rect 5261 22593 5273 22627
rect 5307 22624 5319 22627
rect 5534 22624 5540 22636
rect 5307 22596 5540 22624
rect 5307 22593 5319 22596
rect 5261 22587 5319 22593
rect 5534 22584 5540 22596
rect 5592 22584 5598 22636
rect 7098 22584 7104 22636
rect 7156 22584 7162 22636
rect 10502 22584 10508 22636
rect 10560 22584 10566 22636
rect 11716 22633 11744 22664
rect 11701 22627 11759 22633
rect 10628 22596 11652 22624
rect 4617 22559 4675 22565
rect 4617 22525 4629 22559
rect 4663 22556 4675 22559
rect 4890 22556 4896 22568
rect 4663 22528 4896 22556
rect 4663 22525 4675 22528
rect 4617 22519 4675 22525
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 6546 22516 6552 22568
rect 6604 22556 6610 22568
rect 7469 22559 7527 22565
rect 7469 22556 7481 22559
rect 6604 22528 7481 22556
rect 6604 22516 6610 22528
rect 7469 22525 7481 22528
rect 7515 22525 7527 22559
rect 7469 22519 7527 22525
rect 7745 22559 7803 22565
rect 7745 22525 7757 22559
rect 7791 22556 7803 22559
rect 9122 22556 9128 22568
rect 7791 22528 9128 22556
rect 7791 22525 7803 22528
rect 7745 22519 7803 22525
rect 9122 22516 9128 22528
rect 9180 22516 9186 22568
rect 9217 22559 9275 22565
rect 9217 22525 9229 22559
rect 9263 22556 9275 22559
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 9263 22528 9781 22556
rect 9263 22525 9275 22528
rect 9217 22519 9275 22525
rect 9769 22525 9781 22528
rect 9815 22556 9827 22559
rect 10628 22556 10656 22596
rect 9815 22528 10656 22556
rect 9815 22525 9827 22528
rect 9769 22519 9827 22525
rect 10778 22516 10784 22568
rect 10836 22516 10842 22568
rect 11624 22556 11652 22596
rect 11701 22593 11713 22627
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22593 11943 22627
rect 11885 22587 11943 22593
rect 11900 22556 11928 22587
rect 11624 22528 11928 22556
rect 11992 22556 12020 22664
rect 12084 22633 12112 22732
rect 12345 22729 12357 22763
rect 12391 22760 12403 22763
rect 12434 22760 12440 22772
rect 12391 22732 12440 22760
rect 12391 22729 12403 22732
rect 12345 22723 12403 22729
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 16853 22763 16911 22769
rect 16853 22760 16865 22763
rect 12928 22732 15976 22760
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 12805 22627 12863 22633
rect 12805 22593 12817 22627
rect 12851 22624 12863 22627
rect 12928 22624 12956 22732
rect 12986 22652 12992 22704
rect 13044 22692 13050 22704
rect 13633 22695 13691 22701
rect 13633 22692 13645 22695
rect 13044 22664 13645 22692
rect 13044 22652 13050 22664
rect 13633 22661 13645 22664
rect 13679 22661 13691 22695
rect 13633 22655 13691 22661
rect 13722 22652 13728 22704
rect 13780 22692 13786 22704
rect 14826 22692 14832 22704
rect 13780 22664 14832 22692
rect 13780 22652 13786 22664
rect 14826 22652 14832 22664
rect 14884 22652 14890 22704
rect 15562 22692 15568 22704
rect 15120 22664 15568 22692
rect 12851 22596 12956 22624
rect 12851 22593 12863 22596
rect 12805 22587 12863 22593
rect 12820 22556 12848 22587
rect 13078 22584 13084 22636
rect 13136 22584 13142 22636
rect 13170 22584 13176 22636
rect 13228 22584 13234 22636
rect 13449 22627 13507 22633
rect 13449 22624 13461 22627
rect 13372 22596 13461 22624
rect 11992 22528 12848 22556
rect 13096 22556 13124 22584
rect 13265 22559 13323 22565
rect 13265 22556 13277 22559
rect 13096 22528 13277 22556
rect 5169 22491 5227 22497
rect 5169 22457 5181 22491
rect 5215 22488 5227 22491
rect 5537 22491 5595 22497
rect 5537 22488 5549 22491
rect 5215 22460 5549 22488
rect 5215 22457 5227 22460
rect 5169 22451 5227 22457
rect 5537 22457 5549 22460
rect 5583 22457 5595 22491
rect 5537 22451 5595 22457
rect 5718 22380 5724 22432
rect 5776 22380 5782 22432
rect 10134 22380 10140 22432
rect 10192 22420 10198 22432
rect 10413 22423 10471 22429
rect 10413 22420 10425 22423
rect 10192 22392 10425 22420
rect 10192 22380 10198 22392
rect 10413 22389 10425 22392
rect 10459 22389 10471 22423
rect 11900 22420 11928 22528
rect 13265 22525 13277 22528
rect 13311 22525 13323 22559
rect 13265 22519 13323 22525
rect 12618 22448 12624 22500
rect 12676 22488 12682 22500
rect 13372 22488 13400 22596
rect 13449 22593 13461 22596
rect 13495 22624 13507 22627
rect 13998 22624 14004 22636
rect 13495 22596 14004 22624
rect 13495 22593 13507 22596
rect 13449 22587 13507 22593
rect 13998 22584 14004 22596
rect 14056 22584 14062 22636
rect 14369 22627 14427 22633
rect 14369 22593 14381 22627
rect 14415 22593 14427 22627
rect 14369 22587 14427 22593
rect 14384 22556 14412 22587
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 14918 22584 14924 22636
rect 14976 22624 14982 22636
rect 15120 22633 15148 22664
rect 15562 22652 15568 22664
rect 15620 22652 15626 22704
rect 15948 22692 15976 22732
rect 16592 22732 16865 22760
rect 16592 22704 16620 22732
rect 16853 22729 16865 22732
rect 16899 22760 16911 22763
rect 18322 22760 18328 22772
rect 16899 22732 18328 22760
rect 16899 22729 16911 22732
rect 16853 22723 16911 22729
rect 18322 22720 18328 22732
rect 18380 22720 18386 22772
rect 20901 22763 20959 22769
rect 20901 22760 20913 22763
rect 20088 22732 20913 22760
rect 16390 22692 16396 22704
rect 15948 22664 16396 22692
rect 16390 22652 16396 22664
rect 16448 22652 16454 22704
rect 16574 22652 16580 22704
rect 16632 22652 16638 22704
rect 16669 22695 16727 22701
rect 16669 22661 16681 22695
rect 16715 22692 16727 22695
rect 19334 22692 19340 22704
rect 16715 22664 19340 22692
rect 16715 22661 16727 22664
rect 16669 22655 16727 22661
rect 16868 22636 16896 22664
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 15013 22627 15071 22633
rect 15013 22624 15025 22627
rect 14976 22596 15025 22624
rect 14976 22584 14982 22596
rect 15013 22593 15025 22596
rect 15059 22593 15071 22627
rect 15013 22587 15071 22593
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22624 15531 22627
rect 15654 22624 15660 22636
rect 15519 22596 15660 22624
rect 15519 22593 15531 22596
rect 15473 22587 15531 22593
rect 14660 22556 14688 22584
rect 15028 22556 15056 22587
rect 15654 22584 15660 22596
rect 15712 22584 15718 22636
rect 15749 22627 15807 22633
rect 15749 22593 15761 22627
rect 15795 22624 15807 22627
rect 15795 22596 16804 22624
rect 15795 22593 15807 22596
rect 15749 22587 15807 22593
rect 15565 22559 15623 22565
rect 15565 22556 15577 22559
rect 14384 22528 14964 22556
rect 15028 22528 15577 22556
rect 14936 22488 14964 22528
rect 15565 22525 15577 22528
rect 15611 22525 15623 22559
rect 15565 22519 15623 22525
rect 16574 22488 16580 22500
rect 12676 22460 13400 22488
rect 13464 22460 14596 22488
rect 14936 22460 16580 22488
rect 12676 22448 12682 22460
rect 13464 22420 13492 22460
rect 14568 22432 14596 22460
rect 16574 22448 16580 22460
rect 16632 22448 16638 22500
rect 16776 22488 16804 22596
rect 16850 22584 16856 22636
rect 16908 22584 16914 22636
rect 16942 22584 16948 22636
rect 17000 22584 17006 22636
rect 18138 22584 18144 22636
rect 18196 22584 18202 22636
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22624 18291 22627
rect 18506 22624 18512 22636
rect 18279 22596 18512 22624
rect 18279 22593 18291 22596
rect 18233 22587 18291 22593
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 18598 22584 18604 22636
rect 18656 22624 18662 22636
rect 18693 22627 18751 22633
rect 18693 22624 18705 22627
rect 18656 22596 18705 22624
rect 18656 22584 18662 22596
rect 18693 22593 18705 22596
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 18782 22584 18788 22636
rect 18840 22624 18846 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18840 22596 18889 22624
rect 18840 22584 18846 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 18156 22556 18184 22584
rect 18322 22556 18328 22568
rect 18156 22528 18328 22556
rect 18322 22516 18328 22528
rect 18380 22516 18386 22568
rect 18892 22556 18920 22587
rect 18966 22584 18972 22636
rect 19024 22624 19030 22636
rect 19061 22627 19119 22633
rect 19061 22624 19073 22627
rect 19024 22596 19073 22624
rect 19024 22584 19030 22596
rect 19061 22593 19073 22596
rect 19107 22624 19119 22627
rect 19981 22627 20039 22633
rect 19981 22624 19993 22627
rect 19107 22596 19993 22624
rect 19107 22593 19119 22596
rect 19061 22587 19119 22593
rect 19981 22593 19993 22596
rect 20027 22593 20039 22627
rect 19981 22587 20039 22593
rect 19886 22556 19892 22568
rect 18892 22528 19892 22556
rect 19886 22516 19892 22528
rect 19944 22516 19950 22568
rect 20088 22565 20116 22732
rect 20901 22729 20913 22732
rect 20947 22729 20959 22763
rect 20901 22723 20959 22729
rect 22002 22720 22008 22772
rect 22060 22760 22066 22772
rect 24121 22763 24179 22769
rect 24121 22760 24133 22763
rect 22060 22732 24133 22760
rect 22060 22720 22066 22732
rect 24121 22729 24133 22732
rect 24167 22729 24179 22763
rect 24121 22723 24179 22729
rect 28442 22720 28448 22772
rect 28500 22720 28506 22772
rect 29273 22763 29331 22769
rect 29273 22729 29285 22763
rect 29319 22760 29331 22763
rect 30466 22760 30472 22772
rect 29319 22732 30472 22760
rect 29319 22729 29331 22732
rect 29273 22723 29331 22729
rect 30466 22720 30472 22732
rect 30524 22720 30530 22772
rect 34514 22720 34520 22772
rect 34572 22760 34578 22772
rect 34609 22763 34667 22769
rect 34609 22760 34621 22763
rect 34572 22732 34621 22760
rect 34572 22720 34578 22732
rect 34609 22729 34621 22732
rect 34655 22729 34667 22763
rect 34609 22723 34667 22729
rect 34698 22720 34704 22772
rect 34756 22720 34762 22772
rect 20162 22652 20168 22704
rect 20220 22652 20226 22704
rect 20272 22664 21036 22692
rect 20073 22559 20131 22565
rect 20073 22525 20085 22559
rect 20119 22525 20131 22559
rect 20180 22556 20208 22652
rect 20272 22633 20300 22664
rect 20250 22627 20308 22633
rect 20250 22593 20262 22627
rect 20296 22593 20308 22627
rect 20250 22587 20308 22593
rect 20346 22584 20352 22636
rect 20404 22624 20410 22636
rect 20533 22627 20591 22633
rect 20533 22624 20545 22627
rect 20404 22596 20545 22624
rect 20404 22584 20410 22596
rect 20533 22593 20545 22596
rect 20579 22593 20591 22627
rect 20533 22587 20591 22593
rect 20714 22584 20720 22636
rect 20772 22584 20778 22636
rect 21008 22624 21036 22664
rect 21818 22652 21824 22704
rect 21876 22652 21882 22704
rect 23658 22652 23664 22704
rect 23716 22652 23722 22704
rect 24026 22652 24032 22704
rect 24084 22652 24090 22704
rect 28460 22692 28488 22720
rect 28460 22664 29868 22692
rect 22278 22624 22284 22636
rect 21008 22596 22284 22624
rect 22278 22584 22284 22596
rect 22336 22624 22342 22636
rect 23845 22627 23903 22633
rect 23845 22624 23857 22627
rect 22336 22596 23857 22624
rect 22336 22584 22342 22596
rect 23845 22593 23857 22596
rect 23891 22593 23903 22627
rect 24044 22624 24072 22652
rect 24302 22624 24308 22636
rect 24044 22596 24308 22624
rect 23845 22587 23903 22593
rect 24302 22584 24308 22596
rect 24360 22584 24366 22636
rect 24486 22584 24492 22636
rect 24544 22584 24550 22636
rect 26602 22584 26608 22636
rect 26660 22584 26666 22636
rect 28994 22584 29000 22636
rect 29052 22624 29058 22636
rect 29457 22627 29515 22633
rect 29457 22624 29469 22627
rect 29052 22596 29469 22624
rect 29052 22584 29058 22596
rect 29457 22593 29469 22596
rect 29503 22593 29515 22627
rect 29457 22587 29515 22593
rect 29549 22627 29607 22633
rect 29549 22593 29561 22627
rect 29595 22593 29607 22627
rect 29549 22587 29607 22593
rect 24029 22559 24087 22565
rect 24029 22556 24041 22559
rect 20180 22528 24041 22556
rect 20073 22519 20131 22525
rect 24029 22525 24041 22528
rect 24075 22525 24087 22559
rect 24029 22519 24087 22525
rect 24581 22559 24639 22565
rect 24581 22525 24593 22559
rect 24627 22556 24639 22559
rect 26620 22556 26648 22584
rect 24627 22528 26648 22556
rect 24627 22525 24639 22528
rect 24581 22519 24639 22525
rect 20088 22488 20116 22519
rect 29178 22516 29184 22568
rect 29236 22556 29242 22568
rect 29564 22556 29592 22587
rect 29730 22584 29736 22636
rect 29788 22584 29794 22636
rect 29840 22633 29868 22664
rect 30374 22652 30380 22704
rect 30432 22692 30438 22704
rect 31110 22692 31116 22704
rect 30432 22664 31116 22692
rect 30432 22652 30438 22664
rect 31110 22652 31116 22664
rect 31168 22652 31174 22704
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22593 29883 22627
rect 29825 22587 29883 22593
rect 29914 22584 29920 22636
rect 29972 22584 29978 22636
rect 34716 22624 34744 22720
rect 36998 22652 37004 22704
rect 37056 22692 37062 22704
rect 37056 22664 38042 22692
rect 37056 22652 37062 22664
rect 34793 22627 34851 22633
rect 34793 22624 34805 22627
rect 34716 22596 34805 22624
rect 34793 22593 34805 22596
rect 34839 22593 34851 22627
rect 34793 22587 34851 22593
rect 29932 22556 29960 22584
rect 29236 22528 29960 22556
rect 37277 22559 37335 22565
rect 29236 22516 29242 22528
rect 37277 22525 37289 22559
rect 37323 22525 37335 22559
rect 37277 22519 37335 22525
rect 22094 22488 22100 22500
rect 16776 22460 20116 22488
rect 20456 22460 22100 22488
rect 11900 22392 13492 22420
rect 10413 22383 10471 22389
rect 14274 22380 14280 22432
rect 14332 22420 14338 22432
rect 14461 22423 14519 22429
rect 14461 22420 14473 22423
rect 14332 22392 14473 22420
rect 14332 22380 14338 22392
rect 14461 22389 14473 22392
rect 14507 22389 14519 22423
rect 14461 22383 14519 22389
rect 14550 22380 14556 22432
rect 14608 22380 14614 22432
rect 15102 22380 15108 22432
rect 15160 22380 15166 22432
rect 15286 22380 15292 22432
rect 15344 22380 15350 22432
rect 15470 22380 15476 22432
rect 15528 22380 15534 22432
rect 15930 22380 15936 22432
rect 15988 22380 15994 22432
rect 16666 22380 16672 22432
rect 16724 22380 16730 22432
rect 18230 22380 18236 22432
rect 18288 22380 18294 22432
rect 18598 22380 18604 22432
rect 18656 22380 18662 22432
rect 19426 22380 19432 22432
rect 19484 22420 19490 22432
rect 19981 22423 20039 22429
rect 19981 22420 19993 22423
rect 19484 22392 19993 22420
rect 19484 22380 19490 22392
rect 19981 22389 19993 22392
rect 20027 22389 20039 22423
rect 19981 22383 20039 22389
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 20456 22429 20484 22460
rect 22094 22448 22100 22460
rect 22152 22448 22158 22500
rect 23290 22448 23296 22500
rect 23348 22488 23354 22500
rect 23348 22460 29592 22488
rect 23348 22448 23354 22460
rect 29564 22432 29592 22460
rect 32306 22448 32312 22500
rect 32364 22488 32370 22500
rect 35802 22488 35808 22500
rect 32364 22460 35808 22488
rect 32364 22448 32370 22460
rect 35802 22448 35808 22460
rect 35860 22448 35866 22500
rect 20441 22423 20499 22429
rect 20441 22420 20453 22423
rect 20128 22392 20453 22420
rect 20128 22380 20134 22392
rect 20441 22389 20453 22392
rect 20487 22389 20499 22423
rect 20441 22383 20499 22389
rect 24026 22380 24032 22432
rect 24084 22420 24090 22432
rect 24578 22420 24584 22432
rect 24084 22392 24584 22420
rect 24084 22380 24090 22392
rect 24578 22380 24584 22392
rect 24636 22380 24642 22432
rect 29546 22380 29552 22432
rect 29604 22380 29610 22432
rect 37292 22420 37320 22519
rect 37550 22516 37556 22568
rect 37608 22516 37614 22568
rect 39298 22516 39304 22568
rect 39356 22516 39362 22568
rect 38286 22420 38292 22432
rect 37292 22392 38292 22420
rect 38286 22380 38292 22392
rect 38344 22380 38350 22432
rect 1104 22330 41400 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 41400 22330
rect 1104 22256 41400 22278
rect 1854 22176 1860 22228
rect 1912 22216 1918 22228
rect 2501 22219 2559 22225
rect 2501 22216 2513 22219
rect 1912 22188 2513 22216
rect 1912 22176 1918 22188
rect 2501 22185 2513 22188
rect 2547 22185 2559 22219
rect 2501 22179 2559 22185
rect 5534 22176 5540 22228
rect 5592 22176 5598 22228
rect 7374 22176 7380 22228
rect 7432 22216 7438 22228
rect 12986 22216 12992 22228
rect 7432 22188 12992 22216
rect 7432 22176 7438 22188
rect 12986 22176 12992 22188
rect 13044 22176 13050 22228
rect 13446 22216 13452 22228
rect 13096 22188 13452 22216
rect 10962 22148 10968 22160
rect 9968 22120 10968 22148
rect 3789 22083 3847 22089
rect 3789 22080 3801 22083
rect 2240 22052 3801 22080
rect 2240 22024 2268 22052
rect 3789 22049 3801 22052
rect 3835 22080 3847 22083
rect 4062 22080 4068 22092
rect 3835 22052 4068 22080
rect 3835 22049 3847 22052
rect 3789 22043 3847 22049
rect 4062 22040 4068 22052
rect 4120 22080 4126 22092
rect 5350 22080 5356 22092
rect 4120 22052 5356 22080
rect 4120 22040 4126 22052
rect 5350 22040 5356 22052
rect 5408 22040 5414 22092
rect 8110 22040 8116 22092
rect 8168 22080 8174 22092
rect 8168 22052 8524 22080
rect 8168 22040 8174 22052
rect 2222 21972 2228 22024
rect 2280 21972 2286 22024
rect 2317 22015 2375 22021
rect 2317 21981 2329 22015
rect 2363 22012 2375 22015
rect 7837 22015 7895 22021
rect 2363 21984 2774 22012
rect 2363 21981 2375 21984
rect 2317 21975 2375 21981
rect 2746 21876 2774 21984
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 8021 22015 8079 22021
rect 8021 21981 8033 22015
rect 8067 22012 8079 22015
rect 8496 22012 8524 22052
rect 8570 22040 8576 22092
rect 8628 22040 8634 22092
rect 9766 22012 9772 22024
rect 8067 21984 8432 22012
rect 8496 21984 9772 22012
rect 8067 21981 8079 21984
rect 8021 21975 8079 21981
rect 4065 21947 4123 21953
rect 4065 21913 4077 21947
rect 4111 21944 4123 21947
rect 4111 21916 4476 21944
rect 4111 21913 4123 21916
rect 4065 21907 4123 21913
rect 4448 21888 4476 21916
rect 4522 21904 4528 21956
rect 4580 21904 4586 21956
rect 7852 21944 7880 21975
rect 8202 21944 8208 21956
rect 7852 21916 8208 21944
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 8404 21953 8432 21984
rect 9766 21972 9772 21984
rect 9824 22012 9830 22024
rect 9861 22015 9919 22021
rect 9861 22012 9873 22015
rect 9824 21984 9873 22012
rect 9824 21972 9830 21984
rect 9861 21981 9873 21984
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 8389 21947 8447 21953
rect 8389 21913 8401 21947
rect 8435 21944 8447 21947
rect 9968 21944 9996 22120
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 11885 22083 11943 22089
rect 11885 22080 11897 22083
rect 10060 22052 11897 22080
rect 10060 22021 10088 22052
rect 11885 22049 11897 22052
rect 11931 22049 11943 22083
rect 12618 22080 12624 22092
rect 11885 22043 11943 22049
rect 12176 22052 12624 22080
rect 10045 22015 10103 22021
rect 10045 21981 10057 22015
rect 10091 21981 10103 22015
rect 10045 21975 10103 21981
rect 10134 21972 10140 22024
rect 10192 21972 10198 22024
rect 10226 21972 10232 22024
rect 10284 21972 10290 22024
rect 10594 21972 10600 22024
rect 10652 21972 10658 22024
rect 11514 21972 11520 22024
rect 11572 22012 11578 22024
rect 12176 22021 12204 22052
rect 12618 22040 12624 22052
rect 12676 22040 12682 22092
rect 13096 22080 13124 22188
rect 13446 22176 13452 22188
rect 13504 22176 13510 22228
rect 13998 22176 14004 22228
rect 14056 22176 14062 22228
rect 15749 22219 15807 22225
rect 15749 22185 15761 22219
rect 15795 22216 15807 22219
rect 15838 22216 15844 22228
rect 15795 22188 15844 22216
rect 15795 22185 15807 22188
rect 15749 22179 15807 22185
rect 15838 22176 15844 22188
rect 15896 22176 15902 22228
rect 17497 22219 17555 22225
rect 17497 22185 17509 22219
rect 17543 22216 17555 22219
rect 18138 22216 18144 22228
rect 17543 22188 18144 22216
rect 17543 22185 17555 22188
rect 17497 22179 17555 22185
rect 18138 22176 18144 22188
rect 18196 22176 18202 22228
rect 18601 22219 18659 22225
rect 18601 22185 18613 22219
rect 18647 22216 18659 22219
rect 20070 22216 20076 22228
rect 18647 22188 20076 22216
rect 18647 22185 18659 22188
rect 18601 22179 18659 22185
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 20622 22176 20628 22228
rect 20680 22216 20686 22228
rect 21450 22216 21456 22228
rect 20680 22188 21456 22216
rect 20680 22176 20686 22188
rect 21450 22176 21456 22188
rect 21508 22176 21514 22228
rect 23106 22176 23112 22228
rect 23164 22176 23170 22228
rect 23661 22219 23719 22225
rect 23661 22185 23673 22219
rect 23707 22216 23719 22219
rect 25222 22216 25228 22228
rect 23707 22188 25228 22216
rect 23707 22185 23719 22188
rect 23661 22179 23719 22185
rect 25222 22176 25228 22188
rect 25280 22176 25286 22228
rect 25866 22176 25872 22228
rect 25924 22176 25930 22228
rect 26142 22176 26148 22228
rect 26200 22216 26206 22228
rect 28994 22216 29000 22228
rect 26200 22188 29000 22216
rect 26200 22176 26206 22188
rect 28994 22176 29000 22188
rect 29052 22176 29058 22228
rect 37550 22176 37556 22228
rect 37608 22216 37614 22228
rect 37921 22219 37979 22225
rect 37921 22216 37933 22219
rect 37608 22188 37933 22216
rect 37608 22176 37614 22188
rect 37921 22185 37933 22188
rect 37967 22185 37979 22219
rect 37921 22179 37979 22185
rect 13354 22108 13360 22160
rect 13412 22148 13418 22160
rect 13633 22151 13691 22157
rect 13633 22148 13645 22151
rect 13412 22120 13645 22148
rect 13412 22108 13418 22120
rect 13633 22117 13645 22120
rect 13679 22117 13691 22151
rect 14016 22148 14044 22176
rect 16022 22148 16028 22160
rect 14016 22120 16028 22148
rect 13633 22111 13691 22117
rect 16022 22108 16028 22120
rect 16080 22148 16086 22160
rect 17773 22151 17831 22157
rect 16080 22120 17540 22148
rect 16080 22108 16086 22120
rect 12728 22052 13124 22080
rect 11701 22015 11759 22021
rect 11701 22012 11713 22015
rect 11572 21984 11713 22012
rect 11572 21972 11578 21984
rect 11701 21981 11713 21984
rect 11747 22012 11759 22015
rect 11977 22015 12035 22021
rect 11977 22012 11989 22015
rect 11747 21984 11989 22012
rect 11747 21981 11759 21984
rect 11701 21975 11759 21981
rect 11977 21981 11989 21984
rect 12023 21981 12035 22015
rect 11977 21975 12035 21981
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 8435 21916 9996 21944
rect 10249 21944 10277 21972
rect 10870 21944 10876 21956
rect 10249 21916 10876 21944
rect 8435 21913 8447 21916
rect 8389 21907 8447 21913
rect 10870 21904 10876 21916
rect 10928 21904 10934 21956
rect 11333 21947 11391 21953
rect 11333 21944 11345 21947
rect 11164 21916 11345 21944
rect 2958 21876 2964 21888
rect 2746 21848 2964 21876
rect 2958 21836 2964 21848
rect 3016 21836 3022 21888
rect 4430 21836 4436 21888
rect 4488 21836 4494 21888
rect 5534 21836 5540 21888
rect 5592 21876 5598 21888
rect 5810 21876 5816 21888
rect 5592 21848 5816 21876
rect 5592 21836 5598 21848
rect 5810 21836 5816 21848
rect 5868 21836 5874 21888
rect 7926 21836 7932 21888
rect 7984 21836 7990 21888
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 10413 21879 10471 21885
rect 10413 21876 10425 21879
rect 9180 21848 10425 21876
rect 9180 21836 9186 21848
rect 10413 21845 10425 21848
rect 10459 21845 10471 21879
rect 10413 21839 10471 21845
rect 10502 21836 10508 21888
rect 10560 21876 10566 21888
rect 11164 21876 11192 21916
rect 11333 21913 11345 21916
rect 11379 21913 11391 21947
rect 11333 21907 11391 21913
rect 11609 21947 11667 21953
rect 11609 21913 11621 21947
rect 11655 21944 11667 21947
rect 12176 21944 12204 21975
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 12728 22021 12756 22052
rect 14458 22040 14464 22092
rect 14516 22040 14522 22092
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 21981 12771 22015
rect 12713 21975 12771 21981
rect 12989 22015 13047 22021
rect 12989 21981 13001 22015
rect 13035 21981 13047 22015
rect 12989 21975 13047 21981
rect 11655 21916 12204 21944
rect 11655 21913 11667 21916
rect 11609 21907 11667 21913
rect 10560 21848 11192 21876
rect 10560 21836 10566 21848
rect 11238 21836 11244 21888
rect 11296 21836 11302 21888
rect 11348 21876 11376 21907
rect 12342 21904 12348 21956
rect 12400 21944 12406 21956
rect 12400 21916 12848 21944
rect 12400 21904 12406 21916
rect 12820 21888 12848 21916
rect 11422 21876 11428 21888
rect 11348 21848 11428 21876
rect 11422 21836 11428 21848
rect 11480 21836 11486 21888
rect 11514 21836 11520 21888
rect 11572 21836 11578 21888
rect 12066 21836 12072 21888
rect 12124 21836 12130 21888
rect 12621 21879 12679 21885
rect 12621 21845 12633 21879
rect 12667 21876 12679 21879
rect 12710 21876 12716 21888
rect 12667 21848 12716 21876
rect 12667 21845 12679 21848
rect 12621 21839 12679 21845
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 12802 21836 12808 21888
rect 12860 21836 12866 21888
rect 13004 21876 13032 21975
rect 13170 21972 13176 22024
rect 13228 21972 13234 22024
rect 13262 21972 13268 22024
rect 13320 22012 13326 22024
rect 13633 22015 13691 22021
rect 13633 22012 13645 22015
rect 13320 21984 13645 22012
rect 13320 21972 13326 21984
rect 13633 21981 13645 21984
rect 13679 22012 13691 22015
rect 13814 22012 13820 22024
rect 13679 21984 13820 22012
rect 13679 21981 13691 21984
rect 13633 21975 13691 21981
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 14369 22015 14427 22021
rect 14369 22012 14381 22015
rect 14292 21984 14381 22012
rect 13188 21944 13216 21972
rect 14292 21956 14320 21984
rect 14369 21981 14381 21984
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 14550 21972 14556 22024
rect 14608 22012 14614 22024
rect 17405 22015 17463 22021
rect 14608 21984 15608 22012
rect 14608 21972 14614 21984
rect 13446 21944 13452 21956
rect 13188 21916 13452 21944
rect 13446 21904 13452 21916
rect 13504 21904 13510 21956
rect 14274 21904 14280 21956
rect 14332 21944 14338 21956
rect 15580 21953 15608 21984
rect 17405 21981 17417 22015
rect 17451 21981 17463 22015
rect 17512 22012 17540 22120
rect 17773 22117 17785 22151
rect 17819 22148 17831 22151
rect 17819 22120 18736 22148
rect 17819 22117 17831 22120
rect 17773 22111 17831 22117
rect 17972 22052 18460 22080
rect 17681 22015 17739 22021
rect 17681 22012 17693 22015
rect 17512 21984 17693 22012
rect 17405 21975 17463 21981
rect 17681 21981 17693 21984
rect 17727 21981 17739 22015
rect 17681 21975 17739 21981
rect 15381 21947 15439 21953
rect 15381 21944 15393 21947
rect 14332 21916 15393 21944
rect 14332 21904 14338 21916
rect 15381 21913 15393 21916
rect 15427 21913 15439 21947
rect 15381 21907 15439 21913
rect 15565 21947 15623 21953
rect 15565 21913 15577 21947
rect 15611 21944 15623 21947
rect 15654 21944 15660 21956
rect 15611 21916 15660 21944
rect 15611 21913 15623 21916
rect 15565 21907 15623 21913
rect 15654 21904 15660 21916
rect 15712 21904 15718 21956
rect 17218 21904 17224 21956
rect 17276 21904 17282 21956
rect 17420 21944 17448 21975
rect 17770 21972 17776 22024
rect 17828 22012 17834 22024
rect 17972 22021 18000 22052
rect 17957 22015 18015 22021
rect 17957 22012 17969 22015
rect 17828 21984 17969 22012
rect 17828 21972 17834 21984
rect 17957 21981 17969 21984
rect 18003 21981 18015 22015
rect 18322 22012 18328 22024
rect 17957 21975 18015 21981
rect 18064 21984 18328 22012
rect 18064 21944 18092 21984
rect 18322 21972 18328 21984
rect 18380 21972 18386 22024
rect 17420 21916 18092 21944
rect 18141 21947 18199 21953
rect 18141 21913 18153 21947
rect 18187 21913 18199 21947
rect 18141 21907 18199 21913
rect 15286 21876 15292 21888
rect 13004 21848 15292 21876
rect 15286 21836 15292 21848
rect 15344 21836 15350 21888
rect 17236 21876 17264 21904
rect 17770 21876 17776 21888
rect 17236 21848 17776 21876
rect 17770 21836 17776 21848
rect 17828 21876 17834 21888
rect 18156 21876 18184 21907
rect 17828 21848 18184 21876
rect 18432 21876 18460 22052
rect 18506 22040 18512 22092
rect 18564 22040 18570 22092
rect 18708 22080 18736 22120
rect 18782 22108 18788 22160
rect 18840 22108 18846 22160
rect 20165 22151 20223 22157
rect 18984 22120 19656 22148
rect 18984 22080 19012 22120
rect 18708 22052 19012 22080
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 21981 18659 22015
rect 18601 21975 18659 21981
rect 18877 22015 18935 22021
rect 18877 21981 18889 22015
rect 18923 22012 18935 22015
rect 18984 22012 19012 22052
rect 19168 22052 19472 22080
rect 18923 21984 19012 22012
rect 18923 21981 18935 21984
rect 18877 21975 18935 21981
rect 18616 21944 18644 21975
rect 19058 21972 19064 22024
rect 19116 21972 19122 22024
rect 18969 21947 19027 21953
rect 18969 21944 18981 21947
rect 18616 21916 18981 21944
rect 18969 21913 18981 21916
rect 19015 21913 19027 21947
rect 18969 21907 19027 21913
rect 19168 21876 19196 22052
rect 19242 21972 19248 22024
rect 19300 21972 19306 22024
rect 19334 21972 19340 22024
rect 19392 21972 19398 22024
rect 19444 22021 19472 22052
rect 19518 22040 19524 22092
rect 19576 22080 19582 22092
rect 19628 22080 19656 22120
rect 20165 22117 20177 22151
rect 20211 22148 20223 22151
rect 20714 22148 20720 22160
rect 20211 22120 20720 22148
rect 20211 22117 20223 22120
rect 20165 22111 20223 22117
rect 20714 22108 20720 22120
rect 20772 22108 20778 22160
rect 21082 22108 21088 22160
rect 21140 22108 21146 22160
rect 22278 22108 22284 22160
rect 22336 22148 22342 22160
rect 22557 22151 22615 22157
rect 22557 22148 22569 22151
rect 22336 22120 22569 22148
rect 22336 22108 22342 22120
rect 22557 22117 22569 22120
rect 22603 22117 22615 22151
rect 24946 22148 24952 22160
rect 22557 22111 22615 22117
rect 23216 22120 24952 22148
rect 21910 22080 21916 22092
rect 19576 22052 19656 22080
rect 19720 22052 20484 22080
rect 19576 22040 19582 22052
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19610 21972 19616 22024
rect 19668 22012 19674 22024
rect 19720 22012 19748 22052
rect 19668 21984 19748 22012
rect 19668 21972 19674 21984
rect 20070 21972 20076 22024
rect 20128 22012 20134 22024
rect 20456 22021 20484 22052
rect 20732 22052 21916 22080
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 20128 21984 20361 22012
rect 20128 21972 20134 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 20441 22015 20499 22021
rect 20441 21981 20453 22015
rect 20487 21981 20499 22015
rect 20441 21975 20499 21981
rect 20622 21972 20628 22024
rect 20680 21972 20686 22024
rect 20732 22021 20760 22052
rect 21910 22040 21916 22052
rect 21968 22040 21974 22092
rect 22925 22083 22983 22089
rect 22925 22080 22937 22083
rect 22674 22052 22937 22080
rect 20717 22015 20775 22021
rect 20717 21981 20729 22015
rect 20763 21981 20775 22015
rect 20717 21975 20775 21981
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 21981 20867 22015
rect 20809 21975 20867 21981
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 22674 22012 22702 22052
rect 22925 22049 22937 22052
rect 22971 22080 22983 22083
rect 23216 22080 23244 22120
rect 24946 22108 24952 22120
rect 25004 22108 25010 22160
rect 23382 22080 23388 22092
rect 22971 22052 23244 22080
rect 23308 22052 23388 22080
rect 22971 22049 22983 22052
rect 22925 22043 22983 22049
rect 20993 21975 21051 21981
rect 21284 21984 22702 22012
rect 19352 21944 19380 21972
rect 20162 21944 20168 21956
rect 19352 21916 20168 21944
rect 20162 21904 20168 21916
rect 20220 21904 20226 21956
rect 18432 21848 19196 21876
rect 17828 21836 17834 21848
rect 19334 21836 19340 21888
rect 19392 21836 19398 21888
rect 19886 21836 19892 21888
rect 19944 21876 19950 21888
rect 20824 21876 20852 21975
rect 21008 21944 21036 21975
rect 21284 21944 21312 21984
rect 22738 21972 22744 22024
rect 22796 21972 22802 22024
rect 23014 21972 23020 22024
rect 23072 21972 23078 22024
rect 23308 22021 23336 22052
rect 23382 22040 23388 22052
rect 23440 22040 23446 22092
rect 23477 22083 23535 22089
rect 23477 22049 23489 22083
rect 23523 22080 23535 22083
rect 23750 22080 23756 22092
rect 23523 22052 23756 22080
rect 23523 22049 23535 22052
rect 23477 22043 23535 22049
rect 23750 22040 23756 22052
rect 23808 22040 23814 22092
rect 24118 22040 24124 22092
rect 24176 22040 24182 22092
rect 24394 22080 24400 22092
rect 24228 22052 24400 22080
rect 24228 22024 24256 22052
rect 24394 22040 24400 22052
rect 24452 22080 24458 22092
rect 24765 22083 24823 22089
rect 24765 22080 24777 22083
rect 24452 22052 24777 22080
rect 24452 22040 24458 22052
rect 24765 22049 24777 22052
rect 24811 22049 24823 22083
rect 24765 22043 24823 22049
rect 24854 22040 24860 22092
rect 24912 22040 24918 22092
rect 25884 22080 25912 22176
rect 28902 22148 28908 22160
rect 28736 22120 28908 22148
rect 28736 22089 28764 22120
rect 28902 22108 28908 22120
rect 28960 22108 28966 22160
rect 29546 22108 29552 22160
rect 29604 22148 29610 22160
rect 37734 22148 37740 22160
rect 29604 22120 37740 22148
rect 29604 22108 29610 22120
rect 37734 22108 37740 22120
rect 37792 22108 37798 22160
rect 25148 22052 25912 22080
rect 28721 22083 28779 22089
rect 23293 22015 23351 22021
rect 23293 21981 23305 22015
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 22012 23627 22015
rect 23658 22012 23664 22024
rect 23615 21984 23664 22012
rect 23615 21981 23627 21984
rect 23569 21975 23627 21981
rect 23658 21972 23664 21984
rect 23716 21972 23722 22024
rect 23842 21972 23848 22024
rect 23900 21972 23906 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 21008 21916 21312 21944
rect 21358 21904 21364 21956
rect 21416 21904 21422 21956
rect 22094 21904 22100 21956
rect 22152 21944 22158 21956
rect 24044 21944 24072 21975
rect 24210 21972 24216 22024
rect 24268 21972 24274 22024
rect 24302 21972 24308 22024
rect 24360 22012 24366 22024
rect 25148 22021 25176 22052
rect 28721 22049 28733 22083
rect 28767 22049 28779 22083
rect 28721 22043 28779 22049
rect 24673 22015 24731 22021
rect 24673 22012 24685 22015
rect 24360 21984 24685 22012
rect 24360 21972 24366 21984
rect 24673 21981 24685 21984
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 25133 22015 25191 22021
rect 25133 21981 25145 22015
rect 25179 21981 25191 22015
rect 28445 22015 28503 22021
rect 25133 21975 25191 21981
rect 25608 21984 27752 22012
rect 25148 21944 25176 21975
rect 22152 21916 24072 21944
rect 24136 21916 25176 21944
rect 22152 21904 22158 21916
rect 24136 21876 24164 21916
rect 25608 21888 25636 21984
rect 27522 21904 27528 21956
rect 27580 21904 27586 21956
rect 19944 21848 24164 21876
rect 19944 21836 19950 21848
rect 24394 21836 24400 21888
rect 24452 21836 24458 21888
rect 25590 21836 25596 21888
rect 25648 21836 25654 21888
rect 26326 21836 26332 21888
rect 26384 21876 26390 21888
rect 27430 21876 27436 21888
rect 26384 21848 27436 21876
rect 26384 21836 26390 21848
rect 27430 21836 27436 21848
rect 27488 21876 27494 21888
rect 27617 21879 27675 21885
rect 27617 21876 27629 21879
rect 27488 21848 27629 21876
rect 27488 21836 27494 21848
rect 27617 21845 27629 21848
rect 27663 21845 27675 21879
rect 27724 21876 27752 21984
rect 28445 21981 28457 22015
rect 28491 22012 28503 22015
rect 28626 22012 28632 22024
rect 28491 21984 28632 22012
rect 28491 21981 28503 21984
rect 28445 21975 28503 21981
rect 28626 21972 28632 21984
rect 28684 21972 28690 22024
rect 29564 22021 29592 22108
rect 35434 22040 35440 22092
rect 35492 22080 35498 22092
rect 35621 22083 35679 22089
rect 35621 22080 35633 22083
rect 35492 22052 35633 22080
rect 35492 22040 35498 22052
rect 35621 22049 35633 22052
rect 35667 22049 35679 22083
rect 35621 22043 35679 22049
rect 36081 22083 36139 22089
rect 36081 22049 36093 22083
rect 36127 22080 36139 22083
rect 36127 22052 36860 22080
rect 36127 22049 36139 22052
rect 36081 22043 36139 22049
rect 29549 22015 29607 22021
rect 29549 21981 29561 22015
rect 29595 21981 29607 22015
rect 29549 21975 29607 21981
rect 35342 21972 35348 22024
rect 35400 22012 35406 22024
rect 35713 22015 35771 22021
rect 35713 22012 35725 22015
rect 35400 21984 35725 22012
rect 35400 21972 35406 21984
rect 35713 21981 35725 21984
rect 35759 22012 35771 22015
rect 36630 22012 36636 22024
rect 35759 21984 36636 22012
rect 35759 21981 35771 21984
rect 35713 21975 35771 21981
rect 36630 21972 36636 21984
rect 36688 21972 36694 22024
rect 30006 21904 30012 21956
rect 30064 21944 30070 21956
rect 30285 21947 30343 21953
rect 30285 21944 30297 21947
rect 30064 21916 30297 21944
rect 30064 21904 30070 21916
rect 30285 21913 30297 21916
rect 30331 21913 30343 21947
rect 30285 21907 30343 21913
rect 36832 21888 36860 22052
rect 37642 22040 37648 22092
rect 37700 22040 37706 22092
rect 39298 22080 39304 22092
rect 37752 22052 39304 22080
rect 37550 21972 37556 22024
rect 37608 22012 37614 22024
rect 37752 22012 37780 22052
rect 39298 22040 39304 22052
rect 39356 22040 39362 22092
rect 37608 21984 37780 22012
rect 38105 22015 38163 22021
rect 37608 21972 37614 21984
rect 38105 21981 38117 22015
rect 38151 21981 38163 22015
rect 38105 21975 38163 21981
rect 38120 21944 38148 21975
rect 37108 21916 38148 21944
rect 28077 21879 28135 21885
rect 28077 21876 28089 21879
rect 27724 21848 28089 21876
rect 27617 21839 27675 21845
rect 28077 21845 28089 21848
rect 28123 21845 28135 21879
rect 28077 21839 28135 21845
rect 28258 21836 28264 21888
rect 28316 21876 28322 21888
rect 28537 21879 28595 21885
rect 28537 21876 28549 21879
rect 28316 21848 28549 21876
rect 28316 21836 28322 21848
rect 28537 21845 28549 21848
rect 28583 21845 28595 21879
rect 28537 21839 28595 21845
rect 36814 21836 36820 21888
rect 36872 21836 36878 21888
rect 37108 21885 37136 21916
rect 37093 21879 37151 21885
rect 37093 21845 37105 21879
rect 37139 21845 37151 21879
rect 37093 21839 37151 21845
rect 37458 21836 37464 21888
rect 37516 21836 37522 21888
rect 1104 21786 41400 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 41400 21786
rect 1104 21712 41400 21734
rect 6564 21644 7972 21672
rect 6564 21616 6592 21644
rect 5350 21564 5356 21616
rect 5408 21604 5414 21616
rect 6546 21604 6552 21616
rect 5408 21576 6552 21604
rect 5408 21564 5414 21576
rect 4062 21496 4068 21548
rect 4120 21536 4126 21548
rect 4522 21536 4528 21548
rect 4120 21508 4528 21536
rect 4120 21496 4126 21508
rect 4522 21496 4528 21508
rect 4580 21496 4586 21548
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21536 4675 21539
rect 4798 21536 4804 21548
rect 4663 21508 4804 21536
rect 4663 21505 4675 21508
rect 4617 21499 4675 21505
rect 4798 21496 4804 21508
rect 4856 21536 4862 21548
rect 5166 21536 5172 21548
rect 4856 21508 5172 21536
rect 4856 21496 4862 21508
rect 5166 21496 5172 21508
rect 5224 21496 5230 21548
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21505 5687 21539
rect 5629 21499 5687 21505
rect 1394 21428 1400 21480
rect 1452 21468 1458 21480
rect 2222 21468 2228 21480
rect 1452 21440 2228 21468
rect 1452 21428 1458 21440
rect 2222 21428 2228 21440
rect 2280 21468 2286 21480
rect 2685 21471 2743 21477
rect 2685 21468 2697 21471
rect 2280 21440 2697 21468
rect 2280 21428 2286 21440
rect 2685 21437 2697 21440
rect 2731 21437 2743 21471
rect 2685 21431 2743 21437
rect 2958 21428 2964 21480
rect 3016 21468 3022 21480
rect 4433 21471 4491 21477
rect 3016 21440 4384 21468
rect 3016 21428 3022 21440
rect 4356 21400 4384 21440
rect 4433 21437 4445 21471
rect 4479 21468 4491 21471
rect 4890 21468 4896 21480
rect 4479 21440 4896 21468
rect 4479 21437 4491 21440
rect 4433 21431 4491 21437
rect 4890 21428 4896 21440
rect 4948 21468 4954 21480
rect 5644 21468 5672 21499
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 6380 21545 6408 21576
rect 6546 21564 6552 21576
rect 6604 21564 6610 21616
rect 7098 21564 7104 21616
rect 7156 21564 7162 21616
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 7944 21536 7972 21644
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 10229 21675 10287 21681
rect 9824 21644 10088 21672
rect 9824 21632 9830 21644
rect 9214 21564 9220 21616
rect 9272 21564 9278 21616
rect 7944 21508 8248 21536
rect 6365 21499 6423 21505
rect 4948 21440 5672 21468
rect 4948 21428 4954 21440
rect 6638 21428 6644 21480
rect 6696 21428 6702 21480
rect 7006 21428 7012 21480
rect 7064 21468 7070 21480
rect 8110 21468 8116 21480
rect 7064 21440 8116 21468
rect 7064 21428 7070 21440
rect 8110 21428 8116 21440
rect 8168 21428 8174 21480
rect 8220 21468 8248 21508
rect 8386 21496 8392 21548
rect 8444 21496 8450 21548
rect 10060 21536 10088 21644
rect 10229 21641 10241 21675
rect 10275 21672 10287 21675
rect 10594 21672 10600 21684
rect 10275 21644 10600 21672
rect 10275 21641 10287 21644
rect 10229 21635 10287 21641
rect 10594 21632 10600 21644
rect 10652 21672 10658 21684
rect 10652 21644 10824 21672
rect 10652 21632 10658 21644
rect 10594 21536 10600 21548
rect 10060 21508 10600 21536
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 10686 21496 10692 21548
rect 10744 21496 10750 21548
rect 8481 21471 8539 21477
rect 8481 21468 8493 21471
rect 8220 21440 8493 21468
rect 8481 21437 8493 21440
rect 8527 21437 8539 21471
rect 8481 21431 8539 21437
rect 8757 21471 8815 21477
rect 8757 21437 8769 21471
rect 8803 21468 8815 21471
rect 10796 21468 10824 21644
rect 11238 21632 11244 21684
rect 11296 21632 11302 21684
rect 14734 21672 14740 21684
rect 12406 21644 14740 21672
rect 10965 21607 11023 21613
rect 10965 21573 10977 21607
rect 11011 21604 11023 21607
rect 11256 21604 11284 21632
rect 12066 21604 12072 21616
rect 11011 21576 11284 21604
rect 11348 21576 12072 21604
rect 11011 21573 11023 21576
rect 10965 21567 11023 21573
rect 10870 21496 10876 21548
rect 10928 21536 10934 21548
rect 11057 21539 11115 21545
rect 11057 21536 11069 21539
rect 10928 21508 11069 21536
rect 10928 21496 10934 21508
rect 11057 21505 11069 21508
rect 11103 21536 11115 21539
rect 11348 21536 11376 21576
rect 12066 21564 12072 21576
rect 12124 21564 12130 21616
rect 11103 21508 11376 21536
rect 11517 21539 11575 21545
rect 11103 21505 11115 21508
rect 11057 21499 11115 21505
rect 11517 21505 11529 21539
rect 11563 21536 11575 21539
rect 12406 21536 12434 21644
rect 14734 21632 14740 21644
rect 14792 21632 14798 21684
rect 16390 21632 16396 21684
rect 16448 21632 16454 21684
rect 17218 21632 17224 21684
rect 17276 21632 17282 21684
rect 20070 21672 20076 21684
rect 17604 21644 20076 21672
rect 13280 21576 13676 21604
rect 13280 21545 13308 21576
rect 13648 21548 13676 21576
rect 13814 21564 13820 21616
rect 13872 21604 13878 21616
rect 14001 21607 14059 21613
rect 14001 21604 14013 21607
rect 13872 21576 14013 21604
rect 13872 21564 13878 21576
rect 14001 21573 14013 21576
rect 14047 21573 14059 21607
rect 14001 21567 14059 21573
rect 11563 21508 12434 21536
rect 13265 21539 13323 21545
rect 11563 21505 11575 21508
rect 11517 21499 11575 21505
rect 13265 21505 13277 21539
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 13446 21496 13452 21548
rect 13504 21496 13510 21548
rect 13630 21496 13636 21548
rect 13688 21496 13694 21548
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21536 13783 21539
rect 15930 21536 15936 21548
rect 13771 21508 15936 21536
rect 13771 21505 13783 21508
rect 13725 21499 13783 21505
rect 15930 21496 15936 21508
rect 15988 21496 15994 21548
rect 16408 21536 16436 21632
rect 17604 21604 17632 21644
rect 20070 21632 20076 21644
rect 20128 21632 20134 21684
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 21453 21675 21511 21681
rect 21453 21672 21465 21675
rect 20496 21644 21465 21672
rect 20496 21632 20502 21644
rect 21453 21641 21465 21644
rect 21499 21641 21511 21675
rect 21453 21635 21511 21641
rect 21634 21632 21640 21684
rect 21692 21672 21698 21684
rect 23014 21672 23020 21684
rect 21692 21644 23020 21672
rect 21692 21632 21698 21644
rect 23014 21632 23020 21644
rect 23072 21632 23078 21684
rect 24394 21632 24400 21684
rect 24452 21632 24458 21684
rect 25498 21632 25504 21684
rect 25556 21672 25562 21684
rect 30006 21672 30012 21684
rect 25556 21644 26004 21672
rect 25556 21632 25562 21644
rect 17052 21576 17632 21604
rect 17052 21545 17080 21576
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 16408 21508 17049 21536
rect 17037 21505 17049 21508
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 17221 21539 17279 21545
rect 17221 21505 17233 21539
rect 17267 21536 17279 21539
rect 17497 21539 17555 21545
rect 17267 21534 17356 21536
rect 17497 21534 17509 21539
rect 17267 21508 17509 21534
rect 17267 21505 17279 21508
rect 17328 21506 17509 21508
rect 17221 21499 17279 21505
rect 17497 21505 17509 21506
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 14274 21468 14280 21480
rect 8803 21440 10456 21468
rect 10796 21440 14280 21468
rect 8803 21437 8815 21440
rect 8757 21431 8815 21437
rect 10428 21409 10456 21440
rect 14274 21428 14280 21440
rect 14332 21468 14338 21480
rect 17236 21468 17264 21499
rect 14332 21440 17264 21468
rect 17313 21471 17371 21477
rect 14332 21428 14338 21440
rect 17313 21437 17325 21471
rect 17359 21468 17371 21471
rect 17604 21468 17632 21576
rect 18138 21564 18144 21616
rect 18196 21604 18202 21616
rect 18196 21576 18736 21604
rect 18196 21564 18202 21576
rect 17770 21496 17776 21548
rect 17828 21496 17834 21548
rect 17862 21496 17868 21548
rect 17920 21496 17926 21548
rect 18233 21539 18291 21545
rect 18233 21505 18245 21539
rect 18279 21505 18291 21539
rect 18233 21499 18291 21505
rect 17359 21440 17632 21468
rect 17788 21468 17816 21496
rect 17788 21440 17954 21468
rect 17359 21437 17371 21440
rect 17313 21431 17371 21437
rect 10413 21403 10471 21409
rect 4356 21372 5856 21400
rect 5828 21344 5856 21372
rect 9784 21372 10364 21400
rect 5810 21292 5816 21344
rect 5868 21292 5874 21344
rect 5902 21292 5908 21344
rect 5960 21332 5966 21344
rect 9784 21332 9812 21372
rect 5960 21304 9812 21332
rect 10336 21332 10364 21372
rect 10413 21369 10425 21403
rect 10459 21369 10471 21403
rect 13814 21400 13820 21412
rect 10413 21363 10471 21369
rect 10520 21372 13820 21400
rect 10520 21332 10548 21372
rect 13814 21360 13820 21372
rect 13872 21360 13878 21412
rect 14001 21403 14059 21409
rect 14001 21369 14013 21403
rect 14047 21400 14059 21403
rect 14090 21400 14096 21412
rect 14047 21372 14096 21400
rect 14047 21369 14059 21372
rect 14001 21363 14059 21369
rect 14090 21360 14096 21372
rect 14148 21360 14154 21412
rect 17770 21360 17776 21412
rect 17828 21360 17834 21412
rect 17926 21400 17954 21440
rect 18138 21428 18144 21480
rect 18196 21468 18202 21480
rect 18254 21468 18282 21499
rect 18414 21496 18420 21548
rect 18472 21496 18478 21548
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21526 18567 21539
rect 18598 21526 18604 21548
rect 18555 21505 18604 21526
rect 18509 21499 18604 21505
rect 18524 21498 18604 21499
rect 18598 21496 18604 21498
rect 18656 21496 18662 21548
rect 18196 21440 18282 21468
rect 18708 21468 18736 21576
rect 18800 21576 20392 21604
rect 18800 21545 18828 21576
rect 20364 21548 20392 21576
rect 20622 21564 20628 21616
rect 20680 21604 20686 21616
rect 20680 21576 22692 21604
rect 20680 21564 20686 21576
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 19058 21496 19064 21548
rect 19116 21496 19122 21548
rect 20346 21496 20352 21548
rect 20404 21496 20410 21548
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 21542 21536 21548 21548
rect 21131 21508 21548 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 21542 21496 21548 21508
rect 21600 21536 21606 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21600 21508 21833 21536
rect 21600 21496 21606 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 21910 21496 21916 21548
rect 21968 21536 21974 21548
rect 22664 21545 22692 21576
rect 23474 21564 23480 21616
rect 23532 21564 23538 21616
rect 24412 21604 24440 21632
rect 23676 21576 24440 21604
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 21968 21508 22201 21536
rect 21968 21496 21974 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21505 22707 21539
rect 22649 21499 22707 21505
rect 18877 21471 18935 21477
rect 18877 21468 18889 21471
rect 18708 21440 18889 21468
rect 18196 21428 18202 21440
rect 18877 21437 18889 21440
rect 18923 21437 18935 21471
rect 18877 21431 18935 21437
rect 18969 21471 19027 21477
rect 18969 21437 18981 21471
rect 19015 21437 19027 21471
rect 18969 21431 19027 21437
rect 18984 21400 19012 21431
rect 20162 21428 20168 21480
rect 20220 21468 20226 21480
rect 21177 21471 21235 21477
rect 21177 21468 21189 21471
rect 20220 21440 21189 21468
rect 20220 21428 20226 21440
rect 21177 21437 21189 21440
rect 21223 21437 21235 21471
rect 21177 21431 21235 21437
rect 21634 21428 21640 21480
rect 21692 21428 21698 21480
rect 23676 21477 23704 21576
rect 25222 21564 25228 21616
rect 25280 21604 25286 21616
rect 25976 21613 26004 21644
rect 26988 21644 30012 21672
rect 25961 21607 26019 21613
rect 25280 21576 25912 21604
rect 25280 21564 25286 21576
rect 25884 21548 25912 21576
rect 25961 21573 25973 21607
rect 26007 21573 26019 21607
rect 25961 21567 26019 21573
rect 23750 21496 23756 21548
rect 23808 21536 23814 21548
rect 23845 21539 23903 21545
rect 23845 21536 23857 21539
rect 23808 21508 23857 21536
rect 23808 21496 23814 21508
rect 23845 21505 23857 21508
rect 23891 21505 23903 21539
rect 23845 21499 23903 21505
rect 25590 21496 25596 21548
rect 25648 21496 25654 21548
rect 25682 21496 25688 21548
rect 25740 21496 25746 21548
rect 25866 21496 25872 21548
rect 25924 21496 25930 21548
rect 26142 21545 26148 21548
rect 26099 21539 26148 21545
rect 26099 21505 26111 21539
rect 26145 21505 26148 21539
rect 26099 21499 26148 21505
rect 26142 21496 26148 21499
rect 26200 21496 26206 21548
rect 26326 21496 26332 21548
rect 26384 21496 26390 21548
rect 23661 21471 23719 21477
rect 23661 21437 23673 21471
rect 23707 21437 23719 21471
rect 23661 21431 23719 21437
rect 26602 21428 26608 21480
rect 26660 21428 26666 21480
rect 26786 21428 26792 21480
rect 26844 21468 26850 21480
rect 26988 21477 27016 21644
rect 30006 21632 30012 21644
rect 30064 21632 30070 21684
rect 31478 21672 31484 21684
rect 30668 21644 31484 21672
rect 28626 21564 28632 21616
rect 28684 21604 28690 21616
rect 29273 21607 29331 21613
rect 29273 21604 29285 21607
rect 28684 21576 29285 21604
rect 28684 21564 28690 21576
rect 29273 21573 29285 21576
rect 29319 21573 29331 21607
rect 29273 21567 29331 21573
rect 30558 21564 30564 21616
rect 30616 21604 30622 21616
rect 30668 21604 30696 21644
rect 31144 21613 31172 21644
rect 31478 21632 31484 21644
rect 31536 21632 31542 21684
rect 31570 21632 31576 21684
rect 31628 21632 31634 21684
rect 32214 21632 32220 21684
rect 32272 21632 32278 21684
rect 37001 21675 37059 21681
rect 36004 21644 36768 21672
rect 30955 21607 31013 21613
rect 30955 21604 30967 21607
rect 30616 21576 30696 21604
rect 30616 21564 30622 21576
rect 30668 21545 30696 21576
rect 30944 21573 30967 21604
rect 31001 21573 31013 21607
rect 30944 21567 31013 21573
rect 31129 21607 31187 21613
rect 31129 21573 31141 21607
rect 31175 21573 31187 21607
rect 31389 21607 31447 21613
rect 31389 21604 31401 21607
rect 31129 21567 31187 21573
rect 31220 21576 31401 21604
rect 30653 21539 30711 21545
rect 28382 21508 28672 21536
rect 26973 21471 27031 21477
rect 26973 21468 26985 21471
rect 26844 21440 26985 21468
rect 26844 21428 26850 21440
rect 26973 21437 26985 21440
rect 27019 21437 27031 21471
rect 27249 21471 27307 21477
rect 27249 21468 27261 21471
rect 26973 21431 27031 21437
rect 27080 21440 27261 21468
rect 17926 21372 19012 21400
rect 19242 21360 19248 21412
rect 19300 21400 19306 21412
rect 21652 21400 21680 21428
rect 19300 21372 21680 21400
rect 19300 21360 19306 21372
rect 22646 21360 22652 21412
rect 22704 21360 22710 21412
rect 23753 21403 23811 21409
rect 23753 21369 23765 21403
rect 23799 21400 23811 21403
rect 23842 21400 23848 21412
rect 23799 21372 23848 21400
rect 23799 21369 23811 21372
rect 23753 21363 23811 21369
rect 23842 21360 23848 21372
rect 23900 21360 23906 21412
rect 26237 21403 26295 21409
rect 26237 21369 26249 21403
rect 26283 21400 26295 21403
rect 27080 21400 27108 21440
rect 27249 21437 27261 21440
rect 27295 21437 27307 21471
rect 27249 21431 27307 21437
rect 28534 21428 28540 21480
rect 28592 21428 28598 21480
rect 26283 21372 27108 21400
rect 26283 21369 26295 21372
rect 26237 21363 26295 21369
rect 10336 21304 10548 21332
rect 11701 21335 11759 21341
rect 5960 21292 5966 21304
rect 11701 21301 11713 21335
rect 11747 21332 11759 21335
rect 12066 21332 12072 21344
rect 11747 21304 12072 21332
rect 11747 21301 11759 21304
rect 11701 21295 11759 21301
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 12526 21292 12532 21344
rect 12584 21332 12590 21344
rect 17954 21332 17960 21344
rect 12584 21304 17960 21332
rect 12584 21292 12590 21304
rect 17954 21292 17960 21304
rect 18012 21292 18018 21344
rect 18049 21335 18107 21341
rect 18049 21301 18061 21335
rect 18095 21332 18107 21335
rect 18506 21332 18512 21344
rect 18095 21304 18512 21332
rect 18095 21301 18107 21304
rect 18049 21295 18107 21301
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 18598 21292 18604 21344
rect 18656 21292 18662 21344
rect 21269 21335 21327 21341
rect 21269 21301 21281 21335
rect 21315 21332 21327 21335
rect 22002 21332 22008 21344
rect 21315 21304 22008 21332
rect 21315 21301 21327 21304
rect 21269 21295 21327 21301
rect 22002 21292 22008 21304
rect 22060 21292 22066 21344
rect 23474 21292 23480 21344
rect 23532 21292 23538 21344
rect 28552 21332 28580 21428
rect 28644 21412 28672 21508
rect 30653 21505 30665 21539
rect 30699 21505 30711 21539
rect 30653 21499 30711 21505
rect 30837 21539 30895 21545
rect 30837 21505 30849 21539
rect 30883 21505 30895 21539
rect 30944 21536 30972 21567
rect 31220 21536 31248 21576
rect 31389 21573 31401 21576
rect 31435 21604 31447 21607
rect 31849 21607 31907 21613
rect 31849 21604 31861 21607
rect 31435 21576 31861 21604
rect 31435 21573 31447 21576
rect 31389 21567 31447 21573
rect 31849 21573 31861 21576
rect 31895 21573 31907 21607
rect 32232 21604 32260 21632
rect 36004 21613 36032 21644
rect 35989 21607 36047 21613
rect 35989 21604 36001 21607
rect 31849 21567 31907 21573
rect 32140 21576 32260 21604
rect 35912 21576 36001 21604
rect 30944 21508 31248 21536
rect 30837 21499 30895 21505
rect 29362 21428 29368 21480
rect 29420 21428 29426 21480
rect 29454 21428 29460 21480
rect 29512 21428 29518 21480
rect 28626 21360 28632 21412
rect 28684 21360 28690 21412
rect 30852 21400 30880 21499
rect 31478 21496 31484 21548
rect 31536 21536 31542 21548
rect 32140 21545 32168 21576
rect 31665 21539 31723 21545
rect 31665 21536 31677 21539
rect 31536 21508 31677 21536
rect 31536 21496 31542 21508
rect 31665 21505 31677 21508
rect 31711 21505 31723 21539
rect 31665 21499 31723 21505
rect 31757 21539 31815 21545
rect 31757 21505 31769 21539
rect 31803 21505 31815 21539
rect 31757 21499 31815 21505
rect 32125 21539 32183 21545
rect 32125 21505 32137 21539
rect 32171 21505 32183 21539
rect 32125 21499 32183 21505
rect 31570 21428 31576 21480
rect 31628 21428 31634 21480
rect 31588 21400 31616 21428
rect 30852 21372 31616 21400
rect 28721 21335 28779 21341
rect 28721 21332 28733 21335
rect 28552 21304 28733 21332
rect 28721 21301 28733 21304
rect 28767 21301 28779 21335
rect 28721 21295 28779 21301
rect 28902 21292 28908 21344
rect 28960 21292 28966 21344
rect 30745 21335 30803 21341
rect 30745 21301 30757 21335
rect 30791 21332 30803 21335
rect 31018 21332 31024 21344
rect 30791 21304 31024 21332
rect 30791 21301 30803 21304
rect 30745 21295 30803 21301
rect 31018 21292 31024 21304
rect 31076 21292 31082 21344
rect 31128 21341 31156 21372
rect 31113 21335 31171 21341
rect 31113 21301 31125 21335
rect 31159 21301 31171 21335
rect 31113 21295 31171 21301
rect 31202 21292 31208 21344
rect 31260 21332 31266 21344
rect 31297 21335 31355 21341
rect 31297 21332 31309 21335
rect 31260 21304 31309 21332
rect 31260 21292 31266 21304
rect 31297 21301 31309 21304
rect 31343 21301 31355 21335
rect 31297 21295 31355 21301
rect 31386 21292 31392 21344
rect 31444 21292 31450 21344
rect 31772 21332 31800 21499
rect 32401 21471 32459 21477
rect 32401 21437 32413 21471
rect 32447 21468 32459 21471
rect 32490 21468 32496 21480
rect 32447 21440 32496 21468
rect 32447 21437 32459 21440
rect 32401 21431 32459 21437
rect 32490 21428 32496 21440
rect 32548 21428 32554 21480
rect 33134 21428 33140 21480
rect 33192 21468 33198 21480
rect 33520 21468 33548 21522
rect 33686 21496 33692 21548
rect 33744 21536 33750 21548
rect 35912 21545 35940 21576
rect 35989 21573 36001 21576
rect 36035 21573 36047 21607
rect 35989 21567 36047 21573
rect 36357 21607 36415 21613
rect 36357 21573 36369 21607
rect 36403 21604 36415 21607
rect 36633 21607 36691 21613
rect 36633 21604 36645 21607
rect 36403 21576 36645 21604
rect 36403 21573 36415 21576
rect 36357 21567 36415 21573
rect 36633 21573 36645 21576
rect 36679 21573 36691 21607
rect 36740 21604 36768 21644
rect 37001 21641 37013 21675
rect 37047 21672 37059 21675
rect 37458 21672 37464 21684
rect 37047 21644 37464 21672
rect 37047 21641 37059 21644
rect 37001 21635 37059 21641
rect 37458 21632 37464 21644
rect 37516 21632 37522 21684
rect 36740 21576 37320 21604
rect 36633 21567 36691 21573
rect 37292 21548 37320 21576
rect 35621 21539 35679 21545
rect 35621 21536 35633 21539
rect 33744 21508 35633 21536
rect 33744 21496 33750 21508
rect 33192 21440 33548 21468
rect 34149 21471 34207 21477
rect 33192 21428 33198 21440
rect 34149 21437 34161 21471
rect 34195 21437 34207 21471
rect 34149 21431 34207 21437
rect 32214 21332 32220 21344
rect 31772 21304 32220 21332
rect 32214 21292 32220 21304
rect 32272 21332 32278 21344
rect 34164 21332 34192 21431
rect 32272 21304 34192 21332
rect 35544 21332 35572 21508
rect 35621 21505 35633 21508
rect 35667 21505 35679 21539
rect 35621 21499 35679 21505
rect 35805 21539 35863 21545
rect 35805 21505 35817 21539
rect 35851 21505 35863 21539
rect 35805 21499 35863 21505
rect 35897 21539 35955 21545
rect 35897 21505 35909 21539
rect 35943 21505 35955 21539
rect 36173 21539 36231 21545
rect 36173 21536 36185 21539
rect 35897 21499 35955 21505
rect 36096 21508 36185 21536
rect 35820 21468 35848 21499
rect 36096 21480 36124 21508
rect 36173 21505 36185 21508
rect 36219 21505 36231 21539
rect 36173 21499 36231 21505
rect 36449 21539 36507 21545
rect 36449 21505 36461 21539
rect 36495 21505 36507 21539
rect 36725 21539 36783 21545
rect 36725 21536 36737 21539
rect 36449 21499 36507 21505
rect 36556 21508 36737 21536
rect 36078 21468 36084 21480
rect 35820 21440 36084 21468
rect 36078 21428 36084 21440
rect 36136 21428 36142 21480
rect 35621 21403 35679 21409
rect 35621 21369 35633 21403
rect 35667 21400 35679 21403
rect 36464 21400 36492 21499
rect 35667 21372 36492 21400
rect 35667 21369 35679 21372
rect 35621 21363 35679 21369
rect 36556 21332 36584 21508
rect 36725 21505 36737 21508
rect 36771 21505 36783 21539
rect 36725 21499 36783 21505
rect 36814 21496 36820 21548
rect 36872 21496 36878 21548
rect 37274 21496 37280 21548
rect 37332 21496 37338 21548
rect 35544 21304 36584 21332
rect 32272 21292 32278 21304
rect 1104 21242 41400 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 41400 21242
rect 1104 21168 41400 21190
rect 4525 21131 4583 21137
rect 4525 21097 4537 21131
rect 4571 21128 4583 21131
rect 4614 21128 4620 21140
rect 4571 21100 4620 21128
rect 4571 21097 4583 21100
rect 4525 21091 4583 21097
rect 4614 21088 4620 21100
rect 4672 21088 4678 21140
rect 5902 21088 5908 21140
rect 5960 21088 5966 21140
rect 6273 21131 6331 21137
rect 6273 21097 6285 21131
rect 6319 21128 6331 21131
rect 6638 21128 6644 21140
rect 6319 21100 6644 21128
rect 6319 21097 6331 21100
rect 6273 21091 6331 21097
rect 6638 21088 6644 21100
rect 6696 21088 6702 21140
rect 6730 21088 6736 21140
rect 6788 21128 6794 21140
rect 7837 21131 7895 21137
rect 7837 21128 7849 21131
rect 6788 21100 7849 21128
rect 6788 21088 6794 21100
rect 7837 21097 7849 21100
rect 7883 21097 7895 21131
rect 7837 21091 7895 21097
rect 7926 21088 7932 21140
rect 7984 21088 7990 21140
rect 10597 21131 10655 21137
rect 10597 21097 10609 21131
rect 10643 21097 10655 21131
rect 10597 21091 10655 21097
rect 4709 20927 4767 20933
rect 4709 20893 4721 20927
rect 4755 20924 4767 20927
rect 5626 20924 5632 20936
rect 4755 20896 5632 20924
rect 4755 20893 4767 20896
rect 4709 20887 4767 20893
rect 5626 20884 5632 20896
rect 5684 20884 5690 20936
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20924 5779 20927
rect 5920 20924 5948 21088
rect 6914 21020 6920 21072
rect 6972 21060 6978 21072
rect 7101 21063 7159 21069
rect 7101 21060 7113 21063
rect 6972 21032 7113 21060
rect 6972 21020 6978 21032
rect 7101 21029 7113 21032
rect 7147 21029 7159 21063
rect 7944 21060 7972 21088
rect 7101 21023 7159 21029
rect 7208 21032 7972 21060
rect 6454 20952 6460 21004
rect 6512 20952 6518 21004
rect 6825 20995 6883 21001
rect 6825 20961 6837 20995
rect 6871 20992 6883 20995
rect 7208 20992 7236 21032
rect 6871 20964 7236 20992
rect 6871 20961 6883 20964
rect 6825 20955 6883 20961
rect 5767 20896 5948 20924
rect 6549 20927 6607 20933
rect 5767 20893 5779 20896
rect 5721 20887 5779 20893
rect 6549 20893 6561 20927
rect 6595 20924 6607 20927
rect 6638 20924 6644 20936
rect 6595 20896 6644 20924
rect 6595 20893 6607 20896
rect 6549 20887 6607 20893
rect 6638 20884 6644 20896
rect 6696 20884 6702 20936
rect 6914 20884 6920 20936
rect 6972 20884 6978 20936
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7208 20924 7236 20964
rect 7469 20995 7527 21001
rect 7469 20961 7481 20995
rect 7515 20992 7527 20995
rect 7558 20992 7564 21004
rect 7515 20964 7564 20992
rect 7515 20961 7527 20964
rect 7469 20955 7527 20961
rect 7147 20896 7236 20924
rect 7285 20927 7343 20933
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 7484 20924 7512 20955
rect 7558 20952 7564 20964
rect 7616 20952 7622 21004
rect 7331 20896 7512 20924
rect 7653 20927 7711 20933
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 7653 20893 7665 20927
rect 7699 20924 7711 20927
rect 7944 20924 7972 21032
rect 9214 21020 9220 21072
rect 9272 21060 9278 21072
rect 10612 21060 10640 21091
rect 10686 21088 10692 21140
rect 10744 21128 10750 21140
rect 10781 21131 10839 21137
rect 10781 21128 10793 21131
rect 10744 21100 10793 21128
rect 10744 21088 10750 21100
rect 10781 21097 10793 21100
rect 10827 21097 10839 21131
rect 10781 21091 10839 21097
rect 11514 21088 11520 21140
rect 11572 21088 11578 21140
rect 13357 21131 13415 21137
rect 13357 21097 13369 21131
rect 13403 21128 13415 21131
rect 13538 21128 13544 21140
rect 13403 21100 13544 21128
rect 13403 21097 13415 21100
rect 13357 21091 13415 21097
rect 11532 21060 11560 21088
rect 13372 21060 13400 21091
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 13814 21088 13820 21140
rect 13872 21128 13878 21140
rect 16114 21128 16120 21140
rect 13872 21100 16120 21128
rect 13872 21088 13878 21100
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 17494 21088 17500 21140
rect 17552 21128 17558 21140
rect 17770 21128 17776 21140
rect 17552 21100 17776 21128
rect 17552 21088 17558 21100
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 18230 21088 18236 21140
rect 18288 21128 18294 21140
rect 18414 21128 18420 21140
rect 18288 21100 18420 21128
rect 18288 21088 18294 21100
rect 18414 21088 18420 21100
rect 18472 21088 18478 21140
rect 18598 21088 18604 21140
rect 18656 21128 18662 21140
rect 18656 21100 22094 21128
rect 18656 21088 18662 21100
rect 9272 21032 10548 21060
rect 10612 21032 11560 21060
rect 12544 21032 13400 21060
rect 9272 21020 9278 21032
rect 9968 21001 9996 21032
rect 9953 20995 10011 21001
rect 9953 20961 9965 20995
rect 9999 20961 10011 20995
rect 9953 20955 10011 20961
rect 10226 20952 10232 21004
rect 10284 20992 10290 21004
rect 10520 20992 10548 21032
rect 12544 21004 12572 21032
rect 13906 21020 13912 21072
rect 13964 21060 13970 21072
rect 18782 21060 18788 21072
rect 13964 21032 18788 21060
rect 13964 21020 13970 21032
rect 18782 21020 18788 21032
rect 18840 21020 18846 21072
rect 22066 21060 22094 21100
rect 23474 21088 23480 21140
rect 23532 21088 23538 21140
rect 28077 21131 28135 21137
rect 28077 21128 28089 21131
rect 25240 21100 28089 21128
rect 23382 21060 23388 21072
rect 22066 21032 23388 21060
rect 23382 21020 23388 21032
rect 23440 21020 23446 21072
rect 10284 20964 10456 20992
rect 10520 20964 11192 20992
rect 10284 20952 10290 20964
rect 10428 20933 10456 20964
rect 11164 20936 11192 20964
rect 12158 20952 12164 21004
rect 12216 20952 12222 21004
rect 12250 20952 12256 21004
rect 12308 20952 12314 21004
rect 12526 20952 12532 21004
rect 12584 20952 12590 21004
rect 12805 20995 12863 21001
rect 12805 20961 12817 20995
rect 12851 20992 12863 20995
rect 13814 20992 13820 21004
rect 12851 20964 13820 20992
rect 12851 20961 12863 20964
rect 12805 20955 12863 20961
rect 13814 20952 13820 20964
rect 13872 20952 13878 21004
rect 16022 20952 16028 21004
rect 16080 20952 16086 21004
rect 16298 20952 16304 21004
rect 16356 20992 16362 21004
rect 17221 20995 17279 21001
rect 17221 20992 17233 20995
rect 16356 20964 17233 20992
rect 16356 20952 16362 20964
rect 17221 20961 17233 20964
rect 17267 20961 17279 20995
rect 23492 20992 23520 21088
rect 24762 21020 24768 21072
rect 24820 21060 24826 21072
rect 25240 21060 25268 21100
rect 28077 21097 28089 21100
rect 28123 21097 28135 21131
rect 28077 21091 28135 21097
rect 24820 21032 25268 21060
rect 24820 21020 24826 21032
rect 25866 21020 25872 21072
rect 25924 21060 25930 21072
rect 27709 21063 27767 21069
rect 27709 21060 27721 21063
rect 25924 21032 27721 21060
rect 25924 21020 25930 21032
rect 27709 21029 27721 21032
rect 27755 21029 27767 21063
rect 28092 21060 28120 21091
rect 28258 21088 28264 21140
rect 28316 21088 28322 21140
rect 28442 21088 28448 21140
rect 28500 21088 28506 21140
rect 29270 21128 29276 21140
rect 28552 21100 29276 21128
rect 28460 21060 28488 21088
rect 28092 21032 28488 21060
rect 27709 21023 27767 21029
rect 17221 20955 17279 20961
rect 19536 20964 23520 20992
rect 7699 20896 7972 20924
rect 9677 20927 9735 20933
rect 7699 20893 7711 20896
rect 7653 20887 7711 20893
rect 9677 20893 9689 20927
rect 9723 20924 9735 20927
rect 10413 20927 10471 20933
rect 9723 20896 10364 20924
rect 9723 20893 9735 20896
rect 9677 20887 9735 20893
rect 5810 20816 5816 20868
rect 5868 20856 5874 20868
rect 10336 20856 10364 20896
rect 10413 20893 10425 20927
rect 10459 20893 10471 20927
rect 10413 20887 10471 20893
rect 10502 20884 10508 20936
rect 10560 20884 10566 20936
rect 11146 20884 11152 20936
rect 11204 20884 11210 20936
rect 12066 20884 12072 20936
rect 12124 20884 12130 20936
rect 12618 20884 12624 20936
rect 12676 20924 12682 20936
rect 12897 20927 12955 20933
rect 12897 20924 12909 20927
rect 12676 20896 12909 20924
rect 12676 20884 12682 20896
rect 12897 20893 12909 20896
rect 12943 20893 12955 20927
rect 15930 20924 15936 20936
rect 12897 20887 12955 20893
rect 13004 20896 15936 20924
rect 12084 20856 12112 20884
rect 13004 20856 13032 20896
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 16390 20884 16396 20936
rect 16448 20884 16454 20936
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 16761 20927 16819 20933
rect 16761 20924 16773 20927
rect 16540 20896 16773 20924
rect 16540 20884 16546 20896
rect 16761 20893 16773 20896
rect 16807 20893 16819 20927
rect 16761 20887 16819 20893
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20924 17003 20927
rect 17126 20924 17132 20936
rect 16991 20896 17132 20924
rect 16991 20893 17003 20896
rect 16945 20887 17003 20893
rect 5868 20828 7052 20856
rect 5868 20816 5874 20828
rect 6733 20791 6791 20797
rect 6733 20757 6745 20791
rect 6779 20788 6791 20791
rect 6914 20788 6920 20800
rect 6779 20760 6920 20788
rect 6779 20757 6791 20760
rect 6733 20751 6791 20757
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 7024 20788 7052 20828
rect 7484 20828 7972 20856
rect 10336 20828 12112 20856
rect 12406 20828 13032 20856
rect 13081 20859 13139 20865
rect 7484 20788 7512 20828
rect 7024 20760 7512 20788
rect 7944 20788 7972 20828
rect 12406 20788 12434 20828
rect 13081 20825 13093 20859
rect 13127 20825 13139 20859
rect 13081 20819 13139 20825
rect 7944 20760 12434 20788
rect 12894 20748 12900 20800
rect 12952 20788 12958 20800
rect 13096 20788 13124 20819
rect 14182 20816 14188 20868
rect 14240 20856 14246 20868
rect 15838 20856 15844 20868
rect 14240 20828 15844 20856
rect 14240 20816 14246 20828
rect 15838 20816 15844 20828
rect 15896 20816 15902 20868
rect 16850 20856 16856 20868
rect 16132 20828 16856 20856
rect 16132 20788 16160 20828
rect 16850 20816 16856 20828
rect 16908 20816 16914 20868
rect 12952 20760 16160 20788
rect 12952 20748 12958 20760
rect 16206 20748 16212 20800
rect 16264 20788 16270 20800
rect 16960 20788 16988 20887
rect 17126 20884 17132 20896
rect 17184 20884 17190 20936
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 18966 20924 18972 20936
rect 18012 20896 18972 20924
rect 18012 20884 18018 20896
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 19536 20933 19564 20964
rect 23934 20952 23940 21004
rect 23992 20992 23998 21004
rect 24673 20995 24731 21001
rect 24673 20992 24685 20995
rect 23992 20964 24685 20992
rect 23992 20952 23998 20964
rect 24673 20961 24685 20964
rect 24719 20961 24731 20995
rect 27154 20992 27160 21004
rect 24673 20955 24731 20961
rect 24780 20964 27160 20992
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20254 20924 20260 20936
rect 20027 20896 20260 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 19812 20856 19840 20887
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 21634 20884 21640 20936
rect 21692 20924 21698 20936
rect 24780 20924 24808 20964
rect 27154 20952 27160 20964
rect 27212 20952 27218 21004
rect 27522 20992 27528 21004
rect 27264 20964 27528 20992
rect 21692 20896 24808 20924
rect 21692 20884 21698 20896
rect 24854 20884 24860 20936
rect 24912 20884 24918 20936
rect 27264 20933 27292 20964
rect 27522 20952 27528 20964
rect 27580 20992 27586 21004
rect 28552 20992 28580 21100
rect 29270 21088 29276 21100
rect 29328 21088 29334 21140
rect 29362 21088 29368 21140
rect 29420 21128 29426 21140
rect 29917 21131 29975 21137
rect 29917 21128 29929 21131
rect 29420 21100 29929 21128
rect 29420 21088 29426 21100
rect 29917 21097 29929 21100
rect 29963 21097 29975 21131
rect 39114 21128 39120 21140
rect 29917 21091 29975 21097
rect 31726 21100 39120 21128
rect 31726 21060 31754 21100
rect 39114 21088 39120 21100
rect 39172 21088 39178 21140
rect 27580 20964 28580 20992
rect 28644 21032 31754 21060
rect 27580 20952 27586 20964
rect 27065 20927 27123 20933
rect 27065 20893 27077 20927
rect 27111 20893 27123 20927
rect 27065 20887 27123 20893
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20893 27307 20927
rect 27249 20887 27307 20893
rect 27080 20856 27108 20887
rect 27430 20884 27436 20936
rect 27488 20924 27494 20936
rect 28644 20924 28672 21032
rect 35802 21020 35808 21072
rect 35860 21060 35866 21072
rect 35860 21032 40724 21060
rect 35860 21020 35866 21032
rect 29546 20952 29552 21004
rect 29604 20992 29610 21004
rect 30282 20992 30288 21004
rect 29604 20964 30288 20992
rect 29604 20952 29610 20964
rect 30282 20952 30288 20964
rect 30340 20952 30346 21004
rect 31294 20992 31300 21004
rect 31036 20964 31300 20992
rect 27488 20896 28672 20924
rect 28721 20927 28779 20933
rect 27488 20884 27494 20896
rect 28721 20893 28733 20927
rect 28767 20924 28779 20927
rect 28902 20924 28908 20936
rect 28767 20896 28908 20924
rect 28767 20893 28779 20896
rect 28721 20887 28779 20893
rect 28902 20884 28908 20896
rect 28960 20884 28966 20936
rect 28994 20884 29000 20936
rect 29052 20884 29058 20936
rect 31036 20933 31064 20964
rect 31294 20952 31300 20964
rect 31352 20952 31358 21004
rect 31941 20995 31999 21001
rect 31941 20961 31953 20995
rect 31987 20992 31999 20995
rect 31987 20964 32168 20992
rect 31987 20961 31999 20964
rect 31941 20955 31999 20961
rect 29733 20927 29791 20933
rect 29733 20893 29745 20927
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 30745 20927 30803 20933
rect 30745 20893 30757 20927
rect 30791 20893 30803 20927
rect 30745 20887 30803 20893
rect 30929 20927 30987 20933
rect 30929 20893 30941 20927
rect 30975 20924 30987 20927
rect 31021 20927 31079 20933
rect 31021 20924 31033 20927
rect 30975 20896 31033 20924
rect 30975 20893 30987 20896
rect 30929 20887 30987 20893
rect 31021 20893 31033 20896
rect 31067 20893 31079 20927
rect 31021 20887 31079 20893
rect 28077 20859 28135 20865
rect 28077 20856 28089 20859
rect 19812 20828 20024 20856
rect 27080 20828 28089 20856
rect 19996 20800 20024 20828
rect 28077 20825 28089 20828
rect 28123 20856 28135 20859
rect 28166 20856 28172 20868
rect 28123 20828 28172 20856
rect 28123 20825 28135 20828
rect 28077 20819 28135 20825
rect 28166 20816 28172 20828
rect 28224 20856 28230 20868
rect 29748 20856 29776 20887
rect 28224 20828 29776 20856
rect 30760 20856 30788 20887
rect 31202 20884 31208 20936
rect 31260 20924 31266 20936
rect 31389 20927 31447 20933
rect 31389 20924 31401 20927
rect 31260 20896 31401 20924
rect 31260 20884 31266 20896
rect 31389 20893 31401 20896
rect 31435 20893 31447 20927
rect 31389 20887 31447 20893
rect 31478 20884 31484 20936
rect 31536 20924 31542 20936
rect 31665 20927 31723 20933
rect 31665 20924 31677 20927
rect 31536 20896 31677 20924
rect 31536 20884 31542 20896
rect 31665 20893 31677 20896
rect 31711 20924 31723 20927
rect 32033 20927 32091 20933
rect 32033 20924 32045 20927
rect 31711 20896 32045 20924
rect 31711 20893 31723 20896
rect 31665 20887 31723 20893
rect 32033 20893 32045 20896
rect 32079 20893 32091 20927
rect 32033 20887 32091 20893
rect 31220 20856 31248 20884
rect 30760 20828 31248 20856
rect 28224 20816 28230 20828
rect 31294 20816 31300 20868
rect 31352 20816 31358 20868
rect 16264 20760 16988 20788
rect 16264 20748 16270 20760
rect 17034 20748 17040 20800
rect 17092 20788 17098 20800
rect 17862 20788 17868 20800
rect 17092 20760 17868 20788
rect 17092 20748 17098 20760
rect 17862 20748 17868 20760
rect 17920 20748 17926 20800
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 19705 20791 19763 20797
rect 19705 20788 19717 20791
rect 18380 20760 19717 20788
rect 18380 20748 18386 20760
rect 19705 20757 19717 20760
rect 19751 20757 19763 20791
rect 19705 20751 19763 20757
rect 19886 20748 19892 20800
rect 19944 20748 19950 20800
rect 19978 20748 19984 20800
rect 20036 20748 20042 20800
rect 25038 20748 25044 20800
rect 25096 20748 25102 20800
rect 25866 20748 25872 20800
rect 25924 20788 25930 20800
rect 26418 20788 26424 20800
rect 25924 20760 26424 20788
rect 25924 20748 25930 20760
rect 26418 20748 26424 20760
rect 26476 20748 26482 20800
rect 27154 20748 27160 20800
rect 27212 20748 27218 20800
rect 28534 20748 28540 20800
rect 28592 20748 28598 20800
rect 28902 20748 28908 20800
rect 28960 20748 28966 20800
rect 30837 20791 30895 20797
rect 30837 20757 30849 20791
rect 30883 20788 30895 20791
rect 32140 20788 32168 20964
rect 34514 20952 34520 21004
rect 34572 20992 34578 21004
rect 34701 20995 34759 21001
rect 34701 20992 34713 20995
rect 34572 20964 34713 20992
rect 34572 20952 34578 20964
rect 34701 20961 34713 20964
rect 34747 20961 34759 20995
rect 34701 20955 34759 20961
rect 35529 20995 35587 21001
rect 35529 20961 35541 20995
rect 35575 20992 35587 20995
rect 35575 20964 35756 20992
rect 35575 20961 35587 20964
rect 35529 20955 35587 20961
rect 35161 20927 35219 20933
rect 35161 20924 35173 20927
rect 34716 20896 35173 20924
rect 34716 20800 34744 20896
rect 35161 20893 35173 20896
rect 35207 20893 35219 20927
rect 35161 20887 35219 20893
rect 35250 20884 35256 20936
rect 35308 20924 35314 20936
rect 35728 20933 35756 20964
rect 35443 20927 35501 20933
rect 35443 20926 35455 20927
rect 35360 20924 35455 20926
rect 35308 20898 35455 20924
rect 35308 20896 35388 20898
rect 35308 20884 35314 20896
rect 35443 20893 35455 20898
rect 35489 20893 35501 20927
rect 35621 20927 35679 20933
rect 35621 20924 35633 20927
rect 35443 20887 35501 20893
rect 35544 20896 35633 20924
rect 35544 20868 35572 20896
rect 35621 20893 35633 20896
rect 35667 20893 35679 20927
rect 35621 20887 35679 20893
rect 35719 20927 35777 20933
rect 35719 20893 35731 20927
rect 35765 20893 35777 20927
rect 35719 20887 35777 20893
rect 35891 20927 35949 20933
rect 35891 20902 35903 20927
rect 35937 20902 35949 20927
rect 35891 20887 35900 20902
rect 35526 20816 35532 20868
rect 35584 20816 35590 20868
rect 35894 20850 35900 20887
rect 35952 20850 35958 20902
rect 35986 20884 35992 20936
rect 36044 20884 36050 20936
rect 40696 20933 40724 21032
rect 36173 20927 36231 20933
rect 36173 20893 36185 20927
rect 36219 20893 36231 20927
rect 36173 20887 36231 20893
rect 40681 20927 40739 20933
rect 40681 20893 40693 20927
rect 40727 20893 40739 20927
rect 40681 20887 40739 20893
rect 36188 20800 36216 20887
rect 37642 20816 37648 20868
rect 37700 20856 37706 20868
rect 38381 20859 38439 20865
rect 38381 20856 38393 20859
rect 37700 20828 38393 20856
rect 37700 20816 37706 20828
rect 38381 20825 38393 20828
rect 38427 20856 38439 20859
rect 38562 20856 38568 20868
rect 38427 20828 38568 20856
rect 38427 20825 38439 20828
rect 38381 20819 38439 20825
rect 38562 20816 38568 20828
rect 38620 20816 38626 20868
rect 38838 20816 38844 20868
rect 38896 20816 38902 20868
rect 39022 20816 39028 20868
rect 39080 20816 39086 20868
rect 30883 20760 32168 20788
rect 30883 20757 30895 20760
rect 30837 20751 30895 20757
rect 32398 20748 32404 20800
rect 32456 20748 32462 20800
rect 34698 20748 34704 20800
rect 34756 20748 34762 20800
rect 34790 20748 34796 20800
rect 34848 20788 34854 20800
rect 34977 20791 35035 20797
rect 34977 20788 34989 20791
rect 34848 20760 34989 20788
rect 34848 20748 34854 20760
rect 34977 20757 34989 20760
rect 35023 20757 35035 20791
rect 34977 20751 35035 20757
rect 35069 20791 35127 20797
rect 35069 20757 35081 20791
rect 35115 20788 35127 20791
rect 35802 20788 35808 20800
rect 35115 20760 35808 20788
rect 35115 20757 35127 20760
rect 35069 20751 35127 20757
rect 35802 20748 35808 20760
rect 35860 20748 35866 20800
rect 36078 20748 36084 20800
rect 36136 20748 36142 20800
rect 36170 20748 36176 20800
rect 36228 20748 36234 20800
rect 36446 20748 36452 20800
rect 36504 20788 36510 20800
rect 37090 20788 37096 20800
rect 36504 20760 37096 20788
rect 36504 20748 36510 20760
rect 37090 20748 37096 20760
rect 37148 20788 37154 20800
rect 38473 20791 38531 20797
rect 38473 20788 38485 20791
rect 37148 20760 38485 20788
rect 37148 20748 37154 20760
rect 38473 20757 38485 20760
rect 38519 20757 38531 20791
rect 38473 20751 38531 20757
rect 39206 20748 39212 20800
rect 39264 20748 39270 20800
rect 40957 20791 41015 20797
rect 40957 20757 40969 20791
rect 41003 20788 41015 20791
rect 41003 20760 41552 20788
rect 41003 20757 41015 20760
rect 40957 20751 41015 20757
rect 41524 20732 41552 20760
rect 1104 20698 41400 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 41400 20698
rect 41506 20680 41512 20732
rect 41564 20680 41570 20732
rect 1104 20624 41400 20646
rect 12710 20584 12716 20596
rect 12406 20556 12716 20584
rect 5077 20519 5135 20525
rect 5077 20485 5089 20519
rect 5123 20516 5135 20519
rect 12406 20516 12434 20556
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 12820 20556 13584 20584
rect 5123 20488 12434 20516
rect 5123 20485 5135 20488
rect 5077 20479 5135 20485
rect 5552 20457 5580 20488
rect 4893 20451 4951 20457
rect 4893 20417 4905 20451
rect 4939 20448 4951 20451
rect 5353 20451 5411 20457
rect 5353 20448 5365 20451
rect 4939 20420 5365 20448
rect 4939 20417 4951 20420
rect 4893 20411 4951 20417
rect 5353 20417 5365 20420
rect 5399 20417 5411 20451
rect 5353 20411 5411 20417
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 5368 20380 5396 20411
rect 8570 20408 8576 20460
rect 8628 20408 8634 20460
rect 12158 20408 12164 20460
rect 12216 20408 12222 20460
rect 12250 20408 12256 20460
rect 12308 20408 12314 20460
rect 12345 20451 12403 20457
rect 12345 20417 12357 20451
rect 12391 20448 12403 20451
rect 12526 20448 12532 20460
rect 12391 20420 12532 20448
rect 12391 20417 12403 20420
rect 12345 20411 12403 20417
rect 12526 20408 12532 20420
rect 12584 20408 12590 20460
rect 12618 20408 12624 20460
rect 12676 20448 12682 20460
rect 12713 20451 12771 20457
rect 12713 20448 12725 20451
rect 12676 20420 12725 20448
rect 12676 20408 12682 20420
rect 12713 20417 12725 20420
rect 12759 20448 12771 20451
rect 12820 20448 12848 20556
rect 12986 20476 12992 20528
rect 13044 20516 13050 20528
rect 13044 20488 13492 20516
rect 13044 20476 13050 20488
rect 12759 20420 12848 20448
rect 12759 20417 12771 20420
rect 12713 20411 12771 20417
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 13464 20457 13492 20488
rect 13556 20460 13584 20556
rect 15010 20544 15016 20596
rect 15068 20544 15074 20596
rect 15930 20544 15936 20596
rect 15988 20584 15994 20596
rect 19429 20587 19487 20593
rect 15988 20556 19334 20584
rect 15988 20544 15994 20556
rect 14645 20519 14703 20525
rect 14645 20485 14657 20519
rect 14691 20516 14703 20519
rect 17129 20519 17187 20525
rect 14691 20488 15056 20516
rect 14691 20485 14703 20488
rect 14645 20479 14703 20485
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 12952 20420 13277 20448
rect 12952 20408 12958 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 14737 20451 14795 20457
rect 14737 20417 14749 20451
rect 14783 20448 14795 20451
rect 14826 20448 14832 20460
rect 14783 20420 14832 20448
rect 14783 20417 14795 20420
rect 14737 20411 14795 20417
rect 8588 20380 8616 20408
rect 5368 20352 8616 20380
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12636 20380 12664 20408
rect 12483 20352 12664 20380
rect 14476 20380 14504 20411
rect 14826 20408 14832 20420
rect 14884 20408 14890 20460
rect 15028 20457 15056 20488
rect 15856 20488 16620 20516
rect 15856 20460 15884 20488
rect 15013 20451 15071 20457
rect 15013 20417 15025 20451
rect 15059 20448 15071 20451
rect 15746 20448 15752 20460
rect 15059 20420 15752 20448
rect 15059 20417 15071 20420
rect 15013 20411 15071 20417
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 15838 20408 15844 20460
rect 15896 20408 15902 20460
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 16482 20448 16488 20460
rect 16163 20420 16488 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 15381 20383 15439 20389
rect 15381 20380 15393 20383
rect 14476 20352 15393 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 15381 20349 15393 20352
rect 15427 20349 15439 20383
rect 15381 20343 15439 20349
rect 4890 20272 4896 20324
rect 4948 20312 4954 20324
rect 5353 20315 5411 20321
rect 5353 20312 5365 20315
rect 4948 20284 5365 20312
rect 4948 20272 4954 20284
rect 5353 20281 5365 20284
rect 5399 20281 5411 20315
rect 5353 20275 5411 20281
rect 11977 20315 12035 20321
rect 11977 20281 11989 20315
rect 12023 20312 12035 20315
rect 14182 20312 14188 20324
rect 12023 20284 14188 20312
rect 12023 20281 12035 20284
rect 11977 20275 12035 20281
rect 14182 20272 14188 20284
rect 14240 20272 14246 20324
rect 15396 20312 15424 20343
rect 16206 20340 16212 20392
rect 16264 20340 16270 20392
rect 16298 20340 16304 20392
rect 16356 20340 16362 20392
rect 16393 20383 16451 20389
rect 16393 20349 16405 20383
rect 16439 20380 16451 20383
rect 16592 20380 16620 20488
rect 17129 20485 17141 20519
rect 17175 20516 17187 20519
rect 17402 20516 17408 20528
rect 17175 20488 17408 20516
rect 17175 20485 17187 20488
rect 17129 20479 17187 20485
rect 17402 20476 17408 20488
rect 17460 20476 17466 20528
rect 19306 20516 19334 20556
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 20438 20584 20444 20596
rect 19475 20556 20444 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 21910 20584 21916 20596
rect 20772 20556 21916 20584
rect 20772 20544 20778 20556
rect 21910 20544 21916 20556
rect 21968 20584 21974 20596
rect 22189 20587 22247 20593
rect 22189 20584 22201 20587
rect 21968 20556 22201 20584
rect 21968 20544 21974 20556
rect 22189 20553 22201 20556
rect 22235 20553 22247 20587
rect 22649 20587 22707 20593
rect 22649 20584 22661 20587
rect 22189 20547 22247 20553
rect 22296 20556 22661 20584
rect 17604 20488 19196 20516
rect 19306 20488 20392 20516
rect 16942 20408 16948 20460
rect 17000 20408 17006 20460
rect 17218 20408 17224 20460
rect 17276 20408 17282 20460
rect 17310 20408 17316 20460
rect 17368 20448 17374 20460
rect 17604 20448 17632 20488
rect 17368 20420 17632 20448
rect 17681 20451 17739 20457
rect 17368 20408 17374 20420
rect 17681 20417 17693 20451
rect 17727 20448 17739 20451
rect 17770 20448 17776 20460
rect 17727 20420 17776 20448
rect 17727 20417 17739 20420
rect 17681 20411 17739 20417
rect 17696 20380 17724 20411
rect 17770 20408 17776 20420
rect 17828 20448 17834 20460
rect 18966 20448 18972 20460
rect 17828 20420 18972 20448
rect 17828 20408 17834 20420
rect 18966 20408 18972 20420
rect 19024 20408 19030 20460
rect 19058 20408 19064 20460
rect 19116 20408 19122 20460
rect 16439 20352 16620 20380
rect 16684 20352 17724 20380
rect 16439 20349 16451 20352
rect 16393 20343 16451 20349
rect 16684 20312 16712 20352
rect 17954 20340 17960 20392
rect 18012 20340 18018 20392
rect 19168 20380 19196 20488
rect 19352 20457 19380 20488
rect 19337 20451 19395 20457
rect 19337 20417 19349 20451
rect 19383 20448 19395 20451
rect 19383 20420 19417 20448
rect 19383 20417 19395 20420
rect 19337 20411 19395 20417
rect 19518 20408 19524 20460
rect 19576 20408 19582 20460
rect 20364 20457 20392 20488
rect 20990 20476 20996 20528
rect 21048 20516 21054 20528
rect 21818 20516 21824 20528
rect 21048 20488 21824 20516
rect 21048 20476 21054 20488
rect 21818 20476 21824 20488
rect 21876 20476 21882 20528
rect 22097 20519 22155 20525
rect 22097 20516 22109 20519
rect 21928 20488 22109 20516
rect 19797 20451 19855 20457
rect 19628 20448 19748 20451
rect 19797 20448 19809 20451
rect 19628 20423 19809 20448
rect 19628 20380 19656 20423
rect 19720 20420 19809 20423
rect 19797 20417 19809 20420
rect 19843 20448 19855 20451
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 19843 20420 20177 20448
rect 19843 20417 19855 20420
rect 19797 20411 19855 20417
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20417 20315 20451
rect 20257 20411 20315 20417
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20622 20448 20628 20460
rect 20579 20420 20628 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 19168 20352 19656 20380
rect 19705 20383 19763 20389
rect 19705 20349 19717 20383
rect 19751 20380 19763 20383
rect 19978 20380 19984 20392
rect 19751 20352 19984 20380
rect 19751 20349 19763 20352
rect 19705 20343 19763 20349
rect 19978 20340 19984 20352
rect 20036 20380 20042 20392
rect 20272 20380 20300 20411
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 21358 20408 21364 20460
rect 21416 20408 21422 20460
rect 21726 20408 21732 20460
rect 21784 20448 21790 20460
rect 21928 20448 21956 20488
rect 22097 20485 22109 20488
rect 22143 20516 22155 20519
rect 22296 20516 22324 20556
rect 22649 20553 22661 20556
rect 22695 20553 22707 20587
rect 22649 20547 22707 20553
rect 25222 20544 25228 20596
rect 25280 20584 25286 20596
rect 25961 20587 26019 20593
rect 25961 20584 25973 20587
rect 25280 20556 25973 20584
rect 25280 20544 25286 20556
rect 25961 20553 25973 20556
rect 26007 20553 26019 20587
rect 25961 20547 26019 20553
rect 26142 20544 26148 20596
rect 26200 20544 26206 20596
rect 32398 20544 32404 20596
rect 32456 20544 32462 20596
rect 32490 20544 32496 20596
rect 32548 20584 32554 20596
rect 32769 20587 32827 20593
rect 32769 20584 32781 20587
rect 32548 20556 32781 20584
rect 32548 20544 32554 20556
rect 32769 20553 32781 20556
rect 32815 20553 32827 20587
rect 32769 20547 32827 20553
rect 35342 20544 35348 20596
rect 35400 20584 35406 20596
rect 35618 20584 35624 20596
rect 35400 20556 35624 20584
rect 35400 20544 35406 20556
rect 35618 20544 35624 20556
rect 35676 20544 35682 20596
rect 36173 20587 36231 20593
rect 36173 20553 36185 20587
rect 36219 20584 36231 20587
rect 38838 20584 38844 20596
rect 36219 20556 38844 20584
rect 36219 20553 36231 20556
rect 36173 20547 36231 20553
rect 38838 20544 38844 20556
rect 38896 20544 38902 20596
rect 39040 20556 40448 20584
rect 22143 20488 22324 20516
rect 22465 20519 22523 20525
rect 22143 20485 22155 20488
rect 22097 20479 22155 20485
rect 22465 20485 22477 20519
rect 22511 20516 22523 20519
rect 22554 20516 22560 20528
rect 22511 20488 22560 20516
rect 22511 20485 22523 20488
rect 22465 20479 22523 20485
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 25038 20476 25044 20528
rect 25096 20516 25102 20528
rect 25133 20519 25191 20525
rect 25133 20516 25145 20519
rect 25096 20488 25145 20516
rect 25096 20476 25102 20488
rect 25133 20485 25145 20488
rect 25179 20485 25191 20519
rect 27154 20516 27160 20528
rect 25133 20479 25191 20485
rect 25240 20488 25452 20516
rect 21784 20420 21956 20448
rect 22005 20451 22063 20457
rect 21784 20408 21790 20420
rect 22005 20417 22017 20451
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20448 22431 20451
rect 23017 20451 23075 20457
rect 23017 20448 23029 20451
rect 22419 20420 23029 20448
rect 22419 20417 22431 20420
rect 22373 20411 22431 20417
rect 23017 20417 23029 20420
rect 23063 20417 23075 20451
rect 25240 20448 25268 20488
rect 23017 20411 23075 20417
rect 25148 20420 25268 20448
rect 25424 20448 25452 20488
rect 26528 20488 27160 20516
rect 26528 20457 26556 20488
rect 27154 20476 27160 20488
rect 27212 20476 27218 20528
rect 28534 20476 28540 20528
rect 28592 20476 28598 20528
rect 30282 20476 30288 20528
rect 30340 20476 30346 20528
rect 32416 20516 32444 20544
rect 32416 20488 32628 20516
rect 26086 20451 26144 20457
rect 26086 20448 26098 20451
rect 25424 20420 26098 20448
rect 20036 20352 20300 20380
rect 22020 20380 22048 20411
rect 25148 20392 25176 20420
rect 26086 20417 26098 20420
rect 26132 20417 26144 20451
rect 26086 20411 26144 20417
rect 26513 20451 26571 20457
rect 26513 20417 26525 20451
rect 26559 20417 26571 20451
rect 26513 20411 26571 20417
rect 26786 20408 26792 20460
rect 26844 20448 26850 20460
rect 28261 20451 28319 20457
rect 28261 20448 28273 20451
rect 26844 20420 28273 20448
rect 26844 20408 26850 20420
rect 28261 20417 28273 20420
rect 28307 20417 28319 20451
rect 29670 20434 30880 20448
rect 28261 20411 28319 20417
rect 29656 20420 30880 20434
rect 22094 20380 22100 20392
rect 22020 20352 22100 20380
rect 20036 20340 20042 20352
rect 22094 20340 22100 20352
rect 22152 20380 22158 20392
rect 22646 20380 22652 20392
rect 22152 20352 22652 20380
rect 22152 20340 22158 20352
rect 22646 20340 22652 20352
rect 22704 20340 22710 20392
rect 25130 20340 25136 20392
rect 25188 20340 25194 20392
rect 26605 20383 26663 20389
rect 26605 20380 26617 20383
rect 25337 20352 26617 20380
rect 15396 20284 16712 20312
rect 17678 20272 17684 20324
rect 17736 20312 17742 20324
rect 19610 20312 19616 20324
rect 17736 20284 19616 20312
rect 17736 20272 17742 20284
rect 19610 20272 19616 20284
rect 19668 20272 19674 20324
rect 5258 20204 5264 20256
rect 5316 20204 5322 20256
rect 13262 20204 13268 20256
rect 13320 20204 13326 20256
rect 14274 20204 14280 20256
rect 14332 20204 14338 20256
rect 15930 20204 15936 20256
rect 15988 20204 15994 20256
rect 16761 20247 16819 20253
rect 16761 20213 16773 20247
rect 16807 20244 16819 20247
rect 16850 20244 16856 20256
rect 16807 20216 16856 20244
rect 16807 20213 16819 20216
rect 16761 20207 16819 20213
rect 16850 20204 16856 20216
rect 16908 20244 16914 20256
rect 19150 20244 19156 20256
rect 16908 20216 19156 20244
rect 16908 20204 16914 20216
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 19794 20244 19800 20256
rect 19392 20216 19800 20244
rect 19392 20204 19398 20216
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 19889 20247 19947 20253
rect 19889 20213 19901 20247
rect 19935 20244 19947 20247
rect 20990 20244 20996 20256
rect 19935 20216 20996 20244
rect 19935 20213 19947 20216
rect 19889 20207 19947 20213
rect 20990 20204 20996 20216
rect 21048 20204 21054 20256
rect 22646 20204 22652 20256
rect 22704 20204 22710 20256
rect 22830 20204 22836 20256
rect 22888 20204 22894 20256
rect 23201 20247 23259 20253
rect 23201 20213 23213 20247
rect 23247 20244 23259 20247
rect 23750 20244 23756 20256
rect 23247 20216 23756 20244
rect 23247 20213 23259 20216
rect 23201 20207 23259 20213
rect 23750 20204 23756 20216
rect 23808 20204 23814 20256
rect 24946 20204 24952 20256
rect 25004 20244 25010 20256
rect 25337 20244 25365 20352
rect 26605 20349 26617 20352
rect 26651 20349 26663 20383
rect 26605 20343 26663 20349
rect 28534 20340 28540 20392
rect 28592 20380 28598 20392
rect 29656 20380 29684 20420
rect 28592 20352 29684 20380
rect 28592 20340 28598 20352
rect 30852 20256 30880 20420
rect 32122 20408 32128 20460
rect 32180 20408 32186 20460
rect 32214 20408 32220 20460
rect 32272 20448 32278 20460
rect 32401 20451 32459 20457
rect 32272 20420 32317 20448
rect 32272 20408 32278 20420
rect 32401 20417 32413 20451
rect 32447 20417 32459 20451
rect 32401 20411 32459 20417
rect 25004 20216 25365 20244
rect 25004 20204 25010 20216
rect 25406 20204 25412 20256
rect 25464 20204 25470 20256
rect 26602 20204 26608 20256
rect 26660 20244 26666 20256
rect 27154 20244 27160 20256
rect 26660 20216 27160 20244
rect 26660 20204 26666 20216
rect 27154 20204 27160 20216
rect 27212 20204 27218 20256
rect 30834 20204 30840 20256
rect 30892 20244 30898 20256
rect 31754 20244 31760 20256
rect 30892 20216 31760 20244
rect 30892 20204 30898 20216
rect 31754 20204 31760 20216
rect 31812 20204 31818 20256
rect 32416 20244 32444 20411
rect 32490 20408 32496 20460
rect 32548 20408 32554 20460
rect 32600 20457 32628 20488
rect 33134 20476 33140 20528
rect 33192 20516 33198 20528
rect 39040 20516 39068 20556
rect 33192 20488 34086 20516
rect 35912 20488 36860 20516
rect 33192 20476 33198 20488
rect 35912 20460 35940 20488
rect 32590 20451 32648 20457
rect 32590 20417 32602 20451
rect 32636 20417 32648 20451
rect 32590 20411 32648 20417
rect 32766 20408 32772 20460
rect 32824 20448 32830 20460
rect 33321 20451 33379 20457
rect 33321 20448 33333 20451
rect 32824 20420 33333 20448
rect 32824 20408 32830 20420
rect 33321 20417 33333 20420
rect 33367 20417 33379 20451
rect 33321 20411 33379 20417
rect 35894 20408 35900 20460
rect 35952 20408 35958 20460
rect 36170 20408 36176 20460
rect 36228 20448 36234 20460
rect 36357 20451 36415 20457
rect 36357 20448 36369 20451
rect 36228 20420 36369 20448
rect 36228 20408 36234 20420
rect 36357 20417 36369 20420
rect 36403 20417 36415 20451
rect 36357 20411 36415 20417
rect 36449 20451 36507 20457
rect 36449 20417 36461 20451
rect 36495 20417 36507 20451
rect 36449 20411 36507 20417
rect 33594 20340 33600 20392
rect 33652 20340 33658 20392
rect 35342 20340 35348 20392
rect 35400 20380 35406 20392
rect 35437 20383 35495 20389
rect 35437 20380 35449 20383
rect 35400 20352 35449 20380
rect 35400 20340 35406 20352
rect 35437 20349 35449 20352
rect 35483 20380 35495 20383
rect 35526 20380 35532 20392
rect 35483 20352 35532 20380
rect 35483 20349 35495 20352
rect 35437 20343 35495 20349
rect 35526 20340 35532 20352
rect 35584 20340 35590 20392
rect 36464 20380 36492 20411
rect 36538 20408 36544 20460
rect 36596 20408 36602 20460
rect 36722 20408 36728 20460
rect 36780 20408 36786 20460
rect 36832 20457 36860 20488
rect 37384 20488 39068 20516
rect 37384 20460 37412 20488
rect 36817 20451 36875 20457
rect 36817 20417 36829 20451
rect 36863 20448 36875 20451
rect 37277 20451 37335 20457
rect 37277 20448 37289 20451
rect 36863 20420 37289 20448
rect 36863 20417 36875 20420
rect 36817 20411 36875 20417
rect 37277 20417 37289 20420
rect 37323 20417 37335 20451
rect 37277 20411 37335 20417
rect 37366 20408 37372 20460
rect 37424 20408 37430 20460
rect 37936 20457 37964 20488
rect 39114 20476 39120 20528
rect 39172 20476 39178 20528
rect 40420 20525 40448 20556
rect 40405 20519 40463 20525
rect 40405 20485 40417 20519
rect 40451 20485 40463 20519
rect 40405 20479 40463 20485
rect 37461 20451 37519 20457
rect 37461 20417 37473 20451
rect 37507 20417 37519 20451
rect 37461 20411 37519 20417
rect 37553 20451 37611 20457
rect 37553 20417 37565 20451
rect 37599 20417 37611 20451
rect 37553 20411 37611 20417
rect 37921 20451 37979 20457
rect 37921 20417 37933 20451
rect 37967 20417 37979 20451
rect 37921 20411 37979 20417
rect 36372 20352 36492 20380
rect 36556 20380 36584 20408
rect 37476 20380 37504 20411
rect 36556 20352 37504 20380
rect 34698 20272 34704 20324
rect 34756 20312 34762 20324
rect 36372 20312 36400 20352
rect 34756 20284 36400 20312
rect 34756 20272 34762 20284
rect 33962 20244 33968 20256
rect 32416 20216 33968 20244
rect 33962 20204 33968 20216
rect 34020 20204 34026 20256
rect 34606 20204 34612 20256
rect 34664 20244 34670 20256
rect 36081 20247 36139 20253
rect 36081 20244 36093 20247
rect 34664 20216 36093 20244
rect 34664 20204 34670 20216
rect 36081 20213 36093 20216
rect 36127 20213 36139 20247
rect 36372 20244 36400 20284
rect 37274 20272 37280 20324
rect 37332 20272 37338 20324
rect 37568 20244 37596 20411
rect 37826 20340 37832 20392
rect 37884 20340 37890 20392
rect 38378 20340 38384 20392
rect 38436 20340 38442 20392
rect 38654 20340 38660 20392
rect 38712 20340 38718 20392
rect 36372 20216 37596 20244
rect 38289 20247 38347 20253
rect 36081 20207 36139 20213
rect 38289 20213 38301 20247
rect 38335 20244 38347 20247
rect 39022 20244 39028 20256
rect 38335 20216 39028 20244
rect 38335 20213 38347 20216
rect 38289 20207 38347 20213
rect 39022 20204 39028 20216
rect 39080 20204 39086 20256
rect 1104 20154 41400 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 41400 20154
rect 1104 20080 41400 20102
rect 6638 20000 6644 20052
rect 6696 20000 6702 20052
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 12069 20043 12127 20049
rect 12069 20040 12081 20043
rect 11379 20012 12081 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 12069 20009 12081 20012
rect 12115 20040 12127 20043
rect 13078 20040 13084 20052
rect 12115 20012 13084 20040
rect 12115 20009 12127 20012
rect 12069 20003 12127 20009
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13262 20000 13268 20052
rect 13320 20000 13326 20052
rect 13538 20000 13544 20052
rect 13596 20040 13602 20052
rect 13596 20012 14044 20040
rect 13596 20000 13602 20012
rect 7190 19972 7196 19984
rect 6564 19944 7196 19972
rect 6564 19848 6592 19944
rect 7190 19932 7196 19944
rect 7248 19932 7254 19984
rect 9582 19932 9588 19984
rect 9640 19972 9646 19984
rect 10042 19972 10048 19984
rect 9640 19944 10048 19972
rect 9640 19932 9646 19944
rect 10042 19932 10048 19944
rect 10100 19972 10106 19984
rect 10318 19972 10324 19984
rect 10100 19944 10324 19972
rect 10100 19932 10106 19944
rect 10318 19932 10324 19944
rect 10376 19932 10382 19984
rect 11606 19932 11612 19984
rect 11664 19932 11670 19984
rect 6914 19864 6920 19916
rect 6972 19904 6978 19916
rect 7101 19907 7159 19913
rect 7101 19904 7113 19907
rect 6972 19876 7113 19904
rect 6972 19864 6978 19876
rect 7101 19873 7113 19876
rect 7147 19904 7159 19907
rect 7837 19907 7895 19913
rect 7837 19904 7849 19907
rect 7147 19876 7849 19904
rect 7147 19873 7159 19876
rect 7101 19867 7159 19873
rect 7837 19873 7849 19876
rect 7883 19873 7895 19907
rect 10594 19904 10600 19916
rect 7837 19867 7895 19873
rect 10336 19876 10600 19904
rect 10336 19848 10364 19876
rect 10594 19864 10600 19876
rect 10652 19904 10658 19916
rect 11624 19904 11652 19932
rect 10652 19876 11652 19904
rect 10652 19864 10658 19876
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19836 4491 19839
rect 4798 19836 4804 19848
rect 4479 19808 4804 19836
rect 4479 19805 4491 19808
rect 4433 19799 4491 19805
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19836 4951 19839
rect 5166 19836 5172 19848
rect 4939 19808 5172 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 6546 19796 6552 19848
rect 6604 19796 6610 19848
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19805 6791 19839
rect 6733 19799 6791 19805
rect 934 19728 940 19780
rect 992 19768 998 19780
rect 1489 19771 1547 19777
rect 1489 19768 1501 19771
rect 992 19740 1501 19768
rect 992 19728 998 19740
rect 1489 19737 1501 19740
rect 1535 19737 1547 19771
rect 1489 19731 1547 19737
rect 1670 19728 1676 19780
rect 1728 19728 1734 19780
rect 6748 19768 6776 19799
rect 6822 19796 6828 19848
rect 6880 19836 6886 19848
rect 7009 19839 7067 19845
rect 7009 19836 7021 19839
rect 6880 19808 7021 19836
rect 6880 19796 6886 19808
rect 7009 19805 7021 19808
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7190 19796 7196 19848
rect 7248 19796 7254 19848
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7374 19836 7380 19848
rect 7331 19808 7380 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 7469 19839 7527 19845
rect 7469 19805 7481 19839
rect 7515 19836 7527 19839
rect 7515 19808 8248 19836
rect 7515 19805 7527 19808
rect 7469 19799 7527 19805
rect 8220 19780 8248 19808
rect 10318 19796 10324 19848
rect 10376 19796 10382 19848
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19836 10563 19839
rect 12529 19839 12587 19845
rect 10551 19808 11376 19836
rect 10551 19805 10563 19808
rect 10505 19799 10563 19805
rect 7653 19771 7711 19777
rect 6748 19740 7236 19768
rect 7208 19712 7236 19740
rect 7653 19737 7665 19771
rect 7699 19737 7711 19771
rect 7653 19731 7711 19737
rect 4706 19660 4712 19712
rect 4764 19660 4770 19712
rect 4801 19703 4859 19709
rect 4801 19669 4813 19703
rect 4847 19700 4859 19703
rect 4982 19700 4988 19712
rect 4847 19672 4988 19700
rect 4847 19669 4859 19672
rect 4801 19663 4859 19669
rect 4982 19660 4988 19672
rect 5040 19660 5046 19712
rect 6822 19660 6828 19712
rect 6880 19660 6886 19712
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 7668 19700 7696 19731
rect 8202 19728 8208 19780
rect 8260 19728 8266 19780
rect 8938 19728 8944 19780
rect 8996 19768 9002 19780
rect 11149 19771 11207 19777
rect 8996 19740 10548 19768
rect 8996 19728 9002 19740
rect 7248 19672 7696 19700
rect 7248 19660 7254 19672
rect 9398 19660 9404 19712
rect 9456 19700 9462 19712
rect 10413 19703 10471 19709
rect 10413 19700 10425 19703
rect 9456 19672 10425 19700
rect 9456 19660 9462 19672
rect 10413 19669 10425 19672
rect 10459 19669 10471 19703
rect 10520 19700 10548 19740
rect 11149 19737 11161 19771
rect 11195 19768 11207 19771
rect 11238 19768 11244 19780
rect 11195 19740 11244 19768
rect 11195 19737 11207 19740
rect 11149 19731 11207 19737
rect 11238 19728 11244 19740
rect 11296 19728 11302 19780
rect 11348 19777 11376 19808
rect 12529 19805 12541 19839
rect 12575 19836 12587 19839
rect 12618 19836 12624 19848
rect 12575 19808 12624 19836
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 12802 19796 12808 19848
rect 12860 19796 12866 19848
rect 12894 19796 12900 19848
rect 12952 19796 12958 19848
rect 13280 19836 13308 20000
rect 13633 19975 13691 19981
rect 13633 19941 13645 19975
rect 13679 19972 13691 19975
rect 13906 19972 13912 19984
rect 13679 19944 13912 19972
rect 13679 19941 13691 19944
rect 13633 19935 13691 19941
rect 13906 19932 13912 19944
rect 13964 19932 13970 19984
rect 14016 19972 14044 20012
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16393 20043 16451 20049
rect 16393 20040 16405 20043
rect 16172 20012 16405 20040
rect 16172 20000 16178 20012
rect 16393 20009 16405 20012
rect 16439 20009 16451 20043
rect 16393 20003 16451 20009
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 16666 20040 16672 20052
rect 16531 20012 16672 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 16850 20000 16856 20052
rect 16908 20000 16914 20052
rect 16960 20012 17724 20040
rect 16868 19972 16896 20000
rect 14016 19944 16896 19972
rect 16960 19916 16988 20012
rect 17144 19944 17448 19972
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13648 19876 14105 19904
rect 13648 19845 13676 19876
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 14274 19864 14280 19916
rect 14332 19864 14338 19916
rect 14921 19907 14979 19913
rect 14921 19904 14933 19907
rect 14384 19876 14933 19904
rect 13633 19839 13691 19845
rect 13633 19836 13645 19839
rect 13280 19808 13645 19836
rect 13633 19805 13645 19808
rect 13679 19805 13691 19839
rect 13633 19799 13691 19805
rect 13814 19796 13820 19848
rect 13872 19796 13878 19848
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 13998 19836 14004 19848
rect 13955 19808 14004 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 13998 19796 14004 19808
rect 14056 19836 14062 19848
rect 14384 19836 14412 19876
rect 14921 19873 14933 19876
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 16114 19864 16120 19916
rect 16172 19904 16178 19916
rect 16942 19904 16948 19916
rect 16172 19876 16948 19904
rect 16172 19864 16178 19876
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 14056 19808 14412 19836
rect 14553 19839 14611 19845
rect 14056 19796 14062 19808
rect 14553 19805 14565 19839
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 11333 19771 11391 19777
rect 11333 19737 11345 19771
rect 11379 19768 11391 19771
rect 11422 19768 11428 19780
rect 11379 19740 11428 19768
rect 11379 19737 11391 19740
rect 11333 19731 11391 19737
rect 11422 19728 11428 19740
rect 11480 19728 11486 19780
rect 11790 19728 11796 19780
rect 11848 19728 11854 19780
rect 12345 19771 12403 19777
rect 12345 19737 12357 19771
rect 12391 19768 12403 19771
rect 12713 19771 12771 19777
rect 12391 19740 12664 19768
rect 12391 19737 12403 19740
rect 12345 19731 12403 19737
rect 11517 19703 11575 19709
rect 11517 19700 11529 19703
rect 10520 19672 11529 19700
rect 10413 19663 10471 19669
rect 11517 19669 11529 19672
rect 11563 19669 11575 19703
rect 12636 19700 12664 19740
rect 12713 19737 12725 19771
rect 12759 19768 12771 19771
rect 12912 19768 12940 19796
rect 12759 19740 12940 19768
rect 13832 19768 13860 19796
rect 14568 19768 14596 19799
rect 16574 19796 16580 19848
rect 16632 19796 16638 19848
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19836 16727 19839
rect 17144 19836 17172 19944
rect 17218 19864 17224 19916
rect 17276 19864 17282 19916
rect 17420 19904 17448 19944
rect 17420 19876 17632 19904
rect 16715 19808 17172 19836
rect 16715 19805 16727 19808
rect 16669 19799 16727 19805
rect 13832 19740 14596 19768
rect 12759 19737 12771 19740
rect 12713 19731 12771 19737
rect 16206 19728 16212 19780
rect 16264 19728 16270 19780
rect 16761 19771 16819 19777
rect 16761 19737 16773 19771
rect 16807 19768 16819 19771
rect 17236 19768 17264 19864
rect 17420 19848 17448 19876
rect 17402 19796 17408 19848
rect 17460 19796 17466 19848
rect 17604 19845 17632 19876
rect 17497 19839 17555 19845
rect 17497 19805 17509 19839
rect 17543 19805 17555 19839
rect 17497 19799 17555 19805
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19805 17647 19839
rect 17696 19836 17724 20012
rect 19058 20000 19064 20052
rect 19116 20000 19122 20052
rect 19150 20000 19156 20052
rect 19208 20040 19214 20052
rect 21177 20043 21235 20049
rect 19208 20012 21128 20040
rect 19208 20000 19214 20012
rect 19076 19972 19104 20000
rect 21100 19972 21128 20012
rect 21177 20009 21189 20043
rect 21223 20040 21235 20043
rect 22278 20040 22284 20052
rect 21223 20012 22284 20040
rect 21223 20009 21235 20012
rect 21177 20003 21235 20009
rect 22278 20000 22284 20012
rect 22336 20040 22342 20052
rect 23661 20043 23719 20049
rect 23661 20040 23673 20043
rect 22336 20012 23673 20040
rect 22336 20000 22342 20012
rect 23661 20009 23673 20012
rect 23707 20009 23719 20043
rect 23661 20003 23719 20009
rect 23842 20000 23848 20052
rect 23900 20040 23906 20052
rect 25363 20043 25421 20049
rect 25363 20040 25375 20043
rect 23900 20012 25375 20040
rect 23900 20000 23906 20012
rect 25363 20009 25375 20012
rect 25409 20040 25421 20043
rect 25498 20040 25504 20052
rect 25409 20012 25504 20040
rect 25409 20009 25421 20012
rect 25363 20003 25421 20009
rect 25498 20000 25504 20012
rect 25556 20000 25562 20052
rect 27246 20000 27252 20052
rect 27304 20040 27310 20052
rect 27522 20040 27528 20052
rect 27304 20012 27528 20040
rect 27304 20000 27310 20012
rect 27522 20000 27528 20012
rect 27580 20000 27586 20052
rect 31478 20000 31484 20052
rect 31536 20000 31542 20052
rect 31754 20000 31760 20052
rect 31812 20040 31818 20052
rect 33134 20040 33140 20052
rect 31812 20012 33140 20040
rect 31812 20000 31818 20012
rect 33134 20000 33140 20012
rect 33192 20000 33198 20052
rect 33594 20000 33600 20052
rect 33652 20040 33658 20052
rect 34149 20043 34207 20049
rect 34149 20040 34161 20043
rect 33652 20012 34161 20040
rect 33652 20000 33658 20012
rect 34149 20009 34161 20012
rect 34195 20009 34207 20043
rect 34149 20003 34207 20009
rect 34698 20000 34704 20052
rect 34756 20040 34762 20052
rect 34974 20040 34980 20052
rect 34756 20012 34980 20040
rect 34756 20000 34762 20012
rect 34974 20000 34980 20012
rect 35032 20000 35038 20052
rect 35713 20043 35771 20049
rect 35713 20009 35725 20043
rect 35759 20040 35771 20043
rect 35894 20040 35900 20052
rect 35759 20012 35900 20040
rect 35759 20009 35771 20012
rect 35713 20003 35771 20009
rect 35894 20000 35900 20012
rect 35952 20000 35958 20052
rect 36170 20000 36176 20052
rect 36228 20000 36234 20052
rect 36633 20043 36691 20049
rect 36633 20009 36645 20043
rect 36679 20040 36691 20043
rect 36722 20040 36728 20052
rect 36679 20012 36728 20040
rect 36679 20009 36691 20012
rect 36633 20003 36691 20009
rect 36722 20000 36728 20012
rect 36780 20000 36786 20052
rect 38289 20043 38347 20049
rect 38289 20009 38301 20043
rect 38335 20040 38347 20043
rect 38654 20040 38660 20052
rect 38335 20012 38660 20040
rect 38335 20009 38347 20012
rect 38289 20003 38347 20009
rect 38654 20000 38660 20012
rect 38712 20000 38718 20052
rect 19076 19944 21036 19972
rect 21100 19944 22094 19972
rect 18322 19904 18328 19916
rect 18156 19876 18328 19904
rect 17773 19839 17831 19845
rect 17773 19836 17785 19839
rect 17696 19808 17785 19836
rect 17589 19799 17647 19805
rect 17773 19805 17785 19808
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 17512 19768 17540 19799
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 18156 19845 18184 19876
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 18966 19864 18972 19916
rect 19024 19904 19030 19916
rect 19024 19876 19385 19904
rect 19024 19864 19030 19876
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 17678 19768 17684 19780
rect 16807 19740 17684 19768
rect 16807 19737 16819 19740
rect 16761 19731 16819 19737
rect 17678 19728 17684 19740
rect 17736 19728 17742 19780
rect 19357 19768 19385 19876
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 19484 19876 19625 19904
rect 19484 19864 19490 19876
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 19613 19867 19671 19873
rect 19705 19907 19763 19913
rect 19705 19873 19717 19907
rect 19751 19904 19763 19907
rect 20162 19904 20168 19916
rect 19751 19876 20168 19904
rect 19751 19873 19763 19876
rect 19705 19867 19763 19873
rect 20162 19864 20168 19876
rect 20220 19904 20226 19916
rect 20530 19904 20536 19916
rect 20220 19876 20536 19904
rect 20220 19864 20226 19876
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 21008 19913 21036 19944
rect 20993 19907 21051 19913
rect 20993 19873 21005 19907
rect 21039 19873 21051 19907
rect 20993 19867 21051 19873
rect 19794 19796 19800 19848
rect 19852 19796 19858 19848
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 19904 19768 19932 19799
rect 19978 19796 19984 19848
rect 20036 19796 20042 19848
rect 20070 19796 20076 19848
rect 20128 19796 20134 19848
rect 19357 19740 19932 19768
rect 19996 19768 20024 19796
rect 20254 19768 20260 19780
rect 19996 19740 20260 19768
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 21008 19768 21036 19867
rect 21726 19864 21732 19916
rect 21784 19864 21790 19916
rect 22066 19904 22094 19944
rect 23750 19932 23756 19984
rect 23808 19972 23814 19984
rect 24486 19972 24492 19984
rect 23808 19944 24492 19972
rect 23808 19932 23814 19944
rect 24486 19932 24492 19944
rect 24544 19972 24550 19984
rect 24544 19944 24808 19972
rect 24544 19932 24550 19944
rect 22066 19876 22310 19904
rect 21453 19839 21511 19845
rect 21453 19805 21465 19839
rect 21499 19836 21511 19839
rect 21910 19836 21916 19848
rect 21499 19808 21916 19836
rect 21499 19805 21511 19808
rect 21453 19799 21511 19805
rect 21910 19796 21916 19808
rect 21968 19796 21974 19848
rect 22094 19796 22100 19848
rect 22152 19796 22158 19848
rect 22554 19796 22560 19848
rect 22612 19796 22618 19848
rect 23474 19796 23480 19848
rect 23532 19796 23538 19848
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 23860 19808 24593 19836
rect 22572 19768 22600 19796
rect 23658 19768 23664 19780
rect 21008 19740 22600 19768
rect 23492 19740 23664 19768
rect 14182 19700 14188 19712
rect 12636 19672 14188 19700
rect 11517 19663 11575 19669
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 14366 19660 14372 19712
rect 14424 19660 14430 19712
rect 17313 19703 17371 19709
rect 17313 19669 17325 19703
rect 17359 19700 17371 19703
rect 17770 19700 17776 19712
rect 17359 19672 17776 19700
rect 17359 19669 17371 19672
rect 17313 19663 17371 19669
rect 17770 19660 17776 19672
rect 17828 19660 17834 19712
rect 17954 19660 17960 19712
rect 18012 19660 18018 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 19429 19703 19487 19709
rect 19429 19700 19441 19703
rect 19392 19672 19441 19700
rect 19392 19660 19398 19672
rect 19429 19669 19441 19672
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 20165 19703 20223 19709
rect 20165 19669 20177 19703
rect 20211 19700 20223 19703
rect 20622 19700 20628 19712
rect 20211 19672 20628 19700
rect 20211 19669 20223 19672
rect 20165 19663 20223 19669
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 21358 19660 21364 19712
rect 21416 19660 21422 19712
rect 22554 19660 22560 19712
rect 22612 19700 22618 19712
rect 22659 19703 22717 19709
rect 22659 19700 22671 19703
rect 22612 19672 22671 19700
rect 22612 19660 22618 19672
rect 22659 19669 22671 19672
rect 22705 19700 22717 19703
rect 23492 19700 23520 19740
rect 23658 19728 23664 19740
rect 23716 19768 23722 19780
rect 23860 19777 23888 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24780 19836 24808 19944
rect 25222 19932 25228 19984
rect 25280 19972 25286 19984
rect 32490 19972 32496 19984
rect 25280 19944 25728 19972
rect 25280 19932 25286 19944
rect 24883 19839 24941 19845
rect 24883 19836 24895 19839
rect 24780 19808 24895 19836
rect 24581 19799 24639 19805
rect 24883 19805 24895 19808
rect 24929 19805 24941 19839
rect 24883 19799 24941 19805
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19805 25099 19839
rect 25041 19799 25099 19805
rect 23845 19771 23903 19777
rect 23845 19768 23857 19771
rect 23716 19740 23857 19768
rect 23716 19728 23722 19740
rect 23845 19737 23857 19740
rect 23891 19737 23903 19771
rect 23845 19731 23903 19737
rect 23934 19728 23940 19780
rect 23992 19768 23998 19780
rect 23992 19740 24532 19768
rect 23992 19728 23998 19740
rect 22705 19672 23520 19700
rect 22705 19669 22717 19672
rect 22659 19663 22717 19669
rect 23566 19660 23572 19712
rect 23624 19660 23630 19712
rect 23750 19660 23756 19712
rect 23808 19700 23814 19712
rect 24397 19703 24455 19709
rect 24397 19700 24409 19703
rect 23808 19672 24409 19700
rect 23808 19660 23814 19672
rect 24397 19669 24409 19672
rect 24443 19669 24455 19703
rect 24504 19700 24532 19740
rect 24670 19728 24676 19780
rect 24728 19728 24734 19780
rect 24762 19728 24768 19780
rect 24820 19728 24826 19780
rect 25056 19768 25084 19799
rect 25130 19796 25136 19848
rect 25188 19836 25194 19848
rect 25225 19839 25283 19845
rect 25225 19836 25237 19839
rect 25188 19808 25237 19836
rect 25188 19796 25194 19808
rect 25225 19805 25237 19808
rect 25271 19805 25283 19839
rect 25225 19799 25283 19805
rect 25498 19796 25504 19848
rect 25556 19796 25562 19848
rect 25700 19845 25728 19944
rect 28966 19944 31754 19972
rect 25777 19907 25835 19913
rect 25777 19873 25789 19907
rect 25823 19904 25835 19907
rect 26786 19904 26792 19916
rect 25823 19876 26792 19904
rect 25823 19873 25835 19876
rect 25777 19867 25835 19873
rect 26786 19864 26792 19876
rect 26844 19864 26850 19916
rect 25685 19839 25743 19845
rect 25685 19805 25697 19839
rect 25731 19805 25743 19839
rect 25685 19799 25743 19805
rect 27154 19796 27160 19848
rect 27212 19836 27218 19848
rect 27212 19808 28580 19836
rect 27212 19796 27218 19808
rect 28552 19780 28580 19808
rect 25593 19771 25651 19777
rect 25056 19740 25176 19768
rect 25148 19700 25176 19740
rect 25593 19737 25605 19771
rect 25639 19768 25651 19771
rect 26053 19771 26111 19777
rect 26053 19768 26065 19771
rect 25639 19740 26065 19768
rect 25639 19737 25651 19740
rect 25593 19731 25651 19737
rect 26053 19737 26065 19740
rect 26099 19737 26111 19771
rect 26053 19731 26111 19737
rect 28534 19728 28540 19780
rect 28592 19728 28598 19780
rect 28966 19700 28994 19944
rect 31389 19839 31447 19845
rect 31389 19805 31401 19839
rect 31435 19805 31447 19839
rect 31389 19799 31447 19805
rect 31404 19712 31432 19799
rect 24504 19672 28994 19700
rect 24397 19663 24455 19669
rect 31386 19660 31392 19712
rect 31444 19660 31450 19712
rect 31726 19700 31754 19944
rect 32048 19944 32496 19972
rect 32048 19848 32076 19944
rect 32490 19932 32496 19944
rect 32548 19972 32554 19984
rect 34514 19972 34520 19984
rect 32548 19944 34520 19972
rect 32548 19932 32554 19944
rect 34514 19932 34520 19944
rect 34572 19972 34578 19984
rect 38930 19972 38936 19984
rect 34572 19944 37688 19972
rect 34572 19932 34578 19944
rect 34701 19907 34759 19913
rect 34701 19904 34713 19907
rect 33520 19876 34713 19904
rect 32030 19796 32036 19848
rect 32088 19796 32094 19848
rect 33520 19845 33548 19876
rect 34701 19873 34713 19876
rect 34747 19873 34759 19907
rect 34701 19867 34759 19873
rect 35161 19907 35219 19913
rect 35161 19873 35173 19907
rect 35207 19904 35219 19907
rect 35802 19904 35808 19916
rect 35207 19876 35808 19904
rect 35207 19873 35219 19876
rect 35161 19867 35219 19873
rect 35802 19864 35808 19876
rect 35860 19864 35866 19916
rect 36078 19904 36084 19916
rect 36004 19876 36084 19904
rect 33686 19845 33692 19848
rect 33505 19839 33563 19845
rect 33505 19805 33517 19839
rect 33551 19805 33563 19839
rect 33505 19799 33563 19805
rect 33653 19839 33692 19845
rect 33653 19805 33665 19839
rect 33653 19799 33692 19805
rect 33686 19796 33692 19799
rect 33744 19796 33750 19848
rect 33962 19796 33968 19848
rect 34020 19845 34026 19848
rect 34020 19836 34028 19845
rect 34020 19808 34065 19836
rect 34020 19799 34028 19808
rect 34020 19796 34026 19799
rect 34606 19796 34612 19848
rect 34664 19796 34670 19848
rect 34790 19796 34796 19848
rect 34848 19836 34854 19848
rect 34885 19839 34943 19845
rect 34885 19836 34897 19839
rect 34848 19808 34897 19836
rect 34848 19796 34854 19808
rect 34885 19805 34897 19808
rect 34931 19805 34943 19839
rect 34885 19799 34943 19805
rect 34974 19796 34980 19848
rect 35032 19836 35038 19848
rect 35069 19839 35127 19845
rect 35069 19836 35081 19839
rect 35032 19808 35081 19836
rect 35032 19796 35038 19808
rect 35069 19805 35081 19808
rect 35115 19805 35127 19839
rect 35069 19799 35127 19805
rect 35342 19796 35348 19848
rect 35400 19796 35406 19848
rect 36004 19845 36032 19876
rect 36078 19864 36084 19876
rect 36136 19904 36142 19916
rect 36265 19907 36323 19913
rect 36265 19904 36277 19907
rect 36136 19876 36277 19904
rect 36136 19864 36142 19876
rect 36265 19873 36277 19876
rect 36311 19904 36323 19907
rect 37550 19904 37556 19916
rect 36311 19876 37556 19904
rect 36311 19873 36323 19876
rect 36265 19867 36323 19873
rect 37550 19864 37556 19876
rect 37608 19864 37614 19916
rect 37660 19904 37688 19944
rect 38488 19944 38936 19972
rect 38488 19913 38516 19944
rect 38930 19932 38936 19944
rect 38988 19972 38994 19984
rect 39025 19975 39083 19981
rect 39025 19972 39037 19975
rect 38988 19944 39037 19972
rect 38988 19932 38994 19944
rect 39025 19941 39037 19944
rect 39071 19941 39083 19975
rect 39025 19935 39083 19941
rect 38473 19907 38531 19913
rect 37660 19876 37964 19904
rect 35529 19839 35587 19845
rect 35529 19805 35541 19839
rect 35575 19805 35587 19839
rect 35529 19799 35587 19805
rect 35989 19839 36047 19845
rect 35989 19805 36001 19839
rect 36035 19805 36047 19839
rect 35989 19799 36047 19805
rect 33226 19700 33232 19712
rect 31726 19672 33232 19700
rect 33226 19660 33232 19672
rect 33284 19660 33290 19712
rect 33318 19660 33324 19712
rect 33376 19700 33382 19712
rect 33704 19700 33732 19796
rect 33778 19728 33784 19780
rect 33836 19728 33842 19780
rect 33873 19771 33931 19777
rect 33873 19737 33885 19771
rect 33919 19768 33931 19771
rect 34624 19768 34652 19796
rect 33919 19740 34652 19768
rect 35544 19768 35572 19799
rect 36354 19796 36360 19848
rect 36412 19836 36418 19848
rect 36449 19839 36507 19845
rect 36449 19836 36461 19839
rect 36412 19808 36461 19836
rect 36412 19796 36418 19808
rect 36449 19805 36461 19808
rect 36495 19836 36507 19839
rect 37274 19836 37280 19848
rect 36495 19808 37280 19836
rect 36495 19805 36507 19808
rect 36449 19799 36507 19805
rect 37274 19796 37280 19808
rect 37332 19836 37338 19848
rect 37826 19836 37832 19848
rect 37332 19808 37832 19836
rect 37332 19796 37338 19808
rect 37826 19796 37832 19808
rect 37884 19796 37890 19848
rect 37936 19836 37964 19876
rect 38473 19873 38485 19907
rect 38519 19873 38531 19907
rect 38473 19867 38531 19873
rect 38565 19907 38623 19913
rect 38565 19873 38577 19907
rect 38611 19904 38623 19907
rect 39206 19904 39212 19916
rect 38611 19876 39212 19904
rect 38611 19873 38623 19876
rect 38565 19867 38623 19873
rect 39206 19864 39212 19876
rect 39264 19864 39270 19916
rect 38657 19839 38715 19845
rect 38657 19836 38669 19839
rect 37936 19808 38669 19836
rect 38657 19805 38669 19808
rect 38703 19805 38715 19839
rect 38657 19799 38715 19805
rect 38749 19839 38807 19845
rect 38749 19805 38761 19839
rect 38795 19805 38807 19839
rect 38749 19799 38807 19805
rect 35805 19771 35863 19777
rect 35805 19768 35817 19771
rect 35544 19740 35817 19768
rect 33919 19737 33931 19740
rect 33873 19731 33931 19737
rect 33376 19672 33732 19700
rect 33376 19660 33382 19672
rect 34238 19660 34244 19712
rect 34296 19700 34302 19712
rect 35544 19700 35572 19740
rect 35805 19737 35817 19740
rect 35851 19737 35863 19771
rect 35805 19731 35863 19737
rect 37642 19728 37648 19780
rect 37700 19768 37706 19780
rect 38764 19768 38792 19799
rect 38838 19796 38844 19848
rect 38896 19836 38902 19848
rect 38933 19839 38991 19845
rect 38933 19836 38945 19839
rect 38896 19808 38945 19836
rect 38896 19796 38902 19808
rect 38933 19805 38945 19808
rect 38979 19805 38991 19839
rect 38933 19799 38991 19805
rect 39022 19796 39028 19848
rect 39080 19836 39086 19848
rect 39117 19839 39175 19845
rect 39117 19836 39129 19839
rect 39080 19808 39129 19836
rect 39080 19796 39086 19808
rect 39117 19805 39129 19808
rect 39163 19805 39175 19839
rect 39117 19799 39175 19805
rect 37700 19740 38792 19768
rect 37700 19728 37706 19740
rect 34296 19672 35572 19700
rect 34296 19660 34302 19672
rect 1104 19610 41400 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 41400 19610
rect 1104 19536 41400 19558
rect 4525 19499 4583 19505
rect 4525 19465 4537 19499
rect 4571 19496 4583 19499
rect 4890 19496 4896 19508
rect 4571 19468 4896 19496
rect 4571 19465 4583 19468
rect 4525 19459 4583 19465
rect 4890 19456 4896 19468
rect 4948 19456 4954 19508
rect 4982 19456 4988 19508
rect 5040 19496 5046 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 5040 19468 5365 19496
rect 5040 19456 5046 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 5353 19459 5411 19465
rect 6822 19456 6828 19508
rect 6880 19456 6886 19508
rect 7009 19499 7067 19505
rect 7009 19465 7021 19499
rect 7055 19496 7067 19499
rect 10134 19496 10140 19508
rect 7055 19468 10140 19496
rect 7055 19465 7067 19468
rect 7009 19459 7067 19465
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 10410 19456 10416 19508
rect 10468 19456 10474 19508
rect 10594 19456 10600 19508
rect 10652 19456 10658 19508
rect 11175 19499 11233 19505
rect 11175 19496 11187 19499
rect 10796 19468 11187 19496
rect 4080 19400 4752 19428
rect 4080 19369 4108 19400
rect 4724 19372 4752 19400
rect 4798 19388 4804 19440
rect 4856 19428 4862 19440
rect 4856 19400 5028 19428
rect 4856 19388 4862 19400
rect 3881 19363 3939 19369
rect 3881 19329 3893 19363
rect 3927 19360 3939 19363
rect 4065 19363 4123 19369
rect 3927 19332 4016 19360
rect 3927 19329 3939 19332
rect 3881 19323 3939 19329
rect 3988 19292 4016 19332
rect 4065 19329 4077 19363
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4338 19292 4344 19304
rect 3988 19264 4344 19292
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 4448 19224 4476 19323
rect 4614 19320 4620 19372
rect 4672 19320 4678 19372
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5000 19369 5028 19400
rect 4893 19363 4951 19369
rect 4893 19360 4905 19363
rect 4764 19332 4905 19360
rect 4764 19320 4770 19332
rect 4893 19329 4905 19332
rect 4939 19329 4951 19363
rect 4893 19323 4951 19329
rect 4985 19363 5043 19369
rect 4985 19329 4997 19363
rect 5031 19360 5043 19363
rect 5442 19360 5448 19372
rect 5031 19332 5448 19360
rect 5031 19329 5043 19332
rect 4985 19323 5043 19329
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 6457 19363 6515 19369
rect 6457 19360 6469 19363
rect 5828 19332 6469 19360
rect 4522 19252 4528 19304
rect 4580 19292 4586 19304
rect 4801 19295 4859 19301
rect 4801 19292 4813 19295
rect 4580 19264 4813 19292
rect 4580 19252 4586 19264
rect 4801 19261 4813 19264
rect 4847 19292 4859 19295
rect 4847 19264 4936 19292
rect 4847 19261 4859 19264
rect 4801 19255 4859 19261
rect 4908 19224 4936 19264
rect 5828 19236 5856 19332
rect 6457 19329 6469 19332
rect 6503 19329 6515 19363
rect 6457 19323 6515 19329
rect 6638 19320 6644 19372
rect 6696 19320 6702 19372
rect 6840 19360 6868 19456
rect 9677 19431 9735 19437
rect 9677 19428 9689 19431
rect 8772 19400 9689 19428
rect 6947 19363 7005 19369
rect 6947 19360 6959 19363
rect 6840 19332 6959 19360
rect 6947 19329 6959 19332
rect 6993 19329 7005 19363
rect 6947 19323 7005 19329
rect 7282 19320 7288 19372
rect 7340 19360 7346 19372
rect 8772 19369 8800 19400
rect 9677 19397 9689 19400
rect 9723 19397 9735 19431
rect 9950 19428 9956 19440
rect 9677 19391 9735 19397
rect 9784 19400 9956 19428
rect 8297 19363 8355 19369
rect 8297 19360 8309 19363
rect 7340 19332 8309 19360
rect 7340 19320 7346 19332
rect 8297 19329 8309 19332
rect 8343 19329 8355 19363
rect 8297 19323 8355 19329
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19360 8999 19363
rect 8987 19332 9260 19360
rect 8987 19329 8999 19332
rect 8941 19323 8999 19329
rect 5994 19252 6000 19304
rect 6052 19292 6058 19304
rect 7469 19295 7527 19301
rect 7469 19292 7481 19295
rect 6052 19264 7481 19292
rect 6052 19252 6058 19264
rect 7469 19261 7481 19264
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 5537 19227 5595 19233
rect 5537 19224 5549 19227
rect 4448 19196 4844 19224
rect 4908 19196 5549 19224
rect 4816 19168 4844 19196
rect 5537 19193 5549 19196
rect 5583 19193 5595 19227
rect 5537 19187 5595 19193
rect 5810 19184 5816 19236
rect 5868 19184 5874 19236
rect 6549 19227 6607 19233
rect 6549 19193 6561 19227
rect 6595 19224 6607 19227
rect 7377 19227 7435 19233
rect 7377 19224 7389 19227
rect 6595 19196 7389 19224
rect 6595 19193 6607 19196
rect 6549 19187 6607 19193
rect 7377 19193 7389 19196
rect 7423 19193 7435 19227
rect 7377 19187 7435 19193
rect 3878 19116 3884 19168
rect 3936 19116 3942 19168
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4614 19156 4620 19168
rect 4203 19128 4620 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 4798 19116 4804 19168
rect 4856 19116 4862 19168
rect 5166 19116 5172 19168
rect 5224 19156 5230 19168
rect 5353 19159 5411 19165
rect 5353 19156 5365 19159
rect 5224 19128 5365 19156
rect 5224 19116 5230 19128
rect 5353 19125 5365 19128
rect 5399 19156 5411 19159
rect 6362 19156 6368 19168
rect 5399 19128 6368 19156
rect 5399 19125 5411 19128
rect 5353 19119 5411 19125
rect 6362 19116 6368 19128
rect 6420 19116 6426 19168
rect 6825 19159 6883 19165
rect 6825 19125 6837 19159
rect 6871 19156 6883 19159
rect 7006 19156 7012 19168
rect 6871 19128 7012 19156
rect 6871 19125 6883 19128
rect 6825 19119 6883 19125
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 7929 19159 7987 19165
rect 7929 19156 7941 19159
rect 7800 19128 7941 19156
rect 7800 19116 7806 19128
rect 7929 19125 7941 19128
rect 7975 19125 7987 19159
rect 8312 19156 8340 19323
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19261 8447 19295
rect 8389 19255 8447 19261
rect 8404 19224 8432 19255
rect 8570 19252 8576 19304
rect 8628 19252 8634 19304
rect 8662 19252 8668 19304
rect 8720 19292 8726 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8720 19264 9045 19292
rect 8720 19252 8726 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 9122 19252 9128 19304
rect 9180 19252 9186 19304
rect 9232 19292 9260 19332
rect 9306 19320 9312 19372
rect 9364 19320 9370 19372
rect 9398 19320 9404 19372
rect 9456 19320 9462 19372
rect 9582 19320 9588 19372
rect 9640 19320 9646 19372
rect 9784 19369 9812 19400
rect 9950 19388 9956 19400
rect 10008 19428 10014 19440
rect 10428 19428 10456 19456
rect 10008 19400 10456 19428
rect 10008 19388 10014 19400
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19329 9827 19363
rect 9769 19323 9827 19329
rect 10229 19363 10287 19369
rect 10229 19329 10241 19363
rect 10275 19360 10287 19363
rect 10318 19360 10324 19372
rect 10275 19332 10324 19360
rect 10275 19329 10287 19332
rect 10229 19323 10287 19329
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 10612 19369 10640 19456
rect 10796 19369 10824 19468
rect 11175 19465 11187 19468
rect 11221 19496 11233 19499
rect 12526 19496 12532 19508
rect 11221 19468 12532 19496
rect 11221 19465 11233 19468
rect 11175 19459 11233 19465
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 16482 19496 16488 19508
rect 12636 19468 16488 19496
rect 10965 19431 11023 19437
rect 10965 19397 10977 19431
rect 11011 19428 11023 19431
rect 11330 19428 11336 19440
rect 11011 19400 11336 19428
rect 11011 19397 11023 19400
rect 10965 19391 11023 19397
rect 11330 19388 11336 19400
rect 11388 19428 11394 19440
rect 11517 19431 11575 19437
rect 11517 19428 11529 19431
rect 11388 19400 11529 19428
rect 11388 19388 11394 19400
rect 11517 19397 11529 19400
rect 11563 19397 11575 19431
rect 11517 19391 11575 19397
rect 11701 19431 11759 19437
rect 11701 19397 11713 19431
rect 11747 19428 11759 19431
rect 12342 19428 12348 19440
rect 11747 19400 12348 19428
rect 11747 19397 11759 19400
rect 11701 19391 11759 19397
rect 10413 19363 10471 19369
rect 10413 19329 10425 19363
rect 10459 19334 10471 19363
rect 10597 19363 10655 19369
rect 10459 19329 10548 19334
rect 10413 19323 10548 19329
rect 10597 19329 10609 19363
rect 10643 19329 10655 19363
rect 10597 19323 10655 19329
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19329 10839 19363
rect 11716 19360 11744 19391
rect 12342 19388 12348 19400
rect 12400 19388 12406 19440
rect 12636 19369 12664 19468
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 17313 19499 17371 19505
rect 17313 19465 17325 19499
rect 17359 19496 17371 19499
rect 17402 19496 17408 19508
rect 17359 19468 17408 19496
rect 17359 19465 17371 19468
rect 17313 19459 17371 19465
rect 17402 19456 17408 19468
rect 17460 19496 17466 19508
rect 17681 19499 17739 19505
rect 17681 19496 17693 19499
rect 17460 19468 17693 19496
rect 17460 19456 17466 19468
rect 17681 19465 17693 19468
rect 17727 19465 17739 19499
rect 20622 19496 20628 19508
rect 17681 19459 17739 19465
rect 17788 19468 20628 19496
rect 13814 19388 13820 19440
rect 13872 19428 13878 19440
rect 14093 19431 14151 19437
rect 14093 19428 14105 19431
rect 13872 19400 14105 19428
rect 13872 19388 13878 19400
rect 14093 19397 14105 19400
rect 14139 19397 14151 19431
rect 14093 19391 14151 19397
rect 14182 19388 14188 19440
rect 14240 19428 14246 19440
rect 14461 19431 14519 19437
rect 14461 19428 14473 19431
rect 14240 19400 14473 19428
rect 14240 19388 14246 19400
rect 14461 19397 14473 19400
rect 14507 19428 14519 19431
rect 14737 19431 14795 19437
rect 14737 19428 14749 19431
rect 14507 19400 14749 19428
rect 14507 19397 14519 19400
rect 14461 19391 14519 19397
rect 14737 19397 14749 19400
rect 14783 19428 14795 19431
rect 14826 19428 14832 19440
rect 14783 19400 14832 19428
rect 14783 19397 14795 19400
rect 14737 19391 14795 19397
rect 14826 19388 14832 19400
rect 14884 19388 14890 19440
rect 14921 19431 14979 19437
rect 14921 19397 14933 19431
rect 14967 19428 14979 19431
rect 15010 19428 15016 19440
rect 14967 19400 15016 19428
rect 14967 19397 14979 19400
rect 14921 19391 14979 19397
rect 15010 19388 15016 19400
rect 15068 19388 15074 19440
rect 17497 19431 17555 19437
rect 17497 19428 17509 19431
rect 17328 19400 17509 19428
rect 12621 19363 12679 19369
rect 12621 19360 12633 19363
rect 10781 19323 10839 19329
rect 10888 19332 11744 19360
rect 11808 19332 12633 19360
rect 9416 19292 9444 19320
rect 10428 19306 10548 19323
rect 9232 19264 9444 19292
rect 10520 19292 10548 19306
rect 10888 19292 10916 19332
rect 10520 19264 10916 19292
rect 10962 19252 10968 19304
rect 11020 19292 11026 19304
rect 11808 19292 11836 19332
rect 12621 19329 12633 19332
rect 12667 19329 12679 19363
rect 12621 19323 12679 19329
rect 12710 19320 12716 19372
rect 12768 19360 12774 19372
rect 12805 19363 12863 19369
rect 12805 19360 12817 19363
rect 12768 19332 12817 19360
rect 12768 19320 12774 19332
rect 12805 19329 12817 19332
rect 12851 19329 12863 19363
rect 12805 19323 12863 19329
rect 12986 19320 12992 19372
rect 13044 19320 13050 19372
rect 13998 19320 14004 19372
rect 14056 19360 14062 19372
rect 14277 19363 14335 19369
rect 14277 19360 14289 19363
rect 14056 19332 14289 19360
rect 14056 19320 14062 19332
rect 14277 19329 14289 19332
rect 14323 19329 14335 19363
rect 14277 19323 14335 19329
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19329 14427 19363
rect 14369 19323 14427 19329
rect 11020 19264 11836 19292
rect 11020 19252 11026 19264
rect 9493 19227 9551 19233
rect 9493 19224 9505 19227
rect 8404 19196 9505 19224
rect 9493 19193 9505 19196
rect 9539 19193 9551 19227
rect 11790 19224 11796 19236
rect 9493 19187 9551 19193
rect 11164 19196 11796 19224
rect 9214 19156 9220 19168
rect 8312 19128 9220 19156
rect 7929 19119 7987 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 9582 19116 9588 19168
rect 9640 19156 9646 19168
rect 10321 19159 10379 19165
rect 10321 19156 10333 19159
rect 9640 19128 10333 19156
rect 9640 19116 9646 19128
rect 10321 19125 10333 19128
rect 10367 19125 10379 19159
rect 10321 19119 10379 19125
rect 10410 19116 10416 19168
rect 10468 19156 10474 19168
rect 11164 19165 11192 19196
rect 10597 19159 10655 19165
rect 10597 19156 10609 19159
rect 10468 19128 10609 19156
rect 10468 19116 10474 19128
rect 10597 19125 10609 19128
rect 10643 19125 10655 19159
rect 10597 19119 10655 19125
rect 11149 19159 11207 19165
rect 11149 19125 11161 19159
rect 11195 19125 11207 19159
rect 11149 19119 11207 19125
rect 11330 19116 11336 19168
rect 11388 19116 11394 19168
rect 11716 19165 11744 19196
rect 11790 19184 11796 19196
rect 11848 19224 11854 19236
rect 11848 19196 12664 19224
rect 11848 19184 11854 19196
rect 12636 19168 12664 19196
rect 14274 19184 14280 19236
rect 14332 19224 14338 19236
rect 14384 19224 14412 19323
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 17328 19360 17356 19400
rect 17497 19397 17509 19400
rect 17543 19397 17555 19431
rect 17497 19391 17555 19397
rect 17000 19332 17356 19360
rect 17405 19363 17463 19369
rect 17000 19320 17006 19332
rect 17405 19329 17417 19363
rect 17451 19360 17463 19363
rect 17678 19360 17684 19372
rect 17451 19332 17684 19360
rect 17451 19329 17463 19332
rect 17405 19323 17463 19329
rect 17678 19320 17684 19332
rect 17736 19360 17742 19372
rect 17788 19369 17816 19468
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 24946 19456 24952 19508
rect 25004 19456 25010 19508
rect 25498 19456 25504 19508
rect 25556 19496 25562 19508
rect 26053 19499 26111 19505
rect 26053 19496 26065 19499
rect 25556 19468 26065 19496
rect 25556 19456 25562 19468
rect 26053 19465 26065 19468
rect 26099 19465 26111 19499
rect 26053 19459 26111 19465
rect 31662 19456 31668 19508
rect 31720 19496 31726 19508
rect 34238 19496 34244 19508
rect 31720 19468 34244 19496
rect 31720 19456 31726 19468
rect 17862 19388 17868 19440
rect 17920 19428 17926 19440
rect 20070 19428 20076 19440
rect 17920 19400 20076 19428
rect 17920 19388 17926 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 24964 19428 24992 19456
rect 25409 19431 25467 19437
rect 25409 19428 25421 19431
rect 21744 19400 23336 19428
rect 24964 19400 25421 19428
rect 21744 19372 21772 19400
rect 17773 19363 17831 19369
rect 17773 19360 17785 19363
rect 17736 19332 17785 19360
rect 17736 19320 17742 19332
rect 17773 19329 17785 19332
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 18322 19320 18328 19372
rect 18380 19320 18386 19372
rect 19150 19320 19156 19372
rect 19208 19360 19214 19372
rect 19208 19332 19380 19360
rect 19208 19320 19214 19332
rect 17034 19252 17040 19304
rect 17092 19252 17098 19304
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19292 17187 19295
rect 18340 19292 18368 19320
rect 17175 19264 18368 19292
rect 19352 19292 19380 19332
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19484 19332 19533 19360
rect 19484 19320 19490 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 20162 19320 20168 19372
rect 20220 19320 20226 19372
rect 20254 19320 20260 19372
rect 20312 19320 20318 19372
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 20364 19332 20637 19360
rect 20364 19292 20392 19332
rect 20625 19329 20637 19332
rect 20671 19360 20683 19363
rect 21634 19360 21640 19372
rect 20671 19332 21640 19360
rect 20671 19329 20683 19332
rect 20625 19323 20683 19329
rect 21634 19320 21640 19332
rect 21692 19320 21698 19372
rect 21726 19320 21732 19372
rect 21784 19320 21790 19372
rect 21818 19320 21824 19372
rect 21876 19320 21882 19372
rect 21910 19320 21916 19372
rect 21968 19360 21974 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21968 19332 22017 19360
rect 21968 19320 21974 19332
rect 22005 19329 22017 19332
rect 22051 19360 22063 19363
rect 22186 19360 22192 19372
rect 22051 19332 22192 19360
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22278 19320 22284 19372
rect 22336 19320 22342 19372
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 23308 19369 23336 19400
rect 25409 19397 25421 19400
rect 25455 19397 25467 19431
rect 27430 19428 27436 19440
rect 25409 19391 25467 19397
rect 25792 19400 27436 19428
rect 23017 19363 23075 19369
rect 23017 19360 23029 19363
rect 22704 19332 23029 19360
rect 22704 19320 22710 19332
rect 23017 19329 23029 19332
rect 23063 19329 23075 19363
rect 23017 19323 23075 19329
rect 23293 19363 23351 19369
rect 23293 19329 23305 19363
rect 23339 19329 23351 19363
rect 23293 19323 23351 19329
rect 23400 19332 24164 19360
rect 19352 19264 20392 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 20901 19295 20959 19301
rect 20901 19292 20913 19295
rect 20772 19264 20913 19292
rect 20772 19252 20778 19264
rect 20901 19261 20913 19264
rect 20947 19261 20959 19295
rect 20901 19255 20959 19261
rect 22370 19252 22376 19304
rect 22428 19292 22434 19304
rect 22428 19264 22692 19292
rect 22428 19252 22434 19264
rect 14332 19196 14412 19224
rect 14332 19184 14338 19196
rect 16390 19184 16396 19236
rect 16448 19224 16454 19236
rect 21726 19224 21732 19236
rect 16448 19196 21732 19224
rect 16448 19184 16454 19196
rect 21726 19184 21732 19196
rect 21784 19184 21790 19236
rect 22278 19184 22284 19236
rect 22336 19224 22342 19236
rect 22557 19227 22615 19233
rect 22557 19224 22569 19227
rect 22336 19196 22569 19224
rect 22336 19184 22342 19196
rect 22557 19193 22569 19196
rect 22603 19193 22615 19227
rect 22664 19224 22692 19264
rect 22830 19252 22836 19304
rect 22888 19292 22894 19304
rect 23400 19292 23428 19332
rect 22888 19264 23428 19292
rect 22888 19252 22894 19264
rect 23474 19252 23480 19304
rect 23532 19292 23538 19304
rect 24026 19292 24032 19304
rect 23532 19264 24032 19292
rect 23532 19252 23538 19264
rect 24026 19252 24032 19264
rect 24084 19252 24090 19304
rect 24136 19292 24164 19332
rect 24946 19320 24952 19372
rect 25004 19360 25010 19372
rect 25792 19369 25820 19400
rect 27430 19388 27436 19400
rect 27488 19388 27494 19440
rect 31754 19428 31760 19440
rect 31418 19400 31760 19428
rect 31754 19388 31760 19400
rect 31812 19388 31818 19440
rect 33226 19388 33232 19440
rect 33284 19388 33290 19440
rect 33888 19437 33916 19468
rect 34238 19456 34244 19468
rect 34296 19456 34302 19508
rect 33873 19431 33931 19437
rect 33873 19397 33885 19431
rect 33919 19397 33931 19431
rect 33873 19391 33931 19397
rect 25777 19363 25835 19369
rect 25004 19332 25728 19360
rect 25004 19320 25010 19332
rect 25038 19292 25044 19304
rect 24136 19264 25044 19292
rect 25038 19252 25044 19264
rect 25096 19252 25102 19304
rect 25700 19292 25728 19332
rect 25777 19329 25789 19363
rect 25823 19329 25835 19363
rect 25777 19323 25835 19329
rect 25869 19363 25927 19369
rect 25869 19329 25881 19363
rect 25915 19360 25927 19363
rect 26510 19360 26516 19372
rect 25915 19332 26516 19360
rect 25915 19329 25927 19332
rect 25869 19323 25927 19329
rect 25884 19292 25912 19323
rect 26510 19320 26516 19332
rect 26568 19320 26574 19372
rect 27341 19363 27399 19369
rect 27341 19329 27353 19363
rect 27387 19360 27399 19363
rect 27706 19360 27712 19372
rect 27387 19332 27712 19360
rect 27387 19329 27399 19332
rect 27341 19323 27399 19329
rect 27706 19320 27712 19332
rect 27764 19360 27770 19372
rect 27764 19332 28488 19360
rect 27764 19320 27770 19332
rect 25700 19264 25912 19292
rect 25958 19252 25964 19304
rect 26016 19252 26022 19304
rect 27525 19295 27583 19301
rect 27525 19261 27537 19295
rect 27571 19261 27583 19295
rect 27525 19255 27583 19261
rect 25976 19224 26004 19252
rect 22664 19196 26004 19224
rect 22557 19187 22615 19193
rect 26694 19184 26700 19236
rect 26752 19224 26758 19236
rect 27540 19224 27568 19255
rect 26752 19196 27568 19224
rect 28460 19224 28488 19332
rect 28626 19320 28632 19372
rect 28684 19360 28690 19372
rect 29178 19360 29184 19372
rect 28684 19332 29184 19360
rect 28684 19320 28690 19332
rect 29178 19320 29184 19332
rect 29236 19320 29242 19372
rect 29917 19363 29975 19369
rect 29917 19360 29929 19363
rect 29288 19332 29929 19360
rect 29288 19304 29316 19332
rect 29917 19329 29929 19332
rect 29963 19329 29975 19363
rect 29917 19323 29975 19329
rect 31478 19320 31484 19372
rect 31536 19360 31542 19372
rect 32125 19363 32183 19369
rect 32125 19360 32137 19363
rect 31536 19332 32137 19360
rect 31536 19320 31542 19332
rect 32125 19329 32137 19332
rect 32171 19329 32183 19363
rect 33244 19360 33272 19388
rect 37366 19360 37372 19372
rect 33244 19332 37372 19360
rect 32125 19323 32183 19329
rect 37366 19320 37372 19332
rect 37424 19320 37430 19372
rect 39114 19320 39120 19372
rect 39172 19360 39178 19372
rect 40034 19360 40040 19372
rect 39172 19332 40040 19360
rect 39172 19320 39178 19332
rect 40034 19320 40040 19332
rect 40092 19320 40098 19372
rect 29270 19252 29276 19304
rect 29328 19252 29334 19304
rect 29546 19252 29552 19304
rect 29604 19252 29610 19304
rect 30190 19252 30196 19304
rect 30248 19252 30254 19304
rect 30282 19252 30288 19304
rect 30340 19292 30346 19304
rect 30340 19264 31754 19292
rect 30340 19252 30346 19264
rect 29564 19224 29592 19252
rect 28460 19196 29592 19224
rect 31726 19224 31754 19264
rect 35986 19252 35992 19304
rect 36044 19292 36050 19304
rect 37274 19292 37280 19304
rect 36044 19264 37280 19292
rect 36044 19252 36050 19264
rect 37274 19252 37280 19264
rect 37332 19252 37338 19304
rect 36078 19224 36084 19236
rect 31726 19196 36084 19224
rect 26752 19184 26758 19196
rect 36078 19184 36084 19196
rect 36136 19184 36142 19236
rect 11701 19159 11759 19165
rect 11701 19125 11713 19159
rect 11747 19125 11759 19159
rect 11701 19119 11759 19125
rect 11882 19116 11888 19168
rect 11940 19116 11946 19168
rect 12618 19116 12624 19168
rect 12676 19116 12682 19168
rect 14642 19116 14648 19168
rect 14700 19116 14706 19168
rect 15105 19159 15163 19165
rect 15105 19125 15117 19159
rect 15151 19156 15163 19159
rect 15562 19156 15568 19168
rect 15151 19128 15568 19156
rect 15151 19125 15163 19128
rect 15105 19119 15163 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16669 19159 16727 19165
rect 16669 19125 16681 19159
rect 16715 19156 16727 19159
rect 16850 19156 16856 19168
rect 16715 19128 16856 19156
rect 16715 19125 16727 19128
rect 16669 19119 16727 19125
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 17494 19116 17500 19168
rect 17552 19116 17558 19168
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18782 19156 18788 19168
rect 18104 19128 18788 19156
rect 18104 19116 18110 19128
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 22189 19159 22247 19165
rect 22189 19125 22201 19159
rect 22235 19156 22247 19159
rect 24670 19156 24676 19168
rect 22235 19128 24676 19156
rect 22235 19125 22247 19128
rect 22189 19119 22247 19125
rect 24670 19116 24676 19128
rect 24728 19116 24734 19168
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 26970 19116 26976 19168
rect 27028 19116 27034 19168
rect 28994 19116 29000 19168
rect 29052 19156 29058 19168
rect 30282 19156 30288 19168
rect 29052 19128 30288 19156
rect 29052 19116 29058 19128
rect 30282 19116 30288 19128
rect 30340 19116 30346 19168
rect 30374 19116 30380 19168
rect 30432 19156 30438 19168
rect 31386 19156 31392 19168
rect 30432 19128 31392 19156
rect 30432 19116 30438 19128
rect 31386 19116 31392 19128
rect 31444 19156 31450 19168
rect 31665 19159 31723 19165
rect 31665 19156 31677 19159
rect 31444 19128 31677 19156
rect 31444 19116 31450 19128
rect 31665 19125 31677 19128
rect 31711 19125 31723 19159
rect 31665 19119 31723 19125
rect 32214 19116 32220 19168
rect 32272 19116 32278 19168
rect 32858 19116 32864 19168
rect 32916 19156 32922 19168
rect 33962 19156 33968 19168
rect 32916 19128 33968 19156
rect 32916 19116 32922 19128
rect 33962 19116 33968 19128
rect 34020 19116 34026 19168
rect 34146 19116 34152 19168
rect 34204 19116 34210 19168
rect 1104 19066 41400 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 41400 19066
rect 1104 18992 41400 19014
rect 4522 18912 4528 18964
rect 4580 18952 4586 18964
rect 6914 18952 6920 18964
rect 4580 18924 6920 18952
rect 4580 18912 4586 18924
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 10229 18955 10287 18961
rect 10229 18952 10241 18955
rect 8680 18924 10241 18952
rect 8680 18896 8708 18924
rect 10229 18921 10241 18924
rect 10275 18921 10287 18955
rect 10229 18915 10287 18921
rect 11514 18912 11520 18964
rect 11572 18952 11578 18964
rect 15194 18952 15200 18964
rect 11572 18924 15200 18952
rect 11572 18912 11578 18924
rect 15194 18912 15200 18924
rect 15252 18912 15258 18964
rect 16022 18912 16028 18964
rect 16080 18952 16086 18964
rect 17405 18955 17463 18961
rect 16080 18924 17356 18952
rect 16080 18912 16086 18924
rect 5810 18884 5816 18896
rect 3896 18856 5034 18884
rect 3896 18828 3924 18856
rect 3878 18776 3884 18828
rect 3936 18776 3942 18828
rect 4522 18776 4528 18828
rect 4580 18776 4586 18828
rect 4890 18776 4896 18828
rect 4948 18776 4954 18828
rect 5006 18816 5034 18856
rect 5644 18856 5816 18884
rect 5169 18819 5227 18825
rect 5169 18816 5181 18819
rect 5006 18788 5181 18816
rect 5169 18785 5181 18788
rect 5215 18785 5227 18819
rect 5169 18779 5227 18785
rect 5350 18776 5356 18828
rect 5408 18776 5414 18828
rect 4338 18708 4344 18760
rect 4396 18708 4402 18760
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18717 5043 18751
rect 4985 18711 5043 18717
rect 5077 18751 5135 18757
rect 5077 18717 5089 18751
rect 5123 18748 5135 18751
rect 5442 18748 5448 18760
rect 5123 18720 5448 18748
rect 5123 18717 5135 18720
rect 5077 18711 5135 18717
rect 4249 18683 4307 18689
rect 4249 18649 4261 18683
rect 4295 18680 4307 18683
rect 5000 18680 5028 18711
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 5534 18708 5540 18760
rect 5592 18708 5598 18760
rect 5644 18680 5672 18856
rect 5810 18844 5816 18856
rect 5868 18884 5874 18896
rect 6273 18887 6331 18893
rect 6273 18884 6285 18887
rect 5868 18856 6285 18884
rect 5868 18844 5874 18856
rect 6273 18853 6285 18856
rect 6319 18853 6331 18887
rect 6273 18847 6331 18853
rect 6822 18844 6828 18896
rect 6880 18884 6886 18896
rect 8202 18884 8208 18896
rect 6880 18856 8208 18884
rect 6880 18844 6886 18856
rect 8202 18844 8208 18856
rect 8260 18884 8266 18896
rect 8662 18884 8668 18896
rect 8260 18856 8668 18884
rect 8260 18844 8266 18856
rect 6362 18816 6368 18828
rect 5828 18788 6368 18816
rect 5828 18757 5856 18788
rect 6362 18776 6368 18788
rect 6420 18776 6426 18828
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7024 18788 7849 18816
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18717 5871 18751
rect 5813 18711 5871 18717
rect 4295 18652 4752 18680
rect 5000 18652 5672 18680
rect 4295 18649 4307 18652
rect 4249 18643 4307 18649
rect 3878 18572 3884 18624
rect 3936 18572 3942 18624
rect 4724 18621 4752 18652
rect 6362 18640 6368 18692
rect 6420 18680 6426 18692
rect 6457 18683 6515 18689
rect 6457 18680 6469 18683
rect 6420 18652 6469 18680
rect 6420 18640 6426 18652
rect 6457 18649 6469 18652
rect 6503 18649 6515 18683
rect 6457 18643 6515 18649
rect 6546 18640 6552 18692
rect 6604 18689 6610 18692
rect 6604 18683 6617 18689
rect 6605 18680 6617 18683
rect 6605 18652 6649 18680
rect 6605 18649 6617 18652
rect 6604 18643 6617 18649
rect 6604 18640 6610 18643
rect 6822 18640 6828 18692
rect 6880 18640 6886 18692
rect 6917 18683 6975 18689
rect 6917 18649 6929 18683
rect 6963 18680 6975 18683
rect 7024 18680 7052 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7282 18748 7288 18760
rect 7147 18720 7288 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 7374 18708 7380 18760
rect 7432 18748 7438 18760
rect 7653 18751 7711 18757
rect 7432 18720 7604 18748
rect 7432 18708 7438 18720
rect 6963 18652 7052 18680
rect 6963 18649 6975 18652
rect 6917 18643 6975 18649
rect 7466 18640 7472 18692
rect 7524 18640 7530 18692
rect 7576 18680 7604 18720
rect 7653 18717 7665 18751
rect 7699 18748 7711 18751
rect 7742 18748 7748 18760
rect 7699 18720 7748 18748
rect 7699 18717 7711 18720
rect 7653 18711 7711 18717
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 7926 18708 7932 18760
rect 7984 18708 7990 18760
rect 8496 18757 8524 18856
rect 8662 18844 8668 18856
rect 8720 18844 8726 18896
rect 9214 18844 9220 18896
rect 9272 18884 9278 18896
rect 9769 18887 9827 18893
rect 9769 18884 9781 18887
rect 9272 18856 9781 18884
rect 9272 18844 9278 18856
rect 9769 18853 9781 18856
rect 9815 18853 9827 18887
rect 9769 18847 9827 18853
rect 9858 18844 9864 18896
rect 9916 18884 9922 18896
rect 17328 18884 17356 18924
rect 17405 18921 17417 18955
rect 17451 18952 17463 18955
rect 17678 18952 17684 18964
rect 17451 18924 17684 18952
rect 17451 18921 17463 18924
rect 17405 18915 17463 18921
rect 17678 18912 17684 18924
rect 17736 18952 17742 18964
rect 18138 18952 18144 18964
rect 17736 18924 18144 18952
rect 17736 18912 17742 18924
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 18690 18912 18696 18964
rect 18748 18912 18754 18964
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 20254 18952 20260 18964
rect 19944 18924 20260 18952
rect 19944 18912 19950 18924
rect 20254 18912 20260 18924
rect 20312 18912 20318 18964
rect 22370 18952 22376 18964
rect 20364 18924 22376 18952
rect 9916 18856 12112 18884
rect 9916 18844 9922 18856
rect 9232 18757 9260 18844
rect 9416 18788 10088 18816
rect 9416 18757 9444 18788
rect 10060 18757 10088 18788
rect 8481 18751 8539 18757
rect 8481 18717 8493 18751
rect 8527 18717 8539 18751
rect 8481 18711 8539 18717
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18748 8631 18751
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8619 18720 8953 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18717 9459 18751
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9401 18711 9459 18717
rect 9600 18720 9873 18748
rect 9306 18680 9312 18692
rect 7576 18652 9312 18680
rect 9306 18640 9312 18652
rect 9364 18640 9370 18692
rect 9490 18640 9496 18692
rect 9548 18680 9554 18692
rect 9600 18689 9628 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18748 10103 18751
rect 10091 18720 12020 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 9585 18683 9643 18689
rect 9585 18680 9597 18683
rect 9548 18652 9597 18680
rect 9548 18640 9554 18652
rect 9585 18649 9597 18652
rect 9631 18649 9643 18683
rect 9585 18643 9643 18649
rect 10410 18640 10416 18692
rect 10468 18640 10474 18692
rect 4709 18615 4767 18621
rect 4709 18581 4721 18615
rect 4755 18581 4767 18615
rect 4709 18575 4767 18581
rect 4982 18572 4988 18624
rect 5040 18612 5046 18624
rect 5721 18615 5779 18621
rect 5721 18612 5733 18615
rect 5040 18584 5733 18612
rect 5040 18572 5046 18584
rect 5721 18581 5733 18584
rect 5767 18612 5779 18615
rect 6641 18615 6699 18621
rect 6641 18612 6653 18615
rect 5767 18584 6653 18612
rect 5767 18581 5779 18584
rect 5721 18575 5779 18581
rect 6641 18581 6653 18584
rect 6687 18612 6699 18615
rect 6730 18612 6736 18624
rect 6687 18584 6736 18612
rect 6687 18581 6699 18584
rect 6641 18575 6699 18581
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 7190 18572 7196 18624
rect 7248 18612 7254 18624
rect 7285 18615 7343 18621
rect 7285 18612 7297 18615
rect 7248 18584 7297 18612
rect 7248 18572 7254 18584
rect 7285 18581 7297 18584
rect 7331 18581 7343 18615
rect 7285 18575 7343 18581
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 10428 18612 10456 18640
rect 11992 18624 12020 18720
rect 10962 18612 10968 18624
rect 8628 18584 10968 18612
rect 8628 18572 8634 18584
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11974 18572 11980 18624
rect 12032 18572 12038 18624
rect 12084 18612 12112 18856
rect 13832 18856 17264 18884
rect 17328 18856 17816 18884
rect 12434 18708 12440 18760
rect 12492 18708 12498 18760
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 13832 18748 13860 18856
rect 16390 18776 16396 18828
rect 16448 18776 16454 18828
rect 16574 18776 16580 18828
rect 16632 18776 16638 18828
rect 16666 18776 16672 18828
rect 16724 18776 16730 18828
rect 16761 18819 16819 18825
rect 16761 18785 16773 18819
rect 16807 18816 16819 18819
rect 17236 18816 17264 18856
rect 17788 18816 17816 18856
rect 17862 18844 17868 18896
rect 17920 18884 17926 18896
rect 20364 18884 20392 18924
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 22462 18912 22468 18964
rect 22520 18952 22526 18964
rect 23017 18955 23075 18961
rect 23017 18952 23029 18955
rect 22520 18924 23029 18952
rect 22520 18912 22526 18924
rect 23017 18921 23029 18924
rect 23063 18921 23075 18955
rect 23017 18915 23075 18921
rect 23290 18912 23296 18964
rect 23348 18912 23354 18964
rect 29273 18955 29331 18961
rect 23400 18924 29224 18952
rect 17920 18856 20392 18884
rect 17920 18844 17926 18856
rect 21542 18844 21548 18896
rect 21600 18884 21606 18896
rect 22922 18884 22928 18896
rect 21600 18856 22928 18884
rect 21600 18844 21606 18856
rect 22922 18844 22928 18856
rect 22980 18844 22986 18896
rect 18785 18819 18843 18825
rect 16807 18788 17172 18816
rect 17236 18788 17724 18816
rect 17788 18788 18736 18816
rect 16807 18785 16819 18788
rect 16761 18779 16819 18785
rect 12676 18720 13860 18748
rect 12676 18708 12682 18720
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 14277 18751 14335 18757
rect 14277 18748 14289 18751
rect 13964 18720 14289 18748
rect 13964 18708 13970 18720
rect 14277 18717 14289 18720
rect 14323 18717 14335 18751
rect 14277 18711 14335 18717
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18717 14795 18751
rect 14737 18711 14795 18717
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 12713 18683 12771 18689
rect 12713 18680 12725 18683
rect 12308 18652 12725 18680
rect 12308 18640 12314 18652
rect 12713 18649 12725 18652
rect 12759 18649 12771 18683
rect 12713 18643 12771 18649
rect 13078 18612 13084 18624
rect 12084 18584 13084 18612
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 14292 18612 14320 18711
rect 14752 18680 14780 18711
rect 14826 18708 14832 18760
rect 14884 18748 14890 18760
rect 14921 18751 14979 18757
rect 14921 18748 14933 18751
rect 14884 18720 14933 18748
rect 14884 18708 14890 18720
rect 14921 18717 14933 18720
rect 14967 18717 14979 18751
rect 14921 18711 14979 18717
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 16206 18748 16212 18760
rect 16163 18720 16212 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 17144 18757 17172 18788
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 17494 18748 17500 18760
rect 17175 18720 17500 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 15028 18680 15056 18708
rect 14752 18652 15056 18680
rect 15286 18640 15292 18692
rect 15344 18640 15350 18692
rect 16224 18680 16252 18708
rect 16868 18680 16896 18711
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18717 17647 18751
rect 17696 18748 17724 18788
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 17696 18720 18521 18748
rect 17589 18711 17647 18717
rect 18509 18717 18521 18720
rect 18555 18717 18567 18751
rect 18708 18748 18736 18788
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 18874 18816 18880 18828
rect 18831 18788 18880 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 18874 18776 18880 18788
rect 18932 18776 18938 18828
rect 21910 18776 21916 18828
rect 21968 18816 21974 18828
rect 23308 18816 23336 18912
rect 23400 18828 23428 18924
rect 23658 18844 23664 18896
rect 23716 18884 23722 18896
rect 24394 18884 24400 18896
rect 23716 18856 24400 18884
rect 23716 18844 23722 18856
rect 24394 18844 24400 18856
rect 24452 18884 24458 18896
rect 24452 18856 25268 18884
rect 24452 18844 24458 18856
rect 21968 18788 23336 18816
rect 21968 18776 21974 18788
rect 23382 18776 23388 18828
rect 23440 18776 23446 18828
rect 23474 18776 23480 18828
rect 23532 18816 23538 18828
rect 23532 18788 23980 18816
rect 23532 18776 23538 18788
rect 19426 18748 19432 18760
rect 18708 18720 19432 18748
rect 18509 18711 18567 18717
rect 17604 18680 17632 18711
rect 16224 18652 16896 18680
rect 17512 18652 17632 18680
rect 18524 18680 18552 18711
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18748 19855 18751
rect 20162 18748 20168 18760
rect 19843 18720 20168 18748
rect 19843 18717 19855 18720
rect 19797 18711 19855 18717
rect 20162 18708 20168 18720
rect 20220 18708 20226 18760
rect 22186 18708 22192 18760
rect 22244 18708 22250 18760
rect 22373 18751 22431 18757
rect 22373 18717 22385 18751
rect 22419 18717 22431 18751
rect 22373 18711 22431 18717
rect 22833 18751 22891 18757
rect 22833 18717 22845 18751
rect 22879 18748 22891 18751
rect 23201 18751 23259 18757
rect 23201 18748 23213 18751
rect 22879 18720 23213 18748
rect 22879 18717 22891 18720
rect 22833 18711 22891 18717
rect 23201 18717 23213 18720
rect 23247 18748 23259 18751
rect 23566 18748 23572 18760
rect 23247 18720 23572 18748
rect 23247 18717 23259 18720
rect 23201 18711 23259 18717
rect 22388 18680 22416 18711
rect 23566 18708 23572 18720
rect 23624 18708 23630 18760
rect 23658 18708 23664 18760
rect 23716 18748 23722 18760
rect 23952 18757 23980 18788
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 23716 18720 23765 18748
rect 23716 18708 23722 18720
rect 23753 18717 23765 18720
rect 23799 18717 23811 18751
rect 23753 18711 23811 18717
rect 23937 18751 23995 18757
rect 23937 18717 23949 18751
rect 23983 18717 23995 18751
rect 23937 18711 23995 18717
rect 24210 18708 24216 18760
rect 24268 18708 24274 18760
rect 24596 18757 24624 18856
rect 25133 18819 25191 18825
rect 25133 18816 25145 18819
rect 24688 18788 25145 18816
rect 24688 18760 24716 18788
rect 25133 18785 25145 18788
rect 25179 18785 25191 18819
rect 25133 18779 25191 18785
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24670 18708 24676 18760
rect 24728 18708 24734 18760
rect 25038 18708 25044 18760
rect 25096 18708 25102 18760
rect 25240 18748 25268 18856
rect 27246 18844 27252 18896
rect 27304 18844 27310 18896
rect 29196 18884 29224 18924
rect 29273 18921 29285 18955
rect 29319 18952 29331 18955
rect 29546 18952 29552 18964
rect 29319 18924 29552 18952
rect 29319 18921 29331 18924
rect 29273 18915 29331 18921
rect 29546 18912 29552 18924
rect 29604 18912 29610 18964
rect 33505 18955 33563 18961
rect 33505 18921 33517 18955
rect 33551 18952 33563 18955
rect 33778 18952 33784 18964
rect 33551 18924 33784 18952
rect 33551 18921 33563 18924
rect 33505 18915 33563 18921
rect 33778 18912 33784 18924
rect 33836 18912 33842 18964
rect 33870 18912 33876 18964
rect 33928 18952 33934 18964
rect 35345 18955 35403 18961
rect 33928 18924 35296 18952
rect 33928 18912 33934 18924
rect 29196 18856 29408 18884
rect 27264 18816 27292 18844
rect 26896 18788 27292 18816
rect 27525 18819 27583 18825
rect 25317 18751 25375 18757
rect 25317 18748 25329 18751
rect 25240 18720 25329 18748
rect 25317 18717 25329 18720
rect 25363 18717 25375 18751
rect 25317 18711 25375 18717
rect 23845 18683 23903 18689
rect 23845 18680 23857 18683
rect 18524 18652 19104 18680
rect 15304 18612 15332 18640
rect 17512 18624 17540 18652
rect 19076 18624 19104 18652
rect 22066 18652 22416 18680
rect 22664 18652 23857 18680
rect 14292 18584 15332 18612
rect 15470 18572 15476 18624
rect 15528 18612 15534 18624
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 15528 18584 15577 18612
rect 15528 18572 15534 18584
rect 15565 18581 15577 18584
rect 15611 18581 15623 18615
rect 15565 18575 15623 18581
rect 16301 18615 16359 18621
rect 16301 18581 16313 18615
rect 16347 18612 16359 18615
rect 17494 18612 17500 18624
rect 16347 18584 17500 18612
rect 16347 18581 16359 18584
rect 16301 18575 16359 18581
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 17770 18572 17776 18624
rect 17828 18572 17834 18624
rect 18046 18572 18052 18624
rect 18104 18612 18110 18624
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 18104 18584 18337 18612
rect 18104 18572 18110 18584
rect 18325 18581 18337 18584
rect 18371 18581 18383 18615
rect 18325 18575 18383 18581
rect 19058 18572 19064 18624
rect 19116 18612 19122 18624
rect 21358 18612 21364 18624
rect 19116 18584 21364 18612
rect 19116 18572 19122 18584
rect 21358 18572 21364 18584
rect 21416 18612 21422 18624
rect 22066 18612 22094 18652
rect 22664 18624 22692 18652
rect 23845 18649 23857 18652
rect 23891 18649 23903 18683
rect 23845 18643 23903 18649
rect 24075 18683 24133 18689
rect 24075 18649 24087 18683
rect 24121 18680 24133 18683
rect 24486 18680 24492 18692
rect 24121 18652 24492 18680
rect 24121 18649 24133 18652
rect 24075 18643 24133 18649
rect 24486 18640 24492 18652
rect 24544 18640 24550 18692
rect 24765 18683 24823 18689
rect 24765 18649 24777 18683
rect 24811 18649 24823 18683
rect 24765 18643 24823 18649
rect 24903 18683 24961 18689
rect 24903 18649 24915 18683
rect 24949 18680 24961 18683
rect 25222 18680 25228 18692
rect 24949 18652 25228 18680
rect 24949 18649 24961 18652
rect 24903 18643 24961 18649
rect 21416 18584 22094 18612
rect 22373 18615 22431 18621
rect 21416 18572 21422 18584
rect 22373 18581 22385 18615
rect 22419 18612 22431 18615
rect 22646 18612 22652 18624
rect 22419 18584 22652 18612
rect 22419 18581 22431 18584
rect 22373 18575 22431 18581
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 23290 18572 23296 18624
rect 23348 18572 23354 18624
rect 23566 18572 23572 18624
rect 23624 18572 23630 18624
rect 24302 18572 24308 18624
rect 24360 18612 24366 18624
rect 24397 18615 24455 18621
rect 24397 18612 24409 18615
rect 24360 18584 24409 18612
rect 24360 18572 24366 18584
rect 24397 18581 24409 18584
rect 24443 18581 24455 18615
rect 24780 18612 24808 18643
rect 25222 18640 25228 18652
rect 25280 18640 25286 18692
rect 26896 18680 26924 18788
rect 27525 18785 27537 18819
rect 27571 18816 27583 18819
rect 29270 18816 29276 18828
rect 27571 18788 29276 18816
rect 27571 18785 27583 18788
rect 27525 18779 27583 18785
rect 29270 18776 29276 18788
rect 29328 18776 29334 18828
rect 26970 18708 26976 18760
rect 27028 18748 27034 18760
rect 27433 18751 27491 18757
rect 27433 18748 27445 18751
rect 27028 18720 27445 18748
rect 27028 18708 27034 18720
rect 27433 18717 27445 18720
rect 27479 18717 27491 18751
rect 29380 18748 29408 18856
rect 30193 18819 30251 18825
rect 30193 18785 30205 18819
rect 30239 18816 30251 18819
rect 30282 18816 30288 18828
rect 30239 18788 30288 18816
rect 30239 18785 30251 18788
rect 30193 18779 30251 18785
rect 30282 18776 30288 18788
rect 30340 18776 30346 18828
rect 33226 18776 33232 18828
rect 33284 18776 33290 18828
rect 33597 18819 33655 18825
rect 33597 18785 33609 18819
rect 33643 18816 33655 18819
rect 33643 18788 34376 18816
rect 33643 18785 33655 18788
rect 33597 18779 33655 18785
rect 29917 18751 29975 18757
rect 29917 18748 29929 18751
rect 29380 18720 29929 18748
rect 27433 18711 27491 18717
rect 29917 18717 29929 18720
rect 29963 18748 29975 18751
rect 30374 18748 30380 18760
rect 29963 18720 30380 18748
rect 29963 18717 29975 18720
rect 29917 18711 29975 18717
rect 30374 18708 30380 18720
rect 30432 18708 30438 18760
rect 31297 18751 31355 18757
rect 31297 18717 31309 18751
rect 31343 18748 31355 18751
rect 31478 18748 31484 18760
rect 31343 18720 31484 18748
rect 31343 18717 31355 18720
rect 31297 18711 31355 18717
rect 31478 18708 31484 18720
rect 31536 18708 31542 18760
rect 32033 18751 32091 18757
rect 32033 18717 32045 18751
rect 32079 18748 32091 18751
rect 32079 18720 32113 18748
rect 32079 18717 32091 18720
rect 32033 18711 32091 18717
rect 27801 18683 27859 18689
rect 27801 18680 27813 18683
rect 25332 18652 26924 18680
rect 27264 18652 27813 18680
rect 25332 18612 25360 18652
rect 24780 18584 25360 18612
rect 25501 18615 25559 18621
rect 24397 18575 24455 18581
rect 25501 18581 25513 18615
rect 25547 18612 25559 18615
rect 27154 18612 27160 18624
rect 25547 18584 27160 18612
rect 25547 18581 25559 18584
rect 25501 18575 25559 18581
rect 27154 18572 27160 18584
rect 27212 18572 27218 18624
rect 27264 18621 27292 18652
rect 27801 18649 27813 18652
rect 27847 18649 27859 18683
rect 27801 18643 27859 18649
rect 28534 18640 28540 18692
rect 28592 18640 28598 18692
rect 32048 18680 32076 18711
rect 32214 18708 32220 18760
rect 32272 18708 32278 18760
rect 33134 18708 33140 18760
rect 33192 18708 33198 18760
rect 33612 18680 33640 18779
rect 34348 18760 34376 18788
rect 33778 18708 33784 18760
rect 33836 18708 33842 18760
rect 33962 18708 33968 18760
rect 34020 18708 34026 18760
rect 34330 18708 34336 18760
rect 34388 18708 34394 18760
rect 35268 18757 35296 18924
rect 35345 18921 35357 18955
rect 35391 18952 35403 18955
rect 35802 18952 35808 18964
rect 35391 18924 35808 18952
rect 35391 18921 35403 18924
rect 35345 18915 35403 18921
rect 35802 18912 35808 18924
rect 35860 18912 35866 18964
rect 36633 18955 36691 18961
rect 36633 18921 36645 18955
rect 36679 18952 36691 18955
rect 37642 18952 37648 18964
rect 36679 18924 37648 18952
rect 36679 18921 36691 18924
rect 36633 18915 36691 18921
rect 37642 18912 37648 18924
rect 37700 18912 37706 18964
rect 38562 18912 38568 18964
rect 38620 18952 38626 18964
rect 38620 18924 39528 18952
rect 38620 18912 38626 18924
rect 38841 18887 38899 18893
rect 38841 18853 38853 18887
rect 38887 18853 38899 18887
rect 38841 18847 38899 18853
rect 37277 18819 37335 18825
rect 37277 18785 37289 18819
rect 37323 18816 37335 18819
rect 37366 18816 37372 18828
rect 37323 18788 37372 18816
rect 37323 18785 37335 18788
rect 37277 18779 37335 18785
rect 37366 18776 37372 18788
rect 37424 18776 37430 18828
rect 35253 18751 35311 18757
rect 35253 18717 35265 18751
rect 35299 18717 35311 18751
rect 35253 18711 35311 18717
rect 35437 18751 35495 18757
rect 35437 18717 35449 18751
rect 35483 18748 35495 18751
rect 36078 18748 36084 18760
rect 35483 18720 36084 18748
rect 35483 18717 35495 18720
rect 35437 18711 35495 18717
rect 36078 18708 36084 18720
rect 36136 18708 36142 18760
rect 36814 18708 36820 18760
rect 36872 18708 36878 18760
rect 38856 18748 38884 18847
rect 39500 18825 39528 18924
rect 39485 18819 39543 18825
rect 39485 18785 39497 18819
rect 39531 18816 39543 18819
rect 39666 18816 39672 18828
rect 39531 18788 39672 18816
rect 39531 18785 39543 18788
rect 39485 18779 39543 18785
rect 39666 18776 39672 18788
rect 39724 18776 39730 18828
rect 40037 18751 40095 18757
rect 40037 18748 40049 18751
rect 38856 18720 40049 18748
rect 40037 18717 40049 18720
rect 40083 18717 40095 18751
rect 40037 18711 40095 18717
rect 31404 18652 33640 18680
rect 33888 18652 36676 18680
rect 27249 18615 27307 18621
rect 27249 18581 27261 18615
rect 27295 18581 27307 18615
rect 27249 18575 27307 18581
rect 29546 18572 29552 18624
rect 29604 18572 29610 18624
rect 29638 18572 29644 18624
rect 29696 18612 29702 18624
rect 30009 18615 30067 18621
rect 30009 18612 30021 18615
rect 29696 18584 30021 18612
rect 29696 18572 29702 18584
rect 30009 18581 30021 18584
rect 30055 18581 30067 18615
rect 30009 18575 30067 18581
rect 30650 18572 30656 18624
rect 30708 18612 30714 18624
rect 31404 18612 31432 18652
rect 30708 18584 31432 18612
rect 31573 18615 31631 18621
rect 30708 18572 30714 18584
rect 31573 18581 31585 18615
rect 31619 18612 31631 18615
rect 31938 18612 31944 18624
rect 31619 18584 31944 18612
rect 31619 18581 31631 18584
rect 31573 18575 31631 18581
rect 31938 18572 31944 18584
rect 31996 18572 32002 18624
rect 32030 18572 32036 18624
rect 32088 18572 32094 18624
rect 33318 18572 33324 18624
rect 33376 18612 33382 18624
rect 33888 18612 33916 18652
rect 33376 18584 33916 18612
rect 33376 18572 33382 18584
rect 34146 18572 34152 18624
rect 34204 18612 34210 18624
rect 35986 18612 35992 18624
rect 34204 18584 35992 18612
rect 34204 18572 34210 18584
rect 35986 18572 35992 18584
rect 36044 18572 36050 18624
rect 36648 18612 36676 18652
rect 36722 18640 36728 18692
rect 36780 18680 36786 18692
rect 36909 18683 36967 18689
rect 36909 18680 36921 18683
rect 36780 18652 36921 18680
rect 36780 18640 36786 18652
rect 36909 18649 36921 18652
rect 36955 18649 36967 18683
rect 36909 18643 36967 18649
rect 37001 18683 37059 18689
rect 37001 18649 37013 18683
rect 37047 18649 37059 18683
rect 37001 18643 37059 18649
rect 37016 18612 37044 18643
rect 37090 18640 37096 18692
rect 37148 18689 37154 18692
rect 37148 18683 37177 18689
rect 37165 18649 37177 18683
rect 37148 18643 37177 18649
rect 37148 18640 37154 18643
rect 39298 18640 39304 18692
rect 39356 18680 39362 18692
rect 39356 18652 41000 18680
rect 39356 18640 39362 18652
rect 40972 18624 41000 18652
rect 36648 18584 37044 18612
rect 38746 18572 38752 18624
rect 38804 18612 38810 18624
rect 39209 18615 39267 18621
rect 39209 18612 39221 18615
rect 38804 18584 39221 18612
rect 38804 18572 38810 18584
rect 39209 18581 39221 18584
rect 39255 18581 39267 18615
rect 39209 18575 39267 18581
rect 39850 18572 39856 18624
rect 39908 18572 39914 18624
rect 40954 18572 40960 18624
rect 41012 18572 41018 18624
rect 1104 18522 41400 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 41400 18522
rect 1104 18448 41400 18470
rect 1486 18368 1492 18420
rect 1544 18408 1550 18420
rect 3145 18411 3203 18417
rect 3145 18408 3157 18411
rect 1544 18380 3157 18408
rect 1544 18368 1550 18380
rect 3145 18377 3157 18380
rect 3191 18377 3203 18411
rect 3145 18371 3203 18377
rect 4062 18368 4068 18420
rect 4120 18368 4126 18420
rect 4982 18368 4988 18420
rect 5040 18368 5046 18420
rect 5166 18368 5172 18420
rect 5224 18368 5230 18420
rect 5534 18408 5540 18420
rect 5368 18380 5540 18408
rect 3050 18340 3056 18352
rect 2898 18312 3056 18340
rect 3050 18300 3056 18312
rect 3108 18340 3114 18352
rect 4080 18340 4108 18368
rect 5000 18340 5028 18368
rect 3108 18312 4108 18340
rect 4724 18312 5028 18340
rect 3108 18300 3114 18312
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 4724 18281 4752 18312
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 4982 18232 4988 18284
rect 5040 18272 5046 18284
rect 5184 18272 5212 18368
rect 5368 18281 5396 18380
rect 5534 18368 5540 18380
rect 5592 18408 5598 18420
rect 5813 18411 5871 18417
rect 5592 18380 5764 18408
rect 5592 18368 5598 18380
rect 5442 18300 5448 18352
rect 5500 18300 5506 18352
rect 5645 18343 5703 18349
rect 5645 18340 5657 18343
rect 5552 18312 5657 18340
rect 5040 18244 5212 18272
rect 5353 18275 5411 18281
rect 5040 18232 5046 18244
rect 5353 18241 5365 18275
rect 5399 18241 5411 18275
rect 5353 18235 5411 18241
rect 5552 18216 5580 18312
rect 5645 18309 5657 18312
rect 5691 18309 5703 18343
rect 5645 18303 5703 18309
rect 5736 18272 5764 18380
rect 5813 18377 5825 18411
rect 5859 18408 5871 18411
rect 5994 18408 6000 18420
rect 5859 18380 6000 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 7193 18411 7251 18417
rect 7193 18377 7205 18411
rect 7239 18408 7251 18411
rect 7926 18408 7932 18420
rect 7239 18380 7932 18408
rect 7239 18377 7251 18380
rect 7193 18371 7251 18377
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 8018 18368 8024 18420
rect 8076 18408 8082 18420
rect 11238 18408 11244 18420
rect 8076 18380 11244 18408
rect 8076 18368 8082 18380
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 11974 18368 11980 18420
rect 12032 18368 12038 18420
rect 12621 18411 12679 18417
rect 12621 18408 12633 18411
rect 12176 18380 12633 18408
rect 7374 18340 7380 18352
rect 7116 18312 7380 18340
rect 7116 18281 7144 18312
rect 7374 18300 7380 18312
rect 7432 18300 7438 18352
rect 11054 18300 11060 18352
rect 11112 18340 11118 18352
rect 11112 18312 11560 18340
rect 11112 18300 11118 18312
rect 7101 18275 7159 18281
rect 7101 18272 7113 18275
rect 5736 18244 7113 18272
rect 7101 18241 7113 18244
rect 7147 18241 7159 18275
rect 7101 18235 7159 18241
rect 7190 18232 7196 18284
rect 7248 18272 7254 18284
rect 7285 18275 7343 18281
rect 7285 18272 7297 18275
rect 7248 18244 7297 18272
rect 7248 18232 7254 18244
rect 7285 18241 7297 18244
rect 7331 18241 7343 18275
rect 7285 18235 7343 18241
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 9122 18272 9128 18284
rect 8444 18244 9128 18272
rect 8444 18232 8450 18244
rect 9122 18232 9128 18244
rect 9180 18272 9186 18284
rect 9582 18272 9588 18284
rect 9180 18244 9588 18272
rect 9180 18232 9186 18244
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 10502 18232 10508 18284
rect 10560 18232 10566 18284
rect 10965 18275 11023 18281
rect 10965 18241 10977 18275
rect 11011 18272 11023 18275
rect 11330 18272 11336 18284
rect 11011 18244 11336 18272
rect 11011 18241 11023 18244
rect 10965 18235 11023 18241
rect 11330 18232 11336 18244
rect 11388 18232 11394 18284
rect 11532 18281 11560 18312
rect 12176 18281 12204 18380
rect 12621 18377 12633 18380
rect 12667 18377 12679 18411
rect 12621 18371 12679 18377
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 14700 18380 14872 18408
rect 14700 18368 14706 18380
rect 14844 18349 14872 18380
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 22925 18411 22983 18417
rect 22925 18408 22937 18411
rect 15528 18380 18460 18408
rect 15528 18368 15534 18380
rect 14829 18343 14887 18349
rect 12360 18312 12756 18340
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 12161 18275 12219 18281
rect 12161 18241 12173 18275
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 12360 18281 12388 18312
rect 12345 18275 12403 18281
rect 12345 18272 12357 18275
rect 12308 18244 12357 18272
rect 12308 18232 12314 18244
rect 12345 18241 12357 18244
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12434 18232 12440 18284
rect 12492 18232 12498 18284
rect 12728 18281 12756 18312
rect 14829 18309 14841 18343
rect 14875 18309 14887 18343
rect 15378 18340 15384 18352
rect 14829 18303 14887 18309
rect 15028 18312 15384 18340
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18241 12771 18275
rect 12713 18235 12771 18241
rect 1670 18164 1676 18216
rect 1728 18164 1734 18216
rect 5077 18207 5135 18213
rect 5077 18173 5089 18207
rect 5123 18204 5135 18207
rect 5534 18204 5540 18216
rect 5123 18176 5540 18204
rect 5123 18173 5135 18176
rect 5077 18167 5135 18173
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 7926 18096 7932 18148
rect 7984 18136 7990 18148
rect 10520 18136 10548 18232
rect 10594 18164 10600 18216
rect 10652 18164 10658 18216
rect 12158 18136 12164 18148
rect 7984 18108 8432 18136
rect 10520 18108 12164 18136
rect 7984 18096 7990 18108
rect 4522 18028 4528 18080
rect 4580 18068 4586 18080
rect 4798 18068 4804 18080
rect 4580 18040 4804 18068
rect 4580 18028 4586 18040
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 5350 18028 5356 18080
rect 5408 18068 5414 18080
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5408 18040 5641 18068
rect 5408 18028 5414 18040
rect 5629 18037 5641 18040
rect 5675 18037 5687 18071
rect 5629 18031 5687 18037
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 8294 18068 8300 18080
rect 7340 18040 8300 18068
rect 7340 18028 7346 18040
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 8404 18068 8432 18108
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 8404 18040 11161 18068
rect 11149 18037 11161 18040
rect 11195 18037 11207 18071
rect 11149 18031 11207 18037
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 11701 18071 11759 18077
rect 11701 18068 11713 18071
rect 11388 18040 11713 18068
rect 11388 18028 11394 18040
rect 11701 18037 11713 18040
rect 11747 18037 11759 18071
rect 12544 18068 12572 18235
rect 14366 18232 14372 18284
rect 14424 18272 14430 18284
rect 15028 18272 15056 18312
rect 15378 18300 15384 18312
rect 15436 18340 15442 18352
rect 15436 18312 15792 18340
rect 15436 18300 15442 18312
rect 14424 18244 15056 18272
rect 14424 18232 14430 18244
rect 15286 18232 15292 18284
rect 15344 18232 15350 18284
rect 15562 18232 15568 18284
rect 15620 18232 15626 18284
rect 15764 18281 15792 18312
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16632 18244 16681 18272
rect 16632 18232 16638 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 16816 18244 17049 18272
rect 16816 18232 16822 18244
rect 17037 18241 17049 18244
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 17678 18232 17684 18284
rect 17736 18232 17742 18284
rect 17770 18232 17776 18284
rect 17828 18232 17834 18284
rect 18230 18232 18236 18284
rect 18288 18232 18294 18284
rect 18432 18281 18460 18380
rect 18524 18380 22937 18408
rect 18524 18281 18552 18380
rect 22925 18377 22937 18380
rect 22971 18408 22983 18411
rect 23382 18408 23388 18420
rect 22971 18380 23388 18408
rect 22971 18377 22983 18380
rect 22925 18371 22983 18377
rect 23382 18368 23388 18380
rect 23440 18368 23446 18420
rect 24026 18368 24032 18420
rect 24084 18368 24090 18420
rect 24578 18368 24584 18420
rect 24636 18408 24642 18420
rect 24636 18380 27108 18408
rect 24636 18368 24642 18380
rect 23106 18340 23112 18352
rect 18708 18312 23112 18340
rect 18417 18275 18475 18281
rect 18417 18241 18429 18275
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 18509 18275 18567 18281
rect 18509 18241 18521 18275
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18616 18204 18644 18235
rect 15120 18176 18644 18204
rect 15120 18148 15148 18176
rect 15102 18096 15108 18148
rect 15160 18096 15166 18148
rect 15565 18139 15623 18145
rect 15565 18105 15577 18139
rect 15611 18136 15623 18139
rect 15746 18136 15752 18148
rect 15611 18108 15752 18136
rect 15611 18105 15623 18108
rect 15565 18099 15623 18105
rect 15746 18096 15752 18108
rect 15804 18096 15810 18148
rect 17126 18096 17132 18148
rect 17184 18136 17190 18148
rect 18049 18139 18107 18145
rect 18049 18136 18061 18139
rect 17184 18108 18061 18136
rect 17184 18096 17190 18108
rect 18049 18105 18061 18108
rect 18095 18105 18107 18139
rect 18049 18099 18107 18105
rect 18322 18096 18328 18148
rect 18380 18136 18386 18148
rect 18708 18136 18736 18312
rect 23106 18300 23112 18312
rect 23164 18300 23170 18352
rect 23216 18312 24256 18340
rect 18874 18232 18880 18284
rect 18932 18232 18938 18284
rect 19058 18232 19064 18284
rect 19116 18232 19122 18284
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 18892 18204 18920 18232
rect 19168 18204 19196 18235
rect 19242 18232 19248 18284
rect 19300 18232 19306 18284
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 19978 18272 19984 18284
rect 19484 18244 19984 18272
rect 19484 18232 19490 18244
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 20070 18232 20076 18284
rect 20128 18272 20134 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 20128 18244 20177 18272
rect 20128 18232 20134 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 18892 18176 19196 18204
rect 20180 18204 20208 18235
rect 20254 18232 20260 18284
rect 20312 18232 20318 18284
rect 20346 18232 20352 18284
rect 20404 18272 20410 18284
rect 20441 18275 20499 18281
rect 20441 18272 20453 18275
rect 20404 18244 20453 18272
rect 20404 18232 20410 18244
rect 20441 18241 20453 18244
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 20640 18204 20668 18235
rect 21542 18232 21548 18284
rect 21600 18232 21606 18284
rect 22278 18232 22284 18284
rect 22336 18272 22342 18284
rect 23014 18272 23020 18284
rect 22336 18244 23020 18272
rect 22336 18232 22342 18244
rect 23014 18232 23020 18244
rect 23072 18232 23078 18284
rect 20180 18176 20668 18204
rect 20809 18207 20867 18213
rect 20809 18173 20821 18207
rect 20855 18204 20867 18207
rect 21450 18204 21456 18216
rect 20855 18176 21456 18204
rect 20855 18173 20867 18176
rect 20809 18167 20867 18173
rect 21450 18164 21456 18176
rect 21508 18164 21514 18216
rect 18380 18108 18736 18136
rect 18877 18139 18935 18145
rect 18380 18096 18386 18108
rect 18877 18105 18889 18139
rect 18923 18136 18935 18139
rect 21560 18136 21588 18232
rect 22738 18164 22744 18216
rect 22796 18204 22802 18216
rect 23216 18204 23244 18312
rect 23290 18232 23296 18284
rect 23348 18232 23354 18284
rect 23566 18232 23572 18284
rect 23624 18272 23630 18284
rect 23753 18275 23811 18281
rect 23753 18272 23765 18275
rect 23624 18244 23765 18272
rect 23624 18232 23630 18244
rect 23753 18241 23765 18244
rect 23799 18241 23811 18275
rect 23753 18235 23811 18241
rect 24026 18232 24032 18284
rect 24084 18272 24090 18284
rect 24121 18275 24179 18281
rect 24121 18272 24133 18275
rect 24084 18244 24133 18272
rect 24084 18232 24090 18244
rect 24121 18241 24133 18244
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 22796 18176 23244 18204
rect 23308 18204 23336 18232
rect 24228 18213 24256 18312
rect 24302 18232 24308 18284
rect 24360 18232 24366 18284
rect 24394 18232 24400 18284
rect 24452 18232 24458 18284
rect 24578 18232 24584 18284
rect 24636 18272 24642 18284
rect 26878 18272 26884 18284
rect 24636 18244 26884 18272
rect 24636 18232 24642 18244
rect 26878 18232 26884 18244
rect 26936 18232 26942 18284
rect 27080 18281 27108 18380
rect 27154 18368 27160 18420
rect 27212 18408 27218 18420
rect 27798 18408 27804 18420
rect 27212 18380 27804 18408
rect 27212 18368 27218 18380
rect 27798 18368 27804 18380
rect 27856 18408 27862 18420
rect 29546 18408 29552 18420
rect 27856 18380 27936 18408
rect 27856 18368 27862 18380
rect 27908 18349 27936 18380
rect 29472 18380 29552 18408
rect 27893 18343 27951 18349
rect 27172 18312 27660 18340
rect 26973 18275 27031 18281
rect 26973 18241 26985 18275
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 27066 18275 27124 18281
rect 27066 18241 27078 18275
rect 27112 18241 27124 18275
rect 27066 18235 27124 18241
rect 23661 18207 23719 18213
rect 23661 18204 23673 18207
rect 23308 18176 23673 18204
rect 22796 18164 22802 18176
rect 23661 18173 23673 18176
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 24213 18207 24271 18213
rect 24213 18173 24225 18207
rect 24259 18173 24271 18207
rect 24213 18167 24271 18173
rect 22462 18136 22468 18148
rect 18923 18108 21588 18136
rect 22204 18108 22468 18136
rect 18923 18105 18935 18108
rect 18877 18099 18935 18105
rect 22204 18080 22232 18108
rect 22462 18096 22468 18108
rect 22520 18136 22526 18148
rect 22557 18139 22615 18145
rect 22557 18136 22569 18139
rect 22520 18108 22569 18136
rect 22520 18096 22526 18108
rect 22557 18105 22569 18108
rect 22603 18105 22615 18139
rect 22557 18099 22615 18105
rect 22649 18139 22707 18145
rect 22649 18105 22661 18139
rect 22695 18136 22707 18139
rect 23566 18136 23572 18148
rect 22695 18108 23572 18136
rect 22695 18105 22707 18108
rect 22649 18099 22707 18105
rect 23566 18096 23572 18108
rect 23624 18096 23630 18148
rect 15654 18068 15660 18080
rect 12544 18040 15660 18068
rect 11701 18031 11759 18037
rect 15654 18028 15660 18040
rect 15712 18028 15718 18080
rect 15930 18028 15936 18080
rect 15988 18028 15994 18080
rect 17034 18028 17040 18080
rect 17092 18068 17098 18080
rect 17402 18068 17408 18080
rect 17092 18040 17408 18068
rect 17092 18028 17098 18040
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 18782 18028 18788 18080
rect 18840 18028 18846 18080
rect 18966 18028 18972 18080
rect 19024 18068 19030 18080
rect 19429 18071 19487 18077
rect 19429 18068 19441 18071
rect 19024 18040 19441 18068
rect 19024 18028 19030 18040
rect 19429 18037 19441 18040
rect 19475 18037 19487 18071
rect 19429 18031 19487 18037
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20162 18068 20168 18080
rect 20036 18040 20168 18068
rect 20036 18028 20042 18040
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 20257 18071 20315 18077
rect 20257 18037 20269 18071
rect 20303 18068 20315 18071
rect 20346 18068 20352 18080
rect 20303 18040 20352 18068
rect 20303 18037 20315 18040
rect 20257 18031 20315 18037
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 22186 18028 22192 18080
rect 22244 18028 22250 18080
rect 22278 18028 22284 18080
rect 22336 18028 22342 18080
rect 22738 18028 22744 18080
rect 22796 18028 22802 18080
rect 23198 18028 23204 18080
rect 23256 18068 23262 18080
rect 23385 18071 23443 18077
rect 23385 18068 23397 18071
rect 23256 18040 23397 18068
rect 23256 18028 23262 18040
rect 23385 18037 23397 18040
rect 23431 18037 23443 18071
rect 23676 18068 23704 18167
rect 23845 18139 23903 18145
rect 23845 18105 23857 18139
rect 23891 18136 23903 18139
rect 24320 18136 24348 18232
rect 26988 18204 27016 18235
rect 27172 18204 27200 18312
rect 27249 18275 27307 18281
rect 27249 18241 27261 18275
rect 27295 18241 27307 18275
rect 27249 18235 27307 18241
rect 26988 18176 27200 18204
rect 23891 18108 24348 18136
rect 24581 18139 24639 18145
rect 23891 18105 23903 18108
rect 23845 18099 23903 18105
rect 24581 18105 24593 18139
rect 24627 18136 24639 18139
rect 24854 18136 24860 18148
rect 24627 18108 24860 18136
rect 24627 18105 24639 18108
rect 24581 18099 24639 18105
rect 24854 18096 24860 18108
rect 24912 18136 24918 18148
rect 27264 18136 27292 18235
rect 27338 18232 27344 18284
rect 27396 18232 27402 18284
rect 27522 18281 27528 18284
rect 27479 18275 27528 18281
rect 27479 18241 27491 18275
rect 27525 18241 27528 18275
rect 27479 18235 27528 18241
rect 27522 18232 27528 18235
rect 27580 18232 27586 18284
rect 27632 18204 27660 18312
rect 27893 18309 27905 18343
rect 27939 18309 27951 18343
rect 27893 18303 27951 18309
rect 27706 18232 27712 18284
rect 27764 18232 27770 18284
rect 27982 18232 27988 18284
rect 28040 18232 28046 18284
rect 28074 18232 28080 18284
rect 28132 18232 28138 18284
rect 27632 18176 28304 18204
rect 28276 18145 28304 18176
rect 28350 18164 28356 18216
rect 28408 18204 28414 18216
rect 29086 18204 29092 18216
rect 28408 18176 29092 18204
rect 28408 18164 28414 18176
rect 29086 18164 29092 18176
rect 29144 18164 29150 18216
rect 29472 18213 29500 18380
rect 29546 18368 29552 18380
rect 29604 18368 29610 18420
rect 29917 18411 29975 18417
rect 29917 18377 29929 18411
rect 29963 18408 29975 18411
rect 30190 18408 30196 18420
rect 29963 18380 30196 18408
rect 29963 18377 29975 18380
rect 29917 18371 29975 18377
rect 30190 18368 30196 18380
rect 30248 18368 30254 18420
rect 31573 18411 31631 18417
rect 31573 18377 31585 18411
rect 31619 18408 31631 18411
rect 32122 18408 32128 18420
rect 31619 18380 32128 18408
rect 31619 18377 31631 18380
rect 31573 18371 31631 18377
rect 32122 18368 32128 18380
rect 32180 18368 32186 18420
rect 33226 18368 33232 18420
rect 33284 18408 33290 18420
rect 33505 18411 33563 18417
rect 33505 18408 33517 18411
rect 33284 18380 33517 18408
rect 33284 18368 33290 18380
rect 33505 18377 33517 18380
rect 33551 18377 33563 18411
rect 33505 18371 33563 18377
rect 34149 18411 34207 18417
rect 34149 18377 34161 18411
rect 34195 18408 34207 18411
rect 34698 18408 34704 18420
rect 34195 18380 34704 18408
rect 34195 18377 34207 18380
rect 34149 18371 34207 18377
rect 34698 18368 34704 18380
rect 34756 18408 34762 18420
rect 34993 18411 35051 18417
rect 34993 18408 35005 18411
rect 34756 18380 35005 18408
rect 34756 18368 34762 18380
rect 34993 18377 35005 18380
rect 35039 18377 35051 18411
rect 34993 18371 35051 18377
rect 35161 18411 35219 18417
rect 35161 18377 35173 18411
rect 35207 18408 35219 18411
rect 35434 18408 35440 18420
rect 35207 18380 35440 18408
rect 35207 18377 35219 18380
rect 35161 18371 35219 18377
rect 35434 18368 35440 18380
rect 35492 18368 35498 18420
rect 36633 18411 36691 18417
rect 36633 18377 36645 18411
rect 36679 18408 36691 18411
rect 36722 18408 36728 18420
rect 36679 18380 36728 18408
rect 36679 18377 36691 18380
rect 36633 18371 36691 18377
rect 36722 18368 36728 18380
rect 36780 18368 36786 18420
rect 36814 18368 36820 18420
rect 36872 18408 36878 18420
rect 37093 18411 37151 18417
rect 37093 18408 37105 18411
rect 36872 18380 37105 18408
rect 36872 18368 36878 18380
rect 37093 18377 37105 18380
rect 37139 18377 37151 18411
rect 37093 18371 37151 18377
rect 37829 18411 37887 18417
rect 37829 18377 37841 18411
rect 37875 18408 37887 18411
rect 38749 18411 38807 18417
rect 38749 18408 38761 18411
rect 37875 18380 38761 18408
rect 37875 18377 37887 18380
rect 37829 18371 37887 18377
rect 38749 18377 38761 18380
rect 38795 18377 38807 18411
rect 39850 18408 39856 18420
rect 38749 18371 38807 18377
rect 39500 18380 39856 18408
rect 32214 18300 32220 18352
rect 32272 18300 32278 18352
rect 33137 18343 33195 18349
rect 33137 18309 33149 18343
rect 33183 18309 33195 18343
rect 33137 18303 33195 18309
rect 33353 18343 33411 18349
rect 33353 18309 33365 18343
rect 33399 18340 33411 18343
rect 33689 18343 33747 18349
rect 33689 18340 33701 18343
rect 33399 18312 33701 18340
rect 33399 18309 33411 18312
rect 33353 18303 33411 18309
rect 33689 18309 33701 18312
rect 33735 18309 33747 18343
rect 33689 18303 33747 18309
rect 29549 18275 29607 18281
rect 29549 18241 29561 18275
rect 29595 18272 29607 18275
rect 30650 18272 30656 18284
rect 29595 18244 30656 18272
rect 29595 18241 29607 18244
rect 29549 18235 29607 18241
rect 30650 18232 30656 18244
rect 30708 18232 30714 18284
rect 31478 18232 31484 18284
rect 31536 18232 31542 18284
rect 31665 18275 31723 18281
rect 31665 18241 31677 18275
rect 31711 18272 31723 18275
rect 31938 18272 31944 18284
rect 31711 18244 31944 18272
rect 31711 18241 31723 18244
rect 31665 18235 31723 18241
rect 31938 18232 31944 18244
rect 31996 18232 32002 18284
rect 33152 18272 33180 18303
rect 34606 18300 34612 18352
rect 34664 18340 34670 18352
rect 34793 18343 34851 18349
rect 34793 18340 34805 18343
rect 34664 18312 34805 18340
rect 34664 18300 34670 18312
rect 34793 18309 34805 18312
rect 34839 18309 34851 18343
rect 36909 18343 36967 18349
rect 36909 18340 36921 18343
rect 34793 18303 34851 18309
rect 36648 18312 36921 18340
rect 33060 18244 33180 18272
rect 29457 18207 29515 18213
rect 29457 18173 29469 18207
rect 29503 18173 29515 18207
rect 29457 18167 29515 18173
rect 24912 18108 27292 18136
rect 28261 18139 28319 18145
rect 24912 18096 24918 18108
rect 28261 18105 28273 18139
rect 28307 18105 28319 18139
rect 33060 18136 33088 18244
rect 33594 18232 33600 18284
rect 33652 18232 33658 18284
rect 33778 18232 33784 18284
rect 33836 18232 33842 18284
rect 33873 18275 33931 18281
rect 33873 18241 33885 18275
rect 33919 18241 33931 18275
rect 33873 18235 33931 18241
rect 33134 18164 33140 18216
rect 33192 18204 33198 18216
rect 33888 18204 33916 18235
rect 33192 18176 33916 18204
rect 33192 18164 33198 18176
rect 34146 18164 34152 18216
rect 34204 18164 34210 18216
rect 34624 18136 34652 18300
rect 36449 18275 36507 18281
rect 36449 18272 36461 18275
rect 35912 18244 36461 18272
rect 35912 18216 35940 18244
rect 36449 18241 36461 18244
rect 36495 18241 36507 18275
rect 36449 18235 36507 18241
rect 35894 18164 35900 18216
rect 35952 18164 35958 18216
rect 36464 18204 36492 18235
rect 36538 18232 36544 18284
rect 36596 18272 36602 18284
rect 36648 18281 36676 18312
rect 36909 18309 36921 18312
rect 36955 18309 36967 18343
rect 36909 18303 36967 18309
rect 38378 18300 38384 18352
rect 38436 18340 38442 18352
rect 39500 18349 39528 18380
rect 39850 18368 39856 18380
rect 39908 18368 39914 18420
rect 40954 18368 40960 18420
rect 41012 18368 41018 18420
rect 39485 18343 39543 18349
rect 38436 18312 39252 18340
rect 38436 18300 38442 18312
rect 36633 18275 36691 18281
rect 36633 18272 36645 18275
rect 36596 18244 36645 18272
rect 36596 18232 36602 18244
rect 36633 18241 36645 18244
rect 36679 18241 36691 18275
rect 36633 18235 36691 18241
rect 36725 18275 36783 18281
rect 36725 18241 36737 18275
rect 36771 18241 36783 18275
rect 36725 18235 36783 18241
rect 36740 18204 36768 18235
rect 37090 18232 37096 18284
rect 37148 18272 37154 18284
rect 37458 18272 37464 18284
rect 37148 18244 37464 18272
rect 37148 18232 37154 18244
rect 37458 18232 37464 18244
rect 37516 18232 37522 18284
rect 38746 18232 38752 18284
rect 38804 18232 38810 18284
rect 39224 18281 39252 18312
rect 39485 18309 39497 18343
rect 39531 18309 39543 18343
rect 39485 18303 39543 18309
rect 40034 18300 40040 18352
rect 40092 18300 40098 18352
rect 39209 18275 39267 18281
rect 39209 18241 39221 18275
rect 39255 18241 39267 18275
rect 39209 18235 39267 18241
rect 36464 18176 36768 18204
rect 37553 18207 37611 18213
rect 37553 18173 37565 18207
rect 37599 18204 37611 18207
rect 37826 18204 37832 18216
rect 37599 18176 37832 18204
rect 37599 18173 37611 18176
rect 37553 18167 37611 18173
rect 37826 18164 37832 18176
rect 37884 18164 37890 18216
rect 33060 18108 34652 18136
rect 38381 18139 38439 18145
rect 28261 18099 28319 18105
rect 38381 18105 38393 18139
rect 38427 18136 38439 18139
rect 38764 18136 38792 18232
rect 38838 18164 38844 18216
rect 38896 18164 38902 18216
rect 39025 18207 39083 18213
rect 39025 18173 39037 18207
rect 39071 18204 39083 18207
rect 39114 18204 39120 18216
rect 39071 18176 39120 18204
rect 39071 18173 39083 18176
rect 39025 18167 39083 18173
rect 39114 18164 39120 18176
rect 39172 18164 39178 18216
rect 38427 18108 38792 18136
rect 38427 18105 38439 18108
rect 38381 18099 38439 18105
rect 26878 18068 26884 18080
rect 23676 18040 26884 18068
rect 23385 18031 23443 18037
rect 26878 18028 26884 18040
rect 26936 18068 26942 18080
rect 27246 18068 27252 18080
rect 26936 18040 27252 18068
rect 26936 18028 26942 18040
rect 27246 18028 27252 18040
rect 27304 18028 27310 18080
rect 27617 18071 27675 18077
rect 27617 18037 27629 18071
rect 27663 18068 27675 18071
rect 27706 18068 27712 18080
rect 27663 18040 27712 18068
rect 27663 18037 27675 18040
rect 27617 18031 27675 18037
rect 27706 18028 27712 18040
rect 27764 18028 27770 18080
rect 30006 18028 30012 18080
rect 30064 18068 30070 18080
rect 30282 18068 30288 18080
rect 30064 18040 30288 18068
rect 30064 18028 30070 18040
rect 30282 18028 30288 18040
rect 30340 18068 30346 18080
rect 32309 18071 32367 18077
rect 32309 18068 32321 18071
rect 30340 18040 32321 18068
rect 30340 18028 30346 18040
rect 32309 18037 32321 18040
rect 32355 18068 32367 18071
rect 33226 18068 33232 18080
rect 32355 18040 33232 18068
rect 32355 18037 32367 18040
rect 32309 18031 32367 18037
rect 33226 18028 33232 18040
rect 33284 18028 33290 18080
rect 33318 18028 33324 18080
rect 33376 18028 33382 18080
rect 33502 18028 33508 18080
rect 33560 18068 33566 18080
rect 33778 18068 33784 18080
rect 33560 18040 33784 18068
rect 33560 18028 33566 18040
rect 33778 18028 33784 18040
rect 33836 18068 33842 18080
rect 33965 18071 34023 18077
rect 33965 18068 33977 18071
rect 33836 18040 33977 18068
rect 33836 18028 33842 18040
rect 33965 18037 33977 18040
rect 34011 18037 34023 18071
rect 33965 18031 34023 18037
rect 34514 18028 34520 18080
rect 34572 18068 34578 18080
rect 34977 18071 35035 18077
rect 34977 18068 34989 18071
rect 34572 18040 34989 18068
rect 34572 18028 34578 18040
rect 34977 18037 34989 18040
rect 35023 18037 35035 18071
rect 34977 18031 35035 18037
rect 1104 17978 41400 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 41400 17978
rect 1104 17904 41400 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2685 17867 2743 17873
rect 2685 17864 2697 17867
rect 1728 17836 2697 17864
rect 1728 17824 1734 17836
rect 2685 17833 2697 17836
rect 2731 17833 2743 17867
rect 2685 17827 2743 17833
rect 9401 17867 9459 17873
rect 9401 17833 9413 17867
rect 9447 17864 9459 17867
rect 9490 17864 9496 17876
rect 9447 17836 9496 17864
rect 9447 17833 9459 17836
rect 9401 17827 9459 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 10134 17824 10140 17876
rect 10192 17824 10198 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 12805 17867 12863 17873
rect 12805 17864 12817 17867
rect 12492 17836 12817 17864
rect 12492 17824 12498 17836
rect 12805 17833 12817 17836
rect 12851 17833 12863 17867
rect 12805 17827 12863 17833
rect 15654 17824 15660 17876
rect 15712 17864 15718 17876
rect 22373 17867 22431 17873
rect 15712 17836 22094 17864
rect 15712 17824 15718 17836
rect 4062 17756 4068 17808
rect 4120 17796 4126 17808
rect 4249 17799 4307 17805
rect 4249 17796 4261 17799
rect 4120 17768 4261 17796
rect 4120 17756 4126 17768
rect 4249 17765 4261 17768
rect 4295 17765 4307 17799
rect 11514 17796 11520 17808
rect 4249 17759 4307 17765
rect 4632 17768 11520 17796
rect 1486 17688 1492 17740
rect 1544 17728 1550 17740
rect 1949 17731 2007 17737
rect 1949 17728 1961 17731
rect 1544 17700 1961 17728
rect 1544 17688 1550 17700
rect 1949 17697 1961 17700
rect 1995 17697 2007 17731
rect 4632 17728 4660 17768
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 12066 17756 12072 17808
rect 12124 17796 12130 17808
rect 13354 17796 13360 17808
rect 12124 17768 13360 17796
rect 12124 17756 12130 17768
rect 13354 17756 13360 17768
rect 13412 17756 13418 17808
rect 22066 17796 22094 17836
rect 22373 17833 22385 17867
rect 22419 17864 22431 17867
rect 22738 17864 22744 17876
rect 22419 17836 22744 17864
rect 22419 17833 22431 17836
rect 22373 17827 22431 17833
rect 22738 17824 22744 17836
rect 22796 17824 22802 17876
rect 23014 17824 23020 17876
rect 23072 17864 23078 17876
rect 24026 17864 24032 17876
rect 23072 17836 24032 17864
rect 23072 17824 23078 17836
rect 24026 17824 24032 17836
rect 24084 17824 24090 17876
rect 26050 17824 26056 17876
rect 26108 17864 26114 17876
rect 27430 17864 27436 17876
rect 26108 17836 27436 17864
rect 26108 17824 26114 17836
rect 27430 17824 27436 17836
rect 27488 17864 27494 17876
rect 30929 17867 30987 17873
rect 27488 17836 30880 17864
rect 27488 17824 27494 17836
rect 30852 17796 30880 17836
rect 30929 17833 30941 17867
rect 30975 17864 30987 17867
rect 31478 17864 31484 17876
rect 30975 17836 31484 17864
rect 30975 17833 30987 17836
rect 30929 17827 30987 17833
rect 31478 17824 31484 17836
rect 31536 17824 31542 17876
rect 33870 17824 33876 17876
rect 33928 17824 33934 17876
rect 35529 17867 35587 17873
rect 35529 17833 35541 17867
rect 35575 17864 35587 17867
rect 35894 17864 35900 17876
rect 35575 17836 35900 17864
rect 35575 17833 35587 17836
rect 35529 17827 35587 17833
rect 35894 17824 35900 17836
rect 35952 17864 35958 17876
rect 35952 17836 37136 17864
rect 35952 17824 35958 17836
rect 33888 17796 33916 17824
rect 13464 17768 21980 17796
rect 22066 17768 28994 17796
rect 30852 17768 33916 17796
rect 36817 17799 36875 17805
rect 5442 17728 5448 17740
rect 1949 17691 2007 17697
rect 2884 17700 4660 17728
rect 4724 17700 5448 17728
rect 2884 17669 2912 17700
rect 4724 17672 4752 17700
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 9582 17728 9588 17740
rect 9324 17700 9588 17728
rect 9324 17672 9352 17700
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 11790 17728 11796 17740
rect 10244 17700 11796 17728
rect 2869 17663 2927 17669
rect 2869 17629 2881 17663
rect 2915 17629 2927 17663
rect 2869 17623 2927 17629
rect 2958 17620 2964 17672
rect 3016 17660 3022 17672
rect 3145 17663 3203 17669
rect 3145 17660 3157 17663
rect 3016 17632 3157 17660
rect 3016 17620 3022 17632
rect 3145 17629 3157 17632
rect 3191 17629 3203 17663
rect 3145 17623 3203 17629
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 2593 17595 2651 17601
rect 2593 17561 2605 17595
rect 2639 17592 2651 17595
rect 3053 17595 3111 17601
rect 3053 17592 3065 17595
rect 2639 17564 3065 17592
rect 2639 17561 2651 17564
rect 2593 17555 2651 17561
rect 3053 17561 3065 17564
rect 3099 17561 3111 17595
rect 4448 17592 4476 17623
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 5350 17620 5356 17672
rect 5408 17620 5414 17672
rect 5534 17620 5540 17672
rect 5592 17620 5598 17672
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 9306 17620 9312 17672
rect 9364 17620 9370 17672
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17629 9551 17663
rect 9493 17623 9551 17629
rect 9508 17592 9536 17623
rect 10042 17620 10048 17672
rect 10100 17620 10106 17672
rect 10244 17669 10272 17700
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 12986 17688 12992 17740
rect 13044 17688 13050 17740
rect 13464 17737 13492 17768
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17697 13507 17731
rect 14550 17728 14556 17740
rect 13449 17691 13507 17697
rect 14108 17700 14556 17728
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 4448 17564 5580 17592
rect 3053 17555 3111 17561
rect 5552 17536 5580 17564
rect 9048 17564 9536 17592
rect 9048 17536 9076 17564
rect 10134 17552 10140 17604
rect 10192 17592 10198 17604
rect 11149 17595 11207 17601
rect 11149 17592 11161 17595
rect 10192 17564 11161 17592
rect 10192 17552 10198 17564
rect 11149 17561 11161 17564
rect 11195 17561 11207 17595
rect 11348 17592 11376 17623
rect 11606 17620 11612 17672
rect 11664 17620 11670 17672
rect 11698 17620 11704 17672
rect 11756 17620 11762 17672
rect 11885 17663 11943 17669
rect 11885 17629 11897 17663
rect 11931 17660 11943 17663
rect 12250 17660 12256 17672
rect 11931 17632 12256 17660
rect 11931 17629 11943 17632
rect 11885 17623 11943 17629
rect 11793 17595 11851 17601
rect 11793 17592 11805 17595
rect 11348 17564 11805 17592
rect 11149 17555 11207 17561
rect 11793 17561 11805 17564
rect 11839 17561 11851 17595
rect 11793 17555 11851 17561
rect 5534 17484 5540 17536
rect 5592 17484 5598 17536
rect 9030 17484 9036 17536
rect 9088 17484 9094 17536
rect 11517 17527 11575 17533
rect 11517 17493 11529 17527
rect 11563 17524 11575 17527
rect 11900 17524 11928 17623
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 13004 17660 13032 17688
rect 13633 17663 13691 17669
rect 13633 17660 13645 17663
rect 13004 17632 13645 17660
rect 13633 17629 13645 17632
rect 13679 17629 13691 17663
rect 13633 17623 13691 17629
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14108 17669 14136 17700
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 15562 17728 15568 17740
rect 14660 17700 15568 17728
rect 14660 17669 14688 17700
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 18782 17728 18788 17740
rect 18248 17700 18788 17728
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13872 17632 14105 17660
rect 13872 17620 13878 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 15102 17620 15108 17672
rect 15160 17660 15166 17672
rect 15286 17660 15292 17672
rect 15160 17632 15292 17660
rect 15160 17620 15166 17632
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 15378 17620 15384 17672
rect 15436 17620 15442 17672
rect 18248 17669 18276 17700
rect 18782 17688 18788 17700
rect 18840 17688 18846 17740
rect 19978 17688 19984 17740
rect 20036 17728 20042 17740
rect 20073 17731 20131 17737
rect 20073 17728 20085 17731
rect 20036 17700 20085 17728
rect 20036 17688 20042 17700
rect 20073 17697 20085 17700
rect 20119 17697 20131 17731
rect 20073 17691 20131 17697
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 18966 17660 18972 17672
rect 18555 17632 18972 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 13170 17552 13176 17604
rect 13228 17592 13234 17604
rect 13725 17595 13783 17601
rect 13725 17592 13737 17595
rect 13228 17564 13737 17592
rect 13228 17552 13234 17564
rect 13725 17561 13737 17564
rect 13771 17561 13783 17595
rect 13725 17555 13783 17561
rect 14826 17552 14832 17604
rect 14884 17592 14890 17604
rect 15933 17595 15991 17601
rect 15933 17592 15945 17595
rect 14884 17564 15945 17592
rect 14884 17552 14890 17564
rect 15933 17561 15945 17564
rect 15979 17592 15991 17595
rect 16298 17592 16304 17604
rect 15979 17564 16304 17592
rect 15979 17561 15991 17564
rect 15933 17555 15991 17561
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 17954 17552 17960 17604
rect 18012 17592 18018 17604
rect 18340 17592 18368 17623
rect 18966 17620 18972 17632
rect 19024 17620 19030 17672
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 20088 17632 20177 17660
rect 20088 17604 20116 17632
rect 20165 17629 20177 17632
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 18012 17564 18368 17592
rect 18012 17552 18018 17564
rect 18782 17552 18788 17604
rect 18840 17592 18846 17604
rect 19150 17592 19156 17604
rect 18840 17564 19156 17592
rect 18840 17552 18846 17564
rect 19150 17552 19156 17564
rect 19208 17592 19214 17604
rect 19208 17564 19334 17592
rect 19208 17552 19214 17564
rect 11563 17496 11928 17524
rect 11563 17493 11575 17496
rect 11517 17487 11575 17493
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 14185 17527 14243 17533
rect 14185 17524 14197 17527
rect 13320 17496 14197 17524
rect 13320 17484 13326 17496
rect 14185 17493 14197 17496
rect 14231 17493 14243 17527
rect 14185 17487 14243 17493
rect 15194 17484 15200 17536
rect 15252 17524 15258 17536
rect 18414 17524 18420 17536
rect 15252 17496 18420 17524
rect 15252 17484 15258 17496
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17524 18751 17527
rect 18966 17524 18972 17536
rect 18739 17496 18972 17524
rect 18739 17493 18751 17496
rect 18693 17487 18751 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19306 17524 19334 17564
rect 20070 17552 20076 17604
rect 20128 17552 20134 17604
rect 21952 17592 21980 17768
rect 22370 17688 22376 17740
rect 22428 17728 22434 17740
rect 23290 17728 23296 17740
rect 22428 17700 22784 17728
rect 22428 17688 22434 17700
rect 22554 17620 22560 17672
rect 22612 17620 22618 17672
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 22756 17669 22784 17700
rect 22894 17700 23296 17728
rect 22894 17672 22922 17700
rect 23290 17688 23296 17700
rect 23348 17688 23354 17740
rect 28966 17728 28994 17768
rect 36817 17765 36829 17799
rect 36863 17765 36875 17799
rect 36817 17759 36875 17765
rect 27172 17700 27752 17728
rect 28966 17700 30604 17728
rect 22741 17663 22799 17669
rect 22741 17629 22753 17663
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 22830 17620 22836 17672
rect 22888 17663 22922 17672
rect 22905 17632 22922 17663
rect 22905 17629 22917 17632
rect 22888 17623 22917 17629
rect 22888 17620 22894 17623
rect 23014 17620 23020 17672
rect 23072 17620 23078 17672
rect 24026 17620 24032 17672
rect 24084 17660 24090 17672
rect 26881 17663 26939 17669
rect 26881 17660 26893 17663
rect 24084 17632 26893 17660
rect 24084 17620 24090 17632
rect 26881 17629 26893 17632
rect 26927 17629 26939 17663
rect 26881 17623 26939 17629
rect 26970 17620 26976 17672
rect 27028 17620 27034 17672
rect 27172 17669 27200 17700
rect 27724 17672 27752 17700
rect 27157 17663 27215 17669
rect 27157 17629 27169 17663
rect 27203 17629 27215 17663
rect 27157 17623 27215 17629
rect 27246 17620 27252 17672
rect 27304 17620 27310 17672
rect 27706 17620 27712 17672
rect 27764 17620 27770 17672
rect 28994 17620 29000 17672
rect 29052 17620 29058 17672
rect 26050 17592 26056 17604
rect 21952 17564 26056 17592
rect 26050 17552 26056 17564
rect 26108 17552 26114 17604
rect 26988 17592 27016 17620
rect 29012 17592 29040 17620
rect 26344 17564 26832 17592
rect 26988 17564 29040 17592
rect 30576 17592 30604 17700
rect 30742 17688 30748 17740
rect 30800 17688 30806 17740
rect 31496 17700 34284 17728
rect 30653 17663 30711 17669
rect 30653 17629 30665 17663
rect 30699 17660 30711 17663
rect 31113 17663 31171 17669
rect 31113 17660 31125 17663
rect 30699 17632 31125 17660
rect 30699 17629 30711 17632
rect 30653 17623 30711 17629
rect 31113 17629 31125 17632
rect 31159 17629 31171 17663
rect 31113 17623 31171 17629
rect 31294 17620 31300 17672
rect 31352 17620 31358 17672
rect 31496 17592 31524 17700
rect 31573 17663 31631 17669
rect 31573 17629 31585 17663
rect 31619 17660 31631 17663
rect 33686 17660 33692 17672
rect 31619 17632 33692 17660
rect 31619 17629 31631 17632
rect 31573 17623 31631 17629
rect 33686 17620 33692 17632
rect 33744 17620 33750 17672
rect 34256 17660 34284 17700
rect 34624 17700 35204 17728
rect 34624 17660 34652 17700
rect 34256 17632 34652 17660
rect 34698 17620 34704 17672
rect 34756 17660 34762 17672
rect 35176 17660 35204 17700
rect 35894 17688 35900 17740
rect 35952 17688 35958 17740
rect 36538 17688 36544 17740
rect 36596 17688 36602 17740
rect 35526 17660 35532 17672
rect 34756 17632 35112 17660
rect 35176 17632 35532 17660
rect 34756 17620 34762 17632
rect 30576 17564 31524 17592
rect 26344 17536 26372 17564
rect 20162 17524 20168 17536
rect 19306 17496 20168 17524
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 20533 17527 20591 17533
rect 20533 17493 20545 17527
rect 20579 17524 20591 17527
rect 21082 17524 21088 17536
rect 20579 17496 21088 17524
rect 20579 17493 20591 17496
rect 20533 17487 20591 17493
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 23842 17484 23848 17536
rect 23900 17524 23906 17536
rect 24118 17524 24124 17536
rect 23900 17496 24124 17524
rect 23900 17484 23906 17496
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 26326 17484 26332 17536
rect 26384 17484 26390 17536
rect 26694 17484 26700 17536
rect 26752 17484 26758 17536
rect 26804 17524 26832 17564
rect 34606 17552 34612 17604
rect 34664 17592 34670 17604
rect 34977 17595 35035 17601
rect 34977 17592 34989 17595
rect 34664 17564 34989 17592
rect 34664 17552 34670 17564
rect 34977 17561 34989 17564
rect 35023 17561 35035 17595
rect 35084 17592 35112 17632
rect 35526 17620 35532 17632
rect 35584 17660 35590 17672
rect 35805 17663 35863 17669
rect 35805 17660 35817 17663
rect 35584 17632 35817 17660
rect 35584 17620 35590 17632
rect 35805 17629 35817 17632
rect 35851 17660 35863 17663
rect 36449 17663 36507 17669
rect 36449 17660 36461 17663
rect 35851 17632 36461 17660
rect 35851 17629 35863 17632
rect 35805 17623 35863 17629
rect 36449 17629 36461 17632
rect 36495 17629 36507 17663
rect 36832 17660 36860 17759
rect 37108 17669 37136 17836
rect 38838 17824 38844 17876
rect 38896 17864 38902 17876
rect 39577 17867 39635 17873
rect 39577 17864 39589 17867
rect 38896 17836 39589 17864
rect 38896 17824 38902 17836
rect 39577 17833 39589 17836
rect 39623 17833 39635 17867
rect 39577 17827 39635 17833
rect 36909 17663 36967 17669
rect 36909 17660 36921 17663
rect 36832 17632 36921 17660
rect 36449 17623 36507 17629
rect 36909 17629 36921 17632
rect 36955 17629 36967 17663
rect 36909 17623 36967 17629
rect 37093 17663 37151 17669
rect 37093 17629 37105 17663
rect 37139 17629 37151 17663
rect 40586 17660 40592 17672
rect 37093 17623 37151 17629
rect 39132 17632 40592 17660
rect 35253 17595 35311 17601
rect 35253 17592 35265 17595
rect 35084 17564 35265 17592
rect 34977 17555 35035 17561
rect 35253 17561 35265 17564
rect 35299 17561 35311 17595
rect 35253 17555 35311 17561
rect 35345 17595 35403 17601
rect 35345 17561 35357 17595
rect 35391 17592 35403 17595
rect 35391 17564 36216 17592
rect 35391 17561 35403 17564
rect 35345 17555 35403 17561
rect 28534 17524 28540 17536
rect 26804 17496 28540 17524
rect 28534 17484 28540 17496
rect 28592 17524 28598 17536
rect 29638 17524 29644 17536
rect 28592 17496 29644 17524
rect 28592 17484 28598 17496
rect 29638 17484 29644 17496
rect 29696 17524 29702 17536
rect 31481 17527 31539 17533
rect 31481 17524 31493 17527
rect 29696 17496 31493 17524
rect 29696 17484 29702 17496
rect 31481 17493 31493 17496
rect 31527 17493 31539 17527
rect 31481 17487 31539 17493
rect 34514 17484 34520 17536
rect 34572 17524 34578 17536
rect 36188 17533 36216 17564
rect 36354 17552 36360 17604
rect 36412 17592 36418 17604
rect 39132 17592 39160 17632
rect 40586 17620 40592 17632
rect 40644 17620 40650 17672
rect 36412 17564 39160 17592
rect 39209 17595 39267 17601
rect 36412 17552 36418 17564
rect 39209 17561 39221 17595
rect 39255 17561 39267 17595
rect 39209 17555 39267 17561
rect 35161 17527 35219 17533
rect 35161 17524 35173 17527
rect 34572 17496 35173 17524
rect 34572 17484 34578 17496
rect 35161 17493 35173 17496
rect 35207 17493 35219 17527
rect 35161 17487 35219 17493
rect 36173 17527 36231 17533
rect 36173 17493 36185 17527
rect 36219 17493 36231 17527
rect 36173 17487 36231 17493
rect 37093 17527 37151 17533
rect 37093 17493 37105 17527
rect 37139 17524 37151 17527
rect 37826 17524 37832 17536
rect 37139 17496 37832 17524
rect 37139 17493 37151 17496
rect 37093 17487 37151 17493
rect 37826 17484 37832 17496
rect 37884 17484 37890 17536
rect 39224 17524 39252 17555
rect 39390 17552 39396 17604
rect 39448 17552 39454 17604
rect 40494 17552 40500 17604
rect 40552 17592 40558 17604
rect 40681 17595 40739 17601
rect 40681 17592 40693 17595
rect 40552 17564 40693 17592
rect 40552 17552 40558 17564
rect 40681 17561 40693 17564
rect 40727 17561 40739 17595
rect 40681 17555 40739 17561
rect 39482 17524 39488 17536
rect 39224 17496 39488 17524
rect 39482 17484 39488 17496
rect 39540 17484 39546 17536
rect 40957 17527 41015 17533
rect 40957 17493 40969 17527
rect 41003 17524 41015 17527
rect 41003 17496 41552 17524
rect 41003 17493 41015 17496
rect 40957 17487 41015 17493
rect 41524 17468 41552 17496
rect 1104 17434 41400 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 41400 17434
rect 41506 17416 41512 17468
rect 41564 17416 41570 17468
rect 1104 17360 41400 17382
rect 4890 17280 4896 17332
rect 4948 17320 4954 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 4948 17292 5457 17320
rect 4948 17280 4954 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5445 17283 5503 17289
rect 6733 17323 6791 17329
rect 6733 17289 6745 17323
rect 6779 17320 6791 17323
rect 7190 17320 7196 17332
rect 6779 17292 7196 17320
rect 6779 17289 6791 17292
rect 6733 17283 6791 17289
rect 7190 17280 7196 17292
rect 7248 17280 7254 17332
rect 10134 17320 10140 17332
rect 9416 17292 10140 17320
rect 9416 17264 9444 17292
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 11664 17292 12541 17320
rect 11664 17280 11670 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 12529 17283 12587 17289
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17320 12955 17323
rect 13170 17320 13176 17332
rect 12943 17292 13176 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 13262 17280 13268 17332
rect 13320 17280 13326 17332
rect 15378 17280 15384 17332
rect 15436 17280 15442 17332
rect 15473 17323 15531 17329
rect 15473 17289 15485 17323
rect 15519 17320 15531 17323
rect 15562 17320 15568 17332
rect 15519 17292 15568 17320
rect 15519 17289 15531 17292
rect 15473 17283 15531 17289
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 15654 17280 15660 17332
rect 15712 17280 15718 17332
rect 17586 17280 17592 17332
rect 17644 17280 17650 17332
rect 18414 17280 18420 17332
rect 18472 17320 18478 17332
rect 26970 17320 26976 17332
rect 18472 17292 26976 17320
rect 18472 17280 18478 17292
rect 26970 17280 26976 17292
rect 27028 17280 27034 17332
rect 29638 17280 29644 17332
rect 29696 17320 29702 17332
rect 30101 17323 30159 17329
rect 30101 17320 30113 17323
rect 29696 17292 30113 17320
rect 29696 17280 29702 17292
rect 30101 17289 30113 17292
rect 30147 17289 30159 17323
rect 30101 17283 30159 17289
rect 30650 17280 30656 17332
rect 30708 17280 30714 17332
rect 30742 17280 30748 17332
rect 30800 17320 30806 17332
rect 30929 17323 30987 17329
rect 30929 17320 30941 17323
rect 30800 17292 30941 17320
rect 30800 17280 30806 17292
rect 30929 17289 30941 17292
rect 30975 17289 30987 17323
rect 30929 17283 30987 17289
rect 33137 17323 33195 17329
rect 33137 17289 33149 17323
rect 33183 17320 33195 17323
rect 33318 17320 33324 17332
rect 33183 17292 33324 17320
rect 33183 17289 33195 17292
rect 33137 17283 33195 17289
rect 33318 17280 33324 17292
rect 33376 17280 33382 17332
rect 37366 17280 37372 17332
rect 37424 17280 37430 17332
rect 39393 17323 39451 17329
rect 39393 17320 39405 17323
rect 38764 17292 39405 17320
rect 5810 17252 5816 17264
rect 4632 17224 5816 17252
rect 4632 17193 4660 17224
rect 5810 17212 5816 17224
rect 5868 17212 5874 17264
rect 6932 17224 8340 17252
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17184 4859 17187
rect 4847 17156 5028 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17085 4767 17119
rect 4709 17079 4767 17085
rect 4724 17048 4752 17079
rect 4890 17076 4896 17128
rect 4948 17076 4954 17128
rect 5000 17116 5028 17156
rect 5074 17144 5080 17196
rect 5132 17144 5138 17196
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17184 5319 17187
rect 5350 17184 5356 17196
rect 5307 17156 5356 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 6932 17193 6960 17224
rect 6917 17190 6975 17193
rect 6840 17187 6975 17190
rect 6840 17184 6929 17187
rect 6788 17162 6929 17184
rect 6788 17156 6868 17162
rect 6788 17144 6794 17156
rect 6917 17153 6929 17162
rect 6963 17153 6975 17187
rect 6917 17147 6975 17153
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17184 7895 17187
rect 7926 17184 7932 17196
rect 7883 17156 7932 17184
rect 7883 17153 7895 17156
rect 7837 17147 7895 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8036 17193 8064 17224
rect 8312 17193 8340 17224
rect 8478 17212 8484 17264
rect 8536 17212 8542 17264
rect 8941 17255 8999 17261
rect 8941 17221 8953 17255
rect 8987 17252 8999 17255
rect 9306 17252 9312 17264
rect 8987 17224 9312 17252
rect 8987 17221 8999 17224
rect 8941 17215 8999 17221
rect 9306 17212 9312 17224
rect 9364 17212 9370 17264
rect 9398 17212 9404 17264
rect 9456 17212 9462 17264
rect 11514 17212 11520 17264
rect 11572 17252 11578 17264
rect 11882 17252 11888 17264
rect 11572 17224 11888 17252
rect 11572 17212 11578 17224
rect 11882 17212 11888 17224
rect 11940 17252 11946 17264
rect 12989 17255 13047 17261
rect 11940 17224 12940 17252
rect 11940 17212 11946 17224
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 8297 17187 8355 17193
rect 8297 17153 8309 17187
rect 8343 17184 8355 17187
rect 8754 17184 8760 17196
rect 8343 17156 8760 17184
rect 8343 17153 8355 17156
rect 8297 17147 8355 17153
rect 5534 17116 5540 17128
rect 5000 17088 5540 17116
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 6012 17048 6040 17144
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17085 7251 17119
rect 8220 17116 8248 17147
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 8846 17144 8852 17196
rect 8904 17144 8910 17196
rect 9030 17144 9036 17196
rect 9088 17144 9094 17196
rect 9122 17144 9128 17196
rect 9180 17193 9186 17196
rect 9180 17187 9209 17193
rect 9197 17153 9209 17187
rect 9180 17147 9209 17153
rect 9180 17144 9186 17147
rect 9582 17144 9588 17196
rect 9640 17144 9646 17196
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17184 11759 17187
rect 12250 17184 12256 17196
rect 11747 17156 12256 17184
rect 11747 17153 11759 17156
rect 11701 17147 11759 17153
rect 12250 17144 12256 17156
rect 12308 17144 12314 17196
rect 12912 17184 12940 17224
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 13280 17252 13308 17280
rect 13035 17224 13308 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 14182 17212 14188 17264
rect 14240 17212 14246 17264
rect 15396 17252 15424 17280
rect 15120 17224 15424 17252
rect 17604 17252 17632 17280
rect 17604 17224 18920 17252
rect 14200 17184 14228 17212
rect 12912 17156 14228 17184
rect 14826 17144 14832 17196
rect 14884 17144 14890 17196
rect 15120 17193 15148 17224
rect 14922 17187 14980 17193
rect 14922 17153 14934 17187
rect 14968 17153 14980 17187
rect 14922 17147 14980 17153
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 9306 17116 9312 17128
rect 8220 17088 9312 17116
rect 7193 17079 7251 17085
rect 4724 17020 6040 17048
rect 7208 17048 7236 17079
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 13170 17076 13176 17128
rect 13228 17076 13234 17128
rect 7374 17048 7380 17060
rect 7208 17020 7380 17048
rect 7374 17008 7380 17020
rect 7432 17048 7438 17060
rect 8478 17048 8484 17060
rect 7432 17020 8484 17048
rect 7432 17008 7438 17020
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 8846 17008 8852 17060
rect 8904 17048 8910 17060
rect 10042 17048 10048 17060
rect 8904 17020 10048 17048
rect 8904 17008 8910 17020
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 12158 17008 12164 17060
rect 12216 17048 12222 17060
rect 14937 17048 14965 17147
rect 15194 17144 15200 17196
rect 15252 17144 15258 17196
rect 15286 17144 15292 17196
rect 15344 17193 15350 17196
rect 15344 17184 15352 17193
rect 16117 17187 16175 17193
rect 16117 17184 16129 17187
rect 15344 17156 15389 17184
rect 15488 17156 16129 17184
rect 15344 17147 15352 17156
rect 15344 17144 15350 17147
rect 12216 17020 14965 17048
rect 12216 17008 12222 17020
rect 3418 16940 3424 16992
rect 3476 16980 3482 16992
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 3476 16952 4445 16980
rect 3476 16940 3482 16952
rect 4433 16949 4445 16952
rect 4479 16949 4491 16983
rect 4433 16943 4491 16949
rect 7101 16983 7159 16989
rect 7101 16949 7113 16983
rect 7147 16980 7159 16983
rect 7466 16980 7472 16992
rect 7147 16952 7472 16980
rect 7147 16949 7159 16952
rect 7101 16943 7159 16949
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 7929 16983 7987 16989
rect 7929 16949 7941 16983
rect 7975 16980 7987 16983
rect 8110 16980 8116 16992
rect 7975 16952 8116 16980
rect 7975 16949 7987 16952
rect 7929 16943 7987 16949
rect 8110 16940 8116 16952
rect 8168 16940 8174 16992
rect 8662 16940 8668 16992
rect 8720 16940 8726 16992
rect 9766 16940 9772 16992
rect 9824 16940 9830 16992
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 11756 16952 11897 16980
rect 11756 16940 11762 16952
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 11885 16943 11943 16949
rect 14274 16940 14280 16992
rect 14332 16980 14338 16992
rect 15488 16980 15516 17156
rect 16117 17153 16129 17156
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 17218 17144 17224 17196
rect 17276 17144 17282 17196
rect 18046 17144 18052 17196
rect 18104 17144 18110 17196
rect 18340 17193 18368 17224
rect 18325 17187 18383 17193
rect 18325 17153 18337 17187
rect 18371 17153 18383 17187
rect 18325 17147 18383 17153
rect 18509 17187 18567 17193
rect 18509 17153 18521 17187
rect 18555 17184 18567 17187
rect 18690 17184 18696 17196
rect 18555 17156 18696 17184
rect 18555 17153 18567 17156
rect 18509 17147 18567 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 18785 17187 18843 17193
rect 18785 17153 18797 17187
rect 18831 17182 18843 17187
rect 18892 17182 18920 17224
rect 18966 17212 18972 17264
rect 19024 17252 19030 17264
rect 20530 17252 20536 17264
rect 19024 17224 20536 17252
rect 19024 17212 19030 17224
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 20717 17255 20775 17261
rect 20717 17221 20729 17255
rect 20763 17252 20775 17255
rect 20901 17255 20959 17261
rect 20763 17224 20797 17252
rect 20763 17221 20775 17224
rect 20717 17215 20775 17221
rect 20901 17221 20913 17255
rect 20947 17252 20959 17255
rect 20990 17252 20996 17264
rect 20947 17224 20996 17252
rect 20947 17221 20959 17224
rect 20901 17215 20959 17221
rect 18831 17154 18920 17182
rect 20073 17187 20131 17193
rect 18831 17153 18843 17154
rect 18785 17147 18843 17153
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 15562 17076 15568 17128
rect 15620 17076 15626 17128
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17116 15899 17119
rect 16758 17116 16764 17128
rect 15887 17088 16764 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 17236 17116 17264 17144
rect 17586 17116 17592 17128
rect 17236 17088 17592 17116
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 18064 17116 18092 17144
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 18064 17088 18613 17116
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 18969 17119 19027 17125
rect 18969 17085 18981 17119
rect 19015 17116 19027 17119
rect 19978 17116 19984 17128
rect 19015 17088 19984 17116
rect 19015 17085 19027 17088
rect 18969 17079 19027 17085
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 15580 17048 15608 17076
rect 16025 17051 16083 17057
rect 16025 17048 16037 17051
rect 15580 17020 16037 17048
rect 16025 17017 16037 17020
rect 16071 17017 16083 17051
rect 16025 17011 16083 17017
rect 16114 17008 16120 17060
rect 16172 17048 16178 17060
rect 18138 17048 18144 17060
rect 16172 17020 18144 17048
rect 16172 17008 16178 17020
rect 18138 17008 18144 17020
rect 18196 17008 18202 17060
rect 18325 17051 18383 17057
rect 18325 17017 18337 17051
rect 18371 17048 18383 17051
rect 19426 17048 19432 17060
rect 18371 17020 19432 17048
rect 18371 17017 18383 17020
rect 18325 17011 18383 17017
rect 19426 17008 19432 17020
rect 19484 17008 19490 17060
rect 20088 16992 20116 17147
rect 20162 17144 20168 17196
rect 20220 17184 20226 17196
rect 20257 17187 20315 17193
rect 20257 17184 20269 17187
rect 20220 17156 20269 17184
rect 20220 17144 20226 17156
rect 20257 17153 20269 17156
rect 20303 17153 20315 17187
rect 20257 17147 20315 17153
rect 20438 17144 20444 17196
rect 20496 17184 20502 17196
rect 20732 17184 20760 17215
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 21266 17212 21272 17264
rect 21324 17252 21330 17264
rect 21726 17252 21732 17264
rect 21324 17224 21732 17252
rect 21324 17212 21330 17224
rect 21726 17212 21732 17224
rect 21784 17252 21790 17264
rect 21784 17224 22048 17252
rect 21784 17212 21790 17224
rect 21818 17184 21824 17196
rect 20496 17156 21824 17184
rect 20496 17144 20502 17156
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 22020 17184 22048 17224
rect 22094 17212 22100 17264
rect 22152 17252 22158 17264
rect 26513 17255 26571 17261
rect 26513 17252 26525 17255
rect 22152 17224 24348 17252
rect 22152 17212 22158 17224
rect 23106 17184 23112 17196
rect 22020 17156 23112 17184
rect 23106 17144 23112 17156
rect 23164 17144 23170 17196
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17184 23351 17187
rect 23934 17184 23940 17196
rect 23339 17156 23940 17184
rect 23339 17153 23351 17156
rect 23293 17147 23351 17153
rect 23934 17144 23940 17156
rect 23992 17144 23998 17196
rect 24026 17144 24032 17196
rect 24084 17144 24090 17196
rect 24320 17193 24348 17224
rect 25332 17224 26525 17252
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 24305 17187 24363 17193
rect 24305 17153 24317 17187
rect 24351 17153 24363 17187
rect 24305 17147 24363 17153
rect 24765 17187 24823 17193
rect 24765 17153 24777 17187
rect 24811 17153 24823 17187
rect 24765 17147 24823 17153
rect 24949 17187 25007 17193
rect 24949 17153 24961 17187
rect 24995 17153 25007 17187
rect 24949 17147 25007 17153
rect 23124 17116 23152 17144
rect 24228 17116 24256 17147
rect 24780 17116 24808 17147
rect 23124 17088 24256 17116
rect 20162 17008 20168 17060
rect 20220 17048 20226 17060
rect 20714 17048 20720 17060
rect 20220 17020 20720 17048
rect 20220 17008 20226 17020
rect 20714 17008 20720 17020
rect 20772 17008 20778 17060
rect 20806 17008 20812 17060
rect 20864 17048 20870 17060
rect 21634 17048 21640 17060
rect 20864 17020 21640 17048
rect 20864 17008 20870 17020
rect 21634 17008 21640 17020
rect 21692 17048 21698 17060
rect 23658 17048 23664 17060
rect 21692 17020 23664 17048
rect 21692 17008 21698 17020
rect 23658 17008 23664 17020
rect 23716 17008 23722 17060
rect 14332 16952 15516 16980
rect 14332 16940 14338 16952
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 20070 16980 20076 16992
rect 17368 16952 20076 16980
rect 17368 16940 17374 16952
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20254 16940 20260 16992
rect 20312 16980 20318 16992
rect 20898 16980 20904 16992
rect 20312 16952 20904 16980
rect 20312 16940 20318 16952
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 21085 16983 21143 16989
rect 21085 16949 21097 16983
rect 21131 16980 21143 16983
rect 21726 16980 21732 16992
rect 21131 16952 21732 16980
rect 21131 16949 21143 16952
rect 21085 16943 21143 16949
rect 21726 16940 21732 16952
rect 21784 16940 21790 16992
rect 22462 16940 22468 16992
rect 22520 16980 22526 16992
rect 23014 16980 23020 16992
rect 22520 16952 23020 16980
rect 22520 16940 22526 16952
rect 23014 16940 23020 16952
rect 23072 16940 23078 16992
rect 23474 16940 23480 16992
rect 23532 16940 23538 16992
rect 24228 16980 24256 17088
rect 24320 17088 24808 17116
rect 24320 17057 24348 17088
rect 24305 17051 24363 17057
rect 24305 17017 24317 17051
rect 24351 17017 24363 17051
rect 24305 17011 24363 17017
rect 24394 17008 24400 17060
rect 24452 17048 24458 17060
rect 24964 17048 24992 17147
rect 25038 17144 25044 17196
rect 25096 17144 25102 17196
rect 25332 17193 25360 17224
rect 26513 17221 26525 17224
rect 26559 17221 26571 17255
rect 26513 17215 26571 17221
rect 29917 17255 29975 17261
rect 29917 17221 29929 17255
rect 29963 17252 29975 17255
rect 36630 17252 36636 17264
rect 29963 17224 30880 17252
rect 29963 17221 29975 17224
rect 29917 17215 29975 17221
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 26421 17187 26479 17193
rect 26421 17153 26433 17187
rect 26467 17184 26479 17187
rect 27430 17184 27436 17196
rect 26467 17156 27436 17184
rect 26467 17153 26479 17156
rect 26421 17147 26479 17153
rect 27430 17144 27436 17156
rect 27488 17144 27494 17196
rect 29730 17144 29736 17196
rect 29788 17184 29794 17196
rect 29932 17184 29960 17215
rect 29788 17156 29960 17184
rect 29788 17144 29794 17156
rect 30098 17144 30104 17196
rect 30156 17184 30162 17196
rect 30377 17187 30435 17193
rect 30377 17184 30389 17187
rect 30156 17156 30389 17184
rect 30156 17144 30162 17156
rect 30377 17153 30389 17156
rect 30423 17153 30435 17187
rect 30377 17147 30435 17153
rect 30650 17144 30656 17196
rect 30708 17144 30714 17196
rect 30852 17193 30880 17224
rect 31726 17224 36636 17252
rect 30837 17187 30895 17193
rect 30837 17153 30849 17187
rect 30883 17153 30895 17187
rect 30837 17147 30895 17153
rect 30926 17144 30932 17196
rect 30984 17184 30990 17196
rect 31021 17187 31079 17193
rect 31021 17184 31033 17187
rect 30984 17156 31033 17184
rect 30984 17144 30990 17156
rect 31021 17153 31033 17156
rect 31067 17153 31079 17187
rect 31021 17147 31079 17153
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24452 17020 24992 17048
rect 25056 17088 25145 17116
rect 24452 17008 24458 17020
rect 25056 16980 25084 17088
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 30024 17088 31340 17116
rect 29549 17051 29607 17057
rect 29549 17017 29561 17051
rect 29595 17017 29607 17051
rect 29549 17011 29607 17017
rect 24228 16952 25084 16980
rect 25498 16940 25504 16992
rect 25556 16940 25562 16992
rect 26602 16940 26608 16992
rect 26660 16980 26666 16992
rect 26970 16980 26976 16992
rect 26660 16952 26976 16980
rect 26660 16940 26666 16952
rect 26970 16940 26976 16952
rect 27028 16940 27034 16992
rect 29454 16940 29460 16992
rect 29512 16980 29518 16992
rect 29564 16980 29592 17011
rect 29512 16952 29592 16980
rect 29512 16940 29518 16952
rect 29914 16940 29920 16992
rect 29972 16980 29978 16992
rect 30024 16980 30052 17088
rect 31312 17060 31340 17088
rect 31294 17008 31300 17060
rect 31352 17008 31358 17060
rect 29972 16952 30052 16980
rect 29972 16940 29978 16952
rect 31202 16940 31208 16992
rect 31260 16980 31266 16992
rect 31726 16980 31754 17224
rect 36630 17212 36636 17224
rect 36688 17212 36694 17264
rect 37384 17252 37412 17280
rect 38764 17261 38792 17292
rect 39393 17289 39405 17292
rect 39439 17289 39451 17323
rect 39393 17283 39451 17289
rect 38749 17255 38807 17261
rect 37384 17224 38700 17252
rect 33413 17187 33471 17193
rect 33413 17153 33425 17187
rect 33459 17184 33471 17187
rect 33459 17156 33824 17184
rect 33459 17153 33471 17156
rect 33413 17147 33471 17153
rect 33796 17128 33824 17156
rect 33870 17144 33876 17196
rect 33928 17184 33934 17196
rect 37918 17184 37924 17196
rect 33928 17156 37924 17184
rect 33928 17144 33934 17156
rect 37918 17144 37924 17156
rect 37976 17144 37982 17196
rect 38470 17144 38476 17196
rect 38528 17144 38534 17196
rect 38672 17193 38700 17224
rect 38749 17221 38761 17255
rect 38795 17221 38807 17255
rect 39206 17252 39212 17264
rect 38749 17215 38807 17221
rect 38979 17221 39037 17227
rect 38657 17187 38715 17193
rect 38657 17153 38669 17187
rect 38703 17153 38715 17187
rect 38657 17147 38715 17153
rect 33134 17076 33140 17128
rect 33192 17116 33198 17128
rect 33321 17119 33379 17125
rect 33321 17116 33333 17119
rect 33192 17088 33333 17116
rect 33192 17076 33198 17088
rect 33321 17085 33333 17088
rect 33367 17085 33379 17119
rect 33321 17079 33379 17085
rect 33502 17076 33508 17128
rect 33560 17076 33566 17128
rect 33597 17119 33655 17125
rect 33597 17085 33609 17119
rect 33643 17116 33655 17119
rect 33686 17116 33692 17128
rect 33643 17088 33692 17116
rect 33643 17085 33655 17088
rect 33597 17079 33655 17085
rect 33686 17076 33692 17088
rect 33744 17076 33750 17128
rect 33778 17076 33784 17128
rect 33836 17076 33842 17128
rect 38764 17060 38792 17215
rect 38979 17187 38991 17221
rect 39025 17187 39037 17221
rect 38979 17184 39037 17187
rect 39132 17224 39212 17252
rect 39132 17184 39160 17224
rect 39206 17212 39212 17224
rect 39264 17252 39270 17264
rect 39264 17224 39306 17252
rect 39264 17212 39270 17224
rect 39485 17187 39543 17193
rect 39485 17184 39497 17187
rect 38979 17181 39160 17184
rect 38980 17156 39160 17181
rect 39224 17156 39497 17184
rect 39224 17116 39252 17156
rect 39485 17153 39497 17156
rect 39531 17153 39543 17187
rect 39485 17147 39543 17153
rect 38948 17088 39252 17116
rect 39316 17088 39528 17116
rect 32950 17008 32956 17060
rect 33008 17048 33014 17060
rect 38565 17051 38623 17057
rect 33008 17020 34284 17048
rect 33008 17008 33014 17020
rect 34256 16992 34284 17020
rect 38565 17017 38577 17051
rect 38611 17048 38623 17051
rect 38746 17048 38752 17060
rect 38611 17020 38752 17048
rect 38611 17017 38623 17020
rect 38565 17011 38623 17017
rect 38746 17008 38752 17020
rect 38804 17008 38810 17060
rect 38948 16992 38976 17088
rect 39117 17051 39175 17057
rect 39117 17017 39129 17051
rect 39163 17048 39175 17051
rect 39316 17048 39344 17088
rect 39500 17060 39528 17088
rect 40494 17076 40500 17128
rect 40552 17076 40558 17128
rect 39163 17020 39344 17048
rect 39163 17017 39175 17020
rect 39117 17011 39175 17017
rect 39482 17008 39488 17060
rect 39540 17008 39546 17060
rect 31260 16952 31754 16980
rect 31260 16940 31266 16952
rect 33410 16940 33416 16992
rect 33468 16980 33474 16992
rect 34146 16980 34152 16992
rect 33468 16952 34152 16980
rect 33468 16940 33474 16952
rect 34146 16940 34152 16952
rect 34204 16940 34210 16992
rect 34238 16940 34244 16992
rect 34296 16980 34302 16992
rect 36262 16980 36268 16992
rect 34296 16952 36268 16980
rect 34296 16940 34302 16952
rect 36262 16940 36268 16952
rect 36320 16940 36326 16992
rect 38930 16940 38936 16992
rect 38988 16940 38994 16992
rect 39209 16983 39267 16989
rect 39209 16949 39221 16983
rect 39255 16980 39267 16983
rect 39390 16980 39396 16992
rect 39255 16952 39396 16980
rect 39255 16949 39267 16952
rect 39209 16943 39267 16949
rect 39390 16940 39396 16952
rect 39448 16940 39454 16992
rect 41046 16940 41052 16992
rect 41104 16940 41110 16992
rect 1104 16890 41400 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 41400 16890
rect 1104 16816 41400 16838
rect 8662 16736 8668 16788
rect 8720 16736 8726 16788
rect 8754 16736 8760 16788
rect 8812 16776 8818 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8812 16748 9137 16776
rect 8812 16736 8818 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 9306 16736 9312 16788
rect 9364 16776 9370 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 9364 16748 9413 16776
rect 9364 16736 9370 16748
rect 9401 16745 9413 16748
rect 9447 16745 9459 16779
rect 9401 16739 9459 16745
rect 15194 16736 15200 16788
rect 15252 16776 15258 16788
rect 15381 16779 15439 16785
rect 15381 16776 15393 16779
rect 15252 16748 15393 16776
rect 15252 16736 15258 16748
rect 15381 16745 15393 16748
rect 15427 16776 15439 16779
rect 16022 16776 16028 16788
rect 15427 16748 16028 16776
rect 15427 16745 15439 16748
rect 15381 16739 15439 16745
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 16114 16736 16120 16788
rect 16172 16736 16178 16788
rect 17770 16736 17776 16788
rect 17828 16736 17834 16788
rect 21450 16736 21456 16788
rect 21508 16776 21514 16788
rect 21508 16748 23060 16776
rect 21508 16736 21514 16748
rect 5074 16708 5080 16720
rect 4264 16680 5080 16708
rect 4264 16640 4292 16680
rect 5074 16668 5080 16680
rect 5132 16708 5138 16720
rect 5353 16711 5411 16717
rect 5353 16708 5365 16711
rect 5132 16680 5365 16708
rect 5132 16668 5138 16680
rect 5353 16677 5365 16680
rect 5399 16677 5411 16711
rect 5353 16671 5411 16677
rect 7929 16711 7987 16717
rect 7929 16677 7941 16711
rect 7975 16708 7987 16711
rect 8389 16711 8447 16717
rect 8389 16708 8401 16711
rect 7975 16680 8401 16708
rect 7975 16677 7987 16680
rect 7929 16671 7987 16677
rect 8389 16677 8401 16680
rect 8435 16677 8447 16711
rect 8389 16671 8447 16677
rect 4706 16640 4712 16652
rect 3988 16612 4292 16640
rect 3786 16532 3792 16584
rect 3844 16572 3850 16584
rect 3988 16572 4016 16612
rect 3844 16544 4016 16572
rect 3844 16532 3850 16544
rect 4062 16532 4068 16584
rect 4120 16532 4126 16584
rect 4264 16581 4292 16612
rect 4448 16612 4712 16640
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4172 16504 4200 16535
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4448 16581 4476 16612
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 8021 16643 8079 16649
rect 4908 16612 5580 16640
rect 4433 16575 4491 16581
rect 4433 16572 4445 16575
rect 4396 16544 4445 16572
rect 4396 16532 4402 16544
rect 4433 16541 4445 16544
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 4908 16581 4936 16612
rect 4893 16575 4951 16581
rect 4893 16541 4905 16575
rect 4939 16541 4951 16575
rect 4893 16535 4951 16541
rect 4982 16532 4988 16584
rect 5040 16572 5046 16584
rect 5077 16575 5135 16581
rect 5077 16572 5089 16575
rect 5040 16544 5089 16572
rect 5040 16532 5046 16544
rect 5077 16541 5089 16544
rect 5123 16572 5135 16575
rect 5445 16575 5503 16581
rect 5445 16572 5457 16575
rect 5123 16544 5457 16572
rect 5123 16541 5135 16544
rect 5077 16535 5135 16541
rect 5445 16541 5457 16544
rect 5491 16541 5503 16575
rect 5552 16559 5580 16612
rect 8021 16609 8033 16643
rect 8067 16640 8079 16643
rect 8680 16640 8708 16736
rect 11514 16668 11520 16720
rect 11572 16708 11578 16720
rect 16132 16708 16160 16736
rect 11572 16680 16160 16708
rect 11572 16668 11578 16680
rect 16298 16668 16304 16720
rect 16356 16708 16362 16720
rect 19242 16708 19248 16720
rect 16356 16680 19248 16708
rect 16356 16668 16362 16680
rect 8067 16612 8708 16640
rect 8067 16609 8079 16612
rect 8021 16603 8079 16609
rect 9398 16600 9404 16652
rect 9456 16600 9462 16652
rect 9582 16640 9588 16652
rect 9508 16612 9588 16640
rect 5445 16535 5503 16541
rect 5535 16553 5593 16559
rect 4632 16504 4660 16532
rect 4172 16476 4660 16504
rect 5169 16507 5227 16513
rect 5169 16473 5181 16507
rect 5215 16504 5227 16507
rect 5258 16504 5264 16516
rect 5215 16476 5264 16504
rect 5215 16473 5227 16476
rect 5169 16467 5227 16473
rect 5258 16464 5264 16476
rect 5316 16464 5322 16516
rect 3789 16439 3847 16445
rect 3789 16405 3801 16439
rect 3835 16436 3847 16439
rect 4522 16436 4528 16448
rect 3835 16408 4528 16436
rect 3835 16405 3847 16408
rect 3789 16399 3847 16405
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 5460 16436 5488 16535
rect 5535 16519 5547 16553
rect 5581 16519 5593 16553
rect 7282 16532 7288 16584
rect 7340 16572 7346 16584
rect 7837 16575 7895 16581
rect 7837 16572 7849 16575
rect 7340 16544 7849 16572
rect 7340 16532 7346 16544
rect 7837 16541 7849 16544
rect 7883 16572 7895 16575
rect 7926 16572 7932 16584
rect 7883 16544 7932 16572
rect 7883 16541 7895 16544
rect 7837 16535 7895 16541
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 8110 16532 8116 16584
rect 8168 16532 8174 16584
rect 8294 16532 8300 16584
rect 8352 16532 8358 16584
rect 8386 16532 8392 16584
rect 8444 16532 8450 16584
rect 8478 16532 8484 16584
rect 8536 16572 8542 16584
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 8536 16544 8585 16572
rect 8536 16532 8542 16544
rect 8573 16541 8585 16544
rect 8619 16541 8631 16575
rect 8573 16535 8631 16541
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16572 9367 16575
rect 9416 16572 9444 16600
rect 9508 16581 9536 16612
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10778 16600 10784 16652
rect 10836 16640 10842 16652
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 10836 16612 11897 16640
rect 10836 16600 10842 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 11992 16612 12480 16640
rect 9355 16544 9444 16572
rect 9493 16575 9551 16581
rect 9355 16541 9367 16544
rect 9309 16535 9367 16541
rect 9493 16541 9505 16575
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 5535 16516 5593 16519
rect 5534 16464 5540 16516
rect 5592 16464 5598 16516
rect 8956 16504 8984 16535
rect 9766 16532 9772 16584
rect 9824 16532 9830 16584
rect 11422 16532 11428 16584
rect 11480 16532 11486 16584
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 11698 16572 11704 16584
rect 11655 16544 11704 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 9784 16504 9812 16532
rect 8956 16476 9812 16504
rect 11532 16504 11560 16535
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 11790 16532 11796 16584
rect 11848 16572 11854 16584
rect 11992 16572 12020 16612
rect 11848 16544 12020 16572
rect 12069 16575 12127 16581
rect 11848 16532 11854 16544
rect 12069 16541 12081 16575
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12250 16572 12256 16584
rect 12207 16544 12256 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 12084 16504 12112 16535
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 12342 16532 12348 16584
rect 12400 16532 12406 16584
rect 12452 16581 12480 16612
rect 13078 16600 13084 16652
rect 13136 16600 13142 16652
rect 13814 16600 13820 16652
rect 13872 16600 13878 16652
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 12897 16575 12955 16581
rect 12897 16541 12909 16575
rect 12943 16572 12955 16575
rect 12986 16572 12992 16584
rect 12943 16544 12992 16572
rect 12943 16541 12955 16544
rect 12897 16535 12955 16541
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 13446 16504 13452 16516
rect 11532 16476 12434 16504
rect 5626 16436 5632 16448
rect 5460 16408 5632 16436
rect 5626 16396 5632 16408
rect 5684 16396 5690 16448
rect 5718 16396 5724 16448
rect 5776 16436 5782 16448
rect 7374 16436 7380 16448
rect 5776 16408 7380 16436
rect 5776 16396 5782 16408
rect 7374 16396 7380 16408
rect 7432 16396 7438 16448
rect 7650 16396 7656 16448
rect 7708 16396 7714 16448
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 11149 16439 11207 16445
rect 11149 16436 11161 16439
rect 10928 16408 11161 16436
rect 10928 16396 10934 16408
rect 11149 16405 11161 16408
rect 11195 16405 11207 16439
rect 12406 16436 12434 16476
rect 13004 16476 13452 16504
rect 13004 16445 13032 16476
rect 13446 16464 13452 16476
rect 13504 16504 13510 16516
rect 13832 16504 13860 16600
rect 15378 16532 15384 16584
rect 15436 16572 15442 16584
rect 15565 16575 15623 16581
rect 15565 16572 15577 16575
rect 15436 16544 15577 16572
rect 15436 16532 15442 16544
rect 15565 16541 15577 16544
rect 15611 16541 15623 16575
rect 15565 16535 15623 16541
rect 13504 16476 13860 16504
rect 15580 16504 15608 16535
rect 15654 16532 15660 16584
rect 15712 16532 15718 16584
rect 15838 16532 15844 16584
rect 15896 16532 15902 16584
rect 16316 16581 16344 16668
rect 17236 16652 17264 16680
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 20438 16708 20444 16720
rect 20088 16680 20444 16708
rect 16666 16600 16672 16652
rect 16724 16600 16730 16652
rect 17218 16600 17224 16652
rect 17276 16600 17282 16652
rect 17586 16600 17592 16652
rect 17644 16640 17650 16652
rect 17644 16612 18184 16640
rect 17644 16600 17650 16612
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16572 15991 16575
rect 16025 16575 16083 16581
rect 16025 16572 16037 16575
rect 15979 16544 16037 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 16025 16541 16037 16544
rect 16071 16541 16083 16575
rect 16025 16535 16083 16541
rect 16209 16575 16267 16581
rect 16209 16541 16221 16575
rect 16255 16541 16267 16575
rect 16209 16535 16267 16541
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16541 16359 16575
rect 16301 16535 16359 16541
rect 16393 16575 16451 16581
rect 16393 16541 16405 16575
rect 16439 16572 16451 16575
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16439 16544 16957 16572
rect 16439 16541 16451 16544
rect 16393 16535 16451 16541
rect 16945 16541 16957 16544
rect 16991 16572 17003 16575
rect 17034 16572 17040 16584
rect 16991 16544 17040 16572
rect 16991 16541 17003 16544
rect 16945 16535 17003 16541
rect 15580 16476 16068 16504
rect 13504 16464 13510 16476
rect 16040 16448 16068 16476
rect 12529 16439 12587 16445
rect 12529 16436 12541 16439
rect 12406 16408 12541 16436
rect 11149 16399 11207 16405
rect 12529 16405 12541 16408
rect 12575 16405 12587 16439
rect 12529 16399 12587 16405
rect 12989 16439 13047 16445
rect 12989 16405 13001 16439
rect 13035 16405 13047 16439
rect 12989 16399 13047 16405
rect 13262 16396 13268 16448
rect 13320 16436 13326 16448
rect 15194 16436 15200 16448
rect 13320 16408 15200 16436
rect 13320 16396 13326 16408
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 16022 16396 16028 16448
rect 16080 16396 16086 16448
rect 16224 16436 16252 16535
rect 17034 16532 17040 16544
rect 17092 16572 17098 16584
rect 17092 16544 17448 16572
rect 17092 16532 17098 16544
rect 16482 16464 16488 16516
rect 16540 16513 16546 16516
rect 16540 16507 16569 16513
rect 16557 16473 16569 16507
rect 16540 16467 16569 16473
rect 16540 16464 16546 16467
rect 16758 16464 16764 16516
rect 16816 16504 16822 16516
rect 17129 16507 17187 16513
rect 17129 16504 17141 16507
rect 16816 16476 17141 16504
rect 16816 16464 16822 16476
rect 17129 16473 17141 16476
rect 17175 16504 17187 16507
rect 17310 16504 17316 16516
rect 17175 16476 17316 16504
rect 17175 16473 17187 16476
rect 17129 16467 17187 16473
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 17420 16504 17448 16544
rect 17494 16532 17500 16584
rect 17552 16532 17558 16584
rect 18046 16532 18052 16584
rect 18104 16532 18110 16584
rect 18156 16572 18184 16612
rect 18340 16612 19334 16640
rect 18340 16572 18368 16612
rect 18156 16544 18368 16572
rect 18064 16504 18092 16532
rect 17420 16476 18092 16504
rect 17957 16439 18015 16445
rect 17957 16436 17969 16439
rect 16224 16408 17969 16436
rect 17957 16405 17969 16408
rect 18003 16405 18015 16439
rect 19306 16436 19334 16612
rect 20088 16581 20116 16680
rect 20438 16668 20444 16680
rect 20496 16668 20502 16720
rect 20898 16668 20904 16720
rect 20956 16708 20962 16720
rect 20956 16680 21496 16708
rect 20956 16668 20962 16680
rect 20533 16643 20591 16649
rect 20533 16609 20545 16643
rect 20579 16640 20591 16643
rect 21358 16640 21364 16652
rect 20579 16612 21364 16640
rect 20579 16609 20591 16612
rect 20533 16603 20591 16609
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16541 20131 16575
rect 20073 16535 20131 16541
rect 19904 16504 19932 16535
rect 20162 16532 20168 16584
rect 20220 16532 20226 16584
rect 20254 16532 20260 16584
rect 20312 16532 20318 16584
rect 20346 16532 20352 16584
rect 20404 16532 20410 16584
rect 20806 16532 20812 16584
rect 20864 16532 20870 16584
rect 21174 16532 21180 16584
rect 21232 16532 21238 16584
rect 21468 16581 21496 16680
rect 21818 16668 21824 16720
rect 21876 16708 21882 16720
rect 21876 16680 21956 16708
rect 21876 16668 21882 16680
rect 21634 16600 21640 16652
rect 21692 16640 21698 16652
rect 21729 16643 21787 16649
rect 21729 16640 21741 16643
rect 21692 16612 21741 16640
rect 21692 16600 21698 16612
rect 21729 16609 21741 16612
rect 21775 16609 21787 16643
rect 21729 16603 21787 16609
rect 21928 16581 21956 16680
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 21453 16575 21511 16581
rect 21453 16541 21465 16575
rect 21499 16541 21511 16575
rect 21453 16535 21511 16541
rect 21913 16575 21971 16581
rect 21913 16541 21925 16575
rect 21959 16541 21971 16575
rect 21913 16535 21971 16541
rect 20180 16504 20208 16532
rect 19904 16476 20208 16504
rect 20272 16436 20300 16532
rect 19306 16408 20300 16436
rect 20364 16436 20392 16532
rect 20441 16507 20499 16513
rect 20441 16473 20453 16507
rect 20487 16504 20499 16507
rect 20530 16504 20536 16516
rect 20487 16476 20536 16504
rect 20487 16473 20499 16476
rect 20441 16467 20499 16473
rect 20530 16464 20536 16476
rect 20588 16464 20594 16516
rect 20898 16464 20904 16516
rect 20956 16504 20962 16516
rect 21284 16504 21312 16535
rect 22002 16532 22008 16584
rect 22060 16572 22066 16584
rect 22373 16575 22431 16581
rect 22373 16572 22385 16575
rect 22060 16544 22385 16572
rect 22060 16532 22066 16544
rect 22373 16541 22385 16544
rect 22419 16541 22431 16575
rect 22373 16535 22431 16541
rect 22557 16575 22615 16581
rect 22557 16541 22569 16575
rect 22603 16572 22615 16575
rect 22922 16572 22928 16584
rect 22603 16544 22928 16572
rect 22603 16541 22615 16544
rect 22557 16535 22615 16541
rect 22922 16532 22928 16544
rect 22980 16532 22986 16584
rect 23032 16572 23060 16748
rect 23106 16736 23112 16788
rect 23164 16776 23170 16788
rect 23569 16779 23627 16785
rect 23569 16776 23581 16779
rect 23164 16748 23581 16776
rect 23164 16736 23170 16748
rect 23569 16745 23581 16748
rect 23615 16745 23627 16779
rect 23569 16739 23627 16745
rect 25498 16736 25504 16788
rect 25556 16736 25562 16788
rect 25590 16736 25596 16788
rect 25648 16776 25654 16788
rect 25648 16748 26372 16776
rect 25648 16736 25654 16748
rect 25516 16708 25544 16736
rect 26234 16708 26240 16720
rect 25516 16680 26240 16708
rect 23842 16640 23848 16652
rect 23308 16612 23848 16640
rect 23308 16581 23336 16612
rect 23842 16600 23848 16612
rect 23900 16640 23906 16652
rect 24026 16640 24032 16652
rect 23900 16612 24032 16640
rect 23900 16600 23906 16612
rect 24026 16600 24032 16612
rect 24084 16640 24090 16652
rect 24394 16640 24400 16652
rect 24084 16612 24400 16640
rect 24084 16600 24090 16612
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 25608 16649 25636 16680
rect 26234 16668 26240 16680
rect 26292 16668 26298 16720
rect 25593 16643 25651 16649
rect 25593 16609 25605 16643
rect 25639 16609 25651 16643
rect 25593 16603 25651 16609
rect 25685 16643 25743 16649
rect 25685 16609 25697 16643
rect 25731 16609 25743 16643
rect 26344 16640 26372 16748
rect 26510 16736 26516 16788
rect 26568 16776 26574 16788
rect 26568 16748 27568 16776
rect 26568 16736 26574 16748
rect 26789 16643 26847 16649
rect 26789 16640 26801 16643
rect 26344 16612 26801 16640
rect 25685 16603 25743 16609
rect 26789 16609 26801 16612
rect 26835 16609 26847 16643
rect 26789 16603 26847 16609
rect 23293 16575 23351 16581
rect 23293 16572 23305 16575
rect 23032 16544 23305 16572
rect 23293 16541 23305 16544
rect 23339 16541 23351 16575
rect 23293 16535 23351 16541
rect 23382 16532 23388 16584
rect 23440 16572 23446 16584
rect 23661 16575 23719 16581
rect 23440 16544 23485 16572
rect 23440 16532 23446 16544
rect 23661 16541 23673 16575
rect 23707 16541 23719 16575
rect 23661 16535 23719 16541
rect 21358 16504 21364 16516
rect 20956 16476 21220 16504
rect 21284 16476 21364 16504
rect 20956 16464 20962 16476
rect 20993 16439 21051 16445
rect 20993 16436 21005 16439
rect 20364 16408 21005 16436
rect 17957 16399 18015 16405
rect 20993 16405 21005 16408
rect 21039 16405 21051 16439
rect 21192 16436 21220 16476
rect 21358 16464 21364 16476
rect 21416 16504 21422 16516
rect 22189 16507 22247 16513
rect 22189 16504 22201 16507
rect 21416 16476 22201 16504
rect 21416 16464 21422 16476
rect 22189 16473 22201 16476
rect 22235 16473 22247 16507
rect 23676 16504 23704 16535
rect 24302 16532 24308 16584
rect 24360 16572 24366 16584
rect 25700 16572 25728 16603
rect 26970 16600 26976 16652
rect 27028 16640 27034 16652
rect 27433 16643 27491 16649
rect 27433 16640 27445 16643
rect 27028 16612 27445 16640
rect 27028 16600 27034 16612
rect 27433 16609 27445 16612
rect 27479 16609 27491 16643
rect 27540 16640 27568 16748
rect 29104 16748 29408 16776
rect 28721 16643 28779 16649
rect 27540 16612 28488 16640
rect 27433 16603 27491 16609
rect 24360 16544 25728 16572
rect 26145 16575 26203 16581
rect 24360 16532 24366 16544
rect 26145 16541 26157 16575
rect 26191 16572 26203 16575
rect 26326 16572 26332 16584
rect 26191 16544 26332 16572
rect 26191 16541 26203 16544
rect 26145 16535 26203 16541
rect 26326 16532 26332 16544
rect 26384 16532 26390 16584
rect 26510 16532 26516 16584
rect 26568 16532 26574 16584
rect 26694 16532 26700 16584
rect 26752 16532 26758 16584
rect 27525 16575 27583 16581
rect 27525 16541 27537 16575
rect 27571 16541 27583 16575
rect 27525 16535 27583 16541
rect 24210 16504 24216 16516
rect 22189 16467 22247 16473
rect 22756 16476 23520 16504
rect 23676 16476 24216 16504
rect 22756 16436 22784 16476
rect 23492 16448 23520 16476
rect 24210 16464 24216 16476
rect 24268 16504 24274 16516
rect 26712 16504 26740 16532
rect 27540 16504 27568 16535
rect 27706 16532 27712 16584
rect 27764 16532 27770 16584
rect 28460 16581 28488 16612
rect 28721 16609 28733 16643
rect 28767 16640 28779 16643
rect 28810 16640 28816 16652
rect 28767 16612 28816 16640
rect 28767 16609 28779 16612
rect 28721 16603 28779 16609
rect 28810 16600 28816 16612
rect 28868 16640 28874 16652
rect 29104 16649 29132 16748
rect 29380 16720 29408 16748
rect 29454 16736 29460 16788
rect 29512 16776 29518 16788
rect 30745 16779 30803 16785
rect 30745 16776 30757 16779
rect 29512 16748 30757 16776
rect 29512 16736 29518 16748
rect 30745 16745 30757 16748
rect 30791 16745 30803 16779
rect 30745 16739 30803 16745
rect 30929 16779 30987 16785
rect 30929 16745 30941 16779
rect 30975 16776 30987 16779
rect 33134 16776 33140 16788
rect 30975 16748 33140 16776
rect 30975 16745 30987 16748
rect 30929 16739 30987 16745
rect 29362 16668 29368 16720
rect 29420 16668 29426 16720
rect 29546 16668 29552 16720
rect 29604 16708 29610 16720
rect 29733 16711 29791 16717
rect 29733 16708 29745 16711
rect 29604 16680 29745 16708
rect 29604 16668 29610 16680
rect 29733 16677 29745 16680
rect 29779 16677 29791 16711
rect 29733 16671 29791 16677
rect 30469 16711 30527 16717
rect 30469 16677 30481 16711
rect 30515 16708 30527 16711
rect 30515 16680 32352 16708
rect 30515 16677 30527 16680
rect 30469 16671 30527 16677
rect 28997 16643 29055 16649
rect 28997 16640 29009 16643
rect 28868 16612 29009 16640
rect 28868 16600 28874 16612
rect 28997 16609 29009 16612
rect 29043 16609 29055 16643
rect 28997 16603 29055 16609
rect 29089 16643 29147 16649
rect 29089 16609 29101 16643
rect 29135 16609 29147 16643
rect 29089 16603 29147 16609
rect 29273 16609 29331 16615
rect 28445 16575 28503 16581
rect 28445 16541 28457 16575
rect 28491 16541 28503 16575
rect 28445 16535 28503 16541
rect 24268 16476 26188 16504
rect 26712 16476 27568 16504
rect 24268 16464 24274 16476
rect 21192 16408 22784 16436
rect 20993 16399 21051 16405
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 23109 16439 23167 16445
rect 23109 16436 23121 16439
rect 22888 16408 23121 16436
rect 22888 16396 22894 16408
rect 23109 16405 23121 16408
rect 23155 16405 23167 16439
rect 23109 16399 23167 16405
rect 23474 16396 23480 16448
rect 23532 16396 23538 16448
rect 25130 16396 25136 16448
rect 25188 16396 25194 16448
rect 25501 16439 25559 16445
rect 25501 16405 25513 16439
rect 25547 16436 25559 16439
rect 25590 16436 25596 16448
rect 25547 16408 25596 16436
rect 25547 16405 25559 16408
rect 25501 16399 25559 16405
rect 25590 16396 25596 16408
rect 25648 16396 25654 16448
rect 26050 16396 26056 16448
rect 26108 16396 26114 16448
rect 26160 16436 26188 16476
rect 28166 16464 28172 16516
rect 28224 16464 28230 16516
rect 28460 16504 28488 16535
rect 28534 16532 28540 16584
rect 28592 16572 28598 16584
rect 29181 16575 29239 16581
rect 28592 16544 28637 16572
rect 28592 16532 28598 16544
rect 29181 16541 29193 16575
rect 29227 16541 29239 16575
rect 29273 16575 29285 16609
rect 29319 16575 29331 16609
rect 29638 16600 29644 16652
rect 29696 16600 29702 16652
rect 29748 16640 29776 16671
rect 30098 16640 30104 16652
rect 29748 16612 30104 16640
rect 30098 16600 30104 16612
rect 30156 16600 30162 16652
rect 30190 16600 30196 16652
rect 30248 16640 30254 16652
rect 31021 16643 31079 16649
rect 31021 16640 31033 16643
rect 30248 16612 31033 16640
rect 30248 16600 30254 16612
rect 31021 16609 31033 16612
rect 31067 16609 31079 16643
rect 31021 16603 31079 16609
rect 31294 16600 31300 16652
rect 31352 16640 31358 16652
rect 31389 16643 31447 16649
rect 31389 16640 31401 16643
rect 31352 16612 31401 16640
rect 31352 16600 31358 16612
rect 31389 16609 31401 16612
rect 31435 16609 31447 16643
rect 31389 16603 31447 16609
rect 29273 16574 29331 16575
rect 29273 16569 29408 16574
rect 29656 16572 29684 16600
rect 30926 16572 30932 16584
rect 29288 16562 29408 16569
rect 29564 16562 29684 16572
rect 29288 16546 29684 16562
rect 30806 16547 30932 16572
rect 29181 16535 29239 16541
rect 29380 16544 29684 16546
rect 30791 16544 30932 16547
rect 28460 16476 28948 16504
rect 26786 16436 26792 16448
rect 26160 16408 26792 16436
rect 26786 16396 26792 16408
rect 26844 16396 26850 16448
rect 28718 16396 28724 16448
rect 28776 16436 28782 16448
rect 28813 16439 28871 16445
rect 28813 16436 28825 16439
rect 28776 16408 28825 16436
rect 28776 16396 28782 16408
rect 28813 16405 28825 16408
rect 28859 16405 28871 16439
rect 28920 16436 28948 16476
rect 28994 16436 29000 16448
rect 28920 16408 29000 16436
rect 28813 16399 28871 16405
rect 28994 16396 29000 16408
rect 29052 16396 29058 16448
rect 29196 16436 29224 16535
rect 29380 16534 29592 16544
rect 30791 16541 30849 16544
rect 29733 16507 29791 16513
rect 29733 16504 29745 16507
rect 29472 16476 29745 16504
rect 29472 16448 29500 16476
rect 29733 16473 29745 16476
rect 29779 16473 29791 16507
rect 29733 16467 29791 16473
rect 30098 16464 30104 16516
rect 30156 16504 30162 16516
rect 30561 16507 30619 16513
rect 30561 16504 30573 16507
rect 30156 16476 30573 16504
rect 30156 16464 30162 16476
rect 30561 16473 30573 16476
rect 30607 16473 30619 16507
rect 30791 16507 30803 16541
rect 30837 16507 30849 16541
rect 30926 16532 30932 16544
rect 30984 16532 30990 16584
rect 31202 16532 31208 16584
rect 31260 16532 31266 16584
rect 32324 16581 32352 16680
rect 32968 16640 32996 16748
rect 33134 16736 33140 16748
rect 33192 16736 33198 16788
rect 33229 16779 33287 16785
rect 33229 16745 33241 16779
rect 33275 16776 33287 16779
rect 34514 16776 34520 16788
rect 33275 16748 34520 16776
rect 33275 16745 33287 16748
rect 33229 16739 33287 16745
rect 34514 16736 34520 16748
rect 34572 16736 34578 16788
rect 38470 16776 38476 16788
rect 37752 16748 38476 16776
rect 33045 16711 33103 16717
rect 33045 16677 33057 16711
rect 33091 16708 33103 16711
rect 34606 16708 34612 16720
rect 33091 16680 34612 16708
rect 33091 16677 33103 16680
rect 33045 16671 33103 16677
rect 33505 16643 33563 16649
rect 32968 16612 33088 16640
rect 31481 16575 31539 16581
rect 31481 16541 31493 16575
rect 31527 16541 31539 16575
rect 31481 16535 31539 16541
rect 32309 16575 32367 16581
rect 32309 16541 32321 16575
rect 32355 16541 32367 16575
rect 32309 16535 32367 16541
rect 32769 16575 32827 16581
rect 32769 16541 32781 16575
rect 32815 16541 32827 16575
rect 32769 16535 32827 16541
rect 30791 16501 30849 16507
rect 30561 16467 30619 16473
rect 31018 16464 31024 16516
rect 31076 16504 31082 16516
rect 31496 16504 31524 16535
rect 31076 16476 31524 16504
rect 31076 16464 31082 16476
rect 32324 16448 32352 16535
rect 32401 16507 32459 16513
rect 32401 16473 32413 16507
rect 32447 16504 32459 16507
rect 32784 16504 32812 16535
rect 32950 16532 32956 16584
rect 33008 16532 33014 16584
rect 32447 16476 32812 16504
rect 33060 16504 33088 16612
rect 33505 16609 33517 16643
rect 33551 16640 33563 16643
rect 33594 16640 33600 16652
rect 33551 16612 33600 16640
rect 33551 16609 33563 16612
rect 33505 16603 33563 16609
rect 33594 16600 33600 16612
rect 33652 16600 33658 16652
rect 33410 16581 33416 16584
rect 33137 16575 33195 16581
rect 33137 16541 33149 16575
rect 33183 16572 33195 16575
rect 33401 16575 33416 16581
rect 33401 16572 33413 16575
rect 33183 16544 33413 16572
rect 33183 16541 33195 16544
rect 33137 16535 33195 16541
rect 33401 16541 33413 16544
rect 33401 16535 33416 16541
rect 33410 16532 33416 16535
rect 33468 16532 33474 16584
rect 33873 16575 33931 16581
rect 33873 16572 33885 16575
rect 33612 16544 33885 16572
rect 33612 16504 33640 16544
rect 33873 16541 33885 16544
rect 33919 16572 33931 16575
rect 33962 16572 33968 16584
rect 33919 16544 33968 16572
rect 33919 16541 33931 16544
rect 33873 16535 33931 16541
rect 33962 16532 33968 16544
rect 34020 16532 34026 16584
rect 34072 16572 34100 16680
rect 34606 16668 34612 16680
rect 34664 16668 34670 16720
rect 34241 16575 34299 16581
rect 34241 16572 34253 16575
rect 34072 16544 34253 16572
rect 34241 16541 34253 16544
rect 34287 16541 34299 16575
rect 34241 16535 34299 16541
rect 34425 16575 34483 16581
rect 34425 16541 34437 16575
rect 34471 16541 34483 16575
rect 34425 16535 34483 16541
rect 35897 16575 35955 16581
rect 35897 16541 35909 16575
rect 35943 16572 35955 16575
rect 35986 16572 35992 16584
rect 35943 16544 35992 16572
rect 35943 16541 35955 16544
rect 35897 16535 35955 16541
rect 34440 16504 34468 16535
rect 35986 16532 35992 16544
rect 36044 16572 36050 16584
rect 37752 16581 37780 16748
rect 38470 16736 38476 16748
rect 38528 16776 38534 16788
rect 38838 16776 38844 16788
rect 38528 16748 38844 16776
rect 38528 16736 38534 16748
rect 38838 16736 38844 16748
rect 38896 16736 38902 16788
rect 38930 16736 38936 16788
rect 38988 16736 38994 16788
rect 39206 16736 39212 16788
rect 39264 16736 39270 16788
rect 39298 16736 39304 16788
rect 39356 16736 39362 16788
rect 37918 16668 37924 16720
rect 37976 16708 37982 16720
rect 38654 16708 38660 16720
rect 37976 16680 38660 16708
rect 37976 16668 37982 16680
rect 38654 16668 38660 16680
rect 38712 16668 38718 16720
rect 38948 16640 38976 16736
rect 39316 16640 39344 16736
rect 38764 16612 38976 16640
rect 39132 16612 39344 16640
rect 37737 16575 37795 16581
rect 37737 16572 37749 16575
rect 36044 16544 37749 16572
rect 36044 16532 36050 16544
rect 37737 16541 37749 16544
rect 37783 16541 37795 16575
rect 37737 16535 37795 16541
rect 38565 16575 38623 16581
rect 38565 16541 38577 16575
rect 38611 16572 38623 16575
rect 38654 16572 38660 16584
rect 38611 16544 38660 16572
rect 38611 16541 38623 16544
rect 38565 16535 38623 16541
rect 38654 16532 38660 16544
rect 38712 16532 38718 16584
rect 38764 16572 38792 16612
rect 38841 16575 38899 16581
rect 38841 16572 38853 16575
rect 38764 16544 38853 16572
rect 38841 16541 38853 16544
rect 38887 16541 38899 16575
rect 38841 16535 38899 16541
rect 38930 16532 38936 16584
rect 38988 16532 38994 16584
rect 39132 16581 39160 16612
rect 39574 16600 39580 16652
rect 39632 16640 39638 16652
rect 40497 16643 40555 16649
rect 40497 16640 40509 16643
rect 39632 16612 40509 16640
rect 39632 16600 39638 16612
rect 40497 16609 40509 16612
rect 40543 16609 40555 16643
rect 40497 16603 40555 16609
rect 40586 16600 40592 16652
rect 40644 16600 40650 16652
rect 39117 16575 39175 16581
rect 39117 16541 39129 16575
rect 39163 16541 39175 16575
rect 39117 16535 39175 16541
rect 39209 16575 39267 16581
rect 39209 16541 39221 16575
rect 39255 16572 39267 16575
rect 39255 16544 39344 16572
rect 39255 16541 39267 16544
rect 39209 16535 39267 16541
rect 39316 16516 39344 16544
rect 39390 16532 39396 16584
rect 39448 16532 39454 16584
rect 39669 16575 39727 16581
rect 39669 16541 39681 16575
rect 39715 16572 39727 16575
rect 40405 16575 40463 16581
rect 39715 16544 40080 16572
rect 39715 16541 39727 16544
rect 39669 16535 39727 16541
rect 33060 16476 33640 16504
rect 33888 16476 34468 16504
rect 38749 16507 38807 16513
rect 32447 16473 32459 16476
rect 32401 16467 32459 16473
rect 33888 16448 33916 16476
rect 38749 16473 38761 16507
rect 38795 16473 38807 16507
rect 38749 16467 38807 16473
rect 29454 16436 29460 16448
rect 29196 16408 29460 16436
rect 29454 16396 29460 16408
rect 29512 16396 29518 16448
rect 29638 16396 29644 16448
rect 29696 16436 29702 16448
rect 30285 16439 30343 16445
rect 30285 16436 30297 16439
rect 29696 16408 30297 16436
rect 29696 16396 29702 16408
rect 30285 16405 30297 16408
rect 30331 16405 30343 16439
rect 30285 16399 30343 16405
rect 31294 16396 31300 16448
rect 31352 16436 31358 16448
rect 31662 16436 31668 16448
rect 31352 16408 31668 16436
rect 31352 16396 31358 16408
rect 31662 16396 31668 16408
rect 31720 16396 31726 16448
rect 32306 16396 32312 16448
rect 32364 16396 32370 16448
rect 33502 16396 33508 16448
rect 33560 16436 33566 16448
rect 33597 16439 33655 16445
rect 33597 16436 33609 16439
rect 33560 16408 33609 16436
rect 33560 16396 33566 16408
rect 33597 16405 33609 16408
rect 33643 16405 33655 16439
rect 33597 16399 33655 16405
rect 33778 16396 33784 16448
rect 33836 16396 33842 16448
rect 33870 16396 33876 16448
rect 33928 16396 33934 16448
rect 34422 16396 34428 16448
rect 34480 16396 34486 16448
rect 34514 16396 34520 16448
rect 34572 16436 34578 16448
rect 35894 16436 35900 16448
rect 34572 16408 35900 16436
rect 34572 16396 34578 16408
rect 35894 16396 35900 16408
rect 35952 16436 35958 16448
rect 35989 16439 36047 16445
rect 35989 16436 36001 16439
rect 35952 16408 36001 16436
rect 35952 16396 35958 16408
rect 35989 16405 36001 16408
rect 36035 16405 36047 16439
rect 35989 16399 36047 16405
rect 36538 16396 36544 16448
rect 36596 16436 36602 16448
rect 37734 16436 37740 16448
rect 36596 16408 37740 16436
rect 36596 16396 36602 16408
rect 37734 16396 37740 16408
rect 37792 16396 37798 16448
rect 37921 16439 37979 16445
rect 37921 16405 37933 16439
rect 37967 16436 37979 16439
rect 38470 16436 38476 16448
rect 37967 16408 38476 16436
rect 37967 16405 37979 16408
rect 37921 16399 37979 16405
rect 38470 16396 38476 16408
rect 38528 16396 38534 16448
rect 38654 16396 38660 16448
rect 38712 16445 38718 16448
rect 38712 16399 38721 16445
rect 38764 16436 38792 16467
rect 39298 16464 39304 16516
rect 39356 16464 39362 16516
rect 38838 16436 38844 16448
rect 38764 16408 38844 16436
rect 38712 16396 38718 16399
rect 38838 16396 38844 16408
rect 38896 16396 38902 16448
rect 39025 16439 39083 16445
rect 39025 16405 39037 16439
rect 39071 16436 39083 16439
rect 39408 16436 39436 16532
rect 39071 16408 39436 16436
rect 39071 16405 39083 16408
rect 39025 16399 39083 16405
rect 39482 16396 39488 16448
rect 39540 16396 39546 16448
rect 40052 16445 40080 16544
rect 40405 16541 40417 16575
rect 40451 16572 40463 16575
rect 41046 16572 41052 16584
rect 40451 16544 41052 16572
rect 40451 16541 40463 16544
rect 40405 16535 40463 16541
rect 41046 16532 41052 16544
rect 41104 16532 41110 16584
rect 40037 16439 40095 16445
rect 40037 16405 40049 16439
rect 40083 16405 40095 16439
rect 40037 16399 40095 16405
rect 1104 16346 41400 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 41400 16346
rect 1104 16272 41400 16294
rect 4338 16232 4344 16244
rect 3896 16204 4344 16232
rect 1394 16056 1400 16108
rect 1452 16056 1458 16108
rect 3786 16056 3792 16108
rect 3844 16056 3850 16108
rect 3896 16105 3924 16204
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 5258 16192 5264 16244
rect 5316 16192 5322 16244
rect 5902 16192 5908 16244
rect 5960 16232 5966 16244
rect 5960 16204 6040 16232
rect 5960 16192 5966 16204
rect 6012 16173 6040 16204
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 7558 16232 7564 16244
rect 7432 16204 7564 16232
rect 7432 16192 7438 16204
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 7650 16192 7656 16244
rect 7708 16192 7714 16244
rect 9401 16235 9459 16241
rect 9401 16201 9413 16235
rect 9447 16232 9459 16235
rect 9582 16232 9588 16244
rect 9447 16204 9588 16232
rect 9447 16201 9459 16204
rect 9401 16195 9459 16201
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 11885 16235 11943 16241
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 12342 16232 12348 16244
rect 11931 16204 12348 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 15194 16192 15200 16244
rect 15252 16232 15258 16244
rect 15470 16232 15476 16244
rect 15252 16204 15476 16232
rect 15252 16192 15258 16204
rect 5077 16167 5135 16173
rect 3988 16136 4292 16164
rect 3881 16099 3939 16105
rect 3881 16065 3893 16099
rect 3927 16065 3939 16099
rect 3881 16059 3939 16065
rect 3605 16031 3663 16037
rect 3605 15997 3617 16031
rect 3651 16028 3663 16031
rect 3988 16028 4016 16136
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 3651 16000 4016 16028
rect 4080 16028 4108 16059
rect 4154 16056 4160 16108
rect 4212 16056 4218 16108
rect 4264 16105 4292 16136
rect 5077 16133 5089 16167
rect 5123 16164 5135 16167
rect 5997 16167 6055 16173
rect 5997 16164 6009 16167
rect 5123 16136 6009 16164
rect 5123 16133 5135 16136
rect 5077 16127 5135 16133
rect 5997 16133 6009 16136
rect 6043 16133 6055 16167
rect 7668 16164 7696 16192
rect 5997 16127 6055 16133
rect 6748 16136 7696 16164
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16065 4307 16099
rect 4614 16096 4620 16108
rect 4249 16059 4307 16065
rect 4356 16068 4620 16096
rect 4356 16028 4384 16068
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16096 5319 16099
rect 5353 16099 5411 16105
rect 5307 16065 5320 16096
rect 5261 16059 5320 16065
rect 5353 16065 5365 16099
rect 5399 16096 5411 16099
rect 5718 16096 5724 16108
rect 5399 16068 5724 16096
rect 5399 16065 5411 16068
rect 5353 16059 5411 16065
rect 4080 16000 4384 16028
rect 3651 15997 3663 16000
rect 3605 15991 3663 15997
rect 4522 15988 4528 16040
rect 4580 15988 4586 16040
rect 4890 15960 4896 15972
rect 4632 15932 4896 15960
rect 4632 15904 4660 15932
rect 4890 15920 4896 15932
rect 4948 15920 4954 15972
rect 5292 15960 5320 16059
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 5905 16099 5963 16105
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 6546 16096 6552 16108
rect 5951 16068 6552 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 5537 16031 5595 16037
rect 5537 15997 5549 16031
rect 5583 16028 5595 16031
rect 5626 16028 5632 16040
rect 5583 16000 5632 16028
rect 5583 15997 5595 16000
rect 5537 15991 5595 15997
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 5920 15960 5948 16059
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 6748 16105 6776 16136
rect 9030 16124 9036 16176
rect 9088 16164 9094 16176
rect 14550 16164 14556 16176
rect 9088 16136 11100 16164
rect 9088 16124 9094 16136
rect 9232 16108 9260 16136
rect 11072 16108 11100 16136
rect 11900 16136 14556 16164
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 15997 6883 16031
rect 7208 16028 7236 16059
rect 7466 16056 7472 16108
rect 7524 16056 7530 16108
rect 7558 16056 7564 16108
rect 7616 16056 7622 16108
rect 9214 16056 9220 16108
rect 9272 16056 9278 16108
rect 9398 16056 9404 16108
rect 9456 16056 9462 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11149 16099 11207 16105
rect 11149 16096 11161 16099
rect 11112 16068 11161 16096
rect 11112 16056 11118 16068
rect 11149 16065 11161 16068
rect 11195 16096 11207 16099
rect 11330 16096 11336 16108
rect 11195 16068 11336 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 11422 16056 11428 16108
rect 11480 16096 11486 16108
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 11480 16068 11529 16096
rect 11480 16056 11486 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16065 11759 16099
rect 11900 16096 11928 16136
rect 14550 16124 14556 16136
rect 14608 16124 14614 16176
rect 15396 16173 15424 16204
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 15749 16235 15807 16241
rect 15749 16201 15761 16235
rect 15795 16232 15807 16235
rect 15838 16232 15844 16244
rect 15795 16204 15844 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 15930 16192 15936 16244
rect 15988 16232 15994 16244
rect 16482 16232 16488 16244
rect 15988 16204 16488 16232
rect 15988 16192 15994 16204
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 17037 16235 17095 16241
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 17218 16232 17224 16244
rect 17083 16204 17224 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 17218 16192 17224 16204
rect 17276 16232 17282 16244
rect 17402 16232 17408 16244
rect 17276 16204 17408 16232
rect 17276 16192 17282 16204
rect 17402 16192 17408 16204
rect 17460 16192 17466 16244
rect 18138 16192 18144 16244
rect 18196 16232 18202 16244
rect 18325 16235 18383 16241
rect 18325 16232 18337 16235
rect 18196 16204 18337 16232
rect 18196 16192 18202 16204
rect 18325 16201 18337 16204
rect 18371 16201 18383 16235
rect 18325 16195 18383 16201
rect 20346 16192 20352 16244
rect 20404 16192 20410 16244
rect 20625 16235 20683 16241
rect 20625 16201 20637 16235
rect 20671 16232 20683 16235
rect 20898 16232 20904 16244
rect 20671 16204 20904 16232
rect 20671 16201 20683 16204
rect 20625 16195 20683 16201
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 22388 16204 24716 16232
rect 15381 16167 15439 16173
rect 15381 16133 15393 16167
rect 15427 16133 15439 16167
rect 20364 16164 20392 16192
rect 20717 16167 20775 16173
rect 20717 16164 20729 16167
rect 20364 16136 20729 16164
rect 15381 16127 15439 16133
rect 20717 16133 20729 16136
rect 20763 16133 20775 16167
rect 21177 16167 21235 16173
rect 21177 16164 21189 16167
rect 20717 16127 20775 16133
rect 20824 16136 21189 16164
rect 20824 16108 20852 16136
rect 21177 16133 21189 16136
rect 21223 16133 21235 16167
rect 21177 16127 21235 16133
rect 21358 16124 21364 16176
rect 21416 16124 21422 16176
rect 11977 16099 12035 16105
rect 11977 16096 11989 16099
rect 11900 16068 11989 16096
rect 11701 16059 11759 16065
rect 11977 16065 11989 16068
rect 12023 16065 12035 16099
rect 11977 16059 12035 16065
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 7837 16031 7895 16037
rect 7208 16000 7788 16028
rect 6825 15991 6883 15997
rect 5292 15932 5948 15960
rect 6454 15920 6460 15972
rect 6512 15960 6518 15972
rect 6638 15960 6644 15972
rect 6512 15932 6644 15960
rect 6512 15920 6518 15932
rect 6638 15920 6644 15932
rect 6696 15960 6702 15972
rect 6840 15960 6868 15991
rect 7193 15963 7251 15969
rect 7193 15960 7205 15963
rect 6696 15932 6868 15960
rect 6932 15932 7205 15960
rect 6696 15920 6702 15932
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 992 15864 1593 15892
rect 992 15852 998 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 4614 15852 4620 15904
rect 4672 15852 4678 15904
rect 4798 15852 4804 15904
rect 4856 15852 4862 15904
rect 6932 15901 6960 15932
rect 7193 15929 7205 15932
rect 7239 15929 7251 15963
rect 7193 15923 7251 15929
rect 7466 15920 7472 15972
rect 7524 15960 7530 15972
rect 7760 15969 7788 16000
rect 7837 15997 7849 16031
rect 7883 16028 7895 16031
rect 11716 16028 11744 16059
rect 11882 16028 11888 16040
rect 7883 16000 8156 16028
rect 11716 16000 11888 16028
rect 7883 15997 7895 16000
rect 7837 15991 7895 15997
rect 7653 15963 7711 15969
rect 7653 15960 7665 15963
rect 7524 15932 7665 15960
rect 7524 15920 7530 15932
rect 7653 15929 7665 15932
rect 7699 15929 7711 15963
rect 7653 15923 7711 15929
rect 7745 15963 7803 15969
rect 7745 15929 7757 15963
rect 7791 15929 7803 15963
rect 7745 15923 7803 15929
rect 8128 15904 8156 16000
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 11241 15963 11299 15969
rect 11241 15929 11253 15963
rect 11287 15960 11299 15963
rect 12176 15960 12204 16059
rect 12250 16056 12256 16108
rect 12308 16056 12314 16108
rect 12342 16056 12348 16108
rect 12400 16056 12406 16108
rect 13998 16056 14004 16108
rect 14056 16096 14062 16108
rect 15197 16099 15255 16105
rect 15197 16096 15209 16099
rect 14056 16068 15209 16096
rect 14056 16056 14062 16068
rect 15197 16065 15209 16068
rect 15243 16096 15255 16099
rect 15286 16096 15292 16108
rect 15243 16068 15292 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15470 16056 15476 16108
rect 15528 16056 15534 16108
rect 15565 16099 15623 16105
rect 15565 16065 15577 16099
rect 15611 16096 15623 16099
rect 15746 16096 15752 16108
rect 15611 16068 15752 16096
rect 15611 16065 15623 16068
rect 15565 16059 15623 16065
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16096 16727 16099
rect 17770 16096 17776 16108
rect 16715 16068 17776 16096
rect 16715 16065 16727 16068
rect 16669 16059 16727 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 18138 16056 18144 16108
rect 18196 16094 18202 16108
rect 18196 16066 18239 16094
rect 18196 16056 18202 16066
rect 20530 16056 20536 16108
rect 20588 16096 20594 16108
rect 20806 16096 20812 16108
rect 20588 16068 20812 16096
rect 20588 16056 20594 16068
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 20898 16056 20904 16108
rect 20956 16056 20962 16108
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21082 16096 21088 16108
rect 21039 16068 21088 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 21082 16056 21088 16068
rect 21140 16096 21146 16108
rect 21376 16096 21404 16124
rect 22388 16108 22416 16204
rect 23293 16167 23351 16173
rect 23293 16164 23305 16167
rect 22940 16136 23305 16164
rect 21140 16068 21404 16096
rect 21140 16056 21146 16068
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 22738 16056 22744 16108
rect 22796 16096 22802 16108
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22796 16068 22845 16096
rect 22796 16056 22802 16068
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 17310 15988 17316 16040
rect 17368 16028 17374 16040
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 17368 16000 17969 16028
rect 17368 15988 17374 16000
rect 17957 15997 17969 16000
rect 18003 16028 18015 16031
rect 18003 16000 18276 16028
rect 18003 15997 18015 16000
rect 17957 15991 18015 15997
rect 11287 15932 12204 15960
rect 11287 15929 11299 15932
rect 11241 15923 11299 15929
rect 18248 15904 18276 16000
rect 18414 15988 18420 16040
rect 18472 16028 18478 16040
rect 20714 16028 20720 16040
rect 18472 16000 20720 16028
rect 18472 15988 18478 16000
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 20916 16028 20944 16056
rect 22940 16040 22968 16136
rect 23293 16133 23305 16136
rect 23339 16133 23351 16167
rect 23293 16127 23351 16133
rect 23509 16167 23567 16173
rect 23509 16133 23521 16167
rect 23555 16164 23567 16167
rect 23658 16164 23664 16176
rect 23555 16136 23664 16164
rect 23555 16133 23567 16136
rect 23509 16127 23567 16133
rect 23658 16124 23664 16136
rect 23716 16164 23722 16176
rect 24688 16173 24716 16204
rect 25130 16192 25136 16244
rect 25188 16192 25194 16244
rect 26234 16192 26240 16244
rect 26292 16192 26298 16244
rect 26326 16192 26332 16244
rect 26384 16232 26390 16244
rect 26697 16235 26755 16241
rect 26697 16232 26709 16235
rect 26384 16204 26709 16232
rect 26384 16192 26390 16204
rect 26697 16201 26709 16204
rect 26743 16201 26755 16235
rect 26697 16195 26755 16201
rect 26786 16192 26792 16244
rect 26844 16232 26850 16244
rect 39206 16232 39212 16244
rect 26844 16204 39212 16232
rect 26844 16192 26850 16204
rect 24489 16167 24547 16173
rect 24489 16164 24501 16167
rect 23716 16136 24501 16164
rect 23716 16124 23722 16136
rect 24489 16133 24501 16136
rect 24535 16133 24547 16167
rect 24489 16127 24547 16133
rect 24673 16167 24731 16173
rect 24673 16133 24685 16167
rect 24719 16133 24731 16167
rect 25148 16164 25176 16192
rect 25148 16136 25912 16164
rect 24673 16127 24731 16133
rect 23106 16056 23112 16108
rect 23164 16096 23170 16108
rect 23382 16096 23388 16108
rect 23164 16068 23388 16096
rect 23164 16056 23170 16068
rect 23382 16056 23388 16068
rect 23440 16056 23446 16108
rect 21174 16028 21180 16040
rect 20916 16000 21180 16028
rect 21174 15988 21180 16000
rect 21232 15988 21238 16040
rect 21361 16031 21419 16037
rect 21361 15997 21373 16031
rect 21407 16028 21419 16031
rect 21407 16000 22877 16028
rect 21407 15997 21419 16000
rect 21361 15991 21419 15997
rect 20180 15932 20852 15960
rect 20180 15904 20208 15932
rect 6917 15895 6975 15901
rect 6917 15861 6929 15895
rect 6963 15861 6975 15895
rect 6917 15855 6975 15861
rect 7098 15852 7104 15904
rect 7156 15852 7162 15904
rect 8110 15852 8116 15904
rect 8168 15852 8174 15904
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 11977 15895 12035 15901
rect 11977 15892 11989 15895
rect 11848 15864 11989 15892
rect 11848 15852 11854 15864
rect 11977 15861 11989 15864
rect 12023 15861 12035 15895
rect 11977 15855 12035 15861
rect 17034 15852 17040 15904
rect 17092 15852 17098 15904
rect 17218 15852 17224 15904
rect 17276 15852 17282 15904
rect 18230 15852 18236 15904
rect 18288 15852 18294 15904
rect 20162 15852 20168 15904
rect 20220 15852 20226 15904
rect 20254 15852 20260 15904
rect 20312 15852 20318 15904
rect 20824 15892 20852 15932
rect 20898 15920 20904 15972
rect 20956 15960 20962 15972
rect 21910 15960 21916 15972
rect 20956 15932 21916 15960
rect 20956 15920 20962 15932
rect 21910 15920 21916 15932
rect 21968 15920 21974 15972
rect 22849 15960 22877 16000
rect 22922 15988 22928 16040
rect 22980 15988 22986 16040
rect 23017 16031 23075 16037
rect 23017 15997 23029 16031
rect 23063 16028 23075 16031
rect 24026 16028 24032 16040
rect 23063 16000 24032 16028
rect 23063 15997 23075 16000
rect 23017 15991 23075 15997
rect 23032 15960 23060 15991
rect 24026 15988 24032 16000
rect 24084 16028 24090 16040
rect 24302 16028 24308 16040
rect 24084 16000 24308 16028
rect 24084 15988 24090 16000
rect 24302 15988 24308 16000
rect 24360 15988 24366 16040
rect 24504 16028 24532 16127
rect 24762 16056 24768 16108
rect 24820 16096 24826 16108
rect 25501 16099 25559 16105
rect 25501 16096 25513 16099
rect 24820 16068 25513 16096
rect 24820 16056 24826 16068
rect 25501 16065 25513 16068
rect 25547 16065 25559 16099
rect 25501 16059 25559 16065
rect 25682 16056 25688 16108
rect 25740 16056 25746 16108
rect 25884 16105 25912 16136
rect 25869 16099 25927 16105
rect 25869 16065 25881 16099
rect 25915 16065 25927 16099
rect 26252 16096 26280 16192
rect 26421 16167 26479 16173
rect 26421 16133 26433 16167
rect 26467 16164 26479 16167
rect 27341 16167 27399 16173
rect 27341 16164 27353 16167
rect 26467 16136 27353 16164
rect 26467 16133 26479 16136
rect 26421 16127 26479 16133
rect 27341 16133 27353 16136
rect 27387 16133 27399 16167
rect 27341 16127 27399 16133
rect 28905 16167 28963 16173
rect 28905 16133 28917 16167
rect 28951 16164 28963 16167
rect 29086 16164 29092 16176
rect 28951 16136 29092 16164
rect 28951 16133 28963 16136
rect 28905 16127 28963 16133
rect 29086 16124 29092 16136
rect 29144 16124 29150 16176
rect 29178 16124 29184 16176
rect 29236 16164 29242 16176
rect 29365 16167 29423 16173
rect 29365 16164 29377 16167
rect 29236 16136 29377 16164
rect 29236 16124 29242 16136
rect 29365 16133 29377 16136
rect 29411 16133 29423 16167
rect 29822 16164 29828 16176
rect 29365 16127 29423 16133
rect 29656 16136 29828 16164
rect 26329 16099 26387 16105
rect 26329 16096 26341 16099
rect 26252 16068 26341 16096
rect 25869 16059 25927 16065
rect 26329 16065 26341 16068
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 26605 16099 26663 16105
rect 26605 16065 26617 16099
rect 26651 16096 26663 16099
rect 26694 16096 26700 16108
rect 26651 16068 26700 16096
rect 26651 16065 26663 16068
rect 26605 16059 26663 16065
rect 26694 16056 26700 16068
rect 26752 16056 26758 16108
rect 26786 16056 26792 16108
rect 26844 16056 26850 16108
rect 26973 16099 27031 16105
rect 26973 16065 26985 16099
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 27066 16099 27124 16105
rect 27066 16065 27078 16099
rect 27112 16065 27124 16099
rect 27066 16059 27124 16065
rect 25593 16031 25651 16037
rect 24504 16000 25544 16028
rect 22849 15932 23060 15960
rect 22370 15892 22376 15904
rect 20824 15864 22376 15892
rect 22370 15852 22376 15864
rect 22428 15852 22434 15904
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 22649 15895 22707 15901
rect 22649 15892 22661 15895
rect 22612 15864 22661 15892
rect 22612 15852 22618 15864
rect 22649 15861 22661 15864
rect 22695 15861 22707 15895
rect 22649 15855 22707 15861
rect 22738 15852 22744 15904
rect 22796 15892 22802 15904
rect 23477 15895 23535 15901
rect 23477 15892 23489 15895
rect 22796 15864 23489 15892
rect 22796 15852 22802 15864
rect 23477 15861 23489 15864
rect 23523 15861 23535 15895
rect 23477 15855 23535 15861
rect 23658 15852 23664 15904
rect 23716 15852 23722 15904
rect 24302 15852 24308 15904
rect 24360 15892 24366 15904
rect 24762 15892 24768 15904
rect 24360 15864 24768 15892
rect 24360 15852 24366 15864
rect 24762 15852 24768 15864
rect 24820 15892 24826 15904
rect 24857 15895 24915 15901
rect 24857 15892 24869 15895
rect 24820 15864 24869 15892
rect 24820 15852 24826 15864
rect 24857 15861 24869 15864
rect 24903 15861 24915 15895
rect 25516 15892 25544 16000
rect 25593 15997 25605 16031
rect 25639 16028 25651 16031
rect 26988 16028 27016 16059
rect 25639 16000 27016 16028
rect 25639 15997 25651 16000
rect 25593 15991 25651 15997
rect 25961 15963 26019 15969
rect 25961 15929 25973 15963
rect 26007 15960 26019 15963
rect 26602 15960 26608 15972
rect 26007 15932 26608 15960
rect 26007 15929 26019 15932
rect 25961 15923 26019 15929
rect 26602 15920 26608 15932
rect 26660 15920 26666 15972
rect 26694 15920 26700 15972
rect 26752 15960 26758 15972
rect 27080 15960 27108 16059
rect 27246 16056 27252 16108
rect 27304 16056 27310 16108
rect 27438 16099 27496 16105
rect 27438 16096 27450 16099
rect 27356 16068 27450 16096
rect 26752 15932 27108 15960
rect 26752 15920 26758 15932
rect 27356 15892 27384 16068
rect 27438 16065 27450 16068
rect 27484 16065 27496 16099
rect 27438 16059 27496 16065
rect 28534 16056 28540 16108
rect 28592 16096 28598 16108
rect 28813 16099 28871 16105
rect 28813 16096 28825 16099
rect 28592 16068 28825 16096
rect 28592 16056 28598 16068
rect 28813 16065 28825 16068
rect 28859 16065 28871 16099
rect 28813 16059 28871 16065
rect 28994 16056 29000 16108
rect 29052 16056 29058 16108
rect 29656 16105 29684 16136
rect 29822 16124 29828 16136
rect 29880 16164 29886 16176
rect 30650 16164 30656 16176
rect 29880 16136 30656 16164
rect 29880 16124 29886 16136
rect 30650 16124 30656 16136
rect 30708 16164 30714 16176
rect 34514 16164 34520 16176
rect 30708 16136 34520 16164
rect 30708 16124 30714 16136
rect 33612 16108 33640 16136
rect 34514 16124 34520 16136
rect 34572 16124 34578 16176
rect 36909 16167 36967 16173
rect 35728 16136 36860 16164
rect 29532 16099 29590 16105
rect 29532 16096 29544 16099
rect 29472 16068 29544 16096
rect 29472 16028 29500 16068
rect 29532 16065 29544 16068
rect 29578 16065 29590 16099
rect 29532 16059 29590 16065
rect 29642 16099 29700 16105
rect 29642 16065 29654 16099
rect 29688 16065 29700 16099
rect 29642 16059 29700 16065
rect 29730 16056 29736 16108
rect 29788 16056 29794 16108
rect 29914 16056 29920 16108
rect 29972 16056 29978 16108
rect 32571 16099 32629 16105
rect 32571 16065 32583 16099
rect 32617 16096 32629 16099
rect 32766 16096 32772 16108
rect 32617 16068 32772 16096
rect 32617 16065 32629 16068
rect 32571 16059 32629 16065
rect 32766 16056 32772 16068
rect 32824 16056 32830 16108
rect 33505 16099 33563 16105
rect 33505 16096 33517 16099
rect 32876 16068 33517 16096
rect 29748 16028 29776 16056
rect 29472 16000 29776 16028
rect 30926 15988 30932 16040
rect 30984 15988 30990 16040
rect 32306 15988 32312 16040
rect 32364 16028 32370 16040
rect 32401 16031 32459 16037
rect 32401 16028 32413 16031
rect 32364 16000 32413 16028
rect 32364 15988 32370 16000
rect 32401 15997 32413 16000
rect 32447 15997 32459 16031
rect 32401 15991 32459 15997
rect 29638 15960 29644 15972
rect 27632 15932 29644 15960
rect 27632 15901 27660 15932
rect 29638 15920 29644 15932
rect 29696 15920 29702 15972
rect 29825 15963 29883 15969
rect 29825 15929 29837 15963
rect 29871 15960 29883 15963
rect 30944 15960 30972 15988
rect 32876 15969 32904 16068
rect 33505 16065 33517 16068
rect 33551 16065 33563 16099
rect 33505 16059 33563 16065
rect 33594 16056 33600 16108
rect 33652 16056 33658 16108
rect 33870 16056 33876 16108
rect 33928 16056 33934 16108
rect 33962 16056 33968 16108
rect 34020 16056 34026 16108
rect 34149 16099 34207 16105
rect 34149 16065 34161 16099
rect 34195 16096 34207 16099
rect 34238 16096 34244 16108
rect 34195 16068 34244 16096
rect 34195 16065 34207 16068
rect 34149 16059 34207 16065
rect 34238 16056 34244 16068
rect 34296 16056 34302 16108
rect 34422 16056 34428 16108
rect 34480 16056 34486 16108
rect 34609 16099 34667 16105
rect 34609 16065 34621 16099
rect 34655 16065 34667 16099
rect 34609 16059 34667 16065
rect 33410 15988 33416 16040
rect 33468 16028 33474 16040
rect 33888 16028 33916 16056
rect 33468 16000 33916 16028
rect 34440 16028 34468 16056
rect 34517 16031 34575 16037
rect 34517 16028 34529 16031
rect 34440 16000 34529 16028
rect 33468 15988 33474 16000
rect 34517 15997 34529 16000
rect 34563 15997 34575 16031
rect 34517 15991 34575 15997
rect 29871 15932 30972 15960
rect 32861 15963 32919 15969
rect 29871 15929 29883 15932
rect 29825 15923 29883 15929
rect 32861 15929 32873 15963
rect 32907 15929 32919 15963
rect 32861 15923 32919 15929
rect 25516 15864 27384 15892
rect 27617 15895 27675 15901
rect 24857 15855 24915 15861
rect 27617 15861 27629 15895
rect 27663 15861 27675 15895
rect 27617 15855 27675 15861
rect 28810 15852 28816 15904
rect 28868 15892 28874 15904
rect 29840 15892 29868 15923
rect 34238 15920 34244 15972
rect 34296 15960 34302 15972
rect 34624 15960 34652 16059
rect 34698 16056 34704 16108
rect 34756 16056 34762 16108
rect 34716 16028 34744 16056
rect 35728 16028 35756 16136
rect 36832 16108 36860 16136
rect 36909 16133 36921 16167
rect 36955 16164 36967 16167
rect 36955 16136 37780 16164
rect 36955 16133 36967 16136
rect 36909 16127 36967 16133
rect 36449 16099 36507 16105
rect 36449 16065 36461 16099
rect 36495 16065 36507 16099
rect 36449 16059 36507 16065
rect 34716 16000 35756 16028
rect 36464 16028 36492 16059
rect 36814 16056 36820 16108
rect 36872 16056 36878 16108
rect 37001 16099 37059 16105
rect 37001 16065 37013 16099
rect 37047 16065 37059 16099
rect 37001 16059 37059 16065
rect 37010 16028 37038 16059
rect 37090 16056 37096 16108
rect 37148 16096 37154 16108
rect 37752 16105 37780 16136
rect 37461 16099 37519 16105
rect 37461 16096 37473 16099
rect 37148 16068 37473 16096
rect 37148 16056 37154 16068
rect 37461 16065 37473 16068
rect 37507 16065 37519 16099
rect 37461 16059 37519 16065
rect 37737 16099 37795 16105
rect 37737 16065 37749 16099
rect 37783 16065 37795 16099
rect 37737 16059 37795 16065
rect 37826 16056 37832 16108
rect 37884 16056 37890 16108
rect 38470 16056 38476 16108
rect 38528 16096 38534 16108
rect 38749 16099 38807 16105
rect 38749 16096 38761 16099
rect 38528 16068 38761 16096
rect 38528 16056 38534 16068
rect 38749 16065 38761 16068
rect 38795 16065 38807 16099
rect 38749 16059 38807 16065
rect 37277 16031 37335 16037
rect 37277 16028 37289 16031
rect 36464 16000 37289 16028
rect 37277 15997 37289 16000
rect 37323 16028 37335 16031
rect 38488 16028 38516 16056
rect 37323 16000 38516 16028
rect 38565 16031 38623 16037
rect 37323 15997 37335 16000
rect 37277 15991 37335 15997
rect 38565 15997 38577 16031
rect 38611 16028 38623 16031
rect 38856 16028 38884 16204
rect 39206 16192 39212 16204
rect 39264 16192 39270 16244
rect 39482 16192 39488 16244
rect 39540 16232 39546 16244
rect 39540 16204 39620 16232
rect 39540 16192 39546 16204
rect 39592 16173 39620 16204
rect 40494 16192 40500 16244
rect 40552 16232 40558 16244
rect 41049 16235 41107 16241
rect 41049 16232 41061 16235
rect 40552 16204 41061 16232
rect 40552 16192 40558 16204
rect 41049 16201 41061 16204
rect 41095 16201 41107 16235
rect 41049 16195 41107 16201
rect 39577 16167 39635 16173
rect 39577 16133 39589 16167
rect 39623 16133 39635 16167
rect 39577 16127 39635 16133
rect 40034 16124 40040 16176
rect 40092 16124 40098 16176
rect 38611 16000 38884 16028
rect 38611 15997 38623 16000
rect 38565 15991 38623 15997
rect 39022 15988 39028 16040
rect 39080 16028 39086 16040
rect 39301 16031 39359 16037
rect 39301 16028 39313 16031
rect 39080 16000 39313 16028
rect 39080 15988 39086 16000
rect 39301 15997 39313 16000
rect 39347 15997 39359 16031
rect 39301 15991 39359 15997
rect 34296 15932 34652 15960
rect 34296 15920 34302 15932
rect 36630 15920 36636 15972
rect 36688 15920 36694 15972
rect 37366 15920 37372 15972
rect 37424 15960 37430 15972
rect 38105 15963 38163 15969
rect 38105 15960 38117 15963
rect 37424 15932 38117 15960
rect 37424 15920 37430 15932
rect 38105 15929 38117 15932
rect 38151 15929 38163 15963
rect 38105 15923 38163 15929
rect 28868 15864 29868 15892
rect 33321 15895 33379 15901
rect 28868 15852 28874 15864
rect 33321 15861 33333 15895
rect 33367 15892 33379 15895
rect 33594 15892 33600 15904
rect 33367 15864 33600 15892
rect 33367 15861 33379 15864
rect 33321 15855 33379 15861
rect 33594 15852 33600 15864
rect 33652 15852 33658 15904
rect 33781 15895 33839 15901
rect 33781 15861 33793 15895
rect 33827 15892 33839 15895
rect 33965 15895 34023 15901
rect 33965 15892 33977 15895
rect 33827 15864 33977 15892
rect 33827 15861 33839 15864
rect 33781 15855 33839 15861
rect 33965 15861 33977 15864
rect 34011 15861 34023 15895
rect 33965 15855 34023 15861
rect 34977 15895 35035 15901
rect 34977 15861 34989 15895
rect 35023 15892 35035 15895
rect 35342 15892 35348 15904
rect 35023 15864 35348 15892
rect 35023 15861 35035 15864
rect 34977 15855 35035 15861
rect 35342 15852 35348 15864
rect 35400 15852 35406 15904
rect 37645 15895 37703 15901
rect 37645 15861 37657 15895
rect 37691 15892 37703 15895
rect 37737 15895 37795 15901
rect 37737 15892 37749 15895
rect 37691 15864 37749 15892
rect 37691 15861 37703 15864
rect 37645 15855 37703 15861
rect 37737 15861 37749 15864
rect 37783 15861 37795 15895
rect 37737 15855 37795 15861
rect 38933 15895 38991 15901
rect 38933 15861 38945 15895
rect 38979 15892 38991 15895
rect 39298 15892 39304 15904
rect 38979 15864 39304 15892
rect 38979 15861 38991 15864
rect 38933 15855 38991 15861
rect 39298 15852 39304 15864
rect 39356 15852 39362 15904
rect 1104 15802 41400 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 41400 15802
rect 1104 15728 41400 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1452 15660 1593 15688
rect 1452 15648 1458 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 2028 15691 2086 15697
rect 2028 15657 2040 15691
rect 2074 15688 2086 15691
rect 2074 15660 4016 15688
rect 2074 15657 2086 15660
rect 2028 15651 2086 15657
rect 3988 15620 4016 15660
rect 7098 15648 7104 15700
rect 7156 15648 7162 15700
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 13998 15688 14004 15700
rect 7616 15660 14004 15688
rect 7616 15648 7622 15660
rect 13998 15648 14004 15660
rect 14056 15648 14062 15700
rect 14090 15648 14096 15700
rect 14148 15648 14154 15700
rect 15654 15648 15660 15700
rect 15712 15648 15718 15700
rect 17586 15648 17592 15700
rect 17644 15648 17650 15700
rect 17957 15691 18015 15697
rect 17957 15657 17969 15691
rect 18003 15688 18015 15691
rect 18138 15688 18144 15700
rect 18003 15660 18144 15688
rect 18003 15657 18015 15660
rect 17957 15651 18015 15657
rect 18138 15648 18144 15660
rect 18196 15688 18202 15700
rect 18414 15688 18420 15700
rect 18196 15660 18420 15688
rect 18196 15648 18202 15660
rect 18414 15648 18420 15660
rect 18472 15648 18478 15700
rect 20898 15688 20904 15700
rect 18616 15660 20904 15688
rect 5261 15623 5319 15629
rect 5261 15620 5273 15623
rect 3988 15592 5273 15620
rect 5261 15589 5273 15592
rect 5307 15589 5319 15623
rect 5261 15583 5319 15589
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 2682 15552 2688 15564
rect 1811 15524 2688 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 1780 15484 1808 15515
rect 2682 15512 2688 15524
rect 2740 15512 2746 15564
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15521 3571 15555
rect 3513 15515 3571 15521
rect 1443 15456 1808 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 3050 15444 3056 15496
rect 3108 15484 3114 15496
rect 3528 15484 3556 15515
rect 4798 15512 4804 15564
rect 4856 15512 4862 15564
rect 7116 15552 7144 15648
rect 10778 15580 10784 15632
rect 10836 15580 10842 15632
rect 11974 15620 11980 15632
rect 11164 15592 11980 15620
rect 4908 15524 7144 15552
rect 10413 15555 10471 15561
rect 3970 15484 3976 15496
rect 3108 15456 3174 15484
rect 3528 15456 3976 15484
rect 3108 15444 3114 15456
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 4816 15484 4844 15512
rect 4908 15493 4936 15524
rect 10413 15521 10425 15555
rect 10459 15552 10471 15555
rect 10870 15552 10876 15564
rect 10459 15524 10876 15552
rect 10459 15521 10471 15524
rect 10413 15515 10471 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 4755 15456 4844 15484
rect 4893 15487 4951 15493
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 4893 15447 4951 15453
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 5442 15484 5448 15496
rect 5132 15456 5448 15484
rect 5132 15444 5138 15456
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 11164 15493 11192 15592
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 14108 15552 14136 15648
rect 15672 15620 15700 15648
rect 18616 15620 18644 15660
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 21726 15648 21732 15700
rect 21784 15688 21790 15700
rect 22002 15688 22008 15700
rect 21784 15660 22008 15688
rect 21784 15648 21790 15660
rect 22002 15648 22008 15660
rect 22060 15688 22066 15700
rect 22830 15688 22836 15700
rect 22060 15660 22836 15688
rect 22060 15648 22066 15660
rect 22830 15648 22836 15660
rect 22888 15648 22894 15700
rect 29638 15648 29644 15700
rect 29696 15688 29702 15700
rect 32214 15688 32220 15700
rect 29696 15660 32220 15688
rect 29696 15648 29702 15660
rect 32214 15648 32220 15660
rect 32272 15648 32278 15700
rect 33410 15648 33416 15700
rect 33468 15648 33474 15700
rect 34698 15688 34704 15700
rect 33520 15660 34704 15688
rect 15672 15592 18644 15620
rect 18693 15623 18751 15629
rect 18693 15589 18705 15623
rect 18739 15589 18751 15623
rect 22646 15620 22652 15632
rect 18693 15583 18751 15589
rect 21284 15592 22652 15620
rect 11940 15524 14136 15552
rect 11940 15512 11946 15524
rect 17402 15512 17408 15564
rect 17460 15512 17466 15564
rect 18708 15552 18736 15583
rect 17604 15524 18736 15552
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10888 15456 10977 15484
rect 4985 15419 5043 15425
rect 4985 15385 4997 15419
rect 5031 15385 5043 15419
rect 4985 15379 5043 15385
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15348 4675 15351
rect 5000 15348 5028 15379
rect 4663 15320 5028 15348
rect 4663 15317 4675 15320
rect 4617 15311 4675 15317
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 10888 15357 10916 15456
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15484 11207 15487
rect 11238 15484 11244 15496
rect 11195 15456 11244 15484
rect 11195 15453 11207 15456
rect 11149 15447 11207 15453
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 13354 15444 13360 15496
rect 13412 15444 13418 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 13906 15484 13912 15496
rect 13771 15456 13912 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 10873 15351 10931 15357
rect 10873 15348 10885 15351
rect 10284 15320 10885 15348
rect 10284 15308 10290 15320
rect 10873 15317 10885 15320
rect 10919 15317 10931 15351
rect 10873 15311 10931 15317
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 11333 15351 11391 15357
rect 11333 15348 11345 15351
rect 11204 15320 11345 15348
rect 11204 15308 11210 15320
rect 11333 15317 11345 15320
rect 11379 15317 11391 15351
rect 13372 15348 13400 15444
rect 13817 15419 13875 15425
rect 13817 15385 13829 15419
rect 13863 15416 13875 15419
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 13863 15388 14381 15416
rect 13863 15385 13875 15388
rect 13817 15379 13875 15385
rect 14369 15385 14381 15388
rect 14415 15385 14427 15419
rect 14642 15416 14648 15428
rect 14369 15379 14427 15385
rect 14476 15388 14648 15416
rect 14476 15348 14504 15388
rect 14642 15376 14648 15388
rect 14700 15416 14706 15428
rect 14700 15388 14858 15416
rect 14700 15376 14706 15388
rect 17218 15376 17224 15428
rect 17276 15416 17282 15428
rect 17420 15416 17448 15512
rect 17604 15493 17632 15524
rect 20162 15512 20168 15564
rect 20220 15552 20226 15564
rect 21284 15561 21312 15592
rect 22646 15580 22652 15592
rect 22704 15580 22710 15632
rect 24210 15580 24216 15632
rect 24268 15620 24274 15632
rect 33520 15620 33548 15660
rect 34698 15648 34704 15660
rect 34756 15648 34762 15700
rect 35342 15648 35348 15700
rect 35400 15648 35406 15700
rect 33686 15620 33692 15632
rect 24268 15592 33548 15620
rect 33612 15592 33692 15620
rect 24268 15580 24274 15592
rect 20349 15555 20407 15561
rect 20349 15552 20361 15555
rect 20220 15524 20361 15552
rect 20220 15512 20226 15524
rect 20349 15521 20361 15524
rect 20395 15521 20407 15555
rect 20349 15515 20407 15521
rect 21269 15555 21327 15561
rect 21269 15521 21281 15555
rect 21315 15521 21327 15555
rect 21269 15515 21327 15521
rect 21376 15524 22324 15552
rect 17589 15487 17647 15493
rect 17589 15453 17601 15487
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 17696 15416 17724 15447
rect 18138 15444 18144 15496
rect 18196 15444 18202 15496
rect 18414 15444 18420 15496
rect 18472 15444 18478 15496
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15484 18567 15487
rect 18555 15456 18736 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 18046 15416 18052 15428
rect 17276 15388 17724 15416
rect 17788 15388 18052 15416
rect 17276 15376 17282 15388
rect 13372 15320 14504 15348
rect 15841 15351 15899 15357
rect 11333 15311 11391 15317
rect 15841 15317 15853 15351
rect 15887 15348 15899 15351
rect 16298 15348 16304 15360
rect 15887 15320 16304 15348
rect 15887 15317 15899 15320
rect 15841 15311 15899 15317
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 17788 15348 17816 15388
rect 18046 15376 18052 15388
rect 18104 15416 18110 15428
rect 18325 15419 18383 15425
rect 18325 15416 18337 15419
rect 18104 15388 18337 15416
rect 18104 15376 18110 15388
rect 18325 15385 18337 15388
rect 18371 15385 18383 15419
rect 18325 15379 18383 15385
rect 16908 15320 17816 15348
rect 16908 15308 16914 15320
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 18708 15348 18736 15456
rect 18874 15444 18880 15496
rect 18932 15484 18938 15496
rect 19426 15484 19432 15496
rect 18932 15456 19432 15484
rect 18932 15444 18938 15456
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 21376 15484 21404 15524
rect 20027 15456 21404 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 21450 15444 21456 15496
rect 21508 15444 21514 15496
rect 21652 15493 21680 15524
rect 22296 15496 22324 15524
rect 22480 15524 23525 15552
rect 21601 15487 21680 15493
rect 21601 15453 21613 15487
rect 21647 15456 21680 15487
rect 21647 15453 21659 15456
rect 21601 15447 21659 15453
rect 21726 15444 21732 15496
rect 21784 15444 21790 15496
rect 21918 15487 21976 15493
rect 21918 15453 21930 15487
rect 21964 15453 21976 15487
rect 21918 15447 21976 15453
rect 19444 15416 19472 15444
rect 20165 15419 20223 15425
rect 20165 15416 20177 15419
rect 19444 15388 20177 15416
rect 20165 15385 20177 15388
rect 20211 15416 20223 15419
rect 20441 15419 20499 15425
rect 20441 15416 20453 15419
rect 20211 15388 20453 15416
rect 20211 15385 20223 15388
rect 20165 15379 20223 15385
rect 20441 15385 20453 15388
rect 20487 15385 20499 15419
rect 20441 15379 20499 15385
rect 21818 15376 21824 15428
rect 21876 15376 21882 15428
rect 21928 15416 21956 15447
rect 22278 15444 22284 15496
rect 22336 15444 22342 15496
rect 22480 15416 22508 15524
rect 22557 15487 22615 15493
rect 22557 15453 22569 15487
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 21928 15388 22508 15416
rect 22572 15416 22600 15447
rect 22646 15444 22652 15496
rect 22704 15484 22710 15496
rect 22741 15487 22799 15493
rect 22741 15484 22753 15487
rect 22704 15456 22753 15484
rect 22704 15444 22710 15456
rect 22741 15453 22753 15456
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 23497 15493 23525 15524
rect 23750 15512 23756 15564
rect 23808 15552 23814 15564
rect 23934 15552 23940 15564
rect 23808 15524 23940 15552
rect 23808 15512 23814 15524
rect 23934 15512 23940 15524
rect 23992 15512 23998 15564
rect 27246 15552 27252 15564
rect 24044 15524 27252 15552
rect 23017 15487 23075 15493
rect 23017 15484 23029 15487
rect 22980 15456 23029 15484
rect 22980 15444 22986 15456
rect 23017 15453 23029 15456
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 23110 15487 23168 15493
rect 23110 15453 23122 15487
rect 23156 15453 23168 15487
rect 23110 15447 23168 15453
rect 23482 15487 23540 15493
rect 23482 15453 23494 15487
rect 23528 15453 23540 15487
rect 24044 15484 24072 15524
rect 27246 15512 27252 15524
rect 27304 15512 27310 15564
rect 29178 15512 29184 15564
rect 29236 15552 29242 15564
rect 29641 15555 29699 15561
rect 29641 15552 29653 15555
rect 29236 15524 29653 15552
rect 29236 15512 29242 15524
rect 29641 15521 29653 15524
rect 29687 15521 29699 15555
rect 29641 15515 29699 15521
rect 30098 15512 30104 15564
rect 30156 15512 30162 15564
rect 23482 15447 23540 15453
rect 23584 15456 24072 15484
rect 23124 15416 23152 15447
rect 23198 15416 23204 15428
rect 22572 15388 23204 15416
rect 18196 15320 18736 15348
rect 18196 15308 18202 15320
rect 21358 15308 21364 15360
rect 21416 15348 21422 15360
rect 21928 15348 21956 15388
rect 23198 15376 23204 15388
rect 23256 15376 23262 15428
rect 23293 15419 23351 15425
rect 23293 15385 23305 15419
rect 23339 15385 23351 15419
rect 23293 15379 23351 15385
rect 21416 15320 21956 15348
rect 21416 15308 21422 15320
rect 22094 15308 22100 15360
rect 22152 15308 22158 15360
rect 22278 15308 22284 15360
rect 22336 15348 22342 15360
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 22336 15320 22661 15348
rect 22336 15308 22342 15320
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 22649 15311 22707 15317
rect 22830 15308 22836 15360
rect 22888 15348 22894 15360
rect 23308 15348 23336 15379
rect 23382 15376 23388 15428
rect 23440 15376 23446 15428
rect 23584 15348 23612 15456
rect 24118 15444 24124 15496
rect 24176 15444 24182 15496
rect 24394 15444 24400 15496
rect 24452 15444 24458 15496
rect 24578 15493 24584 15496
rect 24545 15487 24584 15493
rect 24545 15453 24557 15487
rect 24545 15447 24584 15453
rect 24578 15444 24584 15447
rect 24636 15444 24642 15496
rect 24854 15444 24860 15496
rect 24912 15493 24918 15496
rect 24912 15484 24920 15493
rect 24912 15456 24957 15484
rect 24912 15447 24920 15456
rect 24912 15444 24918 15447
rect 29454 15444 29460 15496
rect 29512 15484 29518 15496
rect 33612 15493 33640 15592
rect 33686 15580 33692 15592
rect 33744 15620 33750 15632
rect 34606 15620 34612 15632
rect 33744 15592 34612 15620
rect 33744 15580 33750 15592
rect 34606 15580 34612 15592
rect 34664 15580 34670 15632
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29512 15456 29745 15484
rect 29512 15444 29518 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 33597 15487 33655 15493
rect 33597 15453 33609 15487
rect 33643 15453 33655 15487
rect 33597 15447 33655 15453
rect 33873 15487 33931 15493
rect 33873 15453 33885 15487
rect 33919 15484 33931 15487
rect 33962 15484 33968 15496
rect 33919 15456 33968 15484
rect 33919 15453 33931 15456
rect 33873 15447 33931 15453
rect 33962 15444 33968 15456
rect 34020 15444 34026 15496
rect 34054 15444 34060 15496
rect 34112 15444 34118 15496
rect 35360 15484 35388 15648
rect 35529 15487 35587 15493
rect 35529 15484 35541 15487
rect 35360 15456 35541 15484
rect 35529 15453 35541 15456
rect 35575 15453 35587 15487
rect 35529 15447 35587 15453
rect 35713 15487 35771 15493
rect 35713 15453 35725 15487
rect 35759 15453 35771 15487
rect 35713 15447 35771 15453
rect 24136 15416 24164 15444
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 24136 15388 24685 15416
rect 24596 15360 24624 15388
rect 24673 15385 24685 15388
rect 24719 15385 24731 15419
rect 24673 15379 24731 15385
rect 24762 15376 24768 15428
rect 24820 15376 24826 15428
rect 25130 15376 25136 15428
rect 25188 15416 25194 15428
rect 25188 15388 31754 15416
rect 25188 15376 25194 15388
rect 22888 15320 23612 15348
rect 23661 15351 23719 15357
rect 22888 15308 22894 15320
rect 23661 15317 23673 15351
rect 23707 15348 23719 15351
rect 24210 15348 24216 15360
rect 23707 15320 24216 15348
rect 23707 15317 23719 15320
rect 23661 15311 23719 15317
rect 24210 15308 24216 15320
rect 24268 15308 24274 15360
rect 24578 15308 24584 15360
rect 24636 15308 24642 15360
rect 24946 15308 24952 15360
rect 25004 15348 25010 15360
rect 25041 15351 25099 15357
rect 25041 15348 25053 15351
rect 25004 15320 25053 15348
rect 25004 15308 25010 15320
rect 25041 15317 25053 15320
rect 25087 15317 25099 15351
rect 31726 15348 31754 15388
rect 31938 15376 31944 15428
rect 31996 15416 32002 15428
rect 34072 15416 34100 15444
rect 35728 15416 35756 15447
rect 31996 15388 35756 15416
rect 31996 15376 32002 15388
rect 33778 15348 33784 15360
rect 31726 15320 33784 15348
rect 25041 15311 25099 15317
rect 33778 15308 33784 15320
rect 33836 15308 33842 15360
rect 35526 15308 35532 15360
rect 35584 15348 35590 15360
rect 35621 15351 35679 15357
rect 35621 15348 35633 15351
rect 35584 15320 35633 15348
rect 35584 15308 35590 15320
rect 35621 15317 35633 15320
rect 35667 15317 35679 15351
rect 35621 15311 35679 15317
rect 38654 15308 38660 15360
rect 38712 15348 38718 15360
rect 39482 15348 39488 15360
rect 38712 15320 39488 15348
rect 38712 15308 38718 15320
rect 39482 15308 39488 15320
rect 39540 15308 39546 15360
rect 1104 15258 41400 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 41400 15258
rect 1104 15184 41400 15206
rect 5534 15104 5540 15156
rect 5592 15104 5598 15156
rect 6917 15147 6975 15153
rect 6917 15113 6929 15147
rect 6963 15144 6975 15147
rect 7466 15144 7472 15156
rect 6963 15116 7472 15144
rect 6963 15113 6975 15116
rect 6917 15107 6975 15113
rect 7466 15104 7472 15116
rect 7524 15104 7530 15156
rect 9214 15144 9220 15156
rect 8956 15116 9220 15144
rect 6546 15036 6552 15088
rect 6604 15076 6610 15088
rect 8956 15085 8984 15116
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 9861 15147 9919 15153
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 10410 15144 10416 15156
rect 9907 15116 10416 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 10410 15104 10416 15116
rect 10468 15144 10474 15156
rect 10778 15144 10784 15156
rect 10468 15116 10784 15144
rect 10468 15104 10474 15116
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 10870 15104 10876 15156
rect 10928 15104 10934 15156
rect 11698 15104 11704 15156
rect 11756 15104 11762 15156
rect 12406 15116 13584 15144
rect 8941 15079 8999 15085
rect 6604 15048 7512 15076
rect 6604 15036 6610 15048
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 15008 5411 15011
rect 5810 15008 5816 15020
rect 5399 14980 5816 15008
rect 5399 14977 5411 14980
rect 5353 14971 5411 14977
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 6656 15017 6684 15048
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 6730 14968 6736 15020
rect 6788 14968 6794 15020
rect 7282 14968 7288 15020
rect 7340 14968 7346 15020
rect 7484 15017 7512 15048
rect 8941 15045 8953 15079
rect 8987 15045 8999 15079
rect 8941 15039 8999 15045
rect 9033 15079 9091 15085
rect 9033 15045 9045 15079
rect 9079 15076 9091 15079
rect 10888 15076 10916 15104
rect 9079 15048 9444 15076
rect 9079 15045 9091 15048
rect 9033 15039 9091 15045
rect 9416 15020 9444 15048
rect 9692 15048 11284 15076
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 14977 8355 15011
rect 8297 14971 8355 14977
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14940 5227 14943
rect 5902 14940 5908 14952
rect 5215 14912 5908 14940
rect 5215 14909 5227 14912
rect 5169 14903 5227 14909
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 7484 14940 7512 14971
rect 8113 14943 8171 14949
rect 8113 14940 8125 14943
rect 7484 14912 8125 14940
rect 8113 14909 8125 14912
rect 8159 14940 8171 14943
rect 8202 14940 8208 14952
rect 8159 14912 8208 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8312 14940 8340 14971
rect 8846 14968 8852 15020
rect 8904 14968 8910 15020
rect 9122 14968 9128 15020
rect 9180 15017 9186 15020
rect 9180 15011 9209 15017
rect 9197 14977 9209 15011
rect 9180 14971 9209 14977
rect 9180 14968 9186 14971
rect 9398 14968 9404 15020
rect 9456 14968 9462 15020
rect 9692 15017 9720 15048
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9950 14968 9956 15020
rect 10008 14968 10014 15020
rect 10226 14968 10232 15020
rect 10284 14968 10290 15020
rect 10870 14968 10876 15020
rect 10928 14968 10934 15020
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 15008 11023 15011
rect 11146 15008 11152 15020
rect 11011 14980 11152 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 11256 15017 11284 15048
rect 11330 15036 11336 15088
rect 11388 15076 11394 15088
rect 12406 15076 12434 15116
rect 11388 15048 12434 15076
rect 11388 15036 11394 15048
rect 11241 15011 11299 15017
rect 11241 14977 11253 15011
rect 11287 14977 11299 15011
rect 11241 14971 11299 14977
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 15008 11575 15011
rect 11882 15008 11888 15020
rect 11563 14980 11888 15008
rect 11563 14977 11575 14980
rect 11517 14971 11575 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 13556 15008 13584 15116
rect 13906 15104 13912 15156
rect 13964 15144 13970 15156
rect 14093 15147 14151 15153
rect 14093 15144 14105 15147
rect 13964 15116 14105 15144
rect 13964 15104 13970 15116
rect 14093 15113 14105 15116
rect 14139 15113 14151 15147
rect 16482 15144 16488 15156
rect 14093 15107 14151 15113
rect 15672 15116 16488 15144
rect 15672 15088 15700 15116
rect 16482 15104 16488 15116
rect 16540 15144 16546 15156
rect 17221 15147 17279 15153
rect 16540 15116 17080 15144
rect 16540 15104 16546 15116
rect 14461 15079 14519 15085
rect 14461 15045 14473 15079
rect 14507 15076 14519 15079
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 14507 15048 15025 15076
rect 14507 15045 14519 15048
rect 14461 15039 14519 15045
rect 15013 15045 15025 15048
rect 15059 15045 15071 15079
rect 15013 15039 15071 15045
rect 15654 15036 15660 15088
rect 15712 15036 15718 15088
rect 16945 15079 17003 15085
rect 16945 15076 16957 15079
rect 16316 15048 16957 15076
rect 16316 15020 16344 15048
rect 16945 15045 16957 15048
rect 16991 15045 17003 15079
rect 16945 15039 17003 15045
rect 14921 15011 14979 15017
rect 13556 14994 14780 15008
rect 13570 14980 14780 14994
rect 9306 14940 9312 14952
rect 8312 14912 9312 14940
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 9968 14940 9996 14968
rect 10137 14943 10195 14949
rect 10137 14940 10149 14943
rect 9968 14912 10149 14940
rect 10137 14909 10149 14912
rect 10183 14909 10195 14943
rect 10137 14903 10195 14909
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14909 12219 14943
rect 12161 14903 12219 14909
rect 6362 14832 6368 14884
rect 6420 14872 6426 14884
rect 12176 14872 12204 14903
rect 12434 14900 12440 14952
rect 12492 14900 12498 14952
rect 14458 14900 14464 14952
rect 14516 14900 14522 14952
rect 14550 14900 14556 14952
rect 14608 14900 14614 14952
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14909 14703 14943
rect 14752 14940 14780 14980
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 16298 15008 16304 15020
rect 14967 14980 16304 15008
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 16758 15008 16764 15020
rect 16715 14980 16764 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 17052 15017 17080 15116
rect 17221 15113 17233 15147
rect 17267 15144 17279 15147
rect 17954 15144 17960 15156
rect 17267 15116 17960 15144
rect 17267 15113 17279 15116
rect 17221 15107 17279 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18782 15144 18788 15156
rect 18104 15116 18788 15144
rect 18104 15104 18110 15116
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 19521 15147 19579 15153
rect 19521 15113 19533 15147
rect 19567 15144 19579 15147
rect 19794 15144 19800 15156
rect 19567 15116 19800 15144
rect 19567 15113 19579 15116
rect 19521 15107 19579 15113
rect 19794 15104 19800 15116
rect 19852 15104 19858 15156
rect 22833 15147 22891 15153
rect 22833 15113 22845 15147
rect 22879 15144 22891 15147
rect 23382 15144 23388 15156
rect 22879 15116 23388 15144
rect 22879 15113 22891 15116
rect 22833 15107 22891 15113
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 23474 15104 23480 15156
rect 23532 15144 23538 15156
rect 23532 15116 24164 15144
rect 23532 15104 23538 15116
rect 23658 15076 23664 15088
rect 18156 15048 23664 15076
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 14752 14912 15332 14940
rect 14645 14903 14703 14909
rect 6420 14844 12204 14872
rect 14476 14872 14504 14900
rect 14660 14872 14688 14903
rect 15304 14884 15332 14912
rect 15746 14900 15752 14952
rect 15804 14940 15810 14952
rect 16868 14940 16896 14971
rect 17402 14968 17408 15020
rect 17460 15008 17466 15020
rect 18156 15017 18184 15048
rect 23658 15036 23664 15048
rect 23716 15036 23722 15088
rect 24136 15076 24164 15116
rect 24394 15104 24400 15156
rect 24452 15104 24458 15156
rect 26234 15144 26240 15156
rect 24780 15116 26240 15144
rect 24780 15076 24808 15116
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 27706 15104 27712 15156
rect 27764 15144 27770 15156
rect 28350 15144 28356 15156
rect 27764 15116 28356 15144
rect 27764 15104 27770 15116
rect 28350 15104 28356 15116
rect 28408 15104 28414 15156
rect 29917 15147 29975 15153
rect 29917 15113 29929 15147
rect 29963 15144 29975 15147
rect 30006 15144 30012 15156
rect 29963 15116 30012 15144
rect 29963 15113 29975 15116
rect 29917 15107 29975 15113
rect 30006 15104 30012 15116
rect 30064 15104 30070 15156
rect 30098 15104 30104 15156
rect 30156 15104 30162 15156
rect 39758 15144 39764 15156
rect 30208 15116 39764 15144
rect 24136 15048 24808 15076
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 17460 14980 18153 15008
rect 17460 14968 17466 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 19429 15011 19487 15017
rect 19429 15008 19441 15011
rect 19392 14980 19441 15008
rect 19392 14968 19398 14980
rect 19429 14977 19441 14980
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 15804 14912 16896 14940
rect 15804 14900 15810 14912
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18230 14940 18236 14952
rect 18012 14912 18236 14940
rect 18012 14900 18018 14912
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 19444 14940 19472 14971
rect 19518 14968 19524 15020
rect 19576 15008 19582 15020
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 19576 14980 19625 15008
rect 19576 14968 19582 14980
rect 19613 14977 19625 14980
rect 19659 14977 19671 15011
rect 19613 14971 19671 14977
rect 19705 15011 19763 15017
rect 19705 14977 19717 15011
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 19720 14940 19748 14971
rect 20162 14968 20168 15020
rect 20220 14968 20226 15020
rect 20254 14968 20260 15020
rect 20312 15008 20318 15020
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 20312 14980 20453 15008
rect 20312 14968 20318 14980
rect 20441 14977 20453 14980
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 20901 15011 20959 15017
rect 20901 15008 20913 15011
rect 20772 14980 20913 15008
rect 20772 14968 20778 14980
rect 20901 14977 20913 14980
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 21637 15011 21695 15017
rect 21637 14977 21649 15011
rect 21683 14977 21695 15011
rect 21637 14971 21695 14977
rect 22741 15011 22799 15017
rect 22741 14977 22753 15011
rect 22787 15008 22799 15011
rect 22922 15008 22928 15020
rect 22787 14980 22928 15008
rect 22787 14977 22799 14980
rect 22741 14971 22799 14977
rect 19444 14912 19748 14940
rect 20070 14900 20076 14952
rect 20128 14940 20134 14952
rect 21174 14940 21180 14952
rect 20128 14912 21180 14940
rect 20128 14900 20134 14912
rect 21174 14900 21180 14912
rect 21232 14900 21238 14952
rect 21542 14900 21548 14952
rect 21600 14940 21606 14952
rect 21652 14940 21680 14971
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 23106 14968 23112 15020
rect 23164 14968 23170 15020
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 23845 15011 23903 15017
rect 23845 15008 23857 15011
rect 23808 14980 23857 15008
rect 23808 14968 23814 14980
rect 23845 14977 23857 14980
rect 23891 14977 23903 15011
rect 23845 14971 23903 14977
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 14977 24087 15011
rect 24029 14971 24087 14977
rect 23124 14940 23152 14968
rect 21600 14912 23152 14940
rect 21600 14900 21606 14912
rect 14476 14844 14688 14872
rect 6420 14832 6426 14844
rect 15286 14832 15292 14884
rect 15344 14832 15350 14884
rect 16482 14832 16488 14884
rect 16540 14872 16546 14884
rect 18325 14875 18383 14881
rect 18325 14872 18337 14875
rect 16540 14844 18337 14872
rect 16540 14832 16546 14844
rect 18325 14841 18337 14844
rect 18371 14872 18383 14875
rect 18414 14872 18420 14884
rect 18371 14844 18420 14872
rect 18371 14841 18383 14844
rect 18325 14835 18383 14841
rect 18414 14832 18420 14844
rect 18472 14832 18478 14884
rect 19426 14832 19432 14884
rect 19484 14872 19490 14884
rect 19797 14875 19855 14881
rect 19797 14872 19809 14875
rect 19484 14844 19809 14872
rect 19484 14832 19490 14844
rect 19797 14841 19809 14844
rect 19843 14841 19855 14875
rect 24044 14872 24072 14971
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 24228 15017 24256 15048
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 26510 15076 26516 15088
rect 24912 15048 26516 15076
rect 24912 15036 24918 15048
rect 26510 15036 26516 15048
rect 26568 15076 26574 15088
rect 27157 15079 27215 15085
rect 27157 15076 27169 15079
rect 26568 15048 27169 15076
rect 26568 15036 26574 15048
rect 27157 15045 27169 15048
rect 27203 15045 27215 15079
rect 27157 15039 27215 15045
rect 27246 15036 27252 15088
rect 27304 15076 27310 15088
rect 27304 15048 29868 15076
rect 27304 15036 27310 15048
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 25958 14968 25964 15020
rect 26016 15008 26022 15020
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26016 14980 26985 15008
rect 26016 14968 26022 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 15008 27399 15011
rect 27522 15008 27528 15020
rect 27387 14980 27528 15008
rect 27387 14977 27399 14980
rect 27341 14971 27399 14977
rect 26050 14900 26056 14952
rect 26108 14900 26114 14952
rect 26234 14900 26240 14952
rect 26292 14900 26298 14952
rect 26694 14900 26700 14952
rect 26752 14940 26758 14952
rect 27356 14940 27384 14971
rect 27522 14968 27528 14980
rect 27580 14968 27586 15020
rect 27617 15011 27675 15017
rect 27617 14977 27629 15011
rect 27663 15008 27675 15011
rect 27706 15008 27712 15020
rect 27663 14980 27712 15008
rect 27663 14977 27675 14980
rect 27617 14971 27675 14977
rect 27706 14968 27712 14980
rect 27764 14968 27770 15020
rect 27798 14968 27804 15020
rect 27856 14968 27862 15020
rect 27890 14968 27896 15020
rect 27948 14968 27954 15020
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 15008 28043 15011
rect 28074 15008 28080 15020
rect 28031 14980 28080 15008
rect 28031 14977 28043 14980
rect 27985 14971 28043 14977
rect 28000 14940 28028 14971
rect 28074 14968 28080 14980
rect 28132 15008 28138 15020
rect 28258 15008 28264 15020
rect 28132 14980 28264 15008
rect 28132 14968 28138 14980
rect 28258 14968 28264 14980
rect 28316 14968 28322 15020
rect 29733 15011 29791 15017
rect 29733 14977 29745 15011
rect 29779 14977 29791 15011
rect 29733 14971 29791 14977
rect 26752 14912 27384 14940
rect 27540 14912 28028 14940
rect 26752 14900 26758 14912
rect 26068 14872 26096 14900
rect 19797 14835 19855 14841
rect 19996 14844 21128 14872
rect 24044 14844 26096 14872
rect 26252 14872 26280 14900
rect 27540 14872 27568 14912
rect 26252 14844 27568 14872
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7377 14807 7435 14813
rect 7377 14804 7389 14807
rect 7064 14776 7389 14804
rect 7064 14764 7070 14776
rect 7377 14773 7389 14776
rect 7423 14773 7435 14807
rect 7377 14767 7435 14773
rect 8018 14764 8024 14816
rect 8076 14804 8082 14816
rect 8481 14807 8539 14813
rect 8481 14804 8493 14807
rect 8076 14776 8493 14804
rect 8076 14764 8082 14776
rect 8481 14773 8493 14776
rect 8527 14773 8539 14807
rect 8481 14767 8539 14773
rect 8662 14764 8668 14816
rect 8720 14764 8726 14816
rect 9493 14807 9551 14813
rect 9493 14773 9505 14807
rect 9539 14804 9551 14807
rect 9858 14804 9864 14816
rect 9539 14776 9864 14804
rect 9539 14773 9551 14776
rect 9493 14767 9551 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10594 14764 10600 14816
rect 10652 14764 10658 14816
rect 10686 14764 10692 14816
rect 10744 14764 10750 14816
rect 10962 14764 10968 14816
rect 11020 14804 11026 14816
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 11020 14776 11161 14804
rect 11020 14764 11026 14776
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 11149 14767 11207 14773
rect 13906 14764 13912 14816
rect 13964 14804 13970 14816
rect 16758 14804 16764 14816
rect 13964 14776 16764 14804
rect 13964 14764 13970 14776
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 17034 14764 17040 14816
rect 17092 14804 17098 14816
rect 19996 14804 20024 14844
rect 17092 14776 20024 14804
rect 21100 14804 21128 14844
rect 27614 14832 27620 14884
rect 27672 14872 27678 14884
rect 29748 14872 29776 14971
rect 29840 14940 29868 15048
rect 30009 15011 30067 15017
rect 30009 14977 30021 15011
rect 30055 15008 30067 15011
rect 30116 15008 30144 15104
rect 30055 14980 30144 15008
rect 30055 14977 30067 14980
rect 30009 14971 30067 14977
rect 30208 14940 30236 15116
rect 39758 15104 39764 15116
rect 39816 15104 39822 15156
rect 31205 15079 31263 15085
rect 31205 15076 31217 15079
rect 29840 14912 30236 14940
rect 30300 15048 31217 15076
rect 30300 14872 30328 15048
rect 31205 15045 31217 15048
rect 31251 15045 31263 15079
rect 31938 15076 31944 15088
rect 31205 15039 31263 15045
rect 31312 15048 31944 15076
rect 30745 15011 30803 15017
rect 30745 14977 30757 15011
rect 30791 14977 30803 15011
rect 30745 14971 30803 14977
rect 27672 14844 29684 14872
rect 29748 14844 30328 14872
rect 30760 14872 30788 14971
rect 31312 14952 31340 15048
rect 31938 15036 31944 15048
rect 31996 15036 32002 15088
rect 38676 15033 38734 15039
rect 31386 14968 31392 15020
rect 31444 14968 31450 15020
rect 31481 15011 31539 15017
rect 31481 14977 31493 15011
rect 31527 14977 31539 15011
rect 31481 14971 31539 14977
rect 30837 14943 30895 14949
rect 30837 14909 30849 14943
rect 30883 14940 30895 14943
rect 31294 14940 31300 14952
rect 30883 14912 31300 14940
rect 30883 14909 30895 14912
rect 30837 14903 30895 14909
rect 31294 14900 31300 14912
rect 31352 14900 31358 14952
rect 31496 14940 31524 14971
rect 31570 14968 31576 15020
rect 31628 14968 31634 15020
rect 31711 15011 31769 15017
rect 31711 14977 31723 15011
rect 31757 15008 31769 15011
rect 33962 15008 33968 15020
rect 31757 14980 33968 15008
rect 31757 14977 31769 14980
rect 31711 14971 31769 14977
rect 33962 14968 33968 14980
rect 34020 14968 34026 15020
rect 34698 14968 34704 15020
rect 34756 15008 34762 15020
rect 35345 15011 35403 15017
rect 35345 15008 35357 15011
rect 34756 14980 35357 15008
rect 34756 14968 34762 14980
rect 35345 14977 35357 14980
rect 35391 14977 35403 15011
rect 35345 14971 35403 14977
rect 35529 15011 35587 15017
rect 35529 14977 35541 15011
rect 35575 15008 35587 15011
rect 35618 15008 35624 15020
rect 35575 14980 35624 15008
rect 35575 14977 35587 14980
rect 35529 14971 35587 14977
rect 35618 14968 35624 14980
rect 35676 14968 35682 15020
rect 38676 14999 38688 15033
rect 38722 15030 38734 15033
rect 38722 15008 38976 15030
rect 39298 15008 39304 15020
rect 38722 15002 39304 15008
rect 38722 14999 38734 15002
rect 38676 14993 38734 14999
rect 38948 14980 39304 15002
rect 39298 14968 39304 14980
rect 39356 14968 39362 15020
rect 31496 14912 31702 14940
rect 31674 14872 31702 14912
rect 31846 14900 31852 14952
rect 31904 14900 31910 14952
rect 38933 14943 38991 14949
rect 38933 14909 38945 14943
rect 38979 14940 38991 14943
rect 38979 14912 39436 14940
rect 38979 14909 38991 14912
rect 38933 14903 38991 14909
rect 39408 14884 39436 14912
rect 32214 14872 32220 14884
rect 30760 14844 31248 14872
rect 31674 14844 32220 14872
rect 27672 14832 27678 14844
rect 25038 14804 25044 14816
rect 21100 14776 25044 14804
rect 17092 14764 17098 14776
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 27522 14764 27528 14816
rect 27580 14764 27586 14816
rect 28166 14764 28172 14816
rect 28224 14764 28230 14816
rect 29546 14764 29552 14816
rect 29604 14764 29610 14816
rect 29656 14804 29684 14844
rect 30760 14804 30788 14844
rect 29656 14776 30788 14804
rect 31110 14764 31116 14816
rect 31168 14764 31174 14816
rect 31220 14804 31248 14844
rect 32214 14832 32220 14844
rect 32272 14832 32278 14884
rect 35802 14872 35808 14884
rect 34072 14844 35808 14872
rect 31294 14804 31300 14816
rect 31220 14776 31300 14804
rect 31294 14764 31300 14776
rect 31352 14764 31358 14816
rect 31570 14764 31576 14816
rect 31628 14804 31634 14816
rect 32030 14804 32036 14816
rect 31628 14776 32036 14804
rect 31628 14764 31634 14776
rect 32030 14764 32036 14776
rect 32088 14804 32094 14816
rect 34072 14804 34100 14844
rect 35802 14832 35808 14844
rect 35860 14872 35866 14884
rect 35860 14844 39344 14872
rect 35860 14832 35866 14844
rect 32088 14776 34100 14804
rect 32088 14764 32094 14776
rect 35434 14764 35440 14816
rect 35492 14764 35498 14816
rect 38654 14764 38660 14816
rect 38712 14804 38718 14816
rect 38749 14807 38807 14813
rect 38749 14804 38761 14807
rect 38712 14776 38761 14804
rect 38712 14764 38718 14776
rect 38749 14773 38761 14776
rect 38795 14773 38807 14807
rect 38749 14767 38807 14773
rect 38838 14764 38844 14816
rect 38896 14764 38902 14816
rect 39316 14804 39344 14844
rect 39390 14832 39396 14884
rect 39448 14832 39454 14884
rect 39574 14804 39580 14816
rect 39316 14776 39580 14804
rect 39574 14764 39580 14776
rect 39632 14764 39638 14816
rect 1104 14714 41400 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 41400 14714
rect 1104 14640 41400 14662
rect 3418 14560 3424 14612
rect 3476 14560 3482 14612
rect 5629 14603 5687 14609
rect 5629 14569 5641 14603
rect 5675 14600 5687 14603
rect 5718 14600 5724 14612
rect 5675 14572 5724 14600
rect 5675 14569 5687 14572
rect 5629 14563 5687 14569
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 5810 14560 5816 14612
rect 5868 14560 5874 14612
rect 5902 14560 5908 14612
rect 5960 14600 5966 14612
rect 6089 14603 6147 14609
rect 6089 14600 6101 14603
rect 5960 14572 6101 14600
rect 5960 14560 5966 14572
rect 6089 14569 6101 14572
rect 6135 14569 6147 14603
rect 6089 14563 6147 14569
rect 6656 14572 8064 14600
rect 6549 14535 6607 14541
rect 6549 14532 6561 14535
rect 4172 14504 6561 14532
rect 3605 14467 3663 14473
rect 3605 14433 3617 14467
rect 3651 14464 3663 14467
rect 3973 14467 4031 14473
rect 3973 14464 3985 14467
rect 3651 14436 3985 14464
rect 3651 14433 3663 14436
rect 3605 14427 3663 14433
rect 3973 14433 3985 14436
rect 4019 14433 4031 14467
rect 3973 14427 4031 14433
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14396 3387 14399
rect 4062 14396 4068 14408
rect 3375 14368 4068 14396
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 4172 14405 4200 14504
rect 6549 14501 6561 14504
rect 6595 14501 6607 14535
rect 6549 14495 6607 14501
rect 5074 14464 5080 14476
rect 4448 14436 5080 14464
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 4361 14399 4419 14405
rect 4361 14365 4373 14399
rect 4407 14396 4419 14399
rect 4448 14396 4476 14436
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14464 5595 14467
rect 5810 14464 5816 14476
rect 5583 14436 5816 14464
rect 5583 14433 5595 14436
rect 5537 14427 5595 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 6178 14424 6184 14476
rect 6236 14464 6242 14476
rect 6656 14464 6684 14572
rect 8036 14544 8064 14572
rect 8662 14560 8668 14612
rect 8720 14560 8726 14612
rect 9122 14560 9128 14612
rect 9180 14560 9186 14612
rect 9306 14560 9312 14612
rect 9364 14560 9370 14612
rect 10686 14560 10692 14612
rect 10744 14600 10750 14612
rect 10744 14572 10824 14600
rect 10744 14560 10750 14572
rect 6236 14436 6684 14464
rect 6236 14424 6242 14436
rect 4407 14368 4476 14396
rect 4407 14365 4419 14368
rect 4361 14359 4419 14365
rect 4522 14356 4528 14408
rect 4580 14356 4586 14408
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 3973 14331 4031 14337
rect 3973 14297 3985 14331
rect 4019 14297 4031 14331
rect 3973 14291 4031 14297
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14328 4307 14331
rect 5169 14331 5227 14337
rect 5169 14328 5181 14331
rect 4295 14300 5181 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 5169 14297 5181 14300
rect 5215 14297 5227 14331
rect 5169 14291 5227 14297
rect 3602 14220 3608 14272
rect 3660 14220 3666 14272
rect 3988 14260 4016 14291
rect 4614 14260 4620 14272
rect 3988 14232 4620 14260
rect 4614 14220 4620 14232
rect 4672 14220 4678 14272
rect 4890 14220 4896 14272
rect 4948 14260 4954 14272
rect 5460 14260 5488 14359
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 5997 14399 6055 14405
rect 5776 14390 5856 14396
rect 5905 14393 5963 14399
rect 5905 14390 5917 14393
rect 5776 14368 5917 14390
rect 5776 14356 5782 14368
rect 5828 14362 5917 14368
rect 5905 14359 5917 14362
rect 5951 14359 5963 14393
rect 5997 14365 6009 14399
rect 6043 14396 6055 14399
rect 6043 14368 6132 14396
rect 6043 14365 6055 14368
rect 5997 14359 6055 14365
rect 5905 14353 5963 14359
rect 6104 14260 6132 14368
rect 6270 14356 6276 14408
rect 6328 14356 6334 14408
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14396 6515 14399
rect 6656 14396 6684 14436
rect 6748 14504 7052 14532
rect 6748 14405 6776 14504
rect 7024 14464 7052 14504
rect 7282 14492 7288 14544
rect 7340 14532 7346 14544
rect 7340 14504 7972 14532
rect 7340 14492 7346 14504
rect 7653 14467 7711 14473
rect 7653 14464 7665 14467
rect 7024 14436 7665 14464
rect 7653 14433 7665 14436
rect 7699 14433 7711 14467
rect 7944 14464 7972 14504
rect 8018 14492 8024 14544
rect 8076 14492 8082 14544
rect 8680 14464 8708 14560
rect 8938 14492 8944 14544
rect 8996 14532 9002 14544
rect 9140 14532 9168 14560
rect 10796 14532 10824 14572
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 11149 14603 11207 14609
rect 11149 14600 11161 14603
rect 10928 14572 11161 14600
rect 10928 14560 10934 14572
rect 11149 14569 11161 14572
rect 11195 14569 11207 14603
rect 11149 14563 11207 14569
rect 11885 14603 11943 14609
rect 11885 14569 11897 14603
rect 11931 14600 11943 14603
rect 12434 14600 12440 14612
rect 11931 14572 12440 14600
rect 11931 14569 11943 14572
rect 11885 14563 11943 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 15194 14600 15200 14612
rect 15120 14572 15200 14600
rect 8996 14504 10732 14532
rect 10796 14504 11284 14532
rect 8996 14492 9002 14504
rect 7944 14436 8248 14464
rect 7653 14427 7711 14433
rect 6503 14368 6684 14396
rect 6733 14399 6791 14405
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 6733 14365 6745 14399
rect 6779 14365 6791 14399
rect 6733 14359 6791 14365
rect 6822 14356 6828 14408
rect 6880 14356 6886 14408
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14396 7251 14399
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 7239 14368 7757 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 7745 14365 7757 14368
rect 7791 14365 7803 14399
rect 7745 14359 7803 14365
rect 7926 14356 7932 14408
rect 7984 14356 7990 14408
rect 8018 14356 8024 14408
rect 8076 14356 8082 14408
rect 8220 14405 8248 14436
rect 8312 14436 8708 14464
rect 8312 14405 8340 14436
rect 10410 14424 10416 14476
rect 10468 14464 10474 14476
rect 10468 14436 10640 14464
rect 10468 14424 10474 14436
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 8803 14368 9076 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 6638 14288 6644 14340
rect 6696 14328 6702 14340
rect 6917 14331 6975 14337
rect 6917 14328 6929 14331
rect 6696 14300 6929 14328
rect 6696 14288 6702 14300
rect 6917 14297 6929 14300
rect 6963 14297 6975 14331
rect 6917 14291 6975 14297
rect 7006 14288 7012 14340
rect 7064 14337 7070 14340
rect 7064 14331 7093 14337
rect 7081 14297 7093 14331
rect 7064 14291 7093 14297
rect 7285 14331 7343 14337
rect 7285 14297 7297 14331
rect 7331 14297 7343 14331
rect 7285 14291 7343 14297
rect 7469 14331 7527 14337
rect 7469 14297 7481 14331
rect 7515 14328 7527 14331
rect 8036 14328 8064 14356
rect 7515 14300 8064 14328
rect 8220 14328 8248 14359
rect 8478 14328 8484 14340
rect 8220 14300 8484 14328
rect 7515 14297 7527 14300
rect 7469 14291 7527 14297
rect 7064 14288 7070 14291
rect 4948 14232 6132 14260
rect 6457 14263 6515 14269
rect 4948 14220 4954 14232
rect 6457 14229 6469 14263
rect 6503 14260 6515 14263
rect 6656 14260 6684 14288
rect 6503 14232 6684 14260
rect 6503 14229 6515 14232
rect 6457 14223 6515 14229
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 7300 14260 7328 14291
rect 8478 14288 8484 14300
rect 8536 14288 8542 14340
rect 8588 14328 8616 14359
rect 9048 14340 9076 14368
rect 9214 14356 9220 14408
rect 9272 14396 9278 14408
rect 10612 14405 10640 14436
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 9272 14368 10517 14396
rect 9272 14356 9278 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 10598 14399 10656 14405
rect 10598 14365 10610 14399
rect 10644 14365 10656 14399
rect 10598 14359 10656 14365
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 8588 14300 8953 14328
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 8941 14291 8999 14297
rect 6788 14232 7328 14260
rect 6788 14220 6794 14232
rect 8202 14220 8208 14272
rect 8260 14260 8266 14272
rect 8665 14263 8723 14269
rect 8665 14260 8677 14263
rect 8260 14232 8677 14260
rect 8260 14220 8266 14232
rect 8665 14229 8677 14232
rect 8711 14229 8723 14263
rect 8956 14260 8984 14291
rect 9030 14288 9036 14340
rect 9088 14328 9094 14340
rect 9125 14331 9183 14337
rect 9125 14328 9137 14331
rect 9088 14300 9137 14328
rect 9088 14288 9094 14300
rect 9125 14297 9137 14300
rect 9171 14297 9183 14331
rect 10704 14328 10732 14504
rect 10778 14424 10784 14476
rect 10836 14424 10842 14476
rect 10796 14396 10824 14424
rect 11256 14405 11284 14504
rect 12897 14467 12955 14473
rect 12897 14433 12909 14467
rect 12943 14464 12955 14467
rect 13906 14464 13912 14476
rect 12943 14436 13912 14464
rect 12943 14433 12955 14436
rect 12897 14427 12955 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 10970 14399 11028 14405
rect 10970 14396 10982 14399
rect 10796 14368 10982 14396
rect 10970 14365 10982 14368
rect 11016 14365 11028 14399
rect 10970 14359 11028 14365
rect 11241 14399 11299 14405
rect 11241 14365 11253 14399
rect 11287 14365 11299 14399
rect 11241 14359 11299 14365
rect 11330 14356 11336 14408
rect 11388 14356 11394 14408
rect 11747 14399 11805 14405
rect 11747 14365 11759 14399
rect 11793 14396 11805 14399
rect 11882 14396 11888 14408
rect 11793 14368 11888 14396
rect 11793 14365 11805 14368
rect 11747 14359 11805 14365
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 14829 14399 14887 14405
rect 14829 14365 14841 14399
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 10781 14331 10839 14337
rect 10781 14328 10793 14331
rect 10704 14300 10793 14328
rect 9125 14291 9183 14297
rect 10781 14297 10793 14300
rect 10827 14297 10839 14331
rect 10781 14291 10839 14297
rect 10873 14331 10931 14337
rect 10873 14297 10885 14331
rect 10919 14328 10931 14331
rect 11422 14328 11428 14340
rect 10919 14300 11428 14328
rect 10919 14297 10931 14300
rect 10873 14291 10931 14297
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 11517 14331 11575 14337
rect 11517 14297 11529 14331
rect 11563 14297 11575 14331
rect 11517 14291 11575 14297
rect 11609 14331 11667 14337
rect 11609 14297 11621 14331
rect 11655 14328 11667 14331
rect 13449 14331 13507 14337
rect 13449 14328 13461 14331
rect 11655 14300 13461 14328
rect 11655 14297 11667 14300
rect 11609 14291 11667 14297
rect 13449 14297 13461 14300
rect 13495 14297 13507 14331
rect 14844 14328 14872 14359
rect 14918 14356 14924 14408
rect 14976 14396 14982 14408
rect 15120 14405 15148 14572
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 17221 14603 17279 14609
rect 17221 14569 17233 14603
rect 17267 14600 17279 14603
rect 17494 14600 17500 14612
rect 17267 14572 17500 14600
rect 17267 14569 17279 14572
rect 17221 14563 17279 14569
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 17604 14572 19334 14600
rect 17604 14532 17632 14572
rect 15212 14504 17632 14532
rect 17681 14535 17739 14541
rect 15212 14405 15240 14504
rect 17681 14501 17693 14535
rect 17727 14532 17739 14535
rect 17770 14532 17776 14544
rect 17727 14504 17776 14532
rect 17727 14501 17739 14504
rect 17681 14495 17739 14501
rect 17770 14492 17776 14504
rect 17828 14492 17834 14544
rect 18690 14532 18696 14544
rect 18432 14504 18696 14532
rect 16022 14464 16028 14476
rect 15396 14436 16028 14464
rect 15105 14399 15163 14405
rect 14976 14368 15021 14396
rect 14976 14356 14982 14368
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14365 15255 14399
rect 15197 14359 15255 14365
rect 15294 14399 15352 14405
rect 15294 14365 15306 14399
rect 15340 14390 15352 14399
rect 15396 14390 15424 14436
rect 16022 14424 16028 14436
rect 16080 14464 16086 14476
rect 18138 14464 18144 14476
rect 16080 14436 18144 14464
rect 16080 14424 16086 14436
rect 16114 14396 16120 14408
rect 15340 14365 15424 14390
rect 15294 14362 15424 14365
rect 15488 14368 16120 14396
rect 15294 14359 15352 14362
rect 15488 14328 15516 14368
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 16206 14356 16212 14408
rect 16264 14405 16270 14408
rect 16264 14399 16313 14405
rect 16264 14365 16267 14399
rect 16301 14365 16313 14399
rect 16264 14359 16313 14365
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14365 16451 14399
rect 16393 14359 16451 14365
rect 16264 14356 16270 14359
rect 14844 14300 14964 14328
rect 13449 14291 13507 14297
rect 9674 14260 9680 14272
rect 8956 14232 9680 14260
rect 8665 14223 8723 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 10594 14220 10600 14272
rect 10652 14260 10658 14272
rect 11532 14260 11560 14291
rect 14936 14272 14964 14300
rect 15120 14300 15516 14328
rect 15120 14272 15148 14300
rect 15562 14288 15568 14340
rect 15620 14288 15626 14340
rect 16408 14328 16436 14359
rect 17034 14356 17040 14408
rect 17092 14405 17098 14408
rect 17092 14359 17101 14405
rect 17092 14356 17098 14359
rect 17218 14356 17224 14408
rect 17276 14356 17282 14408
rect 18064 14405 18092 14436
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 18432 14405 18460 14504
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 19306 14532 19334 14572
rect 21910 14560 21916 14612
rect 21968 14600 21974 14612
rect 24486 14600 24492 14612
rect 21968 14572 24492 14600
rect 21968 14560 21974 14572
rect 24486 14560 24492 14572
rect 24544 14560 24550 14612
rect 24578 14560 24584 14612
rect 24636 14560 24642 14612
rect 26878 14560 26884 14612
rect 26936 14600 26942 14612
rect 27249 14603 27307 14609
rect 27249 14600 27261 14603
rect 26936 14572 27261 14600
rect 26936 14560 26942 14572
rect 27249 14569 27261 14572
rect 27295 14569 27307 14603
rect 27249 14563 27307 14569
rect 27341 14603 27399 14609
rect 27341 14569 27353 14603
rect 27387 14600 27399 14603
rect 27522 14600 27528 14612
rect 27387 14572 27528 14600
rect 27387 14569 27399 14572
rect 27341 14563 27399 14569
rect 27522 14560 27528 14572
rect 27580 14560 27586 14612
rect 28166 14600 28172 14612
rect 27724 14572 28172 14600
rect 20438 14532 20444 14544
rect 19306 14504 20444 14532
rect 20438 14492 20444 14504
rect 20496 14492 20502 14544
rect 20717 14535 20775 14541
rect 20717 14501 20729 14535
rect 20763 14532 20775 14535
rect 22738 14532 22744 14544
rect 20763 14504 22744 14532
rect 20763 14501 20775 14504
rect 20717 14495 20775 14501
rect 22738 14492 22744 14504
rect 22796 14492 22802 14544
rect 24596 14532 24624 14560
rect 27433 14535 27491 14541
rect 24596 14504 27384 14532
rect 20533 14467 20591 14473
rect 18616 14436 19334 14464
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 18325 14399 18383 14405
rect 18095 14368 18129 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 18325 14365 18337 14399
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 18340 14328 18368 14359
rect 18616 14328 18644 14436
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 18782 14396 18788 14408
rect 18739 14368 18788 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 18874 14356 18880 14408
rect 18932 14356 18938 14408
rect 16408 14300 17172 14328
rect 10652 14232 11560 14260
rect 10652 14220 10658 14232
rect 14918 14220 14924 14272
rect 14976 14220 14982 14272
rect 15102 14220 15108 14272
rect 15160 14220 15166 14272
rect 15473 14263 15531 14269
rect 15473 14229 15485 14263
rect 15519 14260 15531 14263
rect 15930 14260 15936 14272
rect 15519 14232 15936 14260
rect 15519 14229 15531 14232
rect 15473 14223 15531 14229
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 16114 14220 16120 14272
rect 16172 14260 16178 14272
rect 16758 14260 16764 14272
rect 16172 14232 16764 14260
rect 16172 14220 16178 14232
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 17144 14260 17172 14300
rect 17328 14300 17908 14328
rect 18340 14300 18644 14328
rect 19306 14328 19334 14436
rect 20533 14433 20545 14467
rect 20579 14464 20591 14467
rect 20990 14464 20996 14476
rect 20579 14436 20996 14464
rect 20579 14433 20591 14436
rect 20533 14427 20591 14433
rect 20990 14424 20996 14436
rect 21048 14464 21054 14476
rect 21048 14436 21220 14464
rect 21048 14424 21054 14436
rect 19794 14356 19800 14408
rect 19852 14396 19858 14408
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 19852 14368 20269 14396
rect 19852 14356 19858 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20438 14356 20444 14408
rect 20496 14396 20502 14408
rect 20806 14396 20812 14408
rect 20496 14368 20812 14396
rect 20496 14356 20502 14368
rect 20806 14356 20812 14368
rect 20864 14396 20870 14408
rect 21192 14405 21220 14436
rect 21542 14424 21548 14476
rect 21600 14424 21606 14476
rect 22922 14424 22928 14476
rect 22980 14424 22986 14476
rect 23014 14424 23020 14476
rect 23072 14464 23078 14476
rect 24854 14464 24860 14476
rect 23072 14436 24860 14464
rect 23072 14424 23078 14436
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 26142 14424 26148 14476
rect 26200 14464 26206 14476
rect 26602 14464 26608 14476
rect 26200 14436 26608 14464
rect 26200 14424 26206 14436
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20864 14368 20913 14396
rect 20864 14356 20870 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 21177 14399 21235 14405
rect 21177 14365 21189 14399
rect 21223 14396 21235 14399
rect 21560 14396 21588 14424
rect 21223 14368 21588 14396
rect 22097 14399 22155 14405
rect 21223 14365 21235 14368
rect 21177 14359 21235 14365
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22278 14396 22284 14408
rect 22143 14368 22284 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 22278 14356 22284 14368
rect 22336 14356 22342 14408
rect 22646 14356 22652 14408
rect 22704 14396 22710 14408
rect 26160 14396 26188 14424
rect 22704 14368 26188 14396
rect 22704 14356 22710 14368
rect 26326 14356 26332 14408
rect 26384 14356 26390 14408
rect 26510 14356 26516 14408
rect 26568 14356 26574 14408
rect 26694 14356 26700 14408
rect 26752 14356 26758 14408
rect 27062 14356 27068 14408
rect 27120 14396 27126 14408
rect 27356 14396 27384 14504
rect 27433 14501 27445 14535
rect 27479 14532 27491 14535
rect 27724 14532 27752 14572
rect 28166 14560 28172 14572
rect 28224 14560 28230 14612
rect 29546 14560 29552 14612
rect 29604 14560 29610 14612
rect 31294 14560 31300 14612
rect 31352 14560 31358 14612
rect 31386 14560 31392 14612
rect 31444 14600 31450 14612
rect 32033 14603 32091 14609
rect 32033 14600 32045 14603
rect 31444 14572 32045 14600
rect 31444 14560 31450 14572
rect 32033 14569 32045 14572
rect 32079 14569 32091 14603
rect 32033 14563 32091 14569
rect 32214 14560 32220 14612
rect 32272 14560 32278 14612
rect 35250 14560 35256 14612
rect 35308 14600 35314 14612
rect 35345 14603 35403 14609
rect 35345 14600 35357 14603
rect 35308 14572 35357 14600
rect 35308 14560 35314 14572
rect 35345 14569 35357 14572
rect 35391 14569 35403 14603
rect 37182 14600 37188 14612
rect 35345 14563 35403 14569
rect 36096 14572 37188 14600
rect 27479 14504 27752 14532
rect 29564 14532 29592 14560
rect 31312 14532 31340 14560
rect 31846 14532 31852 14544
rect 29564 14504 29684 14532
rect 31312 14504 31852 14532
rect 27479 14501 27491 14504
rect 27433 14495 27491 14501
rect 27724 14436 28212 14464
rect 27724 14405 27752 14436
rect 27712 14399 27770 14405
rect 27712 14396 27724 14399
rect 27120 14368 27292 14396
rect 27356 14368 27724 14396
rect 27120 14356 27126 14368
rect 19306 14300 25268 14328
rect 17328 14260 17356 14300
rect 17144 14232 17356 14260
rect 17402 14220 17408 14272
rect 17460 14220 17466 14272
rect 17880 14260 17908 14300
rect 18782 14260 18788 14272
rect 17880 14232 18788 14260
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 21085 14263 21143 14269
rect 21085 14229 21097 14263
rect 21131 14260 21143 14263
rect 21174 14260 21180 14272
rect 21131 14232 21180 14260
rect 21131 14229 21143 14232
rect 21085 14223 21143 14229
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 22005 14263 22063 14269
rect 22005 14229 22017 14263
rect 22051 14260 22063 14263
rect 22094 14260 22100 14272
rect 22051 14232 22100 14260
rect 22051 14229 22063 14232
rect 22005 14223 22063 14229
rect 22094 14220 22100 14232
rect 22152 14220 22158 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23658 14260 23664 14272
rect 22796 14232 23664 14260
rect 22796 14220 22802 14232
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 25240 14260 25268 14300
rect 25314 14288 25320 14340
rect 25372 14328 25378 14340
rect 26602 14328 26608 14340
rect 25372 14300 26608 14328
rect 25372 14288 25378 14300
rect 26602 14288 26608 14300
rect 26660 14288 26666 14340
rect 27264 14328 27292 14368
rect 27712 14365 27724 14368
rect 27758 14365 27770 14399
rect 27712 14359 27770 14365
rect 27798 14356 27804 14408
rect 27856 14356 27862 14408
rect 28184 14405 28212 14436
rect 29270 14424 29276 14476
rect 29328 14464 29334 14476
rect 29549 14467 29607 14473
rect 29549 14464 29561 14467
rect 29328 14436 29561 14464
rect 29328 14424 29334 14436
rect 29549 14433 29561 14436
rect 29595 14433 29607 14467
rect 29656 14464 29684 14504
rect 31846 14492 31852 14504
rect 31904 14532 31910 14544
rect 32122 14532 32128 14544
rect 31904 14504 32128 14532
rect 31904 14492 31910 14504
rect 32122 14492 32128 14504
rect 32180 14492 32186 14544
rect 33962 14492 33968 14544
rect 34020 14532 34026 14544
rect 36096 14532 36124 14572
rect 37182 14560 37188 14572
rect 37240 14600 37246 14612
rect 37240 14572 38148 14600
rect 37240 14560 37246 14572
rect 34020 14504 36124 14532
rect 34020 14492 34026 14504
rect 29825 14467 29883 14473
rect 29825 14464 29837 14467
rect 29656 14436 29837 14464
rect 29549 14427 29607 14433
rect 29825 14433 29837 14436
rect 29871 14433 29883 14467
rect 33778 14464 33784 14476
rect 29825 14427 29883 14433
rect 30944 14436 33784 14464
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14396 28227 14399
rect 28350 14396 28356 14408
rect 28215 14368 28356 14396
rect 28215 14365 28227 14368
rect 28169 14359 28227 14365
rect 28350 14356 28356 14368
rect 28408 14356 28414 14408
rect 30834 14356 30840 14408
rect 30892 14396 30898 14408
rect 30944 14396 30972 14436
rect 33778 14424 33784 14436
rect 33836 14424 33842 14476
rect 35161 14467 35219 14473
rect 35161 14433 35173 14467
rect 35207 14464 35219 14467
rect 35342 14464 35348 14476
rect 35207 14436 35348 14464
rect 35207 14433 35219 14436
rect 35161 14427 35219 14433
rect 35342 14424 35348 14436
rect 35400 14424 35406 14476
rect 35434 14424 35440 14476
rect 35492 14424 35498 14476
rect 35802 14424 35808 14476
rect 35860 14424 35866 14476
rect 30892 14382 30972 14396
rect 30892 14368 30958 14382
rect 30892 14356 30898 14368
rect 31294 14356 31300 14408
rect 31352 14356 31358 14408
rect 31478 14356 31484 14408
rect 31536 14396 31542 14408
rect 31665 14399 31723 14405
rect 31665 14396 31677 14399
rect 31536 14368 31677 14396
rect 31536 14356 31542 14368
rect 31665 14365 31677 14368
rect 31711 14396 31723 14399
rect 32125 14399 32183 14405
rect 32125 14396 32137 14399
rect 31711 14368 32137 14396
rect 31711 14365 31723 14368
rect 31665 14359 31723 14365
rect 32125 14365 32137 14368
rect 32171 14365 32183 14399
rect 32125 14359 32183 14365
rect 32309 14399 32367 14405
rect 32309 14365 32321 14399
rect 32355 14365 32367 14399
rect 32309 14359 32367 14365
rect 27985 14331 28043 14337
rect 27985 14328 27997 14331
rect 26712 14300 27108 14328
rect 27264 14300 27997 14328
rect 26712 14260 26740 14300
rect 25240 14232 26740 14260
rect 26878 14220 26884 14272
rect 26936 14220 26942 14272
rect 26970 14220 26976 14272
rect 27028 14220 27034 14272
rect 27080 14260 27108 14300
rect 27985 14297 27997 14300
rect 28031 14297 28043 14331
rect 27985 14291 28043 14297
rect 28077 14331 28135 14337
rect 28077 14297 28089 14331
rect 28123 14297 28135 14331
rect 28077 14291 28135 14297
rect 27614 14260 27620 14272
rect 27080 14232 27620 14260
rect 27614 14220 27620 14232
rect 27672 14220 27678 14272
rect 27706 14220 27712 14272
rect 27764 14260 27770 14272
rect 28092 14260 28120 14291
rect 31110 14288 31116 14340
rect 31168 14288 31174 14340
rect 31312 14328 31340 14356
rect 31573 14331 31631 14337
rect 31573 14328 31585 14331
rect 31312 14300 31585 14328
rect 31573 14297 31585 14300
rect 31619 14297 31631 14331
rect 31849 14331 31907 14337
rect 31849 14328 31861 14331
rect 31573 14291 31631 14297
rect 31726 14300 31861 14328
rect 27764 14232 28120 14260
rect 27764 14220 27770 14232
rect 28166 14220 28172 14272
rect 28224 14260 28230 14272
rect 28353 14263 28411 14269
rect 28353 14260 28365 14263
rect 28224 14232 28365 14260
rect 28224 14220 28230 14232
rect 28353 14229 28365 14232
rect 28399 14229 28411 14263
rect 31128 14260 31156 14288
rect 31478 14260 31484 14272
rect 31128 14232 31484 14260
rect 28353 14223 28411 14229
rect 31478 14220 31484 14232
rect 31536 14260 31542 14272
rect 31726 14260 31754 14300
rect 31849 14297 31861 14300
rect 31895 14328 31907 14331
rect 32324 14328 32352 14359
rect 31895 14300 32352 14328
rect 33796 14328 33824 14424
rect 35069 14399 35127 14405
rect 35069 14365 35081 14399
rect 35115 14396 35127 14399
rect 35452 14396 35480 14424
rect 35115 14368 35480 14396
rect 35115 14365 35127 14368
rect 35069 14359 35127 14365
rect 35526 14356 35532 14408
rect 35584 14356 35590 14408
rect 35677 14399 35735 14405
rect 35677 14365 35689 14399
rect 35723 14396 35735 14399
rect 35820 14396 35848 14424
rect 36096 14408 36124 14504
rect 36173 14535 36231 14541
rect 36173 14501 36185 14535
rect 36219 14501 36231 14535
rect 36173 14495 36231 14501
rect 36188 14464 36216 14495
rect 36541 14467 36599 14473
rect 36541 14464 36553 14467
rect 36188 14436 36553 14464
rect 36541 14433 36553 14436
rect 36587 14433 36599 14467
rect 36541 14427 36599 14433
rect 36078 14405 36084 14408
rect 35723 14368 35848 14396
rect 36035 14399 36084 14405
rect 35723 14365 35735 14368
rect 35677 14359 35735 14365
rect 36035 14365 36047 14399
rect 36081 14365 36084 14399
rect 36035 14359 36084 14365
rect 36078 14356 36084 14359
rect 36136 14356 36142 14408
rect 36170 14356 36176 14408
rect 36228 14396 36234 14408
rect 36265 14399 36323 14405
rect 36265 14396 36277 14399
rect 36228 14368 36277 14396
rect 36228 14356 36234 14368
rect 36265 14365 36277 14368
rect 36311 14365 36323 14399
rect 36265 14359 36323 14365
rect 33796 14300 35204 14328
rect 31895 14297 31907 14300
rect 31849 14291 31907 14297
rect 31536 14232 31754 14260
rect 31536 14220 31542 14232
rect 33318 14220 33324 14272
rect 33376 14260 33382 14272
rect 34514 14260 34520 14272
rect 33376 14232 34520 14260
rect 33376 14220 33382 14232
rect 34514 14220 34520 14232
rect 34572 14220 34578 14272
rect 35176 14260 35204 14300
rect 35250 14288 35256 14340
rect 35308 14328 35314 14340
rect 35805 14331 35863 14337
rect 35805 14328 35817 14331
rect 35308 14300 35817 14328
rect 35308 14288 35314 14300
rect 35805 14297 35817 14300
rect 35851 14297 35863 14331
rect 35805 14291 35863 14297
rect 35894 14288 35900 14340
rect 35952 14288 35958 14340
rect 36004 14300 37030 14328
rect 36004 14260 36032 14300
rect 35176 14232 36032 14260
rect 38120 14260 38148 14572
rect 38746 14532 38752 14544
rect 38396 14504 38752 14532
rect 38396 14405 38424 14504
rect 38746 14492 38752 14504
rect 38804 14492 38810 14544
rect 39482 14492 39488 14544
rect 39540 14492 39546 14544
rect 39117 14467 39175 14473
rect 39117 14464 39129 14467
rect 38544 14436 39129 14464
rect 38544 14405 38572 14436
rect 39117 14433 39129 14436
rect 39163 14433 39175 14467
rect 39117 14427 39175 14433
rect 39758 14424 39764 14476
rect 39816 14464 39822 14476
rect 39853 14467 39911 14473
rect 39853 14464 39865 14467
rect 39816 14436 39865 14464
rect 39816 14424 39822 14436
rect 39853 14433 39865 14436
rect 39899 14433 39911 14467
rect 39853 14427 39911 14433
rect 38381 14399 38439 14405
rect 38381 14365 38393 14399
rect 38427 14365 38439 14399
rect 38381 14359 38439 14365
rect 38529 14399 38587 14405
rect 38529 14365 38541 14399
rect 38575 14365 38587 14399
rect 38529 14359 38587 14365
rect 38654 14356 38660 14408
rect 38712 14356 38718 14408
rect 38746 14356 38752 14408
rect 38804 14356 38810 14408
rect 38846 14399 38904 14405
rect 38846 14365 38858 14399
rect 38892 14365 38904 14399
rect 38846 14359 38904 14365
rect 38286 14288 38292 14340
rect 38344 14288 38350 14340
rect 38856 14328 38884 14359
rect 39298 14356 39304 14408
rect 39356 14356 39362 14408
rect 39390 14356 39396 14408
rect 39448 14356 39454 14408
rect 39574 14356 39580 14408
rect 39632 14356 39638 14408
rect 38580 14300 38884 14328
rect 38580 14260 38608 14300
rect 40494 14288 40500 14340
rect 40552 14288 40558 14340
rect 38120 14232 38608 14260
rect 39025 14263 39083 14269
rect 39025 14229 39037 14263
rect 39071 14260 39083 14263
rect 39298 14260 39304 14272
rect 39071 14232 39304 14260
rect 39071 14229 39083 14232
rect 39025 14223 39083 14229
rect 39298 14220 39304 14232
rect 39356 14220 39362 14272
rect 1104 14170 41400 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 41400 14170
rect 1104 14096 41400 14118
rect 3602 14056 3608 14068
rect 2976 14028 3608 14056
rect 2976 13997 3004 14028
rect 3602 14016 3608 14028
rect 3660 14016 3666 14068
rect 4433 14059 4491 14065
rect 4433 14025 4445 14059
rect 4479 14056 4491 14059
rect 4522 14056 4528 14068
rect 4479 14028 4528 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 2961 13991 3019 13997
rect 2961 13957 2973 13991
rect 3007 13957 3019 13991
rect 2961 13951 3019 13957
rect 3050 13948 3056 14000
rect 3108 13988 3114 14000
rect 4448 13988 4476 14019
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 9214 14056 9220 14068
rect 8536 14028 9220 14056
rect 8536 14016 8542 14028
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 9732 14028 11529 14056
rect 9732 14016 9738 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 11977 14059 12035 14065
rect 11977 14025 11989 14059
rect 12023 14056 12035 14059
rect 12066 14056 12072 14068
rect 12023 14028 12072 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 15010 14056 15016 14068
rect 12492 14028 15016 14056
rect 12492 14016 12498 14028
rect 15010 14016 15016 14028
rect 15068 14056 15074 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 15068 14028 15117 14056
rect 15068 14016 15074 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 15105 14019 15163 14025
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 16850 14056 16856 14068
rect 15252 14028 16856 14056
rect 15252 14016 15258 14028
rect 16850 14016 16856 14028
rect 16908 14056 16914 14068
rect 16908 14028 17724 14056
rect 16908 14016 16914 14028
rect 3108 13960 3450 13988
rect 4448 13960 12434 13988
rect 3108 13948 3114 13960
rect 6914 13880 6920 13932
rect 6972 13920 6978 13932
rect 8110 13920 8116 13932
rect 6972 13892 8116 13920
rect 6972 13880 6978 13892
rect 8110 13880 8116 13892
rect 8168 13920 8174 13932
rect 11330 13920 11336 13932
rect 8168 13892 11336 13920
rect 8168 13880 8174 13892
rect 11330 13880 11336 13892
rect 11388 13880 11394 13932
rect 11882 13880 11888 13932
rect 11940 13880 11946 13932
rect 12406 13920 12434 13960
rect 14366 13948 14372 14000
rect 14424 13988 14430 14000
rect 14424 13960 15700 13988
rect 14424 13948 14430 13960
rect 15194 13920 15200 13932
rect 12406 13892 15200 13920
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15562 13880 15568 13932
rect 15620 13880 15626 13932
rect 15672 13929 15700 13960
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 15933 13991 15991 13997
rect 15933 13988 15945 13991
rect 15896 13960 15945 13988
rect 15896 13948 15902 13960
rect 15933 13957 15945 13960
rect 15979 13957 15991 13991
rect 15933 13951 15991 13957
rect 16942 13948 16948 14000
rect 17000 13948 17006 14000
rect 17696 13997 17724 14028
rect 17681 13991 17739 13997
rect 17681 13957 17693 13991
rect 17727 13988 17739 13991
rect 18276 13994 18414 14022
rect 18782 14016 18788 14068
rect 18840 14016 18846 14068
rect 19978 14016 19984 14068
rect 20036 14016 20042 14068
rect 21450 14056 21456 14068
rect 21104 14028 21456 14056
rect 18276 13988 18304 13994
rect 17727 13960 18304 13988
rect 18386 13988 18414 13994
rect 18509 13991 18567 13997
rect 18386 13960 18460 13988
rect 17727 13957 17739 13960
rect 17681 13951 17739 13957
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 16853 13923 16911 13929
rect 15703 13892 16804 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3694 13852 3700 13864
rect 2740 13824 3700 13852
rect 2740 13812 2746 13824
rect 3694 13812 3700 13824
rect 3752 13812 3758 13864
rect 7926 13812 7932 13864
rect 7984 13852 7990 13864
rect 8662 13852 8668 13864
rect 7984 13824 8668 13852
rect 7984 13812 7990 13824
rect 8662 13812 8668 13824
rect 8720 13852 8726 13864
rect 11238 13852 11244 13864
rect 8720 13824 11244 13852
rect 8720 13812 8726 13824
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13852 12219 13855
rect 12342 13852 12348 13864
rect 12207 13824 12348 13852
rect 12207 13821 12219 13824
rect 12161 13815 12219 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 15102 13812 15108 13864
rect 15160 13852 15166 13864
rect 15289 13855 15347 13861
rect 15289 13852 15301 13855
rect 15160 13824 15301 13852
rect 15160 13812 15166 13824
rect 15289 13821 15301 13824
rect 15335 13821 15347 13855
rect 15289 13815 15347 13821
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 15746 13852 15752 13864
rect 15436 13824 15752 13852
rect 15436 13812 15442 13824
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 15930 13812 15936 13864
rect 15988 13812 15994 13864
rect 16114 13812 16120 13864
rect 16172 13852 16178 13864
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16172 13824 16681 13852
rect 16172 13812 16178 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 15473 13787 15531 13793
rect 15473 13753 15485 13787
rect 15519 13784 15531 13787
rect 15948 13784 15976 13812
rect 15519 13756 15976 13784
rect 16776 13784 16804 13892
rect 16853 13889 16865 13923
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 16868 13852 16896 13883
rect 17034 13880 17040 13932
rect 17092 13880 17098 13932
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17221 13923 17279 13929
rect 17221 13920 17233 13923
rect 17184 13892 17233 13920
rect 17184 13880 17190 13892
rect 17221 13889 17233 13892
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 17402 13880 17408 13932
rect 17460 13880 17466 13932
rect 17497 13923 17555 13929
rect 17497 13889 17509 13923
rect 17543 13889 17555 13923
rect 17497 13883 17555 13889
rect 17420 13852 17448 13880
rect 16868 13824 17448 13852
rect 17512 13784 17540 13883
rect 17770 13880 17776 13932
rect 17828 13880 17834 13932
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 17911 13918 18000 13920
rect 18046 13918 18052 13932
rect 17911 13892 18052 13918
rect 17911 13889 17923 13892
rect 17972 13890 18052 13892
rect 17865 13883 17923 13889
rect 18046 13880 18052 13890
rect 18104 13880 18110 13932
rect 18138 13878 18144 13930
rect 18196 13878 18202 13930
rect 18432 13929 18460 13960
rect 18509 13957 18521 13991
rect 18555 13988 18567 13991
rect 19702 13988 19708 14000
rect 18555 13960 19708 13988
rect 18555 13957 18567 13960
rect 18509 13951 18567 13957
rect 19702 13948 19708 13960
rect 19760 13948 19766 14000
rect 19996 13988 20024 14016
rect 19812 13960 20024 13988
rect 18234 13926 18292 13929
rect 18234 13923 18368 13926
rect 18234 13889 18246 13923
rect 18280 13898 18368 13923
rect 18280 13889 18292 13898
rect 18234 13883 18292 13889
rect 17770 13784 17776 13796
rect 16776 13756 17776 13784
rect 15519 13753 15531 13756
rect 15473 13747 15531 13753
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13784 18107 13787
rect 18230 13784 18236 13796
rect 18095 13756 18236 13784
rect 18095 13753 18107 13756
rect 18049 13747 18107 13753
rect 18230 13744 18236 13756
rect 18288 13744 18294 13796
rect 18340 13784 18368 13898
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 18598 13880 18604 13932
rect 18656 13929 18662 13932
rect 19812 13929 19840 13960
rect 18656 13920 18664 13929
rect 19797 13923 19855 13929
rect 18656 13892 18701 13920
rect 18656 13883 18664 13892
rect 19797 13889 19809 13923
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 19981 13923 20039 13929
rect 19981 13889 19993 13923
rect 20027 13920 20039 13923
rect 20070 13920 20076 13932
rect 20027 13892 20076 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 18656 13880 18662 13883
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13920 20407 13923
rect 20438 13920 20444 13932
rect 20395 13892 20444 13920
rect 20395 13889 20407 13892
rect 20349 13883 20407 13889
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20898 13880 20904 13932
rect 20956 13880 20962 13932
rect 21104 13931 21132 14028
rect 21450 14016 21456 14028
rect 21508 14016 21514 14068
rect 22189 14059 22247 14065
rect 22189 14025 22201 14059
rect 22235 14056 22247 14059
rect 22278 14056 22284 14068
rect 22235 14028 22284 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 23474 14016 23480 14068
rect 23532 14016 23538 14068
rect 23842 14016 23848 14068
rect 23900 14016 23906 14068
rect 25582 14028 25824 14056
rect 25582 14022 25610 14028
rect 21174 13948 21180 14000
rect 21232 13988 21238 14000
rect 23492 13988 23520 14016
rect 21232 13960 23152 13988
rect 21232 13948 21238 13960
rect 21089 13925 21147 13931
rect 21089 13891 21101 13925
rect 21135 13891 21147 13925
rect 21089 13885 21147 13891
rect 21266 13880 21272 13932
rect 21324 13880 21330 13932
rect 21450 13880 21456 13932
rect 21508 13880 21514 13932
rect 22187 13923 22245 13929
rect 22187 13889 22199 13923
rect 22233 13920 22245 13923
rect 22370 13920 22376 13932
rect 22233 13892 22376 13920
rect 22233 13889 22245 13892
rect 22187 13883 22245 13889
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 22738 13880 22744 13932
rect 22796 13880 22802 13932
rect 22830 13880 22836 13932
rect 22888 13880 22894 13932
rect 23014 13880 23020 13932
rect 23072 13880 23078 13932
rect 23124 13929 23152 13960
rect 23262 13960 23520 13988
rect 23860 13988 23888 14016
rect 24688 13994 24900 14022
rect 24688 13988 24716 13994
rect 23860 13960 24716 13988
rect 24872 13988 24900 13994
rect 25332 13994 25610 14022
rect 25332 13988 25360 13994
rect 24872 13960 25360 13988
rect 23262 13929 23290 13960
rect 23109 13923 23167 13929
rect 23109 13889 23121 13923
rect 23155 13889 23167 13923
rect 23109 13883 23167 13889
rect 23247 13923 23305 13929
rect 23247 13889 23259 13923
rect 23293 13889 23305 13923
rect 23247 13883 23305 13889
rect 23474 13880 23480 13932
rect 23532 13880 23538 13932
rect 23658 13880 23664 13932
rect 23716 13880 23722 13932
rect 24136 13929 24164 13960
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13889 24179 13923
rect 24121 13883 24179 13889
rect 24305 13923 24363 13929
rect 24305 13889 24317 13923
rect 24351 13920 24363 13923
rect 24394 13920 24400 13932
rect 24351 13892 24400 13920
rect 24351 13889 24363 13892
rect 24305 13883 24363 13889
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 21177 13855 21235 13861
rect 21177 13852 21189 13855
rect 19576 13824 21189 13852
rect 19576 13812 19582 13824
rect 21177 13821 21189 13824
rect 21223 13821 21235 13855
rect 21177 13815 21235 13821
rect 18414 13784 18420 13796
rect 18340 13756 18420 13784
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 20254 13744 20260 13796
rect 20312 13744 20318 13796
rect 21284 13784 21312 13880
rect 21634 13812 21640 13864
rect 21692 13812 21698 13864
rect 22649 13855 22707 13861
rect 22649 13821 22661 13855
rect 22695 13852 22707 13855
rect 23569 13855 23627 13861
rect 23569 13852 23581 13855
rect 22695 13824 23581 13852
rect 22695 13821 22707 13824
rect 22649 13815 22707 13821
rect 23569 13821 23581 13824
rect 23615 13821 23627 13855
rect 23569 13815 23627 13821
rect 23750 13812 23756 13864
rect 23808 13852 23814 13864
rect 23952 13852 23980 13883
rect 23808 13824 23980 13852
rect 23808 13812 23814 13824
rect 24026 13812 24032 13864
rect 24084 13852 24090 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 24084 13824 24225 13852
rect 24084 13812 24090 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 21284 13756 22508 13784
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 15930 13716 15936 13728
rect 14608 13688 15936 13716
rect 14608 13676 14614 13688
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 17954 13716 17960 13728
rect 16080 13688 17960 13716
rect 16080 13676 16086 13688
rect 17954 13676 17960 13688
rect 18012 13676 18018 13728
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 21726 13716 21732 13728
rect 18196 13688 21732 13716
rect 18196 13676 18202 13688
rect 21726 13676 21732 13688
rect 21784 13716 21790 13728
rect 22005 13719 22063 13725
rect 22005 13716 22017 13719
rect 21784 13688 22017 13716
rect 21784 13676 21790 13688
rect 22005 13685 22017 13688
rect 22051 13685 22063 13719
rect 22480 13716 22508 13756
rect 22554 13744 22560 13796
rect 22612 13744 22618 13796
rect 24320 13784 24348 13883
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 24489 13923 24547 13929
rect 24489 13889 24501 13923
rect 24535 13920 24547 13923
rect 24578 13920 24584 13932
rect 24535 13892 24584 13920
rect 24535 13889 24547 13892
rect 24489 13883 24547 13889
rect 24578 13880 24584 13892
rect 24636 13880 24642 13932
rect 24964 13929 24992 13960
rect 25796 13935 25824 14028
rect 25958 14016 25964 14068
rect 26016 14016 26022 14068
rect 27246 14016 27252 14068
rect 27304 14016 27310 14068
rect 27338 14016 27344 14068
rect 27396 14056 27402 14068
rect 27709 14059 27767 14065
rect 27709 14056 27721 14059
rect 27396 14028 27721 14056
rect 27396 14016 27402 14028
rect 27709 14025 27721 14028
rect 27755 14056 27767 14059
rect 27755 14028 28994 14056
rect 27755 14025 27767 14028
rect 27709 14019 27767 14025
rect 24765 13923 24823 13929
rect 24670 13846 24676 13898
rect 24728 13846 24734 13898
rect 24765 13889 24777 13923
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13889 25007 13923
rect 24949 13883 25007 13889
rect 24673 13821 24685 13846
rect 24719 13821 24731 13846
rect 24673 13815 24731 13821
rect 23308 13756 24348 13784
rect 23308 13716 23336 13756
rect 22480 13688 23336 13716
rect 22005 13679 22063 13685
rect 23382 13676 23388 13728
rect 23440 13676 23446 13728
rect 23750 13676 23756 13728
rect 23808 13716 23814 13728
rect 24780 13716 24808 13883
rect 24964 13784 24992 13883
rect 25038 13880 25044 13932
rect 25096 13880 25102 13932
rect 25130 13880 25136 13932
rect 25188 13880 25194 13932
rect 25314 13880 25320 13932
rect 25372 13880 25378 13932
rect 25781 13929 25839 13935
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13889 25651 13923
rect 25781 13895 25793 13929
rect 25827 13895 25839 13929
rect 25781 13889 25839 13895
rect 25869 13923 25927 13929
rect 25869 13889 25881 13923
rect 25915 13920 25927 13923
rect 25976 13920 26004 14016
rect 27264 13988 27292 14016
rect 28077 13991 28135 13997
rect 28077 13988 28089 13991
rect 26160 13960 27292 13988
rect 27724 13960 28089 13988
rect 26160 13929 26188 13960
rect 27724 13932 27752 13960
rect 28077 13957 28089 13960
rect 28123 13957 28135 13991
rect 28077 13951 28135 13957
rect 25915 13892 26004 13920
rect 26145 13923 26203 13929
rect 25915 13889 25927 13892
rect 25593 13883 25651 13889
rect 25869 13883 25927 13889
rect 26145 13889 26157 13923
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 25038 13784 25044 13796
rect 24964 13756 25044 13784
rect 25038 13744 25044 13756
rect 25096 13744 25102 13796
rect 25608 13784 25636 13883
rect 26878 13880 26884 13932
rect 26936 13920 26942 13932
rect 27433 13923 27491 13929
rect 27433 13920 27445 13923
rect 26936 13892 27445 13920
rect 26936 13880 26942 13892
rect 27433 13889 27445 13892
rect 27479 13889 27491 13923
rect 27433 13883 27491 13889
rect 27706 13880 27712 13932
rect 27764 13880 27770 13932
rect 27804 13923 27862 13929
rect 27804 13889 27816 13923
rect 27850 13920 27862 13923
rect 27893 13923 27951 13929
rect 27850 13889 27864 13920
rect 27804 13883 27864 13889
rect 27893 13889 27905 13923
rect 27939 13889 27951 13923
rect 27893 13883 27951 13889
rect 28169 13923 28227 13929
rect 28169 13889 28181 13923
rect 28215 13889 28227 13923
rect 28169 13883 28227 13889
rect 25961 13855 26019 13861
rect 25961 13821 25973 13855
rect 26007 13821 26019 13855
rect 25961 13815 26019 13821
rect 25148 13756 25636 13784
rect 25148 13728 25176 13756
rect 25774 13744 25780 13796
rect 25832 13784 25838 13796
rect 25976 13784 26004 13815
rect 25832 13756 26004 13784
rect 25832 13744 25838 13756
rect 26786 13744 26792 13796
rect 26844 13784 26850 13796
rect 27338 13784 27344 13796
rect 26844 13756 27344 13784
rect 26844 13744 26850 13756
rect 27338 13744 27344 13756
rect 27396 13744 27402 13796
rect 27836 13784 27864 13883
rect 27908 13852 27936 13883
rect 28074 13852 28080 13864
rect 27908 13824 28080 13852
rect 28074 13812 28080 13824
rect 28132 13812 28138 13864
rect 28184 13852 28212 13883
rect 28258 13880 28264 13932
rect 28316 13880 28322 13932
rect 28966 13920 28994 14028
rect 31018 14016 31024 14068
rect 31076 14016 31082 14068
rect 31297 14059 31355 14065
rect 31297 14025 31309 14059
rect 31343 14056 31355 14059
rect 32950 14056 32956 14068
rect 31343 14028 32956 14056
rect 31343 14025 31355 14028
rect 31297 14019 31355 14025
rect 32950 14016 32956 14028
rect 33008 14016 33014 14068
rect 33045 14059 33103 14065
rect 33045 14025 33057 14059
rect 33091 14056 33103 14059
rect 33226 14056 33232 14068
rect 33091 14028 33232 14056
rect 33091 14025 33103 14028
rect 33045 14019 33103 14025
rect 33226 14016 33232 14028
rect 33284 14016 33290 14068
rect 33321 14059 33379 14065
rect 33321 14025 33333 14059
rect 33367 14056 33379 14059
rect 33962 14056 33968 14068
rect 33367 14028 33968 14056
rect 33367 14025 33379 14028
rect 33321 14019 33379 14025
rect 33962 14016 33968 14028
rect 34020 14016 34026 14068
rect 34072 14028 34560 14056
rect 30837 13991 30895 13997
rect 30837 13957 30849 13991
rect 30883 13988 30895 13991
rect 31036 13988 31064 14016
rect 30883 13960 31064 13988
rect 30883 13957 30895 13960
rect 30837 13951 30895 13957
rect 31386 13948 31392 14000
rect 31444 13988 31450 14000
rect 31665 13991 31723 13997
rect 31665 13988 31677 13991
rect 31444 13960 31677 13988
rect 31444 13948 31450 13960
rect 31665 13957 31677 13960
rect 31711 13957 31723 13991
rect 32968 13988 32996 14016
rect 34072 13988 34100 14028
rect 31665 13951 31723 13957
rect 31864 13960 32260 13988
rect 32968 13960 34100 13988
rect 30190 13920 30196 13932
rect 28966 13892 30196 13920
rect 30190 13880 30196 13892
rect 30248 13920 30254 13932
rect 31018 13920 31024 13932
rect 30248 13892 31024 13920
rect 30248 13880 30254 13892
rect 31018 13880 31024 13892
rect 31076 13880 31082 13932
rect 31205 13923 31263 13929
rect 31205 13889 31217 13923
rect 31251 13920 31263 13923
rect 31481 13923 31539 13929
rect 31481 13920 31493 13923
rect 31251 13892 31493 13920
rect 31251 13889 31263 13892
rect 31205 13883 31263 13889
rect 31481 13889 31493 13892
rect 31527 13889 31539 13923
rect 31481 13883 31539 13889
rect 31570 13880 31576 13932
rect 31628 13880 31634 13932
rect 31864 13929 31892 13960
rect 32232 13932 32260 13960
rect 31849 13923 31907 13929
rect 31849 13889 31861 13923
rect 31895 13889 31907 13923
rect 31849 13883 31907 13889
rect 31941 13923 31999 13929
rect 31941 13889 31953 13923
rect 31987 13889 31999 13923
rect 31941 13883 31999 13889
rect 28442 13852 28448 13864
rect 28184 13824 28448 13852
rect 28442 13812 28448 13824
rect 28500 13812 28506 13864
rect 28350 13784 28356 13796
rect 27836 13756 28356 13784
rect 28350 13744 28356 13756
rect 28408 13744 28414 13796
rect 31956 13784 31984 13883
rect 32030 13880 32036 13932
rect 32088 13880 32094 13932
rect 32122 13880 32128 13932
rect 32180 13880 32186 13932
rect 32214 13880 32220 13932
rect 32272 13880 32278 13932
rect 32309 13923 32367 13929
rect 32309 13889 32321 13923
rect 32355 13889 32367 13923
rect 32309 13883 32367 13889
rect 32769 13923 32827 13929
rect 32769 13889 32781 13923
rect 32815 13920 32827 13923
rect 33134 13920 33140 13932
rect 32815 13892 33140 13920
rect 32815 13889 32827 13892
rect 32769 13883 32827 13889
rect 32048 13852 32076 13880
rect 32324 13852 32352 13883
rect 33134 13880 33140 13892
rect 33192 13880 33198 13932
rect 33318 13920 33324 13932
rect 33279 13892 33324 13920
rect 33318 13880 33324 13892
rect 33376 13880 33382 13932
rect 33594 13880 33600 13932
rect 33652 13920 33658 13932
rect 34072 13929 34100 13960
rect 34238 13948 34244 14000
rect 34296 13988 34302 14000
rect 34532 13988 34560 14028
rect 34698 14016 34704 14068
rect 34756 14016 34762 14068
rect 35176 14028 35848 14056
rect 35176 13997 35204 14028
rect 35161 13991 35219 13997
rect 35161 13988 35173 13991
rect 34296 13960 34468 13988
rect 34532 13960 35173 13988
rect 34296 13948 34302 13960
rect 33781 13923 33839 13929
rect 33781 13920 33793 13923
rect 33652 13892 33793 13920
rect 33652 13880 33658 13892
rect 33781 13889 33793 13892
rect 33827 13889 33839 13923
rect 33781 13883 33839 13889
rect 34057 13923 34115 13929
rect 34057 13889 34069 13923
rect 34103 13889 34115 13923
rect 34057 13883 34115 13889
rect 34146 13880 34152 13932
rect 34204 13880 34210 13932
rect 34330 13880 34336 13932
rect 34388 13880 34394 13932
rect 34440 13929 34468 13960
rect 35161 13957 35173 13960
rect 35207 13957 35219 13991
rect 35161 13951 35219 13957
rect 35253 13991 35311 13997
rect 35253 13957 35265 13991
rect 35299 13957 35311 13991
rect 35253 13951 35311 13957
rect 34425 13923 34483 13929
rect 34425 13889 34437 13923
rect 34471 13889 34483 13923
rect 34425 13883 34483 13889
rect 34606 13880 34612 13932
rect 34664 13880 34670 13932
rect 34698 13880 34704 13932
rect 34756 13920 34762 13932
rect 34793 13923 34851 13929
rect 34793 13920 34805 13923
rect 34756 13892 34805 13920
rect 34756 13880 34762 13892
rect 34793 13889 34805 13892
rect 34839 13889 34851 13923
rect 34793 13883 34851 13889
rect 34882 13880 34888 13932
rect 34940 13920 34946 13932
rect 35069 13923 35127 13929
rect 34940 13918 35036 13920
rect 35069 13918 35081 13923
rect 34940 13892 35081 13918
rect 34940 13880 34946 13892
rect 35008 13890 35081 13892
rect 35069 13889 35081 13890
rect 35115 13889 35127 13923
rect 35069 13883 35127 13889
rect 32048 13824 32352 13852
rect 32493 13855 32551 13861
rect 32493 13821 32505 13855
rect 32539 13821 32551 13855
rect 32493 13815 32551 13821
rect 33045 13855 33103 13861
rect 33045 13821 33057 13855
rect 33091 13852 33103 13855
rect 34164 13852 34192 13880
rect 35268 13852 35296 13951
rect 35342 13948 35348 14000
rect 35400 13988 35406 14000
rect 35621 13991 35679 13997
rect 35621 13988 35633 13991
rect 35400 13960 35633 13988
rect 35400 13948 35406 13960
rect 35621 13957 35633 13960
rect 35667 13957 35679 13991
rect 35820 13988 35848 14028
rect 35894 14016 35900 14068
rect 35952 14056 35958 14068
rect 37001 14059 37059 14065
rect 37001 14056 37013 14059
rect 35952 14028 37013 14056
rect 35952 14016 35958 14028
rect 37001 14025 37013 14028
rect 37047 14025 37059 14059
rect 39390 14056 39396 14068
rect 37001 14019 37059 14025
rect 38948 14028 39396 14056
rect 35820 13960 36124 13988
rect 35621 13951 35679 13957
rect 35437 13923 35495 13929
rect 35437 13889 35449 13923
rect 35483 13889 35495 13923
rect 35437 13883 35495 13889
rect 33091 13824 33180 13852
rect 34164 13824 35296 13852
rect 35452 13852 35480 13883
rect 35526 13880 35532 13932
rect 35584 13920 35590 13932
rect 36096 13929 36124 13960
rect 35805 13923 35863 13929
rect 35805 13920 35817 13923
rect 35584 13892 35817 13920
rect 35584 13880 35590 13892
rect 35805 13889 35817 13892
rect 35851 13889 35863 13923
rect 35805 13883 35863 13889
rect 35989 13923 36047 13929
rect 35989 13889 36001 13923
rect 36035 13889 36047 13923
rect 35989 13883 36047 13889
rect 36081 13923 36139 13929
rect 36081 13889 36093 13923
rect 36127 13889 36139 13923
rect 36081 13883 36139 13889
rect 38565 13923 38623 13929
rect 38565 13889 38577 13923
rect 38611 13920 38623 13923
rect 38654 13920 38660 13932
rect 38611 13892 38660 13920
rect 38611 13889 38623 13892
rect 38565 13883 38623 13889
rect 35894 13852 35900 13864
rect 35452 13824 35900 13852
rect 33091 13821 33103 13824
rect 33045 13815 33103 13821
rect 32508 13784 32536 13815
rect 33152 13793 33180 13824
rect 31956 13756 32536 13784
rect 33137 13787 33195 13793
rect 25130 13716 25136 13728
rect 23808 13688 25136 13716
rect 23808 13676 23814 13688
rect 25130 13676 25136 13688
rect 25188 13676 25194 13728
rect 25314 13676 25320 13728
rect 25372 13716 25378 13728
rect 25501 13719 25559 13725
rect 25501 13716 25513 13719
rect 25372 13688 25513 13716
rect 25372 13676 25378 13688
rect 25501 13685 25513 13688
rect 25547 13685 25559 13719
rect 25501 13679 25559 13685
rect 26234 13676 26240 13728
rect 26292 13716 26298 13728
rect 26329 13719 26387 13725
rect 26329 13716 26341 13719
rect 26292 13688 26341 13716
rect 26292 13676 26298 13688
rect 26329 13685 26341 13688
rect 26375 13685 26387 13719
rect 26329 13679 26387 13685
rect 27065 13719 27123 13725
rect 27065 13685 27077 13719
rect 27111 13716 27123 13719
rect 27246 13716 27252 13728
rect 27111 13688 27252 13716
rect 27111 13685 27123 13688
rect 27065 13679 27123 13685
rect 27246 13676 27252 13688
rect 27304 13676 27310 13728
rect 27525 13719 27583 13725
rect 27525 13685 27537 13719
rect 27571 13716 27583 13719
rect 28445 13719 28503 13725
rect 28445 13716 28457 13719
rect 27571 13688 28457 13716
rect 27571 13685 27583 13688
rect 27525 13679 27583 13685
rect 28445 13685 28457 13688
rect 28491 13685 28503 13719
rect 28445 13679 28503 13685
rect 31846 13676 31852 13728
rect 31904 13716 31910 13728
rect 31956 13716 31984 13756
rect 33137 13753 33149 13787
rect 33183 13753 33195 13787
rect 33873 13787 33931 13793
rect 33873 13784 33885 13787
rect 33137 13747 33195 13753
rect 33336 13756 33885 13784
rect 31904 13688 31984 13716
rect 32861 13719 32919 13725
rect 31904 13676 31910 13688
rect 32861 13685 32873 13719
rect 32907 13716 32919 13719
rect 33336 13716 33364 13756
rect 33873 13753 33885 13756
rect 33919 13753 33931 13787
rect 33873 13747 33931 13753
rect 34790 13744 34796 13796
rect 34848 13784 34854 13796
rect 34885 13787 34943 13793
rect 34885 13784 34897 13787
rect 34848 13756 34897 13784
rect 34848 13744 34854 13756
rect 34885 13753 34897 13756
rect 34931 13753 34943 13787
rect 34885 13747 34943 13753
rect 32907 13688 33364 13716
rect 32907 13685 32919 13688
rect 32861 13679 32919 13685
rect 33686 13676 33692 13728
rect 33744 13716 33750 13728
rect 33962 13716 33968 13728
rect 33744 13688 33968 13716
rect 33744 13676 33750 13688
rect 33962 13676 33968 13688
rect 34020 13676 34026 13728
rect 35268 13716 35296 13824
rect 35894 13812 35900 13824
rect 35952 13812 35958 13864
rect 36004 13784 36032 13883
rect 38654 13880 38660 13892
rect 38712 13880 38718 13932
rect 36357 13855 36415 13861
rect 36357 13821 36369 13855
rect 36403 13852 36415 13855
rect 38286 13852 38292 13864
rect 36403 13824 38292 13852
rect 36403 13821 36415 13824
rect 36357 13815 36415 13821
rect 36262 13784 36268 13796
rect 35912 13756 36268 13784
rect 35912 13716 35940 13756
rect 36262 13744 36268 13756
rect 36320 13744 36326 13796
rect 35268 13688 35940 13716
rect 35986 13676 35992 13728
rect 36044 13716 36050 13728
rect 36372 13716 36400 13815
rect 38286 13812 38292 13824
rect 38344 13812 38350 13864
rect 38470 13812 38476 13864
rect 38528 13852 38534 13864
rect 38746 13852 38752 13864
rect 38528 13824 38752 13852
rect 38528 13812 38534 13824
rect 38746 13812 38752 13824
rect 38804 13812 38810 13864
rect 38948 13861 38976 14028
rect 39390 14016 39396 14028
rect 39448 14016 39454 14068
rect 39298 13948 39304 14000
rect 39356 13948 39362 14000
rect 40034 13948 40040 14000
rect 40092 13948 40098 14000
rect 38933 13855 38991 13861
rect 38933 13821 38945 13855
rect 38979 13821 38991 13855
rect 38933 13815 38991 13821
rect 39022 13812 39028 13864
rect 39080 13812 39086 13864
rect 41049 13855 41107 13861
rect 41049 13821 41061 13855
rect 41095 13821 41107 13855
rect 41049 13815 41107 13821
rect 39040 13784 39068 13812
rect 38396 13756 39068 13784
rect 38396 13728 38424 13756
rect 36044 13688 36400 13716
rect 36044 13676 36050 13688
rect 38378 13676 38384 13728
rect 38436 13676 38442 13728
rect 38654 13676 38660 13728
rect 38712 13716 38718 13728
rect 39758 13716 39764 13728
rect 38712 13688 39764 13716
rect 38712 13676 38718 13688
rect 39758 13676 39764 13688
rect 39816 13716 39822 13728
rect 41064 13716 41092 13815
rect 39816 13688 41092 13716
rect 39816 13676 39822 13688
rect 1104 13626 41400 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 41400 13626
rect 1104 13552 41400 13574
rect 5721 13515 5779 13521
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 6270 13512 6276 13524
rect 5767 13484 6276 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 6270 13472 6276 13484
rect 6328 13512 6334 13524
rect 6730 13512 6736 13524
rect 6328 13484 6736 13512
rect 6328 13472 6334 13484
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 10962 13512 10968 13524
rect 8536 13484 10968 13512
rect 8536 13472 8542 13484
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11940 13484 12081 13512
rect 11940 13472 11946 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 16482 13512 16488 13524
rect 12860 13484 16488 13512
rect 12860 13472 12866 13484
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 16853 13515 16911 13521
rect 16853 13481 16865 13515
rect 16899 13512 16911 13515
rect 19334 13512 19340 13524
rect 16899 13484 19340 13512
rect 16899 13481 16911 13484
rect 16853 13475 16911 13481
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 23566 13512 23572 13524
rect 22066 13484 23572 13512
rect 7374 13444 7380 13456
rect 5920 13416 7380 13444
rect 5718 13336 5724 13388
rect 5776 13376 5782 13388
rect 5920 13376 5948 13416
rect 7374 13404 7380 13416
rect 7432 13404 7438 13456
rect 16022 13444 16028 13456
rect 11716 13416 16028 13444
rect 6822 13376 6828 13388
rect 5776 13348 5948 13376
rect 5776 13336 5782 13348
rect 5920 13317 5948 13348
rect 6288 13348 6828 13376
rect 6288 13317 6316 13348
rect 6822 13336 6828 13348
rect 6880 13376 6886 13388
rect 6880 13348 8064 13376
rect 6880 13336 6886 13348
rect 8036 13320 8064 13348
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 6181 13311 6239 13317
rect 6181 13277 6193 13311
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 6196 13240 6224 13271
rect 6730 13240 6736 13252
rect 6196 13212 6736 13240
rect 6730 13200 6736 13212
rect 6788 13200 6794 13252
rect 7944 13240 7972 13271
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 8076 13280 8125 13308
rect 8076 13268 8082 13280
rect 8113 13277 8125 13280
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8386 13240 8392 13252
rect 7944 13212 8392 13240
rect 8386 13200 8392 13212
rect 8444 13200 8450 13252
rect 11716 13184 11744 13416
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 17589 13447 17647 13453
rect 17589 13444 17601 13447
rect 16132 13416 17601 13444
rect 12710 13336 12716 13388
rect 12768 13336 12774 13388
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13376 13415 13379
rect 13446 13376 13452 13388
rect 13403 13348 13452 13376
rect 13403 13345 13415 13348
rect 13357 13339 13415 13345
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13308 12495 13311
rect 12986 13308 12992 13320
rect 12483 13280 12992 13308
rect 12483 13277 12495 13280
rect 12437 13271 12495 13277
rect 12986 13268 12992 13280
rect 13044 13308 13050 13320
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 13044 13280 13277 13308
rect 13044 13268 13050 13280
rect 13265 13277 13277 13280
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 13372 13252 13400 13339
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 13538 13336 13544 13388
rect 13596 13376 13602 13388
rect 13596 13348 15792 13376
rect 13596 13336 13602 13348
rect 12529 13243 12587 13249
rect 12529 13209 12541 13243
rect 12575 13240 12587 13243
rect 13354 13240 13360 13252
rect 12575 13212 13360 13240
rect 12575 13209 12587 13212
rect 12529 13203 12587 13209
rect 13354 13200 13360 13212
rect 13412 13200 13418 13252
rect 6089 13175 6147 13181
rect 6089 13141 6101 13175
rect 6135 13172 6147 13175
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6135 13144 6377 13172
rect 6135 13141 6147 13144
rect 6089 13135 6147 13141
rect 6365 13141 6377 13144
rect 6411 13172 6423 13175
rect 6914 13172 6920 13184
rect 6411 13144 6920 13172
rect 6411 13141 6423 13144
rect 6365 13135 6423 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 8018 13132 8024 13184
rect 8076 13132 8082 13184
rect 11698 13132 11704 13184
rect 11756 13132 11762 13184
rect 12894 13132 12900 13184
rect 12952 13132 12958 13184
rect 15764 13172 15792 13348
rect 15838 13200 15844 13252
rect 15896 13240 15902 13252
rect 16132 13240 16160 13416
rect 17589 13413 17601 13416
rect 17635 13413 17647 13447
rect 17589 13407 17647 13413
rect 20717 13447 20775 13453
rect 20717 13413 20729 13447
rect 20763 13444 20775 13447
rect 20990 13444 20996 13456
rect 20763 13416 20996 13444
rect 20763 13413 20775 13416
rect 20717 13407 20775 13413
rect 20990 13404 20996 13416
rect 21048 13444 21054 13456
rect 21818 13444 21824 13456
rect 21048 13416 21824 13444
rect 21048 13404 21054 13416
rect 21818 13404 21824 13416
rect 21876 13404 21882 13456
rect 17126 13376 17132 13388
rect 16224 13348 17132 13376
rect 16224 13317 16252 13348
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 17218 13336 17224 13388
rect 17276 13336 17282 13388
rect 17402 13336 17408 13388
rect 17460 13376 17466 13388
rect 18046 13376 18052 13388
rect 17460 13348 18052 13376
rect 17460 13336 17466 13348
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 20162 13336 20168 13388
rect 20220 13376 20226 13388
rect 20533 13379 20591 13385
rect 20533 13376 20545 13379
rect 20220 13348 20545 13376
rect 20220 13336 20226 13348
rect 20533 13345 20545 13348
rect 20579 13345 20591 13379
rect 22066 13376 22094 13484
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 24578 13472 24584 13524
rect 24636 13512 24642 13524
rect 30098 13512 30104 13524
rect 24636 13484 30104 13512
rect 24636 13472 24642 13484
rect 22278 13404 22284 13456
rect 22336 13444 22342 13456
rect 22336 13416 24624 13444
rect 22336 13404 22342 13416
rect 20533 13339 20591 13345
rect 20732 13348 22094 13376
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 16298 13268 16304 13320
rect 16356 13268 16362 13320
rect 16715 13311 16773 13317
rect 16715 13277 16727 13311
rect 16761 13308 16773 13311
rect 18230 13308 18236 13320
rect 16761 13280 18236 13308
rect 16761 13277 16773 13280
rect 16715 13271 16773 13277
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 20732 13308 20760 13348
rect 22186 13336 22192 13388
rect 22244 13376 22250 13388
rect 22244 13348 23612 13376
rect 22244 13336 22250 13348
rect 20364 13280 20760 13308
rect 20809 13311 20867 13317
rect 16485 13243 16543 13249
rect 16485 13240 16497 13243
rect 15896 13212 16497 13240
rect 15896 13200 15902 13212
rect 16485 13209 16497 13212
rect 16531 13209 16543 13243
rect 16485 13203 16543 13209
rect 16574 13200 16580 13252
rect 16632 13200 16638 13252
rect 16942 13200 16948 13252
rect 17000 13200 17006 13252
rect 20364 13249 20392 13280
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 21818 13308 21824 13320
rect 20855 13280 21824 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 21818 13268 21824 13280
rect 21876 13268 21882 13320
rect 22278 13268 22284 13320
rect 22336 13268 22342 13320
rect 22572 13317 22600 13348
rect 22373 13311 22431 13317
rect 22373 13277 22385 13311
rect 22419 13277 22431 13311
rect 22373 13271 22431 13277
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13277 22615 13311
rect 22557 13271 22615 13277
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13308 22707 13311
rect 23382 13308 23388 13320
rect 22695 13280 23388 13308
rect 22695 13277 22707 13280
rect 22649 13271 22707 13277
rect 20349 13243 20407 13249
rect 20349 13240 20361 13243
rect 17052 13212 20361 13240
rect 16114 13172 16120 13184
rect 15764 13144 16120 13172
rect 16114 13132 16120 13144
rect 16172 13132 16178 13184
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 17052 13172 17080 13212
rect 20349 13209 20361 13212
rect 20395 13209 20407 13243
rect 20349 13203 20407 13209
rect 21450 13200 21456 13252
rect 21508 13240 21514 13252
rect 22388 13240 22416 13271
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 22738 13240 22744 13252
rect 21508 13212 22744 13240
rect 21508 13200 21514 13212
rect 22738 13200 22744 13212
rect 22796 13200 22802 13252
rect 22833 13243 22891 13249
rect 22833 13209 22845 13243
rect 22879 13240 22891 13243
rect 23474 13240 23480 13252
rect 22879 13212 23480 13240
rect 22879 13209 22891 13212
rect 22833 13203 22891 13209
rect 16816 13144 17080 13172
rect 17313 13175 17371 13181
rect 16816 13132 16822 13144
rect 17313 13141 17325 13175
rect 17359 13172 17371 13175
rect 19058 13172 19064 13184
rect 17359 13144 19064 13172
rect 17359 13141 17371 13144
rect 17313 13135 17371 13141
rect 19058 13132 19064 13144
rect 19116 13172 19122 13184
rect 19242 13172 19248 13184
rect 19116 13144 19248 13172
rect 19116 13132 19122 13144
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 22094 13132 22100 13184
rect 22152 13132 22158 13184
rect 22646 13132 22652 13184
rect 22704 13172 22710 13184
rect 22848 13172 22876 13203
rect 23474 13200 23480 13212
rect 23532 13200 23538 13252
rect 23584 13240 23612 13348
rect 24596 13320 24624 13416
rect 24578 13268 24584 13320
rect 24636 13268 24642 13320
rect 24688 13317 24716 13484
rect 30098 13472 30104 13484
rect 30156 13472 30162 13524
rect 30944 13484 33088 13512
rect 25774 13444 25780 13456
rect 24780 13416 25360 13444
rect 24780 13388 24808 13416
rect 24762 13336 24768 13388
rect 24820 13336 24826 13388
rect 25130 13336 25136 13388
rect 25188 13336 25194 13388
rect 25332 13385 25360 13416
rect 25424 13416 25780 13444
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13345 25375 13379
rect 25317 13339 25375 13345
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13277 24731 13311
rect 24673 13271 24731 13277
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 24872 13240 24900 13271
rect 24946 13268 24952 13320
rect 25004 13268 25010 13320
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13308 25099 13311
rect 25148 13308 25176 13336
rect 25087 13280 25176 13308
rect 25225 13311 25283 13317
rect 25087 13277 25099 13280
rect 25041 13271 25099 13277
rect 25225 13277 25237 13311
rect 25271 13277 25283 13311
rect 25225 13271 25283 13277
rect 25240 13240 25268 13271
rect 23584 13212 24900 13240
rect 25056 13212 25268 13240
rect 25332 13240 25360 13339
rect 25424 13317 25452 13416
rect 25774 13404 25780 13416
rect 25832 13404 25838 13456
rect 25958 13404 25964 13456
rect 26016 13444 26022 13456
rect 27706 13444 27712 13456
rect 26016 13416 27712 13444
rect 26016 13404 26022 13416
rect 27706 13404 27712 13416
rect 27764 13404 27770 13456
rect 27341 13379 27399 13385
rect 27341 13376 27353 13379
rect 25514 13348 26097 13376
rect 25409 13311 25467 13317
rect 25409 13277 25421 13311
rect 25455 13277 25467 13311
rect 25409 13271 25467 13277
rect 25514 13240 25542 13348
rect 25593 13311 25651 13317
rect 25593 13277 25605 13311
rect 25639 13277 25651 13311
rect 25593 13271 25651 13277
rect 25332 13212 25542 13240
rect 25608 13240 25636 13271
rect 25958 13268 25964 13320
rect 26016 13268 26022 13320
rect 26069 13317 26097 13348
rect 26344 13348 27016 13376
rect 26054 13311 26112 13317
rect 26054 13277 26066 13311
rect 26100 13277 26112 13311
rect 26344 13308 26372 13348
rect 26054 13271 26112 13277
rect 26160 13280 26372 13308
rect 26160 13240 26188 13280
rect 26418 13268 26424 13320
rect 26476 13317 26482 13320
rect 26476 13308 26484 13317
rect 26476 13280 26521 13308
rect 26476 13271 26484 13280
rect 26476 13268 26482 13271
rect 26694 13268 26700 13320
rect 26752 13308 26758 13320
rect 26988 13317 27016 13348
rect 27172 13348 27353 13376
rect 26881 13311 26939 13317
rect 26881 13308 26893 13311
rect 26752 13280 26893 13308
rect 26752 13268 26758 13280
rect 26881 13277 26893 13280
rect 26927 13277 26939 13311
rect 26881 13271 26939 13277
rect 26973 13311 27031 13317
rect 26973 13277 26985 13311
rect 27019 13308 27031 13311
rect 27062 13308 27068 13320
rect 27019 13280 27068 13308
rect 27019 13277 27031 13280
rect 26973 13271 27031 13277
rect 27062 13268 27068 13280
rect 27120 13268 27126 13320
rect 27172 13317 27200 13348
rect 27341 13345 27353 13348
rect 27387 13345 27399 13379
rect 30944 13376 30972 13484
rect 31018 13404 31024 13456
rect 31076 13444 31082 13456
rect 31076 13416 31984 13444
rect 31076 13404 31082 13416
rect 27341 13339 27399 13345
rect 27724 13348 30972 13376
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13277 27215 13311
rect 27157 13271 27215 13277
rect 27249 13311 27307 13317
rect 27249 13277 27261 13311
rect 27295 13277 27307 13311
rect 27525 13311 27583 13317
rect 27525 13308 27537 13311
rect 27249 13271 27307 13277
rect 27356 13280 27537 13308
rect 25608 13212 26188 13240
rect 26237 13243 26295 13249
rect 25056 13184 25084 13212
rect 26237 13209 26249 13243
rect 26283 13209 26295 13243
rect 26237 13203 26295 13209
rect 22704 13144 22876 13172
rect 22704 13132 22710 13144
rect 22922 13132 22928 13184
rect 22980 13132 22986 13184
rect 24394 13132 24400 13184
rect 24452 13132 24458 13184
rect 25038 13132 25044 13184
rect 25096 13132 25102 13184
rect 25498 13132 25504 13184
rect 25556 13172 25562 13184
rect 25777 13175 25835 13181
rect 25777 13172 25789 13175
rect 25556 13144 25789 13172
rect 25556 13132 25562 13144
rect 25777 13141 25789 13144
rect 25823 13141 25835 13175
rect 26252 13172 26280 13203
rect 26326 13200 26332 13252
rect 26384 13200 26390 13252
rect 26510 13200 26516 13252
rect 26568 13200 26574 13252
rect 27264 13240 27292 13271
rect 27356 13252 27384 13280
rect 27525 13277 27537 13280
rect 27571 13277 27583 13311
rect 27525 13271 27583 13277
rect 26620 13212 27292 13240
rect 26528 13172 26556 13200
rect 26620 13181 26648 13212
rect 27338 13200 27344 13252
rect 27396 13200 27402 13252
rect 26252 13144 26556 13172
rect 26605 13175 26663 13181
rect 25777 13135 25835 13141
rect 26605 13141 26617 13175
rect 26651 13141 26663 13175
rect 26605 13135 26663 13141
rect 26694 13132 26700 13184
rect 26752 13132 26758 13184
rect 26786 13132 26792 13184
rect 26844 13172 26850 13184
rect 27724 13181 27752 13348
rect 31956 13320 31984 13416
rect 32030 13404 32036 13456
rect 32088 13404 32094 13456
rect 33060 13444 33088 13484
rect 33134 13472 33140 13524
rect 33192 13512 33198 13524
rect 33413 13515 33471 13521
rect 33413 13512 33425 13515
rect 33192 13484 33425 13512
rect 33192 13472 33198 13484
rect 33413 13481 33425 13484
rect 33459 13481 33471 13515
rect 33413 13475 33471 13481
rect 35069 13515 35127 13521
rect 35069 13481 35081 13515
rect 35115 13512 35127 13515
rect 35434 13512 35440 13524
rect 35115 13484 35440 13512
rect 35115 13481 35127 13484
rect 35069 13475 35127 13481
rect 35434 13472 35440 13484
rect 35492 13472 35498 13524
rect 35529 13515 35587 13521
rect 35529 13481 35541 13515
rect 35575 13512 35587 13515
rect 35618 13512 35624 13524
rect 35575 13484 35624 13512
rect 35575 13481 35587 13484
rect 35529 13475 35587 13481
rect 35618 13472 35624 13484
rect 35676 13472 35682 13524
rect 35894 13472 35900 13524
rect 35952 13512 35958 13524
rect 35989 13515 36047 13521
rect 35989 13512 36001 13515
rect 35952 13484 36001 13512
rect 35952 13472 35958 13484
rect 35989 13481 36001 13484
rect 36035 13481 36047 13515
rect 35989 13475 36047 13481
rect 36096 13484 36400 13512
rect 34698 13444 34704 13456
rect 33060 13416 34704 13444
rect 34698 13404 34704 13416
rect 34756 13444 34762 13456
rect 35452 13444 35480 13472
rect 36096 13444 36124 13484
rect 34756 13416 35020 13444
rect 35452 13416 36124 13444
rect 36173 13447 36231 13453
rect 34756 13404 34762 13416
rect 32048 13376 32076 13404
rect 34992 13376 35020 13416
rect 36173 13413 36185 13447
rect 36219 13444 36231 13447
rect 36262 13444 36268 13456
rect 36219 13416 36268 13444
rect 36219 13413 36231 13416
rect 36173 13407 36231 13413
rect 36262 13404 36268 13416
rect 36320 13404 36326 13456
rect 35621 13379 35679 13385
rect 35621 13376 35633 13379
rect 32048 13348 34928 13376
rect 34992 13348 35633 13376
rect 27801 13311 27859 13317
rect 27801 13277 27813 13311
rect 27847 13308 27859 13311
rect 28350 13308 28356 13320
rect 27847 13280 28356 13308
rect 27847 13277 27859 13280
rect 27801 13271 27859 13277
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 31478 13268 31484 13320
rect 31536 13268 31542 13320
rect 31570 13268 31576 13320
rect 31628 13268 31634 13320
rect 31938 13268 31944 13320
rect 31996 13268 32002 13320
rect 32048 13317 32076 13348
rect 32033 13311 32091 13317
rect 32033 13277 32045 13311
rect 32079 13277 32091 13311
rect 32033 13271 32091 13277
rect 32950 13268 32956 13320
rect 33008 13308 33014 13320
rect 33413 13311 33471 13317
rect 33413 13308 33425 13311
rect 33008 13280 33425 13308
rect 33008 13268 33014 13280
rect 33413 13277 33425 13280
rect 33459 13277 33471 13311
rect 33413 13271 33471 13277
rect 33597 13311 33655 13317
rect 33597 13277 33609 13311
rect 33643 13308 33655 13311
rect 34146 13308 34152 13320
rect 33643 13280 34152 13308
rect 33643 13277 33655 13280
rect 33597 13271 33655 13277
rect 34146 13268 34152 13280
rect 34204 13268 34210 13320
rect 34348 13317 34376 13348
rect 34333 13311 34391 13317
rect 34333 13277 34345 13311
rect 34379 13277 34391 13311
rect 34333 13271 34391 13277
rect 34422 13268 34428 13320
rect 34480 13268 34486 13320
rect 34514 13268 34520 13320
rect 34572 13308 34578 13320
rect 34900 13317 34928 13348
rect 35621 13345 35633 13348
rect 35667 13376 35679 13379
rect 35986 13376 35992 13388
rect 35667 13348 35992 13376
rect 35667 13345 35679 13348
rect 35621 13339 35679 13345
rect 35986 13336 35992 13348
rect 36044 13336 36050 13388
rect 34701 13311 34759 13317
rect 34701 13308 34713 13311
rect 34572 13280 34713 13308
rect 34572 13268 34578 13280
rect 34701 13277 34713 13280
rect 34747 13277 34759 13311
rect 34701 13271 34759 13277
rect 34885 13311 34943 13317
rect 34885 13277 34897 13311
rect 34931 13308 34943 13311
rect 35161 13311 35219 13317
rect 35161 13308 35173 13311
rect 34931 13280 35173 13308
rect 34931 13277 34943 13280
rect 34885 13271 34943 13277
rect 35161 13277 35173 13280
rect 35207 13308 35219 13311
rect 35526 13308 35532 13320
rect 35207 13280 35532 13308
rect 35207 13277 35219 13280
rect 35161 13271 35219 13277
rect 35526 13268 35532 13280
rect 35584 13268 35590 13320
rect 35805 13311 35863 13317
rect 35805 13277 35817 13311
rect 35851 13277 35863 13311
rect 35805 13271 35863 13277
rect 28994 13200 29000 13252
rect 29052 13240 29058 13252
rect 35066 13240 35072 13252
rect 29052 13212 35072 13240
rect 29052 13200 29058 13212
rect 35066 13200 35072 13212
rect 35124 13200 35130 13252
rect 35345 13243 35403 13249
rect 35345 13209 35357 13243
rect 35391 13209 35403 13243
rect 35345 13203 35403 13209
rect 27709 13175 27767 13181
rect 27709 13172 27721 13175
rect 26844 13144 27721 13172
rect 26844 13132 26850 13144
rect 27709 13141 27721 13144
rect 27755 13141 27767 13175
rect 27709 13135 27767 13141
rect 31294 13132 31300 13184
rect 31352 13172 31358 13184
rect 31757 13175 31815 13181
rect 31757 13172 31769 13175
rect 31352 13144 31769 13172
rect 31352 13132 31358 13144
rect 31757 13141 31769 13144
rect 31803 13141 31815 13175
rect 31757 13135 31815 13141
rect 32214 13132 32220 13184
rect 32272 13132 32278 13184
rect 34698 13132 34704 13184
rect 34756 13172 34762 13184
rect 35360 13172 35388 13203
rect 35710 13200 35716 13252
rect 35768 13240 35774 13252
rect 35820 13240 35848 13271
rect 35894 13268 35900 13320
rect 35952 13308 35958 13320
rect 36372 13317 36400 13484
rect 38930 13472 38936 13524
rect 38988 13472 38994 13524
rect 38657 13447 38715 13453
rect 38657 13413 38669 13447
rect 38703 13444 38715 13447
rect 38948 13444 38976 13472
rect 38703 13416 38976 13444
rect 38703 13413 38715 13416
rect 38657 13407 38715 13413
rect 38562 13336 38568 13388
rect 38620 13376 38626 13388
rect 38933 13379 38991 13385
rect 38933 13376 38945 13379
rect 38620 13348 38945 13376
rect 38620 13336 38626 13348
rect 38933 13345 38945 13348
rect 38979 13345 38991 13379
rect 39577 13379 39635 13385
rect 39577 13376 39589 13379
rect 38933 13339 38991 13345
rect 39408 13348 39589 13376
rect 39408 13320 39436 13348
rect 39577 13345 39589 13348
rect 39623 13345 39635 13379
rect 39577 13339 39635 13345
rect 36173 13311 36231 13317
rect 36173 13308 36185 13311
rect 35952 13280 36185 13308
rect 35952 13268 35958 13280
rect 36173 13277 36185 13280
rect 36219 13277 36231 13311
rect 36173 13271 36231 13277
rect 36357 13311 36415 13317
rect 36357 13277 36369 13311
rect 36403 13277 36415 13311
rect 38378 13308 38384 13320
rect 36357 13271 36415 13277
rect 36556 13280 38384 13308
rect 35768 13212 35848 13240
rect 35768 13200 35774 13212
rect 36262 13200 36268 13252
rect 36320 13240 36326 13252
rect 36556 13240 36584 13280
rect 38378 13268 38384 13280
rect 38436 13308 38442 13320
rect 38473 13311 38531 13317
rect 38473 13308 38485 13311
rect 38436 13280 38485 13308
rect 38436 13268 38442 13280
rect 38473 13277 38485 13280
rect 38519 13277 38531 13311
rect 38473 13271 38531 13277
rect 38654 13268 38660 13320
rect 38712 13268 38718 13320
rect 38841 13311 38899 13317
rect 38841 13277 38853 13311
rect 38887 13308 38899 13311
rect 39114 13308 39120 13320
rect 38887 13280 39120 13308
rect 38887 13277 38899 13280
rect 38841 13271 38899 13277
rect 39114 13268 39120 13280
rect 39172 13268 39178 13320
rect 39390 13268 39396 13320
rect 39448 13268 39454 13320
rect 39485 13311 39543 13317
rect 39485 13277 39497 13311
rect 39531 13308 39543 13311
rect 39758 13308 39764 13320
rect 39531 13280 39764 13308
rect 39531 13277 39543 13280
rect 39485 13271 39543 13277
rect 39758 13268 39764 13280
rect 39816 13268 39822 13320
rect 39945 13311 40003 13317
rect 39945 13277 39957 13311
rect 39991 13308 40003 13311
rect 40497 13311 40555 13317
rect 40497 13308 40509 13311
rect 39991 13280 40509 13308
rect 39991 13277 40003 13280
rect 39945 13271 40003 13277
rect 40497 13277 40509 13280
rect 40543 13308 40555 13311
rect 40543 13280 41460 13308
rect 40543 13277 40555 13280
rect 40497 13271 40555 13277
rect 36320 13212 36584 13240
rect 36320 13200 36326 13212
rect 36630 13200 36636 13252
rect 36688 13240 36694 13252
rect 37645 13243 37703 13249
rect 37645 13240 37657 13243
rect 36688 13212 37657 13240
rect 36688 13200 36694 13212
rect 37645 13209 37657 13212
rect 37691 13209 37703 13243
rect 37645 13203 37703 13209
rect 38746 13200 38752 13252
rect 38804 13240 38810 13252
rect 39408 13240 39436 13268
rect 38804 13212 39436 13240
rect 38804 13200 38810 13212
rect 34756 13144 35388 13172
rect 39485 13175 39543 13181
rect 34756 13132 34762 13144
rect 39485 13141 39497 13175
rect 39531 13172 39543 13175
rect 39758 13172 39764 13184
rect 39531 13144 39764 13172
rect 39531 13141 39543 13144
rect 39485 13135 39543 13141
rect 39758 13132 39764 13144
rect 39816 13132 39822 13184
rect 39850 13132 39856 13184
rect 39908 13172 39914 13184
rect 40037 13175 40095 13181
rect 40037 13172 40049 13175
rect 39908 13144 40049 13172
rect 39908 13132 39914 13144
rect 40037 13141 40049 13144
rect 40083 13141 40095 13175
rect 40037 13135 40095 13141
rect 41046 13132 41052 13184
rect 41104 13132 41110 13184
rect 1104 13082 41400 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 41400 13082
rect 1104 13008 41400 13030
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 6380 12940 7941 12968
rect 6086 12860 6092 12912
rect 6144 12900 6150 12912
rect 6270 12900 6276 12912
rect 6144 12872 6276 12900
rect 6144 12860 6150 12872
rect 6270 12860 6276 12872
rect 6328 12860 6334 12912
rect 6380 12909 6408 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 7929 12931 7987 12937
rect 8018 12928 8024 12980
rect 8076 12928 8082 12980
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 8754 12968 8760 12980
rect 8628 12940 8760 12968
rect 8628 12928 8634 12940
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12937 9275 12971
rect 10778 12968 10784 12980
rect 9217 12931 9275 12937
rect 9600 12940 10784 12968
rect 6365 12903 6423 12909
rect 6365 12869 6377 12903
rect 6411 12869 6423 12903
rect 6365 12863 6423 12869
rect 6549 12903 6607 12909
rect 6549 12869 6561 12903
rect 6595 12900 6607 12903
rect 6825 12903 6883 12909
rect 6825 12900 6837 12903
rect 6595 12872 6837 12900
rect 6595 12869 6607 12872
rect 6549 12863 6607 12869
rect 6825 12869 6837 12872
rect 6871 12869 6883 12903
rect 6825 12863 6883 12869
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 4908 12696 4936 12795
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 5166 12792 5172 12844
rect 5224 12792 5230 12844
rect 5258 12792 5264 12844
rect 5316 12792 5322 12844
rect 6638 12792 6644 12844
rect 6696 12792 6702 12844
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7374 12792 7380 12844
rect 7432 12792 7438 12844
rect 7834 12792 7840 12844
rect 7892 12792 7898 12844
rect 7926 12792 7932 12844
rect 7984 12792 7990 12844
rect 8036 12832 8064 12928
rect 9232 12900 9260 12931
rect 8220 12872 9260 12900
rect 8220 12841 8248 12872
rect 9600 12844 9628 12940
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 11882 12968 11888 12980
rect 11480 12940 11888 12968
rect 11480 12928 11486 12940
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12345 12971 12403 12977
rect 12345 12937 12357 12971
rect 12391 12937 12403 12971
rect 12345 12931 12403 12937
rect 12713 12971 12771 12977
rect 12713 12937 12725 12971
rect 12759 12968 12771 12971
rect 12894 12968 12900 12980
rect 12759 12940 12900 12968
rect 12759 12937 12771 12940
rect 12713 12931 12771 12937
rect 9953 12903 10011 12909
rect 9953 12900 9965 12903
rect 9692 12872 9965 12900
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 8036 12804 8125 12832
rect 8113 12801 8125 12804
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8205 12835 8263 12841
rect 8205 12801 8217 12835
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 5276 12764 5304 12792
rect 7024 12764 7052 12792
rect 5276 12736 7052 12764
rect 5442 12696 5448 12708
rect 4908 12668 5448 12696
rect 5442 12656 5448 12668
rect 5500 12696 5506 12708
rect 6822 12696 6828 12708
rect 5500 12668 6828 12696
rect 5500 12656 5506 12668
rect 6822 12656 6828 12668
rect 6880 12656 6886 12708
rect 7392 12696 7420 12792
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 7944 12764 7972 12792
rect 7791 12736 7972 12764
rect 8496 12764 8524 12795
rect 8570 12792 8576 12844
rect 8628 12792 8634 12844
rect 8721 12835 8779 12841
rect 8721 12801 8733 12835
rect 8767 12832 8779 12835
rect 8767 12801 8800 12832
rect 8721 12795 8800 12801
rect 8496 12736 8616 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 8588 12696 8616 12736
rect 7392 12668 8616 12696
rect 8772 12696 8800 12795
rect 8846 12792 8852 12844
rect 8904 12792 8910 12844
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 9122 12841 9128 12844
rect 9079 12835 9128 12841
rect 9079 12801 9091 12835
rect 9125 12801 9128 12835
rect 9079 12795 9128 12801
rect 9122 12792 9128 12795
rect 9180 12832 9186 12844
rect 9582 12832 9588 12844
rect 9180 12804 9588 12832
rect 9180 12792 9186 12804
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 9692 12841 9720 12872
rect 9953 12869 9965 12872
rect 9999 12900 10011 12903
rect 12360 12900 12388 12931
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 16485 12971 16543 12977
rect 15212 12940 16436 12968
rect 15212 12900 15240 12940
rect 9999 12872 12388 12900
rect 12728 12872 15240 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 12728 12844 12756 12872
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 16408 12900 16436 12940
rect 16485 12937 16497 12971
rect 16531 12968 16543 12971
rect 16574 12968 16580 12980
rect 16531 12940 16580 12968
rect 16531 12937 16543 12940
rect 16485 12931 16543 12937
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17678 12968 17684 12980
rect 17184 12940 17684 12968
rect 17184 12928 17190 12940
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 19518 12968 19524 12980
rect 18524 12940 19524 12968
rect 18524 12900 18552 12940
rect 19518 12928 19524 12940
rect 19576 12928 19582 12980
rect 19705 12971 19763 12977
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 20714 12968 20720 12980
rect 19751 12940 20720 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 24946 12928 24952 12980
rect 25004 12968 25010 12980
rect 25590 12968 25596 12980
rect 25004 12940 25596 12968
rect 25004 12928 25010 12940
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 31386 12928 31392 12980
rect 31444 12968 31450 12980
rect 31846 12968 31852 12980
rect 31444 12940 31852 12968
rect 31444 12928 31450 12940
rect 31846 12928 31852 12940
rect 31904 12928 31910 12980
rect 36170 12968 36176 12980
rect 33060 12940 36176 12968
rect 15344 12872 15502 12900
rect 16408 12872 18552 12900
rect 15344 12860 15350 12872
rect 18598 12860 18604 12912
rect 18656 12900 18662 12912
rect 18656 12872 19196 12900
rect 18656 12860 18662 12872
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 10778 12832 10784 12844
rect 10183 12804 10784 12832
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12764 9551 12767
rect 9766 12764 9772 12776
rect 9539 12736 9772 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 9766 12724 9772 12736
rect 9824 12764 9830 12776
rect 10152 12764 10180 12795
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 12710 12792 12716 12844
rect 12768 12792 12774 12844
rect 12802 12792 12808 12844
rect 12860 12792 12866 12844
rect 14090 12792 14096 12844
rect 14148 12832 14154 12844
rect 14737 12835 14795 12841
rect 14737 12832 14749 12835
rect 14148 12804 14749 12832
rect 14148 12792 14154 12804
rect 14737 12801 14749 12804
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17862 12832 17868 12844
rect 17000 12804 17868 12832
rect 17000 12792 17006 12804
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 18782 12832 18788 12844
rect 18288 12804 18788 12832
rect 18288 12792 18294 12804
rect 18782 12792 18788 12804
rect 18840 12832 18846 12844
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18840 12804 19073 12832
rect 18840 12792 18846 12804
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 9824 12736 10180 12764
rect 9824 12724 9830 12736
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 11112 12736 11529 12764
rect 11112 12724 11118 12736
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 12618 12764 12624 12776
rect 12400 12736 12624 12764
rect 12400 12724 12406 12736
rect 12618 12724 12624 12736
rect 12676 12764 12682 12776
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12676 12736 12909 12764
rect 12676 12724 12682 12736
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 18012 12736 18981 12764
rect 18012 12724 18018 12736
rect 18969 12733 18981 12736
rect 19015 12764 19027 12767
rect 19168 12764 19196 12872
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 19392 12872 20116 12900
rect 19392 12860 19398 12872
rect 19242 12792 19248 12844
rect 19300 12832 19306 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 19300 12804 19441 12832
rect 19300 12792 19306 12804
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 19521 12835 19579 12841
rect 19521 12801 19533 12835
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 19536 12764 19564 12795
rect 19978 12792 19984 12844
rect 20036 12792 20042 12844
rect 20088 12841 20116 12872
rect 20732 12872 23520 12900
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 20162 12792 20168 12844
rect 20220 12792 20226 12844
rect 20254 12792 20260 12844
rect 20312 12832 20318 12844
rect 20732 12841 20760 12872
rect 23492 12844 23520 12872
rect 23934 12860 23940 12912
rect 23992 12900 23998 12912
rect 24121 12903 24179 12909
rect 24121 12900 24133 12903
rect 23992 12872 24133 12900
rect 23992 12860 23998 12872
rect 24121 12869 24133 12872
rect 24167 12869 24179 12903
rect 24121 12863 24179 12869
rect 24210 12860 24216 12912
rect 24268 12900 24274 12912
rect 25314 12900 25320 12912
rect 24268 12872 25320 12900
rect 24268 12860 24274 12872
rect 25314 12860 25320 12872
rect 25372 12860 25378 12912
rect 25682 12860 25688 12912
rect 25740 12860 25746 12912
rect 28810 12860 28816 12912
rect 28868 12900 28874 12912
rect 28994 12900 29000 12912
rect 28868 12872 29000 12900
rect 28868 12860 28874 12872
rect 28994 12860 29000 12872
rect 29052 12860 29058 12912
rect 29270 12860 29276 12912
rect 29328 12900 29334 12912
rect 29549 12903 29607 12909
rect 29549 12900 29561 12903
rect 29328 12872 29561 12900
rect 29328 12860 29334 12872
rect 29549 12869 29561 12872
rect 29595 12869 29607 12903
rect 29549 12863 29607 12869
rect 30742 12860 30748 12912
rect 30800 12900 30806 12912
rect 31481 12903 31539 12909
rect 31481 12900 31493 12903
rect 30800 12872 31493 12900
rect 30800 12860 30806 12872
rect 31481 12869 31493 12872
rect 31527 12869 31539 12903
rect 32214 12900 32220 12912
rect 31481 12863 31539 12869
rect 31588 12872 32220 12900
rect 20349 12835 20407 12841
rect 20349 12832 20361 12835
rect 20312 12804 20361 12832
rect 20312 12792 20318 12804
rect 20349 12801 20361 12804
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12832 21051 12835
rect 21082 12832 21088 12844
rect 21039 12804 21088 12832
rect 21039 12801 21051 12804
rect 20993 12795 21051 12801
rect 20732 12764 20760 12795
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 23474 12792 23480 12844
rect 23532 12792 23538 12844
rect 23658 12792 23664 12844
rect 23716 12832 23722 12844
rect 23753 12835 23811 12841
rect 23753 12832 23765 12835
rect 23716 12804 23765 12832
rect 23716 12792 23722 12804
rect 23753 12801 23765 12804
rect 23799 12801 23811 12835
rect 23753 12795 23811 12801
rect 23845 12835 23903 12841
rect 23845 12801 23857 12835
rect 23891 12832 23903 12835
rect 24578 12832 24584 12844
rect 23891 12804 24584 12832
rect 23891 12801 23903 12804
rect 23845 12795 23903 12801
rect 24578 12792 24584 12804
rect 24636 12792 24642 12844
rect 25700 12832 25728 12860
rect 24688 12804 25728 12832
rect 31205 12835 31263 12841
rect 19015 12736 19104 12764
rect 19168 12736 19564 12764
rect 20272 12736 20760 12764
rect 19015 12733 19027 12736
rect 18969 12727 19027 12733
rect 19076 12708 19104 12736
rect 9030 12696 9036 12708
rect 8772 12668 9036 12696
rect 4890 12588 4896 12640
rect 4948 12588 4954 12640
rect 6362 12588 6368 12640
rect 6420 12588 6426 12640
rect 8386 12588 8392 12640
rect 8444 12588 8450 12640
rect 8588 12628 8616 12668
rect 9030 12656 9036 12668
rect 9088 12696 9094 12708
rect 9088 12668 9996 12696
rect 9088 12656 9094 12668
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 8588 12600 9873 12628
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 9968 12628 9996 12668
rect 10042 12656 10048 12708
rect 10100 12696 10106 12708
rect 10100 12668 12020 12696
rect 10100 12656 10106 12668
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9968 12600 10333 12628
rect 9861 12591 9919 12597
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 11992 12628 12020 12668
rect 13538 12656 13544 12708
rect 13596 12656 13602 12708
rect 16114 12656 16120 12708
rect 16172 12696 16178 12708
rect 16172 12668 19012 12696
rect 16172 12656 16178 12668
rect 13556 12628 13584 12656
rect 15010 12637 15016 12640
rect 11992 12600 13584 12628
rect 15000 12631 15016 12637
rect 10321 12591 10379 12597
rect 15000 12597 15012 12631
rect 15000 12591 15016 12597
rect 15010 12588 15016 12591
rect 15068 12588 15074 12640
rect 15378 12588 15384 12640
rect 15436 12628 15442 12640
rect 15654 12628 15660 12640
rect 15436 12600 15660 12628
rect 15436 12588 15442 12600
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 18509 12631 18567 12637
rect 18509 12597 18521 12631
rect 18555 12628 18567 12631
rect 18874 12628 18880 12640
rect 18555 12600 18880 12628
rect 18555 12597 18567 12600
rect 18509 12591 18567 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 18984 12628 19012 12668
rect 19058 12656 19064 12708
rect 19116 12656 19122 12708
rect 19150 12656 19156 12708
rect 19208 12696 19214 12708
rect 20272 12696 20300 12736
rect 20806 12724 20812 12776
rect 20864 12724 20870 12776
rect 24688 12764 24716 12804
rect 31205 12801 31217 12835
rect 31251 12801 31263 12835
rect 31205 12795 31263 12801
rect 21192 12736 24716 12764
rect 21192 12705 21220 12736
rect 25038 12724 25044 12776
rect 25096 12764 25102 12776
rect 28626 12764 28632 12776
rect 25096 12736 28632 12764
rect 25096 12724 25102 12736
rect 28626 12724 28632 12736
rect 28684 12724 28690 12776
rect 31220 12764 31248 12795
rect 31294 12792 31300 12844
rect 31352 12792 31358 12844
rect 31588 12841 31616 12872
rect 32214 12860 32220 12872
rect 32272 12860 32278 12912
rect 31573 12835 31631 12841
rect 31573 12801 31585 12835
rect 31619 12801 31631 12835
rect 31573 12795 31631 12801
rect 31754 12792 31760 12844
rect 31812 12792 31818 12844
rect 33060 12841 33088 12940
rect 36170 12928 36176 12940
rect 36228 12928 36234 12980
rect 38654 12968 38660 12980
rect 37844 12940 38660 12968
rect 33226 12860 33232 12912
rect 33284 12900 33290 12912
rect 33321 12903 33379 12909
rect 33321 12900 33333 12903
rect 33284 12872 33333 12900
rect 33284 12860 33290 12872
rect 33321 12869 33333 12872
rect 33367 12869 33379 12903
rect 33321 12863 33379 12869
rect 33778 12860 33784 12912
rect 33836 12860 33842 12912
rect 35066 12860 35072 12912
rect 35124 12900 35130 12912
rect 36630 12900 36636 12912
rect 35124 12872 36636 12900
rect 35124 12860 35130 12872
rect 36630 12860 36636 12872
rect 36688 12860 36694 12912
rect 33045 12835 33103 12841
rect 33045 12801 33057 12835
rect 33091 12801 33103 12835
rect 33045 12795 33103 12801
rect 37458 12792 37464 12844
rect 37516 12792 37522 12844
rect 31386 12764 31392 12776
rect 31220 12736 31392 12764
rect 31386 12724 31392 12736
rect 31444 12724 31450 12776
rect 31481 12767 31539 12773
rect 31481 12733 31493 12767
rect 31527 12764 31539 12767
rect 31662 12764 31668 12776
rect 31527 12736 31668 12764
rect 31527 12733 31539 12736
rect 31481 12727 31539 12733
rect 31662 12724 31668 12736
rect 31720 12724 31726 12776
rect 34514 12724 34520 12776
rect 34572 12764 34578 12776
rect 34793 12767 34851 12773
rect 34793 12764 34805 12767
rect 34572 12736 34805 12764
rect 34572 12724 34578 12736
rect 34793 12733 34805 12736
rect 34839 12733 34851 12767
rect 34793 12727 34851 12733
rect 37366 12724 37372 12776
rect 37424 12724 37430 12776
rect 37844 12773 37872 12940
rect 38654 12928 38660 12940
rect 38712 12928 38718 12980
rect 41049 12971 41107 12977
rect 41049 12937 41061 12971
rect 41095 12968 41107 12971
rect 41432 12968 41460 13280
rect 41095 12940 41460 12968
rect 41095 12937 41107 12940
rect 41049 12931 41107 12937
rect 40034 12860 40040 12912
rect 40092 12860 40098 12912
rect 38378 12792 38384 12844
rect 38436 12832 38442 12844
rect 39301 12835 39359 12841
rect 39301 12832 39313 12835
rect 38436 12804 39313 12832
rect 38436 12792 38442 12804
rect 39301 12801 39313 12804
rect 39347 12801 39359 12835
rect 39301 12795 39359 12801
rect 37829 12767 37887 12773
rect 37829 12733 37841 12767
rect 37875 12733 37887 12767
rect 37829 12727 37887 12733
rect 39574 12724 39580 12776
rect 39632 12724 39638 12776
rect 19208 12668 20300 12696
rect 21177 12699 21235 12705
rect 19208 12656 19214 12668
rect 21177 12665 21189 12699
rect 21223 12665 21235 12699
rect 21177 12659 21235 12665
rect 23474 12656 23480 12708
rect 23532 12696 23538 12708
rect 25056 12696 25084 12724
rect 23532 12668 25084 12696
rect 23532 12656 23538 12668
rect 27062 12656 27068 12708
rect 27120 12696 27126 12708
rect 32214 12696 32220 12708
rect 27120 12668 32220 12696
rect 27120 12656 27126 12668
rect 32214 12656 32220 12668
rect 32272 12656 32278 12708
rect 20714 12628 20720 12640
rect 18984 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 23569 12631 23627 12637
rect 23569 12597 23581 12631
rect 23615 12628 23627 12631
rect 23934 12628 23940 12640
rect 23615 12600 23940 12628
rect 23615 12597 23627 12600
rect 23569 12591 23627 12597
rect 23934 12588 23940 12600
rect 23992 12588 23998 12640
rect 26602 12588 26608 12640
rect 26660 12628 26666 12640
rect 32582 12628 32588 12640
rect 26660 12600 32588 12628
rect 26660 12588 26666 12600
rect 32582 12588 32588 12600
rect 32640 12588 32646 12640
rect 33042 12588 33048 12640
rect 33100 12628 33106 12640
rect 39666 12628 39672 12640
rect 33100 12600 39672 12628
rect 33100 12588 33106 12600
rect 39666 12588 39672 12600
rect 39724 12588 39730 12640
rect 1104 12538 41400 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 41400 12538
rect 1104 12464 41400 12486
rect 6365 12427 6423 12433
rect 2608 12396 5120 12424
rect 2608 12229 2636 12396
rect 5092 12356 5120 12396
rect 6365 12393 6377 12427
rect 6411 12424 6423 12427
rect 6638 12424 6644 12436
rect 6411 12396 6644 12424
rect 6411 12393 6423 12396
rect 6365 12387 6423 12393
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 8662 12424 8668 12436
rect 8260 12396 8668 12424
rect 8260 12384 8266 12396
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 9490 12424 9496 12436
rect 9364 12396 9496 12424
rect 9364 12384 9370 12396
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 10778 12384 10784 12436
rect 10836 12384 10842 12436
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 12986 12424 12992 12436
rect 11756 12396 12992 12424
rect 11756 12384 11762 12396
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13354 12424 13360 12436
rect 13280 12396 13360 12424
rect 5092 12328 10732 12356
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 3752 12260 3801 12288
rect 3752 12248 3758 12260
rect 3789 12257 3801 12260
rect 3835 12288 3847 12291
rect 6086 12288 6092 12300
rect 3835 12260 6092 12288
rect 3835 12257 3847 12260
rect 3789 12251 3847 12257
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 6270 12248 6276 12300
rect 6328 12248 6334 12300
rect 8312 12260 8800 12288
rect 8312 12232 8340 12260
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 2593 12183 2651 12189
rect 2866 12180 2872 12232
rect 2924 12180 2930 12232
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2976 12192 3065 12220
rect 2976 12164 3004 12192
rect 3053 12189 3065 12192
rect 3099 12189 3111 12223
rect 5810 12223 5868 12229
rect 5810 12220 5822 12223
rect 3053 12183 3111 12189
rect 5736 12192 5822 12220
rect 2958 12112 2964 12164
rect 3016 12112 3022 12164
rect 4062 12112 4068 12164
rect 4120 12112 4126 12164
rect 4706 12112 4712 12164
rect 4764 12112 4770 12164
rect 5736 12152 5764 12192
rect 5810 12189 5822 12192
rect 5856 12220 5868 12223
rect 6181 12223 6239 12229
rect 5856 12192 6132 12220
rect 5856 12189 5868 12192
rect 5810 12183 5868 12189
rect 5552 12124 5764 12152
rect 6104 12152 6132 12192
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6365 12223 6423 12229
rect 6227 12192 6316 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6288 12152 6316 12192
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6546 12220 6552 12232
rect 6411 12192 6552 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 6638 12180 6644 12232
rect 6696 12180 6702 12232
rect 7466 12220 7472 12232
rect 6886 12192 7472 12220
rect 6454 12152 6460 12164
rect 6104 12124 6224 12152
rect 6288 12124 6460 12152
rect 2222 12044 2228 12096
rect 2280 12084 2286 12096
rect 5552 12093 5580 12124
rect 6196 12096 6224 12124
rect 6454 12112 6460 12124
rect 6512 12112 6518 12164
rect 6564 12152 6592 12180
rect 6886 12152 6914 12192
rect 7466 12180 7472 12192
rect 7524 12220 7530 12232
rect 8294 12220 8300 12232
rect 7524 12192 8300 12220
rect 7524 12180 7530 12192
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 6564 12124 6914 12152
rect 7834 12112 7840 12164
rect 7892 12152 7898 12164
rect 8404 12152 8432 12183
rect 8478 12180 8484 12232
rect 8536 12180 8542 12232
rect 8570 12180 8576 12232
rect 8628 12180 8634 12232
rect 8772 12229 8800 12260
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10704 12288 10732 12328
rect 12066 12288 12072 12300
rect 9732 12260 9812 12288
rect 10704 12260 12072 12288
rect 9732 12248 9738 12260
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 7892 12124 9168 12152
rect 7892 12112 7898 12124
rect 9140 12096 9168 12124
rect 9232 12096 9260 12183
rect 9306 12180 9312 12232
rect 9364 12180 9370 12232
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12189 9643 12223
rect 9585 12183 9643 12189
rect 9600 12152 9628 12183
rect 9508 12124 9628 12152
rect 9677 12155 9735 12161
rect 2409 12087 2467 12093
rect 2409 12084 2421 12087
rect 2280 12056 2421 12084
rect 2280 12044 2286 12056
rect 2409 12053 2421 12056
rect 2455 12053 2467 12087
rect 2409 12047 2467 12053
rect 2777 12087 2835 12093
rect 2777 12053 2789 12087
rect 2823 12084 2835 12087
rect 3605 12087 3663 12093
rect 3605 12084 3617 12087
rect 2823 12056 3617 12084
rect 2823 12053 2835 12056
rect 2777 12047 2835 12053
rect 3605 12053 3617 12056
rect 3651 12053 3663 12087
rect 3605 12047 3663 12053
rect 5537 12087 5595 12093
rect 5537 12053 5549 12087
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 5626 12044 5632 12096
rect 5684 12044 5690 12096
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 5813 12087 5871 12093
rect 5813 12084 5825 12087
rect 5776 12056 5825 12084
rect 5776 12044 5782 12056
rect 5813 12053 5825 12056
rect 5859 12053 5871 12087
rect 5813 12047 5871 12053
rect 6178 12044 6184 12096
rect 6236 12044 6242 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 6822 12084 6828 12096
rect 6595 12056 6828 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 8113 12087 8171 12093
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 8662 12084 8668 12096
rect 8159 12056 8668 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 9030 12044 9036 12096
rect 9088 12044 9094 12096
rect 9122 12044 9128 12096
rect 9180 12044 9186 12096
rect 9214 12044 9220 12096
rect 9272 12044 9278 12096
rect 9508 12084 9536 12124
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 9784 12152 9812 12260
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12434 12248 12440 12300
rect 12492 12248 12498 12300
rect 12618 12248 12624 12300
rect 12676 12248 12682 12300
rect 13280 12297 13308 12396
rect 13354 12384 13360 12396
rect 13412 12424 13418 12436
rect 13412 12396 14596 12424
rect 13412 12384 13418 12396
rect 14568 12297 14596 12396
rect 15010 12384 15016 12436
rect 15068 12424 15074 12436
rect 15105 12427 15163 12433
rect 15105 12424 15117 12427
rect 15068 12396 15117 12424
rect 15068 12384 15074 12396
rect 15105 12393 15117 12396
rect 15151 12393 15163 12427
rect 15105 12387 15163 12393
rect 15396 12396 19288 12424
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 14553 12291 14611 12297
rect 14553 12257 14565 12291
rect 14599 12257 14611 12291
rect 14553 12251 14611 12257
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 15396 12288 15424 12396
rect 15473 12359 15531 12365
rect 15473 12325 15485 12359
rect 15519 12325 15531 12359
rect 15473 12319 15531 12325
rect 14783 12260 15424 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 10502 12180 10508 12232
rect 10560 12180 10566 12232
rect 10594 12180 10600 12232
rect 10652 12180 10658 12232
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 12952 12192 13185 12220
rect 12952 12180 12958 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 9723 12124 9812 12152
rect 12345 12155 12403 12161
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 12345 12121 12357 12155
rect 12391 12152 12403 12155
rect 13464 12152 13492 12251
rect 15013 12223 15071 12229
rect 15013 12189 15025 12223
rect 15059 12220 15071 12223
rect 15488 12220 15516 12319
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 18138 12356 18144 12368
rect 16448 12328 18144 12356
rect 16448 12316 16454 12328
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 19260 12356 19288 12396
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 19392 12396 19717 12424
rect 19392 12384 19398 12396
rect 19705 12393 19717 12396
rect 19751 12393 19763 12427
rect 22278 12424 22284 12436
rect 19705 12387 19763 12393
rect 20824 12396 22284 12424
rect 20824 12368 20852 12396
rect 22278 12384 22284 12396
rect 22336 12384 22342 12436
rect 23198 12384 23204 12436
rect 23256 12384 23262 12436
rect 27433 12427 27491 12433
rect 27433 12424 27445 12427
rect 24320 12396 27445 12424
rect 20806 12356 20812 12368
rect 19260 12328 20812 12356
rect 20806 12316 20812 12328
rect 20864 12316 20870 12368
rect 21450 12316 21456 12368
rect 21508 12356 21514 12368
rect 21729 12359 21787 12365
rect 21729 12356 21741 12359
rect 21508 12328 21741 12356
rect 21508 12316 21514 12328
rect 21729 12325 21741 12328
rect 21775 12325 21787 12359
rect 23216 12356 23244 12384
rect 23845 12359 23903 12365
rect 23845 12356 23857 12359
rect 23216 12328 23857 12356
rect 21729 12319 21787 12325
rect 23845 12325 23857 12328
rect 23891 12325 23903 12359
rect 23845 12319 23903 12325
rect 15930 12248 15936 12300
rect 15988 12248 15994 12300
rect 16114 12248 16120 12300
rect 16172 12248 16178 12300
rect 16224 12260 16436 12288
rect 16224 12220 16252 12260
rect 15059 12192 15516 12220
rect 15580 12192 16252 12220
rect 15059 12189 15071 12192
rect 15013 12183 15071 12189
rect 15580 12152 15608 12192
rect 16298 12180 16304 12232
rect 16356 12180 16362 12232
rect 16408 12220 16436 12260
rect 19610 12248 19616 12300
rect 19668 12288 19674 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 19668 12260 19809 12288
rect 19668 12248 19674 12260
rect 19797 12257 19809 12260
rect 19843 12288 19855 12291
rect 19978 12288 19984 12300
rect 19843 12260 19984 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 21634 12288 21640 12300
rect 21468 12260 21640 12288
rect 16408 12192 18736 12220
rect 12391 12124 12940 12152
rect 13464 12124 15608 12152
rect 15841 12155 15899 12161
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 9582 12084 9588 12096
rect 9508 12056 9588 12084
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 10376 12056 11989 12084
rect 10376 12044 10382 12056
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 11977 12047 12035 12053
rect 12802 12044 12808 12096
rect 12860 12044 12866 12096
rect 12912 12084 12940 12124
rect 15841 12121 15853 12155
rect 15887 12152 15899 12155
rect 16393 12155 16451 12161
rect 16393 12152 16405 12155
rect 15887 12124 16405 12152
rect 15887 12121 15899 12124
rect 15841 12115 15899 12121
rect 16393 12121 16405 12124
rect 16439 12121 16451 12155
rect 16393 12115 16451 12121
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 18708 12152 18736 12192
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 18932 12192 19533 12220
rect 18932 12180 18938 12192
rect 19521 12189 19533 12192
rect 19567 12220 19579 12223
rect 20162 12220 20168 12232
rect 19567 12192 20168 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 21174 12180 21180 12232
rect 21232 12180 21238 12232
rect 21468 12229 21496 12260
rect 21634 12248 21640 12260
rect 21692 12248 21698 12300
rect 22738 12288 22744 12300
rect 21744 12260 22744 12288
rect 21453 12223 21511 12229
rect 21453 12220 21465 12223
rect 21284 12192 21465 12220
rect 21284 12164 21312 12192
rect 21453 12189 21465 12192
rect 21499 12189 21511 12223
rect 21453 12183 21511 12189
rect 21542 12180 21548 12232
rect 21600 12180 21606 12232
rect 19150 12152 19156 12164
rect 16632 12124 18644 12152
rect 18708 12124 19156 12152
rect 16632 12112 16638 12124
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 12912 12056 14105 12084
rect 14093 12053 14105 12056
rect 14139 12053 14151 12087
rect 14093 12047 14151 12053
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14240 12056 14473 12084
rect 14240 12044 14246 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 15746 12084 15752 12096
rect 15528 12056 15752 12084
rect 15528 12044 15534 12056
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 18506 12084 18512 12096
rect 16356 12056 18512 12084
rect 16356 12044 16362 12056
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 18616 12084 18644 12124
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 19337 12155 19395 12161
rect 19337 12121 19349 12155
rect 19383 12152 19395 12155
rect 20990 12152 20996 12164
rect 19383 12124 20996 12152
rect 19383 12121 19395 12124
rect 19337 12115 19395 12121
rect 20990 12112 20996 12124
rect 21048 12112 21054 12164
rect 21266 12112 21272 12164
rect 21324 12112 21330 12164
rect 21358 12112 21364 12164
rect 21416 12112 21422 12164
rect 21744 12152 21772 12260
rect 22738 12248 22744 12260
rect 22796 12248 22802 12300
rect 23934 12248 23940 12300
rect 23992 12248 23998 12300
rect 21821 12223 21879 12229
rect 21821 12189 21833 12223
rect 21867 12189 21879 12223
rect 21821 12183 21879 12189
rect 21561 12124 21772 12152
rect 21836 12152 21864 12183
rect 22370 12180 22376 12232
rect 22428 12220 22434 12232
rect 23415 12223 23473 12229
rect 23415 12220 23427 12223
rect 22428 12192 23427 12220
rect 22428 12180 22434 12192
rect 23415 12189 23427 12192
rect 23461 12189 23473 12223
rect 24320 12220 24348 12396
rect 27433 12393 27445 12396
rect 27479 12393 27491 12427
rect 27433 12387 27491 12393
rect 28718 12384 28724 12436
rect 28776 12384 28782 12436
rect 28902 12384 28908 12436
rect 28960 12424 28966 12436
rect 30006 12424 30012 12436
rect 28960 12396 30012 12424
rect 28960 12384 28966 12396
rect 30006 12384 30012 12396
rect 30064 12384 30070 12436
rect 30282 12384 30288 12436
rect 30340 12424 30346 12436
rect 30340 12396 31524 12424
rect 30340 12384 30346 12396
rect 24673 12359 24731 12365
rect 24673 12325 24685 12359
rect 24719 12356 24731 12359
rect 24762 12356 24768 12368
rect 24719 12328 24768 12356
rect 24719 12325 24731 12328
rect 24673 12319 24731 12325
rect 24762 12316 24768 12328
rect 24820 12316 24826 12368
rect 25056 12328 26188 12356
rect 25056 12229 25084 12328
rect 26160 12288 26188 12328
rect 28736 12288 28764 12384
rect 29365 12359 29423 12365
rect 29365 12325 29377 12359
rect 29411 12356 29423 12359
rect 29411 12328 30880 12356
rect 29411 12325 29423 12328
rect 29365 12319 29423 12325
rect 28905 12291 28963 12297
rect 28905 12288 28917 12291
rect 26160 12260 27660 12288
rect 28736 12260 28917 12288
rect 26160 12232 26188 12260
rect 24489 12223 24547 12229
rect 24489 12220 24501 12223
rect 23415 12183 23473 12189
rect 23558 12192 24501 12220
rect 23558 12161 23586 12192
rect 24489 12189 24501 12192
rect 24535 12189 24547 12223
rect 24489 12183 24547 12189
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12189 25099 12223
rect 25041 12183 25099 12189
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 23543 12155 23601 12161
rect 21836 12124 23428 12152
rect 21561 12084 21589 12124
rect 18616 12056 21589 12084
rect 21818 12044 21824 12096
rect 21876 12084 21882 12096
rect 21913 12087 21971 12093
rect 21913 12084 21925 12087
rect 21876 12056 21925 12084
rect 21876 12044 21882 12056
rect 21913 12053 21925 12056
rect 21959 12053 21971 12087
rect 21913 12047 21971 12053
rect 22738 12044 22744 12096
rect 22796 12084 22802 12096
rect 23106 12084 23112 12096
rect 22796 12056 23112 12084
rect 22796 12044 22802 12056
rect 23106 12044 23112 12056
rect 23164 12084 23170 12096
rect 23293 12087 23351 12093
rect 23293 12084 23305 12087
rect 23164 12056 23305 12084
rect 23164 12044 23170 12056
rect 23293 12053 23305 12056
rect 23339 12053 23351 12087
rect 23400 12084 23428 12124
rect 23543 12121 23555 12155
rect 23589 12121 23601 12155
rect 23543 12115 23601 12121
rect 23658 12112 23664 12164
rect 23716 12152 23722 12164
rect 25056 12152 25084 12183
rect 23716 12124 25084 12152
rect 25240 12152 25268 12183
rect 25314 12180 25320 12232
rect 25372 12220 25378 12232
rect 25498 12220 25504 12232
rect 25372 12192 25504 12220
rect 25372 12180 25378 12192
rect 25498 12180 25504 12192
rect 25556 12180 25562 12232
rect 26142 12180 26148 12232
rect 26200 12180 26206 12232
rect 26620 12229 26648 12260
rect 26421 12223 26479 12229
rect 26421 12189 26433 12223
rect 26467 12189 26479 12223
rect 26421 12183 26479 12189
rect 26605 12223 26663 12229
rect 26605 12189 26617 12223
rect 26651 12189 26663 12223
rect 26605 12183 26663 12189
rect 26441 12152 26469 12183
rect 26970 12180 26976 12232
rect 27028 12180 27034 12232
rect 27062 12180 27068 12232
rect 27120 12180 27126 12232
rect 27246 12180 27252 12232
rect 27304 12180 27310 12232
rect 27338 12180 27344 12232
rect 27396 12180 27402 12232
rect 27632 12229 27660 12260
rect 28905 12257 28917 12260
rect 28951 12257 28963 12291
rect 28905 12251 28963 12257
rect 30190 12248 30196 12300
rect 30248 12248 30254 12300
rect 30282 12248 30288 12300
rect 30340 12248 30346 12300
rect 27433 12223 27491 12229
rect 27433 12189 27445 12223
rect 27479 12189 27491 12223
rect 27433 12183 27491 12189
rect 27617 12223 27675 12229
rect 27617 12189 27629 12223
rect 27663 12189 27675 12223
rect 27617 12183 27675 12189
rect 28721 12223 28779 12229
rect 28721 12189 28733 12223
rect 28767 12189 28779 12223
rect 28721 12183 28779 12189
rect 28997 12223 29055 12229
rect 28997 12189 29009 12223
rect 29043 12220 29055 12223
rect 29546 12220 29552 12232
rect 29043 12192 29552 12220
rect 29043 12189 29055 12192
rect 28997 12183 29055 12189
rect 26988 12152 27016 12180
rect 25240 12124 25360 12152
rect 26441 12124 27016 12152
rect 27264 12152 27292 12180
rect 27448 12152 27476 12183
rect 27264 12124 27476 12152
rect 28736 12152 28764 12183
rect 29546 12180 29552 12192
rect 29604 12180 29610 12232
rect 30561 12223 30619 12229
rect 30561 12189 30573 12223
rect 30607 12220 30619 12223
rect 30650 12220 30656 12232
rect 30607 12192 30656 12220
rect 30607 12189 30619 12192
rect 30561 12183 30619 12189
rect 30650 12180 30656 12192
rect 30708 12180 30714 12232
rect 30852 12220 30880 12328
rect 31294 12316 31300 12368
rect 31352 12316 31358 12368
rect 31496 12356 31524 12396
rect 31754 12384 31760 12436
rect 31812 12424 31818 12436
rect 31849 12427 31907 12433
rect 31849 12424 31861 12427
rect 31812 12396 31861 12424
rect 31812 12384 31818 12396
rect 31849 12393 31861 12396
rect 31895 12393 31907 12427
rect 31849 12387 31907 12393
rect 39485 12427 39543 12433
rect 39485 12393 39497 12427
rect 39531 12424 39543 12427
rect 39574 12424 39580 12436
rect 39531 12396 39580 12424
rect 39531 12393 39543 12396
rect 39485 12387 39543 12393
rect 39574 12384 39580 12396
rect 39632 12384 39638 12436
rect 33042 12356 33048 12368
rect 31496 12328 33048 12356
rect 33042 12316 33048 12328
rect 33100 12316 33106 12368
rect 31312 12288 31340 12316
rect 31312 12260 31524 12288
rect 30953 12223 31011 12229
rect 30953 12220 30965 12223
rect 30852 12192 30965 12220
rect 30953 12189 30965 12192
rect 30999 12189 31011 12223
rect 30953 12183 31011 12189
rect 31110 12180 31116 12232
rect 31168 12220 31174 12232
rect 31205 12223 31263 12229
rect 31205 12220 31217 12223
rect 31168 12192 31217 12220
rect 31168 12180 31174 12192
rect 31205 12189 31217 12192
rect 31251 12189 31263 12223
rect 31205 12183 31263 12189
rect 31386 12180 31392 12232
rect 31444 12180 31450 12232
rect 31496 12229 31524 12260
rect 31570 12248 31576 12300
rect 31628 12248 31634 12300
rect 33686 12288 33692 12300
rect 31680 12260 33692 12288
rect 31680 12232 31708 12260
rect 33686 12248 33692 12260
rect 33744 12248 33750 12300
rect 35710 12248 35716 12300
rect 35768 12288 35774 12300
rect 40497 12291 40555 12297
rect 40497 12288 40509 12291
rect 35768 12260 40509 12288
rect 35768 12248 35774 12260
rect 40497 12257 40509 12260
rect 40543 12257 40555 12291
rect 40497 12251 40555 12257
rect 40586 12248 40592 12300
rect 40644 12248 40650 12300
rect 31481 12223 31539 12229
rect 31481 12189 31493 12223
rect 31527 12189 31539 12223
rect 31481 12183 31539 12189
rect 31662 12180 31668 12232
rect 31720 12180 31726 12232
rect 31849 12223 31907 12229
rect 31849 12189 31861 12223
rect 31895 12189 31907 12223
rect 31849 12183 31907 12189
rect 30101 12155 30159 12161
rect 28736 12124 29776 12152
rect 23716 12112 23722 12124
rect 23676 12084 23704 12112
rect 23400 12056 23704 12084
rect 23293 12047 23351 12053
rect 24578 12044 24584 12096
rect 24636 12084 24642 12096
rect 24762 12084 24768 12096
rect 24636 12056 24768 12084
rect 24636 12044 24642 12056
rect 24762 12044 24768 12056
rect 24820 12084 24826 12096
rect 25332 12084 25360 12124
rect 24820 12056 25360 12084
rect 24820 12044 24826 12056
rect 26510 12044 26516 12096
rect 26568 12044 26574 12096
rect 26878 12044 26884 12096
rect 26936 12044 26942 12096
rect 28534 12044 28540 12096
rect 28592 12044 28598 12096
rect 29748 12093 29776 12124
rect 30101 12121 30113 12155
rect 30147 12152 30159 12155
rect 30147 12124 30604 12152
rect 30147 12121 30159 12124
rect 30101 12115 30159 12121
rect 29733 12087 29791 12093
rect 29733 12053 29745 12087
rect 29779 12053 29791 12087
rect 30576 12084 30604 12124
rect 30742 12112 30748 12164
rect 30800 12112 30806 12164
rect 30834 12112 30840 12164
rect 30892 12152 30898 12164
rect 31294 12152 31300 12164
rect 30892 12124 31300 12152
rect 30892 12112 30898 12124
rect 31294 12112 31300 12124
rect 31352 12112 31358 12164
rect 31864 12152 31892 12183
rect 32030 12180 32036 12232
rect 32088 12180 32094 12232
rect 32950 12180 32956 12232
rect 33008 12220 33014 12232
rect 34606 12220 34612 12232
rect 33008 12192 34612 12220
rect 33008 12180 33014 12192
rect 34606 12180 34612 12192
rect 34664 12180 34670 12232
rect 38654 12180 38660 12232
rect 38712 12180 38718 12232
rect 39669 12223 39727 12229
rect 39669 12189 39681 12223
rect 39715 12220 39727 12223
rect 40405 12223 40463 12229
rect 39715 12192 40080 12220
rect 39715 12189 39727 12192
rect 39669 12183 39727 12189
rect 32968 12152 32996 12180
rect 31864 12124 32996 12152
rect 31113 12087 31171 12093
rect 31113 12084 31125 12087
rect 30576 12056 31125 12084
rect 29733 12047 29791 12053
rect 31113 12053 31125 12056
rect 31159 12053 31171 12087
rect 31113 12047 31171 12053
rect 38470 12044 38476 12096
rect 38528 12044 38534 12096
rect 40052 12093 40080 12192
rect 40405 12189 40417 12223
rect 40451 12220 40463 12223
rect 41046 12220 41052 12232
rect 40451 12192 41052 12220
rect 40451 12189 40463 12192
rect 40405 12183 40463 12189
rect 41046 12180 41052 12192
rect 41104 12180 41110 12232
rect 40037 12087 40095 12093
rect 40037 12053 40049 12087
rect 40083 12053 40095 12087
rect 40037 12047 40095 12053
rect 1104 11994 41400 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 41400 11994
rect 1104 11920 41400 11942
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 4120 11852 4905 11880
rect 4120 11840 4126 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 5626 11880 5632 11892
rect 4893 11843 4951 11849
rect 5000 11852 5632 11880
rect 1949 11815 2007 11821
rect 1949 11781 1961 11815
rect 1995 11812 2007 11815
rect 2222 11812 2228 11824
rect 1995 11784 2228 11812
rect 1995 11781 2007 11784
rect 1949 11775 2007 11781
rect 2222 11772 2228 11784
rect 2280 11772 2286 11824
rect 3050 11704 3056 11756
rect 3108 11704 3114 11756
rect 3694 11704 3700 11756
rect 3752 11704 3758 11756
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 4663 11747 4721 11753
rect 4663 11713 4675 11747
rect 4709 11744 4721 11747
rect 4890 11744 4896 11756
rect 4709 11716 4896 11744
rect 4709 11713 4721 11716
rect 4663 11707 4721 11713
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 3712 11676 3740 11704
rect 1719 11648 3740 11676
rect 4540 11676 4568 11707
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 5000 11753 5028 11852
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6089 11883 6147 11889
rect 6089 11849 6101 11883
rect 6135 11880 6147 11883
rect 6270 11880 6276 11892
rect 6135 11852 6276 11880
rect 6135 11849 6147 11852
rect 6089 11843 6147 11849
rect 6270 11840 6276 11852
rect 6328 11880 6334 11892
rect 6733 11883 6791 11889
rect 6733 11880 6745 11883
rect 6328 11852 6745 11880
rect 6328 11840 6334 11852
rect 6733 11849 6745 11852
rect 6779 11880 6791 11883
rect 7837 11883 7895 11889
rect 7837 11880 7849 11883
rect 6779 11852 7849 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 7837 11849 7849 11852
rect 7883 11849 7895 11883
rect 7837 11843 7895 11849
rect 8205 11883 8263 11889
rect 8205 11849 8217 11883
rect 8251 11880 8263 11883
rect 8570 11880 8576 11892
rect 8251 11852 8576 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 5077 11815 5135 11821
rect 5077 11781 5089 11815
rect 5123 11781 5135 11815
rect 5077 11775 5135 11781
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11713 5043 11747
rect 5092 11744 5120 11775
rect 5166 11772 5172 11824
rect 5224 11812 5230 11824
rect 5277 11815 5335 11821
rect 5277 11812 5289 11815
rect 5224 11784 5289 11812
rect 5224 11772 5230 11784
rect 5277 11781 5289 11784
rect 5323 11781 5335 11815
rect 5277 11775 5335 11781
rect 5442 11772 5448 11824
rect 5500 11772 5506 11824
rect 5905 11815 5963 11821
rect 5905 11781 5917 11815
rect 5951 11812 5963 11815
rect 7852 11812 7880 11843
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 8754 11880 8760 11892
rect 8680 11852 8760 11880
rect 5951 11784 7788 11812
rect 7852 11784 8524 11812
rect 5951 11781 5963 11784
rect 5905 11775 5963 11781
rect 5460 11744 5488 11772
rect 6564 11753 6592 11784
rect 5092 11716 5488 11744
rect 6181 11747 6239 11753
rect 4985 11707 5043 11713
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6549 11747 6607 11753
rect 6227 11716 6500 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6472 11676 6500 11716
rect 6549 11713 6561 11747
rect 6595 11713 6607 11747
rect 6809 11747 6867 11753
rect 6809 11744 6821 11747
rect 6549 11707 6607 11713
rect 6656 11716 6821 11744
rect 6656 11676 6684 11716
rect 6809 11713 6821 11716
rect 6855 11713 6867 11747
rect 6809 11707 6867 11713
rect 7466 11704 7472 11756
rect 7524 11704 7530 11756
rect 7760 11744 7788 11784
rect 7834 11744 7840 11756
rect 7760 11716 7840 11744
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11713 8079 11747
rect 8021 11707 8079 11713
rect 4540 11648 4660 11676
rect 6472 11648 6776 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 4632 11620 4660 11648
rect 4614 11568 4620 11620
rect 4672 11568 4678 11620
rect 4801 11611 4859 11617
rect 4801 11577 4813 11611
rect 4847 11608 4859 11611
rect 5445 11611 5503 11617
rect 5445 11608 5457 11611
rect 4847 11580 5457 11608
rect 4847 11577 4859 11580
rect 4801 11571 4859 11577
rect 5445 11577 5457 11580
rect 5491 11577 5503 11611
rect 6638 11608 6644 11620
rect 5445 11571 5503 11577
rect 5920 11580 6644 11608
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 2958 11540 2964 11552
rect 1544 11512 2964 11540
rect 1544 11500 1550 11512
rect 2958 11500 2964 11512
rect 3016 11540 3022 11552
rect 3421 11543 3479 11549
rect 3421 11540 3433 11543
rect 3016 11512 3433 11540
rect 3016 11500 3022 11512
rect 3421 11509 3433 11512
rect 3467 11509 3479 11543
rect 3421 11503 3479 11509
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5920 11549 5948 11580
rect 6638 11568 6644 11580
rect 6696 11568 6702 11620
rect 6748 11608 6776 11648
rect 6822 11608 6828 11620
rect 6748 11580 6828 11608
rect 6822 11568 6828 11580
rect 6880 11568 6886 11620
rect 8036 11608 8064 11707
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 8496 11753 8524 11784
rect 8680 11753 8708 11852
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 9030 11840 9036 11892
rect 9088 11840 9094 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9493 11883 9551 11889
rect 9493 11880 9505 11883
rect 9180 11852 9505 11880
rect 9180 11840 9186 11852
rect 9493 11849 9505 11852
rect 9539 11849 9551 11883
rect 9493 11843 9551 11849
rect 10318 11840 10324 11892
rect 10376 11840 10382 11892
rect 12802 11880 12808 11892
rect 11900 11852 12808 11880
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11744 8815 11747
rect 9048 11744 9076 11840
rect 10336 11812 10364 11840
rect 11900 11821 11928 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 12894 11840 12900 11892
rect 12952 11880 12958 11892
rect 13357 11883 13415 11889
rect 13357 11880 13369 11883
rect 12952 11852 13369 11880
rect 12952 11840 12958 11852
rect 13357 11849 13369 11852
rect 13403 11849 13415 11883
rect 13357 11843 13415 11849
rect 11885 11815 11943 11821
rect 9600 11784 10364 11812
rect 10428 11784 11836 11812
rect 9600 11753 9628 11784
rect 10428 11753 10456 11784
rect 8803 11716 9076 11744
rect 9309 11747 9367 11753
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 9309 11713 9321 11747
rect 9355 11744 9367 11747
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9355 11716 9597 11744
rect 9355 11713 9367 11716
rect 9309 11707 9367 11713
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 8312 11676 8340 11704
rect 8680 11676 8708 11707
rect 8312 11648 8708 11676
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9784 11676 9812 11707
rect 10870 11704 10876 11756
rect 10928 11704 10934 11756
rect 9180 11648 9812 11676
rect 9180 11636 9186 11648
rect 9214 11608 9220 11620
rect 8036 11580 9220 11608
rect 9214 11568 9220 11580
rect 9272 11608 9278 11620
rect 9585 11611 9643 11617
rect 9585 11608 9597 11611
rect 9272 11580 9597 11608
rect 9272 11568 9278 11580
rect 9585 11577 9597 11580
rect 9631 11577 9643 11611
rect 9784 11608 9812 11648
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 10502 11676 10508 11688
rect 10275 11648 10508 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 10502 11636 10508 11648
rect 10560 11676 10566 11688
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10560 11648 10701 11676
rect 10560 11636 10566 11648
rect 10689 11645 10701 11648
rect 10735 11676 10747 11679
rect 11054 11676 11060 11688
rect 10735 11648 11060 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 9784 11580 10609 11608
rect 9585 11571 9643 11577
rect 10597 11577 10609 11580
rect 10643 11577 10655 11611
rect 11808 11608 11836 11784
rect 11885 11781 11897 11815
rect 11931 11781 11943 11815
rect 11885 11775 11943 11781
rect 12066 11772 12072 11824
rect 12124 11772 12130 11824
rect 13372 11812 13400 11843
rect 13446 11840 13452 11892
rect 13504 11840 13510 11892
rect 15378 11840 15384 11892
rect 15436 11840 15442 11892
rect 15749 11883 15807 11889
rect 15749 11849 15761 11883
rect 15795 11880 15807 11883
rect 16206 11880 16212 11892
rect 15795 11852 16212 11880
rect 15795 11849 15807 11852
rect 15749 11843 15807 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 17034 11840 17040 11892
rect 17092 11840 17098 11892
rect 17589 11883 17647 11889
rect 17589 11849 17601 11883
rect 17635 11880 17647 11883
rect 18325 11883 18383 11889
rect 18325 11880 18337 11883
rect 17635 11852 18337 11880
rect 17635 11849 17647 11852
rect 17589 11843 17647 11849
rect 18325 11849 18337 11852
rect 18371 11880 18383 11883
rect 18414 11880 18420 11892
rect 18371 11852 18420 11880
rect 18371 11849 18383 11852
rect 18325 11843 18383 11849
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 18506 11840 18512 11892
rect 18564 11880 18570 11892
rect 20346 11880 20352 11892
rect 18564 11852 20352 11880
rect 18564 11840 18570 11852
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 21174 11880 21180 11892
rect 20956 11852 21180 11880
rect 20956 11840 20962 11852
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 21910 11889 21916 11892
rect 21903 11883 21916 11889
rect 21903 11880 21915 11883
rect 21871 11852 21915 11880
rect 21903 11849 21915 11852
rect 21903 11843 21916 11849
rect 21910 11840 21916 11843
rect 21968 11840 21974 11892
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 22373 11883 22431 11889
rect 22373 11880 22385 11883
rect 22152 11852 22385 11880
rect 22152 11840 22158 11852
rect 22373 11849 22385 11852
rect 22419 11849 22431 11883
rect 22373 11843 22431 11849
rect 24210 11840 24216 11892
rect 24268 11880 24274 11892
rect 24268 11852 24808 11880
rect 24268 11840 24274 11852
rect 14182 11812 14188 11824
rect 13372 11784 14188 11812
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 15286 11772 15292 11824
rect 15344 11772 15350 11824
rect 15396 11812 15424 11840
rect 15396 11784 15608 11812
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 14734 11744 14740 11756
rect 13044 11716 14740 11744
rect 13044 11704 13050 11716
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 15194 11704 15200 11756
rect 15252 11704 15258 11756
rect 15304 11744 15332 11772
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 15304 11716 15393 11744
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15580 11753 15608 11784
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 16022 11744 16028 11756
rect 15611 11716 16028 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 17052 11744 17080 11840
rect 20254 11772 20260 11824
rect 20312 11812 20318 11824
rect 20625 11815 20683 11821
rect 20312 11784 20576 11812
rect 20312 11772 20318 11784
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 17052 11716 17141 11744
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 18138 11704 18144 11756
rect 18196 11744 18202 11756
rect 18785 11747 18843 11753
rect 18785 11744 18797 11747
rect 18196 11716 18797 11744
rect 18196 11704 18202 11716
rect 18785 11713 18797 11716
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11713 19119 11747
rect 19061 11707 19119 11713
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11676 12219 11679
rect 12618 11676 12624 11688
rect 12207 11648 12624 11676
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 13630 11636 13636 11688
rect 13688 11636 13694 11688
rect 15212 11676 15240 11704
rect 15212 11648 15608 11676
rect 15580 11620 15608 11648
rect 17218 11636 17224 11688
rect 17276 11676 17282 11688
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 17276 11648 18429 11676
rect 17276 11636 17282 11648
rect 18417 11645 18429 11648
rect 18463 11676 18475 11679
rect 18506 11676 18512 11688
rect 18463 11648 18512 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 18601 11679 18659 11685
rect 18601 11645 18613 11679
rect 18647 11645 18659 11679
rect 18601 11639 18659 11645
rect 15378 11608 15384 11620
rect 11808 11580 15384 11608
rect 10597 11571 10655 11577
rect 15378 11568 15384 11580
rect 15436 11608 15442 11620
rect 15436 11580 15516 11608
rect 15436 11568 15442 11580
rect 5261 11543 5319 11549
rect 5261 11540 5273 11543
rect 5132 11512 5273 11540
rect 5132 11500 5138 11512
rect 5261 11509 5273 11512
rect 5307 11540 5319 11543
rect 5905 11543 5963 11549
rect 5905 11540 5917 11543
rect 5307 11512 5917 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 5905 11509 5917 11512
rect 5951 11509 5963 11543
rect 5905 11503 5963 11509
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 6730 11540 6736 11552
rect 6420 11512 6736 11540
rect 6420 11500 6426 11512
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 7561 11543 7619 11549
rect 7561 11509 7573 11543
rect 7607 11540 7619 11543
rect 8202 11540 8208 11552
rect 7607 11512 8208 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 8996 11512 11069 11540
rect 8996 11500 9002 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 11057 11503 11115 11509
rect 11606 11500 11612 11552
rect 11664 11500 11670 11552
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 12989 11543 13047 11549
rect 12989 11540 13001 11543
rect 12584 11512 13001 11540
rect 12584 11500 12590 11512
rect 12989 11509 13001 11512
rect 13035 11509 13047 11543
rect 15488 11540 15516 11580
rect 15562 11568 15568 11620
rect 15620 11568 15626 11620
rect 16482 11568 16488 11620
rect 16540 11568 16546 11620
rect 17954 11568 17960 11620
rect 18012 11568 18018 11620
rect 18046 11568 18052 11620
rect 18104 11608 18110 11620
rect 18616 11608 18644 11639
rect 18874 11636 18880 11688
rect 18932 11636 18938 11688
rect 19076 11676 19104 11707
rect 20438 11704 20444 11756
rect 20496 11704 20502 11756
rect 20548 11744 20576 11784
rect 20625 11781 20637 11815
rect 20671 11812 20683 11815
rect 21266 11812 21272 11824
rect 20671 11784 21272 11812
rect 20671 11781 20683 11784
rect 20625 11775 20683 11781
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 21450 11772 21456 11824
rect 21508 11772 21514 11824
rect 21637 11815 21695 11821
rect 21637 11781 21649 11815
rect 21683 11812 21695 11815
rect 22002 11812 22008 11824
rect 21683 11784 22008 11812
rect 21683 11781 21695 11784
rect 21637 11775 21695 11781
rect 22002 11772 22008 11784
rect 22060 11812 22066 11824
rect 23474 11812 23480 11824
rect 22060 11784 23480 11812
rect 22060 11772 22066 11784
rect 23474 11772 23480 11784
rect 23532 11772 23538 11824
rect 24302 11812 24308 11824
rect 23768 11784 24308 11812
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20548 11716 20729 11744
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 20809 11747 20867 11753
rect 20809 11713 20821 11747
rect 20855 11744 20867 11747
rect 20898 11744 20904 11756
rect 20855 11716 20904 11744
rect 20855 11713 20867 11716
rect 20809 11707 20867 11713
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 21174 11704 21180 11756
rect 21232 11704 21238 11756
rect 21361 11747 21419 11753
rect 21361 11713 21373 11747
rect 21407 11744 21419 11747
rect 21468 11744 21496 11772
rect 21407 11716 21496 11744
rect 21545 11747 21603 11753
rect 21407 11713 21419 11716
rect 21361 11707 21419 11713
rect 21545 11713 21557 11747
rect 21591 11713 21603 11747
rect 22094 11744 22100 11756
rect 21545 11707 21603 11713
rect 21744 11716 22100 11744
rect 19076 11648 20760 11676
rect 18892 11608 18920 11636
rect 20732 11620 20760 11648
rect 21266 11636 21272 11688
rect 21324 11676 21330 11688
rect 21560 11676 21588 11707
rect 21744 11676 21772 11716
rect 22094 11704 22100 11716
rect 22152 11704 22158 11756
rect 23198 11704 23204 11756
rect 23256 11704 23262 11756
rect 23385 11747 23443 11753
rect 23385 11713 23397 11747
rect 23431 11713 23443 11747
rect 23385 11707 23443 11713
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11744 23627 11747
rect 23658 11744 23664 11756
rect 23615 11716 23664 11744
rect 23615 11713 23627 11716
rect 23569 11707 23627 11713
rect 21324 11648 21772 11676
rect 22281 11679 22339 11685
rect 21324 11636 21330 11648
rect 22281 11645 22293 11679
rect 22327 11645 22339 11679
rect 22281 11639 22339 11645
rect 22465 11679 22523 11685
rect 22465 11645 22477 11679
rect 22511 11676 22523 11679
rect 23216 11676 23244 11704
rect 22511 11648 23244 11676
rect 22511 11645 22523 11648
rect 22465 11639 22523 11645
rect 19886 11608 19892 11620
rect 18104 11580 18828 11608
rect 18892 11580 19892 11608
rect 18104 11568 18110 11580
rect 16500 11540 16528 11568
rect 15488 11512 16528 11540
rect 12989 11503 13047 11509
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 18800 11549 18828 11580
rect 19886 11568 19892 11580
rect 19944 11568 19950 11620
rect 20714 11568 20720 11620
rect 20772 11568 20778 11620
rect 20993 11611 21051 11617
rect 20993 11577 21005 11611
rect 21039 11608 21051 11611
rect 22296 11608 22324 11639
rect 21039 11580 22324 11608
rect 23400 11608 23428 11707
rect 23658 11704 23664 11716
rect 23716 11704 23722 11756
rect 23768 11753 23796 11784
rect 24302 11772 24308 11784
rect 24360 11772 24366 11824
rect 24780 11821 24808 11852
rect 25038 11840 25044 11892
rect 25096 11880 25102 11892
rect 25133 11883 25191 11889
rect 25133 11880 25145 11883
rect 25096 11852 25145 11880
rect 25096 11840 25102 11852
rect 25133 11849 25145 11852
rect 25179 11849 25191 11883
rect 25590 11880 25596 11892
rect 25133 11843 25191 11849
rect 25332 11852 25596 11880
rect 24765 11815 24823 11821
rect 24765 11781 24777 11815
rect 24811 11781 24823 11815
rect 24765 11775 24823 11781
rect 24854 11772 24860 11824
rect 24912 11772 24918 11824
rect 23753 11747 23811 11753
rect 23753 11713 23765 11747
rect 23799 11713 23811 11747
rect 23753 11707 23811 11713
rect 23842 11704 23848 11756
rect 23900 11744 23906 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23900 11716 23949 11744
rect 23900 11704 23906 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 24320 11744 24348 11772
rect 24489 11747 24547 11753
rect 24489 11744 24501 11747
rect 24320 11716 24501 11744
rect 23937 11707 23995 11713
rect 24489 11713 24501 11716
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 25041 11747 25099 11753
rect 25041 11713 25053 11747
rect 25087 11744 25099 11747
rect 25332 11744 25360 11852
rect 25590 11840 25596 11852
rect 25648 11880 25654 11892
rect 26510 11880 26516 11892
rect 25648 11852 26516 11880
rect 25648 11840 25654 11852
rect 26510 11840 26516 11852
rect 26568 11840 26574 11892
rect 26878 11840 26884 11892
rect 26936 11880 26942 11892
rect 28626 11880 28632 11892
rect 26936 11852 28212 11880
rect 26936 11840 26942 11852
rect 27341 11815 27399 11821
rect 27341 11812 27353 11815
rect 26068 11784 27353 11812
rect 25087 11716 25360 11744
rect 25409 11747 25467 11753
rect 25087 11713 25099 11716
rect 25041 11707 25099 11713
rect 25409 11713 25421 11747
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 25593 11747 25651 11753
rect 25593 11713 25605 11747
rect 25639 11744 25651 11747
rect 25682 11744 25688 11756
rect 25639 11716 25688 11744
rect 25639 11713 25651 11716
rect 25593 11707 25651 11713
rect 24397 11679 24455 11685
rect 24397 11645 24409 11679
rect 24443 11676 24455 11679
rect 24762 11676 24768 11688
rect 24443 11648 24768 11676
rect 24443 11645 24455 11648
rect 24397 11639 24455 11645
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 24486 11608 24492 11620
rect 23400 11580 24492 11608
rect 21039 11577 21051 11580
rect 20993 11571 21051 11577
rect 24486 11568 24492 11580
rect 24544 11568 24550 11620
rect 25424 11608 25452 11707
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 26068 11753 26096 11784
rect 27341 11781 27353 11784
rect 27387 11781 27399 11815
rect 27341 11775 27399 11781
rect 26053 11747 26111 11753
rect 26053 11713 26065 11747
rect 26099 11713 26111 11747
rect 26053 11707 26111 11713
rect 26146 11747 26204 11753
rect 26146 11713 26158 11747
rect 26192 11713 26204 11747
rect 26146 11707 26204 11713
rect 26160 11676 26188 11707
rect 26234 11704 26240 11756
rect 26292 11704 26298 11756
rect 26326 11704 26332 11756
rect 26384 11704 26390 11756
rect 26421 11747 26479 11753
rect 26421 11713 26433 11747
rect 26467 11713 26479 11747
rect 26421 11707 26479 11713
rect 26068 11648 26188 11676
rect 26252 11676 26280 11704
rect 26436 11676 26464 11707
rect 26510 11704 26516 11756
rect 26568 11753 26574 11756
rect 26568 11744 26576 11753
rect 26568 11716 26613 11744
rect 26568 11707 26576 11716
rect 26568 11704 26574 11707
rect 26970 11704 26976 11756
rect 27028 11704 27034 11756
rect 27062 11704 27068 11756
rect 27120 11704 27126 11756
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11744 27215 11747
rect 27203 11716 27384 11744
rect 27203 11713 27215 11716
rect 27157 11707 27215 11713
rect 26786 11676 26792 11688
rect 26252 11648 26792 11676
rect 26068 11620 26096 11648
rect 26786 11636 26792 11648
rect 26844 11636 26850 11688
rect 26050 11608 26056 11620
rect 25424 11580 26056 11608
rect 26050 11568 26056 11580
rect 26108 11568 26114 11620
rect 27080 11608 27108 11704
rect 27356 11688 27384 11716
rect 27338 11636 27344 11688
rect 27396 11636 27402 11688
rect 28184 11676 28212 11852
rect 28276 11852 28632 11880
rect 28276 11753 28304 11852
rect 28626 11840 28632 11852
rect 28684 11880 28690 11892
rect 29270 11880 29276 11892
rect 28684 11852 29276 11880
rect 28684 11840 28690 11852
rect 29270 11840 29276 11852
rect 29328 11840 29334 11892
rect 30006 11840 30012 11892
rect 30064 11880 30070 11892
rect 30064 11852 30420 11880
rect 30064 11840 30070 11852
rect 28534 11772 28540 11824
rect 28592 11772 28598 11824
rect 30190 11772 30196 11824
rect 30248 11812 30254 11824
rect 30285 11815 30343 11821
rect 30285 11812 30297 11815
rect 30248 11784 30297 11812
rect 30248 11772 30254 11784
rect 30285 11781 30297 11784
rect 30331 11781 30343 11815
rect 30392 11812 30420 11852
rect 30466 11840 30472 11892
rect 30524 11880 30530 11892
rect 36081 11883 36139 11889
rect 30524 11852 35940 11880
rect 30524 11840 30530 11852
rect 35710 11812 35716 11824
rect 30392 11784 35716 11812
rect 30285 11775 30343 11781
rect 35710 11772 35716 11784
rect 35768 11772 35774 11824
rect 28261 11747 28319 11753
rect 28261 11713 28273 11747
rect 28307 11713 28319 11747
rect 28261 11707 28319 11713
rect 29638 11704 29644 11756
rect 29696 11704 29702 11756
rect 35912 11753 35940 11852
rect 36081 11849 36093 11883
rect 36127 11880 36139 11883
rect 36817 11883 36875 11889
rect 36817 11880 36829 11883
rect 36127 11852 36829 11880
rect 36127 11849 36139 11852
rect 36081 11843 36139 11849
rect 36817 11849 36829 11852
rect 36863 11849 36875 11883
rect 36817 11843 36875 11849
rect 36357 11815 36415 11821
rect 36357 11812 36369 11815
rect 36096 11784 36369 11812
rect 36096 11756 36124 11784
rect 36357 11781 36369 11784
rect 36403 11781 36415 11815
rect 36357 11775 36415 11781
rect 36541 11815 36599 11821
rect 36541 11781 36553 11815
rect 36587 11812 36599 11815
rect 38378 11812 38384 11824
rect 36587 11784 36952 11812
rect 36587 11781 36599 11784
rect 36541 11775 36599 11781
rect 35621 11747 35679 11753
rect 35621 11713 35633 11747
rect 35667 11713 35679 11747
rect 35621 11707 35679 11713
rect 35805 11747 35863 11753
rect 35805 11713 35817 11747
rect 35851 11713 35863 11747
rect 35805 11707 35863 11713
rect 35897 11747 35955 11753
rect 35897 11713 35909 11747
rect 35943 11713 35955 11747
rect 35897 11707 35955 11713
rect 35526 11676 35532 11688
rect 28184 11648 35532 11676
rect 35526 11636 35532 11648
rect 35584 11676 35590 11688
rect 35636 11676 35664 11707
rect 35584 11648 35664 11676
rect 35584 11636 35590 11648
rect 26436 11580 27108 11608
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 17184 11512 17233 11540
rect 17184 11500 17190 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17221 11503 17279 11509
rect 18785 11543 18843 11549
rect 18785 11509 18797 11543
rect 18831 11509 18843 11543
rect 18785 11503 18843 11509
rect 19245 11543 19303 11549
rect 19245 11509 19257 11543
rect 19291 11540 19303 11543
rect 19610 11540 19616 11552
rect 19291 11512 19616 11540
rect 19291 11509 19303 11512
rect 19245 11503 19303 11509
rect 19610 11500 19616 11512
rect 19668 11500 19674 11552
rect 21358 11500 21364 11552
rect 21416 11540 21422 11552
rect 21818 11540 21824 11552
rect 21416 11512 21824 11540
rect 21416 11500 21422 11512
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 23198 11500 23204 11552
rect 23256 11540 23262 11552
rect 23385 11543 23443 11549
rect 23385 11540 23397 11543
rect 23256 11512 23397 11540
rect 23256 11500 23262 11512
rect 23385 11509 23397 11512
rect 23431 11509 23443 11543
rect 23385 11503 23443 11509
rect 23750 11500 23756 11552
rect 23808 11500 23814 11552
rect 24213 11543 24271 11549
rect 24213 11509 24225 11543
rect 24259 11540 24271 11543
rect 26436 11540 26464 11580
rect 33594 11568 33600 11620
rect 33652 11608 33658 11620
rect 35820 11608 35848 11707
rect 35912 11676 35940 11707
rect 36078 11704 36084 11756
rect 36136 11704 36142 11756
rect 36924 11753 36952 11784
rect 38120 11784 38384 11812
rect 38120 11753 38148 11784
rect 38378 11772 38384 11784
rect 38436 11772 38442 11824
rect 38838 11772 38844 11824
rect 38896 11772 38902 11824
rect 36173 11747 36231 11753
rect 36173 11713 36185 11747
rect 36219 11713 36231 11747
rect 36173 11707 36231 11713
rect 36633 11747 36691 11753
rect 36633 11713 36645 11747
rect 36679 11713 36691 11747
rect 36633 11707 36691 11713
rect 36909 11747 36967 11753
rect 36909 11713 36921 11747
rect 36955 11713 36967 11747
rect 36909 11707 36967 11713
rect 38105 11747 38163 11753
rect 38105 11713 38117 11747
rect 38151 11713 38163 11747
rect 38105 11707 38163 11713
rect 36188 11676 36216 11707
rect 35912 11648 36216 11676
rect 36648 11676 36676 11707
rect 37550 11676 37556 11688
rect 36648 11648 37556 11676
rect 33652 11580 35848 11608
rect 36188 11608 36216 11648
rect 37550 11636 37556 11648
rect 37608 11636 37614 11688
rect 38381 11679 38439 11685
rect 38381 11645 38393 11679
rect 38427 11676 38439 11679
rect 38470 11676 38476 11688
rect 38427 11648 38476 11676
rect 38427 11645 38439 11648
rect 38381 11639 38439 11645
rect 38470 11636 38476 11648
rect 38528 11636 38534 11688
rect 37458 11608 37464 11620
rect 36188 11580 37464 11608
rect 33652 11568 33658 11580
rect 24259 11512 26464 11540
rect 26697 11543 26755 11549
rect 24259 11509 24271 11512
rect 24213 11503 24271 11509
rect 26697 11509 26709 11543
rect 26743 11540 26755 11543
rect 26878 11540 26884 11552
rect 26743 11512 26884 11540
rect 26743 11509 26755 11512
rect 26697 11503 26755 11509
rect 26878 11500 26884 11512
rect 26936 11540 26942 11552
rect 30466 11540 30472 11552
rect 26936 11512 30472 11540
rect 26936 11500 26942 11512
rect 30466 11500 30472 11512
rect 30524 11500 30530 11552
rect 35710 11500 35716 11552
rect 35768 11500 35774 11552
rect 35820 11540 35848 11580
rect 37458 11568 37464 11580
rect 37516 11568 37522 11620
rect 35986 11540 35992 11552
rect 35820 11512 35992 11540
rect 35986 11500 35992 11512
rect 36044 11540 36050 11552
rect 36538 11540 36544 11552
rect 36044 11512 36544 11540
rect 36044 11500 36050 11512
rect 36538 11500 36544 11512
rect 36596 11500 36602 11552
rect 36633 11543 36691 11549
rect 36633 11509 36645 11543
rect 36679 11540 36691 11543
rect 36722 11540 36728 11552
rect 36679 11512 36728 11540
rect 36679 11509 36691 11512
rect 36633 11503 36691 11509
rect 36722 11500 36728 11512
rect 36780 11500 36786 11552
rect 39850 11500 39856 11552
rect 39908 11500 39914 11552
rect 1104 11450 41400 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 41400 11450
rect 1104 11376 41400 11398
rect 934 11296 940 11348
rect 992 11336 998 11348
rect 1581 11339 1639 11345
rect 1581 11336 1593 11339
rect 992 11308 1593 11336
rect 992 11296 998 11308
rect 1581 11305 1593 11308
rect 1627 11305 1639 11339
rect 1581 11299 1639 11305
rect 3050 11296 3056 11348
rect 3108 11296 3114 11348
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 4672 11308 5733 11336
rect 4672 11296 4678 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 5721 11299 5779 11305
rect 5828 11308 6914 11336
rect 3068 11268 3096 11296
rect 5828 11268 5856 11308
rect 3068 11240 5856 11268
rect 6886 11268 6914 11308
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9398 11336 9404 11348
rect 9088 11308 9404 11336
rect 9088 11296 9094 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 10928 11308 13492 11336
rect 10928 11296 10934 11308
rect 11698 11268 11704 11280
rect 6886 11240 11704 11268
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 12066 11228 12072 11280
rect 12124 11228 12130 11280
rect 12526 11268 12532 11280
rect 12452 11240 12532 11268
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 5224 11172 5764 11200
rect 5224 11160 5230 11172
rect 1486 11092 1492 11144
rect 1544 11092 1550 11144
rect 5626 11092 5632 11144
rect 5684 11092 5690 11144
rect 5736 11141 5764 11172
rect 8386 11160 8392 11212
rect 8444 11200 8450 11212
rect 9214 11200 9220 11212
rect 8444 11172 9220 11200
rect 8444 11160 8450 11172
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 12452 11209 12480 11240
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11132 5871 11135
rect 6362 11132 6368 11144
rect 5859 11104 6368 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 5644 11064 5672 11092
rect 5828 11064 5856 11095
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 9950 11064 9956 11076
rect 2924 11036 5580 11064
rect 5644 11036 5856 11064
rect 5920 11036 9956 11064
rect 2924 11024 2930 11036
rect 5552 10996 5580 11036
rect 5920 10996 5948 11036
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 12526 11024 12532 11076
rect 12584 11064 12590 11076
rect 13262 11064 13268 11076
rect 12584 11036 13268 11064
rect 12584 11024 12590 11036
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 13464 11064 13492 11308
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 16669 11339 16727 11345
rect 13596 11308 14504 11336
rect 13596 11296 13602 11308
rect 14093 11271 14151 11277
rect 14093 11237 14105 11271
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 14108 11200 14136 11231
rect 14476 11212 14504 11308
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 17034 11336 17040 11348
rect 16715 11308 17040 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 18230 11296 18236 11348
rect 18288 11336 18294 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 18288 11308 18429 11336
rect 18288 11296 18294 11308
rect 18417 11305 18429 11308
rect 18463 11336 18475 11339
rect 18874 11336 18880 11348
rect 18463 11308 18880 11336
rect 18463 11305 18475 11308
rect 18417 11299 18475 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 19426 11296 19432 11348
rect 19484 11296 19490 11348
rect 19797 11339 19855 11345
rect 19797 11336 19809 11339
rect 19536 11308 19809 11336
rect 18046 11228 18052 11280
rect 18104 11268 18110 11280
rect 19536 11268 19564 11308
rect 19797 11305 19809 11308
rect 19843 11305 19855 11339
rect 19797 11299 19855 11305
rect 20806 11296 20812 11348
rect 20864 11296 20870 11348
rect 21634 11296 21640 11348
rect 21692 11336 21698 11348
rect 22370 11336 22376 11348
rect 21692 11308 22376 11336
rect 21692 11296 21698 11308
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 25041 11339 25099 11345
rect 23348 11308 24808 11336
rect 23348 11296 23354 11308
rect 20257 11271 20315 11277
rect 20257 11268 20269 11271
rect 18104 11240 19564 11268
rect 19812 11240 20269 11268
rect 18104 11228 18110 11240
rect 13924 11172 14136 11200
rect 13924 11141 13952 11172
rect 14458 11160 14464 11212
rect 14516 11200 14522 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 14516 11172 14657 11200
rect 14516 11160 14522 11172
rect 14645 11169 14657 11172
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 15068 11172 15301 11200
rect 15068 11160 15074 11172
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 18064 11200 18092 11228
rect 15289 11163 15347 11169
rect 16500 11172 18092 11200
rect 13909 11135 13967 11141
rect 13909 11101 13921 11135
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 14148 11104 16436 11132
rect 14148 11092 14154 11104
rect 14553 11067 14611 11073
rect 14553 11064 14565 11067
rect 13464 11036 14565 11064
rect 14553 11033 14565 11036
rect 14599 11064 14611 11067
rect 14599 11036 14688 11064
rect 14599 11033 14611 11036
rect 14553 11027 14611 11033
rect 5552 10968 5948 10996
rect 6086 10956 6092 11008
rect 6144 10956 6150 11008
rect 6178 10956 6184 11008
rect 6236 10996 6242 11008
rect 9398 10996 9404 11008
rect 6236 10968 9404 10996
rect 6236 10956 6242 10968
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 9582 10956 9588 11008
rect 9640 10996 9646 11008
rect 11882 10996 11888 11008
rect 9640 10968 11888 10996
rect 9640 10956 9646 10968
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 13722 10956 13728 11008
rect 13780 10956 13786 11008
rect 14458 10956 14464 11008
rect 14516 10956 14522 11008
rect 14660 10996 14688 11036
rect 14734 11024 14740 11076
rect 14792 11064 14798 11076
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 14792 11036 15025 11064
rect 14792 11024 14798 11036
rect 15013 11033 15025 11036
rect 15059 11033 15071 11067
rect 15930 11064 15936 11076
rect 15013 11027 15071 11033
rect 15120 11036 15936 11064
rect 15120 10996 15148 11036
rect 15930 11024 15936 11036
rect 15988 11064 15994 11076
rect 16298 11064 16304 11076
rect 15988 11036 16304 11064
rect 15988 11024 15994 11036
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 14660 10968 15148 10996
rect 16408 10996 16436 11104
rect 16500 11073 16528 11172
rect 18782 11160 18788 11212
rect 18840 11200 18846 11212
rect 18840 11172 19012 11200
rect 18840 11160 18846 11172
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 16592 11104 17785 11132
rect 16485 11067 16543 11073
rect 16485 11033 16497 11067
rect 16531 11033 16543 11067
rect 16485 11027 16543 11033
rect 16592 10996 16620 11104
rect 17773 11101 17785 11104
rect 17819 11132 17831 11135
rect 17954 11132 17960 11144
rect 17819 11104 17960 11132
rect 17819 11101 17831 11104
rect 17773 11095 17831 11101
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18138 11092 18144 11144
rect 18196 11132 18202 11144
rect 18196 11104 18460 11132
rect 18196 11092 18202 11104
rect 16669 11067 16727 11073
rect 16669 11033 16681 11067
rect 16715 11064 16727 11067
rect 16715 11036 16988 11064
rect 16715 11033 16727 11036
rect 16669 11027 16727 11033
rect 16408 10968 16620 10996
rect 16850 10956 16856 11008
rect 16908 10956 16914 11008
rect 16960 10996 16988 11036
rect 17034 11024 17040 11076
rect 17092 11064 17098 11076
rect 18322 11064 18328 11076
rect 17092 11036 18328 11064
rect 17092 11024 17098 11036
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 18432 11073 18460 11104
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 18984 11132 19012 11172
rect 19058 11160 19064 11212
rect 19116 11200 19122 11212
rect 19116 11172 19380 11200
rect 19116 11160 19122 11172
rect 19352 11141 19380 11172
rect 19610 11160 19616 11212
rect 19668 11160 19674 11212
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18564 11104 18920 11132
rect 18984 11104 19257 11132
rect 18564 11092 18570 11104
rect 18417 11067 18475 11073
rect 18417 11033 18429 11067
rect 18463 11064 18475 11067
rect 18782 11064 18788 11076
rect 18463 11036 18788 11064
rect 18463 11033 18475 11036
rect 18417 11027 18475 11033
rect 18782 11024 18788 11036
rect 18840 11024 18846 11076
rect 17218 10996 17224 11008
rect 16960 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 18598 10956 18604 11008
rect 18656 10956 18662 11008
rect 18892 10996 18920 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19337 11135 19395 11141
rect 19337 11101 19349 11135
rect 19383 11132 19395 11135
rect 19426 11132 19432 11144
rect 19383 11104 19432 11132
rect 19383 11101 19395 11104
rect 19337 11095 19395 11101
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11132 19579 11135
rect 19812 11132 19840 11240
rect 20257 11237 20269 11240
rect 20303 11237 20315 11271
rect 20257 11231 20315 11237
rect 22830 11228 22836 11280
rect 22888 11228 22894 11280
rect 19886 11160 19892 11212
rect 19944 11160 19950 11212
rect 21358 11160 21364 11212
rect 21416 11160 21422 11212
rect 21450 11160 21456 11212
rect 21508 11200 21514 11212
rect 22925 11203 22983 11209
rect 21508 11172 21956 11200
rect 21508 11160 21514 11172
rect 19567 11104 19840 11132
rect 19567 11101 19579 11104
rect 19521 11095 19579 11101
rect 20070 11092 20076 11144
rect 20128 11092 20134 11144
rect 21542 11092 21548 11144
rect 21600 11092 21606 11144
rect 21634 11092 21640 11144
rect 21692 11092 21698 11144
rect 21821 11135 21879 11141
rect 21821 11101 21833 11135
rect 21867 11101 21879 11135
rect 21821 11095 21879 11101
rect 19797 11067 19855 11073
rect 19797 11064 19809 11067
rect 19444 11036 19809 11064
rect 19444 10996 19472 11036
rect 19797 11033 19809 11036
rect 19843 11033 19855 11067
rect 19797 11027 19855 11033
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 20806 11064 20812 11076
rect 20220 11036 20812 11064
rect 20220 11024 20226 11036
rect 20806 11024 20812 11036
rect 20864 11024 20870 11076
rect 20898 11024 20904 11076
rect 20956 11064 20962 11076
rect 21085 11067 21143 11073
rect 21085 11064 21097 11067
rect 20956 11036 21097 11064
rect 20956 11024 20962 11036
rect 21085 11033 21097 11036
rect 21131 11033 21143 11067
rect 21085 11027 21143 11033
rect 21266 11024 21272 11076
rect 21324 11024 21330 11076
rect 21560 11064 21588 11092
rect 21836 11064 21864 11095
rect 21928 11073 21956 11172
rect 22925 11169 22937 11203
rect 22971 11200 22983 11203
rect 23308 11200 23336 11296
rect 24670 11228 24676 11280
rect 24728 11228 24734 11280
rect 24780 11268 24808 11308
rect 25041 11305 25053 11339
rect 25087 11336 25099 11339
rect 32490 11336 32496 11348
rect 25087 11308 32496 11336
rect 25087 11305 25099 11308
rect 25041 11299 25099 11305
rect 32490 11296 32496 11308
rect 32548 11296 32554 11348
rect 33229 11339 33287 11345
rect 33229 11336 33241 11339
rect 32692 11308 33241 11336
rect 25869 11271 25927 11277
rect 25869 11268 25881 11271
rect 24780 11240 25881 11268
rect 25869 11237 25881 11240
rect 25915 11237 25927 11271
rect 25869 11231 25927 11237
rect 22971 11172 23336 11200
rect 22971 11169 22983 11172
rect 22925 11163 22983 11169
rect 23750 11160 23756 11212
rect 23808 11200 23814 11212
rect 23808 11172 24164 11200
rect 23808 11160 23814 11172
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 22463 11135 22521 11141
rect 22463 11101 22475 11135
rect 22509 11132 22521 11135
rect 23198 11132 23204 11144
rect 22509 11104 23204 11132
rect 22509 11101 22521 11104
rect 22463 11095 22521 11101
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 23474 11092 23480 11144
rect 23532 11092 23538 11144
rect 23658 11092 23664 11144
rect 23716 11092 23722 11144
rect 23842 11092 23848 11144
rect 23900 11092 23906 11144
rect 24136 11132 24164 11172
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 24136 11104 24409 11132
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24486 11092 24492 11144
rect 24544 11132 24550 11144
rect 24688 11132 24716 11228
rect 25590 11160 25596 11212
rect 25648 11200 25654 11212
rect 25884 11200 25912 11231
rect 25958 11228 25964 11280
rect 26016 11268 26022 11280
rect 26142 11268 26148 11280
rect 26016 11240 26148 11268
rect 26016 11228 26022 11240
rect 26142 11228 26148 11240
rect 26200 11228 26206 11280
rect 26510 11228 26516 11280
rect 26568 11268 26574 11280
rect 27525 11271 27583 11277
rect 26568 11240 27389 11268
rect 26568 11228 26574 11240
rect 26697 11203 26755 11209
rect 26697 11200 26709 11203
rect 25648 11172 25820 11200
rect 25884 11172 26709 11200
rect 25648 11160 25654 11172
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 24544 11104 24589 11132
rect 24688 11104 24777 11132
rect 24544 11092 24550 11104
rect 24765 11101 24777 11104
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 24854 11092 24860 11144
rect 24912 11141 24918 11144
rect 24912 11132 24920 11141
rect 25499 11135 25557 11141
rect 24912 11104 24957 11132
rect 24912 11095 24920 11104
rect 25499 11101 25511 11135
rect 25545 11132 25557 11135
rect 25682 11132 25688 11144
rect 25545 11104 25688 11132
rect 25545 11101 25557 11104
rect 25499 11095 25557 11101
rect 24912 11092 24918 11095
rect 25682 11092 25688 11104
rect 25740 11092 25746 11144
rect 21560 11036 21864 11064
rect 21913 11067 21971 11073
rect 21913 11033 21925 11067
rect 21959 11064 21971 11067
rect 22204 11064 22232 11092
rect 22646 11064 22652 11076
rect 21959 11036 22232 11064
rect 22296 11036 22652 11064
rect 21959 11033 21971 11036
rect 21913 11027 21971 11033
rect 22296 11005 22324 11036
rect 22646 11024 22652 11036
rect 22704 11024 22710 11076
rect 23492 11064 23520 11092
rect 24578 11064 24584 11076
rect 23492 11036 24584 11064
rect 24578 11024 24584 11036
rect 24636 11064 24642 11076
rect 24673 11067 24731 11073
rect 24673 11064 24685 11067
rect 24636 11036 24685 11064
rect 24636 11024 24642 11036
rect 24673 11033 24685 11036
rect 24719 11033 24731 11067
rect 24673 11027 24731 11033
rect 18892 10968 19472 10996
rect 22281 10999 22339 11005
rect 22281 10965 22293 10999
rect 22327 10965 22339 10999
rect 22281 10959 22339 10965
rect 22370 10956 22376 11008
rect 22428 10996 22434 11008
rect 22465 10999 22523 11005
rect 22465 10996 22477 10999
rect 22428 10968 22477 10996
rect 22428 10956 22434 10968
rect 22465 10965 22477 10968
rect 22511 10965 22523 10999
rect 22465 10959 22523 10965
rect 23109 10999 23167 11005
rect 23109 10965 23121 10999
rect 23155 10996 23167 10999
rect 23198 10996 23204 11008
rect 23155 10968 23204 10996
rect 23155 10965 23167 10968
rect 23109 10959 23167 10965
rect 23198 10956 23204 10968
rect 23256 10956 23262 11008
rect 25038 10956 25044 11008
rect 25096 10996 25102 11008
rect 25317 10999 25375 11005
rect 25317 10996 25329 10999
rect 25096 10968 25329 10996
rect 25096 10956 25102 10968
rect 25317 10965 25329 10968
rect 25363 10965 25375 10999
rect 25317 10959 25375 10965
rect 25501 10999 25559 11005
rect 25501 10965 25513 10999
rect 25547 10996 25559 10999
rect 25792 10996 25820 11172
rect 26697 11169 26709 11172
rect 26743 11169 26755 11203
rect 26697 11163 26755 11169
rect 25958 11092 25964 11144
rect 26016 11092 26022 11144
rect 26510 11092 26516 11144
rect 26568 11132 26574 11144
rect 26568 11104 26832 11132
rect 26568 11092 26574 11104
rect 26234 11024 26240 11076
rect 26292 11064 26298 11076
rect 26421 11067 26479 11073
rect 26421 11064 26433 11067
rect 26292 11036 26433 11064
rect 26292 11024 26298 11036
rect 26421 11033 26433 11036
rect 26467 11033 26479 11067
rect 26421 11027 26479 11033
rect 26605 11067 26663 11073
rect 26605 11033 26617 11067
rect 26651 11064 26663 11067
rect 26694 11064 26700 11076
rect 26651 11036 26700 11064
rect 26651 11033 26663 11036
rect 26605 11027 26663 11033
rect 26694 11024 26700 11036
rect 26752 11024 26758 11076
rect 26804 11064 26832 11104
rect 26878 11092 26884 11144
rect 26936 11092 26942 11144
rect 26970 11092 26976 11144
rect 27028 11092 27034 11144
rect 27361 11141 27389 11240
rect 27525 11237 27537 11271
rect 27571 11268 27583 11271
rect 32582 11268 32588 11280
rect 27571 11240 32588 11268
rect 27571 11237 27583 11240
rect 27525 11231 27583 11237
rect 32582 11228 32588 11240
rect 32640 11228 32646 11280
rect 32122 11160 32128 11212
rect 32180 11200 32186 11212
rect 32692 11200 32720 11308
rect 33229 11305 33241 11308
rect 33275 11305 33287 11339
rect 33229 11299 33287 11305
rect 35710 11296 35716 11348
rect 35768 11336 35774 11348
rect 36633 11339 36691 11345
rect 36633 11336 36645 11339
rect 35768 11308 36645 11336
rect 35768 11296 35774 11308
rect 36633 11305 36645 11308
rect 36679 11305 36691 11339
rect 36633 11299 36691 11305
rect 38289 11339 38347 11345
rect 38289 11305 38301 11339
rect 38335 11336 38347 11339
rect 38654 11336 38660 11348
rect 38335 11308 38660 11336
rect 38335 11305 38347 11308
rect 38289 11299 38347 11305
rect 38654 11296 38660 11308
rect 38712 11296 38718 11348
rect 39850 11268 39856 11280
rect 32784 11240 39856 11268
rect 32784 11212 32812 11240
rect 32180 11172 32720 11200
rect 32180 11160 32186 11172
rect 32766 11160 32772 11212
rect 32824 11160 32830 11212
rect 33045 11203 33103 11209
rect 33045 11169 33057 11203
rect 33091 11200 33103 11203
rect 33502 11200 33508 11212
rect 33091 11172 33508 11200
rect 33091 11169 33103 11172
rect 33045 11163 33103 11169
rect 33502 11160 33508 11172
rect 33560 11160 33566 11212
rect 34790 11160 34796 11212
rect 34848 11160 34854 11212
rect 35986 11160 35992 11212
rect 36044 11200 36050 11212
rect 36722 11200 36728 11212
rect 36044 11172 36216 11200
rect 36044 11160 36050 11172
rect 27346 11135 27404 11141
rect 27346 11101 27358 11135
rect 27392 11101 27404 11135
rect 27346 11095 27404 11101
rect 32674 11092 32680 11144
rect 32732 11132 32738 11144
rect 32953 11135 33011 11141
rect 32953 11132 32965 11135
rect 32732 11104 32965 11132
rect 32732 11092 32738 11104
rect 32953 11101 32965 11104
rect 32999 11101 33011 11135
rect 32953 11095 33011 11101
rect 34931 11135 34989 11141
rect 34931 11101 34943 11135
rect 34977 11132 34989 11135
rect 36078 11132 36084 11144
rect 34977 11104 36084 11132
rect 34977 11101 34989 11104
rect 34931 11095 34989 11101
rect 27157 11067 27215 11073
rect 27157 11064 27169 11067
rect 26804 11036 27169 11064
rect 27157 11033 27169 11036
rect 27203 11033 27215 11067
rect 27157 11027 27215 11033
rect 27249 11067 27307 11073
rect 27249 11033 27261 11067
rect 27295 11033 27307 11067
rect 27249 11027 27307 11033
rect 25547 10968 25820 10996
rect 25547 10965 25559 10968
rect 25501 10959 25559 10965
rect 25866 10956 25872 11008
rect 25924 10996 25930 11008
rect 27264 10996 27292 11027
rect 25924 10968 27292 10996
rect 25924 10956 25930 10968
rect 30650 10956 30656 11008
rect 30708 10996 30714 11008
rect 33410 10996 33416 11008
rect 30708 10968 33416 10996
rect 30708 10956 30714 10968
rect 33410 10956 33416 10968
rect 33468 10996 33474 11008
rect 34956 10996 34984 11095
rect 36078 11092 36084 11104
rect 36136 11092 36142 11144
rect 36188 11141 36216 11172
rect 36280 11172 36728 11200
rect 36173 11135 36231 11141
rect 36173 11101 36185 11135
rect 36219 11101 36231 11135
rect 36173 11095 36231 11101
rect 35526 11024 35532 11076
rect 35584 11064 35590 11076
rect 35989 11067 36047 11073
rect 35989 11064 36001 11067
rect 35584 11036 36001 11064
rect 35584 11024 35590 11036
rect 35989 11033 36001 11036
rect 36035 11064 36047 11067
rect 36280 11064 36308 11172
rect 36722 11160 36728 11172
rect 36780 11200 36786 11212
rect 37461 11203 37519 11209
rect 37461 11200 37473 11203
rect 36780 11172 37473 11200
rect 36780 11160 36786 11172
rect 37461 11169 37473 11172
rect 37507 11169 37519 11203
rect 37461 11163 37519 11169
rect 37921 11203 37979 11209
rect 37921 11169 37933 11203
rect 37967 11200 37979 11203
rect 38746 11200 38752 11212
rect 37967 11172 38752 11200
rect 37967 11169 37979 11172
rect 37921 11163 37979 11169
rect 38746 11160 38752 11172
rect 38804 11160 38810 11212
rect 36357 11135 36415 11141
rect 36357 11101 36369 11135
rect 36403 11132 36415 11135
rect 37553 11135 37611 11141
rect 36403 11104 36584 11132
rect 36403 11101 36415 11104
rect 36357 11095 36415 11101
rect 36449 11067 36507 11073
rect 36449 11064 36461 11067
rect 36035 11036 36216 11064
rect 36280 11036 36461 11064
rect 36035 11033 36047 11036
rect 35989 11027 36047 11033
rect 33468 10968 34984 10996
rect 33468 10956 33474 10968
rect 35250 10956 35256 11008
rect 35308 10956 35314 11008
rect 36188 10996 36216 11036
rect 36449 11033 36461 11036
rect 36495 11033 36507 11067
rect 36556 11064 36584 11104
rect 37553 11101 37565 11135
rect 37599 11132 37611 11135
rect 38010 11132 38016 11144
rect 37599 11104 38016 11132
rect 37599 11101 37611 11104
rect 37553 11095 37611 11101
rect 36649 11067 36707 11073
rect 36649 11064 36661 11067
rect 36556 11036 36661 11064
rect 36449 11027 36507 11033
rect 36649 11033 36661 11036
rect 36695 11033 36707 11067
rect 37568 11064 37596 11095
rect 38010 11092 38016 11104
rect 38068 11092 38074 11144
rect 36649 11027 36707 11033
rect 36740 11036 37596 11064
rect 38749 11067 38807 11073
rect 36740 10996 36768 11036
rect 38749 11033 38761 11067
rect 38795 11064 38807 11067
rect 38856 11064 38884 11240
rect 39850 11228 39856 11240
rect 39908 11228 39914 11280
rect 38933 11203 38991 11209
rect 38933 11169 38945 11203
rect 38979 11200 38991 11203
rect 39666 11200 39672 11212
rect 38979 11172 39672 11200
rect 38979 11169 38991 11172
rect 38933 11163 38991 11169
rect 39666 11160 39672 11172
rect 39724 11160 39730 11212
rect 39022 11064 39028 11076
rect 38795 11036 39028 11064
rect 38795 11033 38807 11036
rect 38749 11027 38807 11033
rect 39022 11024 39028 11036
rect 39080 11024 39086 11076
rect 36188 10968 36768 10996
rect 36814 10956 36820 11008
rect 36872 10956 36878 11008
rect 38654 10956 38660 11008
rect 38712 10956 38718 11008
rect 1104 10906 41400 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 41400 10906
rect 1104 10832 41400 10854
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 7926 10792 7932 10804
rect 4028 10764 7932 10792
rect 4028 10752 4034 10764
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 9582 10792 9588 10804
rect 8904 10764 9588 10792
rect 8904 10752 8910 10764
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 8570 10656 8576 10668
rect 8251 10628 8576 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8754 10656 8760 10668
rect 8711 10628 8760 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 8956 10665 8984 10764
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10689 10795 10747 10801
rect 10689 10792 10701 10795
rect 9916 10764 10701 10792
rect 9916 10752 9922 10764
rect 10689 10761 10701 10764
rect 10735 10761 10747 10795
rect 13722 10792 13728 10804
rect 10689 10755 10747 10761
rect 13556 10764 13728 10792
rect 13556 10733 13584 10764
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14458 10752 14464 10804
rect 14516 10792 14522 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 14516 10764 15025 10792
rect 14516 10752 14522 10764
rect 15013 10761 15025 10764
rect 15059 10792 15071 10795
rect 15470 10792 15476 10804
rect 15059 10764 15476 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 17589 10795 17647 10801
rect 17589 10761 17601 10795
rect 17635 10792 17647 10795
rect 18230 10792 18236 10804
rect 17635 10764 18236 10792
rect 17635 10761 17647 10764
rect 17589 10755 17647 10761
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 18506 10752 18512 10804
rect 18564 10801 18570 10804
rect 18564 10792 18576 10801
rect 18564 10764 18609 10792
rect 18564 10755 18576 10764
rect 18564 10752 18570 10755
rect 18782 10752 18788 10804
rect 18840 10792 18846 10804
rect 19254 10795 19312 10801
rect 19254 10792 19266 10795
rect 18840 10764 19266 10792
rect 18840 10752 18846 10764
rect 19254 10761 19266 10764
rect 19300 10761 19312 10795
rect 19978 10792 19984 10804
rect 19254 10755 19312 10761
rect 19352 10764 19984 10792
rect 13541 10727 13599 10733
rect 13541 10693 13553 10727
rect 13587 10693 13599 10727
rect 15488 10724 15516 10752
rect 13541 10687 13599 10693
rect 15304 10696 15516 10724
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 8386 10548 8392 10600
rect 8444 10548 8450 10600
rect 8478 10548 8484 10600
rect 8536 10548 8542 10600
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10588 9275 10591
rect 9306 10588 9312 10600
rect 9263 10560 9312 10588
rect 9263 10557 9275 10560
rect 9217 10551 9275 10557
rect 9306 10548 9312 10560
rect 9364 10588 9370 10600
rect 10520 10588 10548 10619
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11112 10628 11529 10656
rect 11112 10616 11118 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 13170 10656 13176 10668
rect 11747 10628 13176 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 15010 10656 15016 10668
rect 14674 10628 15016 10656
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 15304 10665 15332 10696
rect 15562 10684 15568 10736
rect 15620 10684 15626 10736
rect 17126 10684 17132 10736
rect 17184 10684 17190 10736
rect 18046 10684 18052 10736
rect 18104 10724 18110 10736
rect 18141 10727 18199 10733
rect 18141 10724 18153 10727
rect 18104 10696 18153 10724
rect 18104 10684 18110 10696
rect 18141 10693 18153 10696
rect 18187 10724 18199 10727
rect 18877 10727 18935 10733
rect 18877 10724 18889 10727
rect 18187 10696 18889 10724
rect 18187 10693 18199 10696
rect 18141 10687 18199 10693
rect 18877 10693 18889 10696
rect 18923 10693 18935 10727
rect 18877 10687 18935 10693
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10656 15715 10659
rect 16850 10656 16856 10668
rect 15703 10628 16856 10656
rect 15703 10625 15715 10628
rect 15657 10619 15715 10625
rect 13265 10591 13323 10597
rect 9364 10560 10456 10588
rect 10520 10560 11008 10588
rect 9364 10548 9370 10560
rect 8297 10523 8355 10529
rect 8297 10489 8309 10523
rect 8343 10520 8355 10523
rect 8757 10523 8815 10529
rect 8757 10520 8769 10523
rect 8343 10492 8769 10520
rect 8343 10489 8355 10492
rect 8297 10483 8355 10489
rect 8757 10489 8769 10492
rect 8803 10489 8815 10523
rect 10321 10523 10379 10529
rect 10321 10520 10333 10523
rect 8757 10483 8815 10489
rect 8864 10492 10333 10520
rect 8018 10412 8024 10464
rect 8076 10412 8082 10464
rect 8110 10412 8116 10464
rect 8168 10452 8174 10464
rect 8864 10452 8892 10492
rect 10321 10489 10333 10492
rect 10367 10489 10379 10523
rect 10321 10483 10379 10489
rect 8168 10424 8892 10452
rect 9125 10455 9183 10461
rect 8168 10412 8174 10424
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 9582 10452 9588 10464
rect 9171 10424 9588 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 10428 10452 10456 10560
rect 10980 10532 11008 10560
rect 13265 10557 13277 10591
rect 13311 10588 13323 10591
rect 13630 10588 13636 10600
rect 13311 10560 13636 10588
rect 13311 10557 13323 10560
rect 13265 10551 13323 10557
rect 13630 10548 13636 10560
rect 13688 10588 13694 10600
rect 14090 10588 14096 10600
rect 13688 10560 14096 10588
rect 13688 10548 13694 10560
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 15488 10588 15516 10619
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10656 18843 10659
rect 19352 10656 19380 10764
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 26237 10795 26295 10801
rect 22066 10764 23520 10792
rect 19426 10684 19432 10736
rect 19484 10724 19490 10736
rect 19484 10696 19840 10724
rect 19484 10684 19490 10696
rect 19812 10665 19840 10696
rect 20806 10684 20812 10736
rect 20864 10724 20870 10736
rect 21818 10724 21824 10736
rect 20864 10696 21824 10724
rect 20864 10684 20870 10696
rect 21818 10684 21824 10696
rect 21876 10724 21882 10736
rect 22066 10724 22094 10764
rect 23492 10736 23520 10764
rect 25424 10764 25958 10792
rect 23385 10727 23443 10733
rect 23385 10724 23397 10727
rect 21876 10696 22094 10724
rect 23216 10696 23397 10724
rect 21876 10684 21882 10696
rect 23216 10668 23244 10696
rect 23385 10693 23397 10696
rect 23431 10693 23443 10727
rect 23385 10687 23443 10693
rect 23474 10684 23480 10736
rect 23532 10684 23538 10736
rect 23615 10727 23673 10733
rect 23615 10693 23627 10727
rect 23661 10724 23673 10727
rect 24670 10724 24676 10736
rect 23661 10696 24676 10724
rect 23661 10693 23673 10696
rect 23615 10687 23673 10693
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 25222 10684 25228 10736
rect 25280 10684 25286 10736
rect 25424 10733 25452 10764
rect 25409 10727 25467 10733
rect 25409 10693 25421 10727
rect 25455 10693 25467 10727
rect 25930 10724 25958 10764
rect 26237 10761 26249 10795
rect 26283 10792 26295 10795
rect 26510 10792 26516 10804
rect 26283 10764 26516 10792
rect 26283 10761 26295 10764
rect 26237 10755 26295 10761
rect 26510 10752 26516 10764
rect 26568 10752 26574 10804
rect 26789 10795 26847 10801
rect 26789 10761 26801 10795
rect 26835 10792 26847 10795
rect 26878 10792 26884 10804
rect 26835 10764 26884 10792
rect 26835 10761 26847 10764
rect 26789 10755 26847 10761
rect 26878 10752 26884 10764
rect 26936 10752 26942 10804
rect 27430 10752 27436 10804
rect 27488 10752 27494 10804
rect 30101 10795 30159 10801
rect 30101 10761 30113 10795
rect 30147 10792 30159 10795
rect 30929 10795 30987 10801
rect 30929 10792 30941 10795
rect 30147 10764 30941 10792
rect 30147 10761 30159 10764
rect 30101 10755 30159 10761
rect 30929 10761 30941 10764
rect 30975 10761 30987 10795
rect 30929 10755 30987 10761
rect 31297 10795 31355 10801
rect 31297 10761 31309 10795
rect 31343 10792 31355 10795
rect 32122 10792 32128 10804
rect 31343 10764 32128 10792
rect 31343 10761 31355 10764
rect 31297 10755 31355 10761
rect 32122 10752 32128 10764
rect 32180 10752 32186 10804
rect 33226 10792 33232 10804
rect 32416 10764 33232 10792
rect 27338 10724 27344 10736
rect 25930 10696 26193 10724
rect 25409 10687 25467 10693
rect 18831 10628 19380 10656
rect 19613 10659 19671 10665
rect 18831 10625 18843 10628
rect 18785 10619 18843 10625
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10625 19855 10659
rect 19797 10619 19855 10625
rect 15838 10588 15844 10600
rect 15488 10560 15844 10588
rect 15838 10548 15844 10560
rect 15896 10588 15902 10600
rect 16482 10588 16488 10600
rect 15896 10560 16488 10588
rect 15896 10548 15902 10560
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 19628 10588 19656 10619
rect 22830 10616 22836 10668
rect 22888 10656 22894 10668
rect 23109 10659 23167 10665
rect 23109 10656 23121 10659
rect 22888 10628 23121 10656
rect 22888 10616 22894 10628
rect 23109 10625 23121 10628
rect 23155 10625 23167 10659
rect 23109 10619 23167 10625
rect 23198 10616 23204 10668
rect 23256 10616 23262 10668
rect 23293 10659 23351 10665
rect 23293 10625 23305 10659
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 23753 10659 23811 10665
rect 23753 10625 23765 10659
rect 23799 10656 23811 10659
rect 24026 10656 24032 10668
rect 23799 10628 24032 10656
rect 23799 10625 23811 10628
rect 23753 10619 23811 10625
rect 18656 10560 19656 10588
rect 19981 10591 20039 10597
rect 18656 10548 18662 10560
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 20162 10588 20168 10600
rect 20027 10560 20168 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 20254 10548 20260 10600
rect 20312 10588 20318 10600
rect 23308 10588 23336 10619
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 25240 10656 25268 10684
rect 25501 10659 25559 10665
rect 25501 10656 25513 10659
rect 25240 10628 25513 10656
rect 25501 10625 25513 10628
rect 25547 10625 25559 10659
rect 25501 10619 25559 10625
rect 25682 10616 25688 10668
rect 25740 10616 25746 10668
rect 25823 10659 25881 10665
rect 25823 10656 25835 10659
rect 25796 10625 25835 10656
rect 25869 10625 25881 10659
rect 25796 10619 25881 10625
rect 20312 10560 25360 10588
rect 20312 10548 20318 10560
rect 10962 10480 10968 10532
rect 11020 10480 11026 10532
rect 16942 10480 16948 10532
rect 17000 10520 17006 10532
rect 17405 10523 17463 10529
rect 17405 10520 17417 10523
rect 17000 10492 17417 10520
rect 17000 10480 17006 10492
rect 17405 10489 17417 10492
rect 17451 10489 17463 10523
rect 17405 10483 17463 10489
rect 18524 10492 19288 10520
rect 11330 10452 11336 10464
rect 10428 10424 11336 10452
rect 11330 10412 11336 10424
rect 11388 10452 11394 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 11388 10424 11897 10452
rect 11388 10412 11394 10424
rect 11885 10421 11897 10424
rect 11931 10421 11943 10455
rect 11885 10415 11943 10421
rect 15838 10412 15844 10464
rect 15896 10412 15902 10464
rect 18414 10412 18420 10464
rect 18472 10452 18478 10464
rect 18524 10461 18552 10492
rect 19260 10461 19288 10492
rect 21082 10480 21088 10532
rect 21140 10520 21146 10532
rect 24949 10523 25007 10529
rect 24949 10520 24961 10523
rect 21140 10492 24961 10520
rect 21140 10480 21146 10492
rect 24949 10489 24961 10492
rect 24995 10489 25007 10523
rect 24949 10483 25007 10489
rect 18509 10455 18567 10461
rect 18509 10452 18521 10455
rect 18472 10424 18521 10452
rect 18472 10412 18478 10424
rect 18509 10421 18521 10424
rect 18555 10421 18567 10455
rect 18509 10415 18567 10421
rect 19245 10455 19303 10461
rect 19245 10421 19257 10455
rect 19291 10421 19303 10455
rect 19245 10415 19303 10421
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10452 19487 10455
rect 20346 10452 20352 10464
rect 19475 10424 20352 10452
rect 19475 10421 19487 10424
rect 19429 10415 19487 10421
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 25332 10452 25360 10560
rect 25406 10548 25412 10600
rect 25464 10548 25470 10600
rect 25796 10520 25824 10619
rect 25958 10616 25964 10668
rect 26016 10616 26022 10668
rect 26050 10616 26056 10668
rect 26108 10616 26114 10668
rect 26165 10588 26193 10696
rect 26620 10696 27344 10724
rect 26234 10616 26240 10668
rect 26292 10656 26298 10668
rect 26620 10665 26648 10696
rect 27338 10684 27344 10696
rect 27396 10684 27402 10736
rect 27448 10724 27476 10752
rect 30193 10727 30251 10733
rect 30193 10724 30205 10727
rect 27448 10696 30205 10724
rect 30193 10693 30205 10696
rect 30239 10724 30251 10727
rect 30374 10724 30380 10736
rect 30239 10696 30380 10724
rect 30239 10693 30251 10696
rect 30193 10687 30251 10693
rect 30374 10684 30380 10696
rect 30432 10684 30438 10736
rect 26605 10659 26663 10665
rect 26605 10656 26617 10659
rect 26292 10628 26617 10656
rect 26292 10616 26298 10628
rect 26605 10625 26617 10628
rect 26651 10625 26663 10659
rect 26605 10619 26663 10625
rect 26694 10616 26700 10668
rect 26752 10616 26758 10668
rect 26786 10616 26792 10668
rect 26844 10616 26850 10668
rect 32416 10656 32444 10764
rect 33226 10752 33232 10764
rect 33284 10792 33290 10804
rect 33594 10792 33600 10804
rect 33284 10764 33600 10792
rect 33284 10752 33290 10764
rect 33594 10752 33600 10764
rect 33652 10752 33658 10804
rect 34790 10752 34796 10804
rect 34848 10752 34854 10804
rect 35250 10752 35256 10804
rect 35308 10752 35314 10804
rect 38654 10752 38660 10804
rect 38712 10752 38718 10804
rect 38746 10752 38752 10804
rect 38804 10792 38810 10804
rect 39025 10795 39083 10801
rect 39025 10792 39037 10795
rect 38804 10764 39037 10792
rect 38804 10752 38810 10764
rect 39025 10761 39037 10764
rect 39071 10761 39083 10795
rect 39025 10755 39083 10761
rect 32582 10684 32588 10736
rect 32640 10724 32646 10736
rect 32640 10696 34652 10724
rect 32640 10684 32646 10696
rect 32493 10659 32551 10665
rect 32493 10656 32505 10659
rect 32416 10628 32505 10656
rect 32493 10625 32505 10628
rect 32539 10625 32551 10659
rect 32493 10619 32551 10625
rect 26421 10591 26479 10597
rect 26421 10588 26433 10591
rect 26165 10560 26433 10588
rect 26421 10557 26433 10560
rect 26467 10588 26479 10591
rect 26712 10588 26740 10616
rect 26467 10560 26740 10588
rect 26467 10557 26479 10560
rect 26421 10551 26479 10557
rect 26804 10520 26832 10616
rect 30282 10548 30288 10600
rect 30340 10548 30346 10600
rect 31386 10548 31392 10600
rect 31444 10548 31450 10600
rect 32600 10597 32628 10684
rect 34624 10668 34652 10696
rect 33042 10616 33048 10668
rect 33100 10616 33106 10668
rect 33321 10659 33379 10665
rect 33321 10625 33333 10659
rect 33367 10656 33379 10659
rect 33367 10628 33732 10656
rect 33367 10625 33379 10628
rect 33321 10619 33379 10625
rect 31573 10591 31631 10597
rect 31573 10557 31585 10591
rect 31619 10557 31631 10591
rect 31573 10551 31631 10557
rect 32585 10591 32643 10597
rect 32585 10557 32597 10591
rect 32631 10557 32643 10591
rect 32585 10551 32643 10557
rect 25796 10492 26832 10520
rect 31588 10520 31616 10551
rect 32858 10548 32864 10600
rect 32916 10548 32922 10600
rect 33229 10591 33287 10597
rect 33229 10557 33241 10591
rect 33275 10557 33287 10591
rect 33229 10551 33287 10557
rect 31662 10520 31668 10532
rect 31588 10492 31668 10520
rect 31662 10480 31668 10492
rect 31720 10520 31726 10532
rect 32876 10520 32904 10548
rect 31720 10492 32904 10520
rect 33244 10520 33272 10551
rect 33594 10548 33600 10600
rect 33652 10548 33658 10600
rect 33704 10588 33732 10628
rect 33778 10616 33784 10668
rect 33836 10616 33842 10668
rect 34606 10616 34612 10668
rect 34664 10616 34670 10668
rect 34808 10656 34836 10752
rect 35161 10659 35219 10665
rect 34808 10628 35112 10656
rect 35084 10588 35112 10628
rect 35161 10625 35173 10659
rect 35207 10656 35219 10659
rect 35268 10656 35296 10752
rect 35989 10727 36047 10733
rect 35360 10696 35848 10724
rect 35360 10665 35388 10696
rect 35820 10665 35848 10696
rect 35989 10693 36001 10727
rect 36035 10724 36047 10727
rect 36081 10727 36139 10733
rect 36081 10724 36093 10727
rect 36035 10696 36093 10724
rect 36035 10693 36047 10696
rect 35989 10687 36047 10693
rect 36081 10693 36093 10696
rect 36127 10693 36139 10727
rect 36814 10724 36820 10736
rect 36081 10687 36139 10693
rect 36188 10696 36820 10724
rect 35207 10628 35296 10656
rect 35345 10659 35403 10665
rect 35207 10625 35219 10628
rect 35161 10619 35219 10625
rect 35345 10625 35357 10659
rect 35391 10625 35403 10659
rect 35345 10619 35403 10625
rect 35713 10659 35771 10665
rect 35713 10625 35725 10659
rect 35759 10625 35771 10659
rect 35713 10619 35771 10625
rect 35805 10659 35863 10665
rect 35805 10625 35817 10659
rect 35851 10656 35863 10659
rect 36188 10656 36216 10696
rect 36372 10665 36400 10696
rect 36814 10684 36820 10696
rect 36872 10684 36878 10736
rect 35851 10628 36216 10656
rect 36265 10659 36323 10665
rect 35851 10625 35863 10628
rect 35805 10619 35863 10625
rect 36265 10625 36277 10659
rect 36311 10625 36323 10659
rect 36265 10619 36323 10625
rect 36357 10659 36415 10665
rect 36357 10625 36369 10659
rect 36403 10625 36415 10659
rect 36357 10619 36415 10625
rect 35728 10588 35756 10619
rect 33704 10560 34836 10588
rect 35084 10560 35756 10588
rect 33965 10523 34023 10529
rect 33965 10520 33977 10523
rect 33244 10492 33977 10520
rect 31720 10480 31726 10492
rect 33965 10489 33977 10492
rect 34011 10489 34023 10523
rect 33965 10483 34023 10489
rect 34808 10464 34836 10560
rect 35728 10520 35756 10560
rect 35986 10548 35992 10600
rect 36044 10548 36050 10600
rect 36280 10520 36308 10619
rect 39114 10548 39120 10600
rect 39172 10548 39178 10600
rect 39298 10548 39304 10600
rect 39356 10548 39362 10600
rect 35728 10492 36308 10520
rect 25958 10452 25964 10464
rect 25332 10424 25964 10452
rect 25958 10412 25964 10424
rect 26016 10412 26022 10464
rect 29730 10412 29736 10464
rect 29788 10412 29794 10464
rect 32769 10455 32827 10461
rect 32769 10421 32781 10455
rect 32815 10452 32827 10455
rect 33045 10455 33103 10461
rect 33045 10452 33057 10455
rect 32815 10424 33057 10452
rect 32815 10421 32827 10424
rect 32769 10415 32827 10421
rect 33045 10421 33057 10424
rect 33091 10452 33103 10455
rect 33134 10452 33140 10464
rect 33091 10424 33140 10452
rect 33091 10421 33103 10424
rect 33045 10415 33103 10421
rect 33134 10412 33140 10424
rect 33192 10412 33198 10464
rect 33502 10412 33508 10464
rect 33560 10412 33566 10464
rect 34790 10412 34796 10464
rect 34848 10452 34854 10464
rect 35253 10455 35311 10461
rect 35253 10452 35265 10455
rect 34848 10424 35265 10452
rect 34848 10412 34854 10424
rect 35253 10421 35265 10424
rect 35299 10421 35311 10455
rect 35253 10415 35311 10421
rect 36078 10412 36084 10464
rect 36136 10412 36142 10464
rect 38654 10412 38660 10464
rect 38712 10452 38718 10464
rect 39316 10452 39344 10548
rect 38712 10424 39344 10452
rect 38712 10412 38718 10424
rect 1104 10362 41400 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 41400 10362
rect 1104 10288 41400 10310
rect 4893 10251 4951 10257
rect 4893 10217 4905 10251
rect 4939 10248 4951 10251
rect 5166 10248 5172 10260
rect 4939 10220 5172 10248
rect 4939 10217 4951 10220
rect 4893 10211 4951 10217
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5644 10220 7144 10248
rect 5184 10112 5212 10208
rect 5537 10115 5595 10121
rect 5537 10112 5549 10115
rect 5184 10084 5549 10112
rect 5537 10081 5549 10084
rect 5583 10081 5595 10115
rect 5537 10075 5595 10081
rect 4798 10004 4804 10056
rect 4856 10004 4862 10056
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 4614 9936 4620 9988
rect 4672 9936 4678 9988
rect 4908 9976 4936 10007
rect 5166 10004 5172 10056
rect 5224 10004 5230 10056
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5644 10044 5672 10220
rect 6549 10183 6607 10189
rect 6549 10149 6561 10183
rect 6595 10180 6607 10183
rect 6730 10180 6736 10192
rect 6595 10152 6736 10180
rect 6595 10149 6607 10152
rect 6549 10143 6607 10149
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 6822 10140 6828 10192
rect 6880 10140 6886 10192
rect 6840 10112 6868 10140
rect 7116 10124 7144 10220
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 8444 10220 8769 10248
rect 8444 10208 8450 10220
rect 8757 10217 8769 10220
rect 8803 10217 8815 10251
rect 8757 10211 8815 10217
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 11606 10248 11612 10260
rect 9640 10220 11612 10248
rect 9640 10208 9646 10220
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 12066 10208 12072 10260
rect 12124 10208 12130 10260
rect 15838 10208 15844 10260
rect 15896 10208 15902 10260
rect 18874 10208 18880 10260
rect 18932 10208 18938 10260
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 22373 10251 22431 10257
rect 22373 10248 22385 10251
rect 20772 10220 22385 10248
rect 20772 10208 20778 10220
rect 22373 10217 22385 10220
rect 22419 10217 22431 10251
rect 22373 10211 22431 10217
rect 23293 10251 23351 10257
rect 23293 10217 23305 10251
rect 23339 10248 23351 10251
rect 23842 10248 23848 10260
rect 23339 10220 23848 10248
rect 23339 10217 23351 10220
rect 23293 10211 23351 10217
rect 23842 10208 23848 10220
rect 23900 10208 23906 10260
rect 24026 10208 24032 10260
rect 24084 10208 24090 10260
rect 24946 10208 24952 10260
rect 25004 10248 25010 10260
rect 25498 10248 25504 10260
rect 25004 10220 25504 10248
rect 25004 10208 25010 10220
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 25958 10208 25964 10260
rect 26016 10208 26022 10260
rect 26329 10251 26387 10257
rect 26329 10217 26341 10251
rect 26375 10248 26387 10251
rect 26418 10248 26424 10260
rect 26375 10220 26424 10248
rect 26375 10217 26387 10220
rect 26329 10211 26387 10217
rect 26418 10208 26424 10220
rect 26476 10208 26482 10260
rect 29730 10208 29736 10260
rect 29788 10208 29794 10260
rect 30929 10251 30987 10257
rect 30929 10217 30941 10251
rect 30975 10248 30987 10251
rect 31386 10248 31392 10260
rect 30975 10220 31392 10248
rect 30975 10217 30987 10220
rect 30929 10211 30987 10217
rect 31386 10208 31392 10220
rect 31444 10208 31450 10260
rect 32861 10251 32919 10257
rect 32861 10217 32873 10251
rect 32907 10248 32919 10251
rect 33042 10248 33048 10260
rect 32907 10220 33048 10248
rect 32907 10217 32919 10220
rect 32861 10211 32919 10217
rect 33042 10208 33048 10220
rect 33100 10208 33106 10260
rect 35986 10248 35992 10260
rect 33244 10220 35992 10248
rect 8110 10180 8116 10192
rect 8036 10152 8116 10180
rect 5736 10084 6868 10112
rect 5736 10053 5764 10084
rect 5491 10016 5672 10044
rect 5721 10047 5779 10053
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10044 5963 10047
rect 6270 10044 6276 10056
rect 5951 10016 6276 10044
rect 5951 10013 5963 10016
rect 5905 10007 5963 10013
rect 5626 9976 5632 9988
rect 4908 9948 5632 9976
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 5736 9976 5764 10007
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6840 10053 6868 10084
rect 7098 10072 7104 10124
rect 7156 10072 7162 10124
rect 8036 10053 8064 10152
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 11330 10180 11336 10192
rect 10520 10152 11336 10180
rect 8220 10112 8248 10140
rect 9122 10112 9128 10124
rect 8128 10084 8248 10112
rect 8496 10084 9128 10112
rect 8128 10053 8156 10084
rect 8496 10053 8524 10084
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6472 10016 6684 10044
rect 6783 10016 6837 10044
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 5736 9948 6101 9976
rect 6089 9945 6101 9948
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 5074 9868 5080 9920
rect 5132 9868 5138 9920
rect 6288 9908 6316 10004
rect 6472 9985 6500 10016
rect 6457 9979 6515 9985
rect 6457 9945 6469 9979
rect 6503 9945 6515 9979
rect 6457 9939 6515 9945
rect 6546 9936 6552 9988
rect 6604 9936 6610 9988
rect 6656 9976 6684 10016
rect 6825 10013 6837 10016
rect 6871 10044 6883 10047
rect 7561 10047 7619 10053
rect 7561 10044 7573 10047
rect 6871 10016 7573 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7561 10013 7573 10016
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 8206 10047 8264 10053
rect 8206 10013 8218 10047
rect 8252 10013 8264 10047
rect 8206 10007 8264 10013
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 8619 10047 8677 10053
rect 8619 10013 8631 10047
rect 8665 10044 8677 10047
rect 9490 10044 9496 10056
rect 8665 10016 9496 10044
rect 8665 10013 8677 10016
rect 8619 10007 8677 10013
rect 6914 9976 6920 9988
rect 6656 9948 6920 9976
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 7760 9976 7788 10007
rect 8220 9976 8248 10007
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 9582 10004 9588 10056
rect 9640 10004 9646 10056
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10044 10379 10047
rect 10520 10044 10548 10152
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 10980 10084 11713 10112
rect 10980 10053 11008 10084
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 11974 10072 11980 10124
rect 12032 10072 12038 10124
rect 12084 10112 12112 10208
rect 12084 10084 12480 10112
rect 11146 10053 11152 10056
rect 10367 10016 10548 10044
rect 10965 10047 11023 10053
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 10965 10013 10977 10047
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11113 10047 11152 10053
rect 11113 10013 11125 10047
rect 11113 10007 11152 10013
rect 11146 10004 11152 10007
rect 11204 10004 11210 10056
rect 11330 10004 11336 10056
rect 11388 10004 11394 10056
rect 11422 10004 11428 10056
rect 11480 10053 11486 10056
rect 11480 10007 11488 10053
rect 11480 10004 11486 10007
rect 11882 10004 11888 10056
rect 11940 10004 11946 10056
rect 11992 10044 12020 10072
rect 12452 10053 12480 10084
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 11992 10016 12173 10044
rect 12161 10013 12173 10016
rect 12207 10044 12219 10047
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 12207 10016 12265 10044
rect 12207 10013 12219 10016
rect 12161 10007 12219 10013
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 15657 10047 15715 10053
rect 15657 10013 15669 10047
rect 15703 10013 15715 10047
rect 15856 10044 15884 10208
rect 23474 10140 23480 10192
rect 23532 10140 23538 10192
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 21450 10112 21456 10124
rect 16439 10084 21456 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 22370 10072 22376 10124
rect 22428 10112 22434 10124
rect 22428 10084 23336 10112
rect 22428 10072 22434 10084
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 15856 10016 16589 10044
rect 15657 10007 15715 10013
rect 16577 10013 16589 10016
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 8294 9976 8300 9988
rect 7760 9948 8300 9976
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 8386 9936 8392 9988
rect 8444 9936 8450 9988
rect 11241 9979 11299 9985
rect 11241 9976 11253 9979
rect 8588 9948 9982 9976
rect 10612 9948 11253 9976
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 6288 9880 6745 9908
rect 6733 9877 6745 9880
rect 6779 9877 6791 9911
rect 6733 9871 6791 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 7929 9911 7987 9917
rect 7929 9908 7941 9911
rect 7800 9880 7941 9908
rect 7800 9868 7806 9880
rect 7929 9877 7941 9880
rect 7975 9908 7987 9911
rect 8588 9908 8616 9948
rect 7975 9880 8616 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 10612 9908 10640 9948
rect 11241 9945 11253 9948
rect 11287 9945 11299 9979
rect 12621 9979 12679 9985
rect 12621 9976 12633 9979
rect 11241 9939 11299 9945
rect 11348 9948 12633 9976
rect 9272 9880 10640 9908
rect 9272 9868 9278 9880
rect 10962 9868 10968 9920
rect 11020 9908 11026 9920
rect 11348 9908 11376 9948
rect 12621 9945 12633 9948
rect 12667 9945 12679 9979
rect 12621 9939 12679 9945
rect 11020 9880 11376 9908
rect 11020 9868 11026 9880
rect 11606 9868 11612 9920
rect 11664 9868 11670 9920
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 15672 9908 15700 10007
rect 16761 9979 16819 9985
rect 16761 9976 16773 9979
rect 15856 9948 16773 9976
rect 15856 9908 15884 9948
rect 16761 9945 16773 9948
rect 16807 9945 16819 9979
rect 16868 9976 16896 10007
rect 18598 10004 18604 10056
rect 18656 10004 18662 10056
rect 18874 10004 18880 10056
rect 18932 10004 18938 10056
rect 21726 10004 21732 10056
rect 21784 10004 21790 10056
rect 22281 10047 22339 10053
rect 22281 10013 22293 10047
rect 22327 10044 22339 10047
rect 22462 10044 22468 10056
rect 22327 10016 22468 10044
rect 22327 10013 22339 10016
rect 22281 10007 22339 10013
rect 22462 10004 22468 10016
rect 22520 10004 22526 10056
rect 23198 10044 23204 10056
rect 22756 10016 23204 10044
rect 18892 9976 18920 10004
rect 19242 9976 19248 9988
rect 16868 9948 19248 9976
rect 16761 9939 16819 9945
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 22002 9936 22008 9988
rect 22060 9936 22066 9988
rect 22756 9920 22784 10016
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 15528 9880 15884 9908
rect 15528 9868 15534 9880
rect 16298 9868 16304 9920
rect 16356 9868 16362 9920
rect 22738 9868 22744 9920
rect 22796 9868 22802 9920
rect 23308 9908 23336 10084
rect 23385 10047 23443 10053
rect 23385 10013 23397 10047
rect 23431 10044 23443 10047
rect 23492 10044 23520 10140
rect 24044 10112 24072 10208
rect 25682 10112 25688 10124
rect 24044 10084 25688 10112
rect 25682 10072 25688 10084
rect 25740 10112 25746 10124
rect 25740 10084 25820 10112
rect 25740 10072 25746 10084
rect 25222 10044 25228 10056
rect 23431 10016 25228 10044
rect 23431 10013 23443 10016
rect 23385 10007 23443 10013
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 25314 10004 25320 10056
rect 25372 10004 25378 10056
rect 25792 10053 25820 10084
rect 25777 10047 25835 10053
rect 25777 10013 25789 10047
rect 25823 10013 25835 10047
rect 25976 10044 26004 10208
rect 26053 10047 26111 10053
rect 26053 10044 26065 10047
rect 25976 10016 26065 10044
rect 25777 10007 25835 10013
rect 26053 10013 26065 10016
rect 26099 10013 26111 10047
rect 26053 10007 26111 10013
rect 26145 10047 26203 10053
rect 26145 10013 26157 10047
rect 26191 10044 26203 10047
rect 26970 10044 26976 10056
rect 26191 10016 26976 10044
rect 26191 10013 26203 10016
rect 26145 10007 26203 10013
rect 26970 10004 26976 10016
rect 27028 10004 27034 10056
rect 27982 10004 27988 10056
rect 28040 10004 28046 10056
rect 29365 10047 29423 10053
rect 29365 10013 29377 10047
rect 29411 10044 29423 10047
rect 29748 10044 29776 10208
rect 32582 10140 32588 10192
rect 32640 10180 32646 10192
rect 33137 10183 33195 10189
rect 33137 10180 33149 10183
rect 32640 10152 33149 10180
rect 32640 10140 32646 10152
rect 33137 10149 33149 10152
rect 33183 10149 33195 10183
rect 33137 10143 33195 10149
rect 30745 10115 30803 10121
rect 30745 10081 30757 10115
rect 30791 10112 30803 10115
rect 31110 10112 31116 10124
rect 30791 10084 31116 10112
rect 30791 10081 30803 10084
rect 30745 10075 30803 10081
rect 31110 10072 31116 10084
rect 31168 10072 31174 10124
rect 31294 10072 31300 10124
rect 31352 10112 31358 10124
rect 32769 10115 32827 10121
rect 32769 10112 32781 10115
rect 31352 10084 32781 10112
rect 31352 10072 31358 10084
rect 32769 10081 32781 10084
rect 32815 10112 32827 10115
rect 33244 10112 33272 10220
rect 35986 10208 35992 10220
rect 36044 10208 36050 10260
rect 39114 10208 39120 10260
rect 39172 10248 39178 10260
rect 40313 10251 40371 10257
rect 40313 10248 40325 10251
rect 39172 10220 40325 10248
rect 39172 10208 39178 10220
rect 40313 10217 40325 10220
rect 40359 10217 40371 10251
rect 40313 10211 40371 10217
rect 34698 10140 34704 10192
rect 34756 10180 34762 10192
rect 35161 10183 35219 10189
rect 35161 10180 35173 10183
rect 34756 10152 35173 10180
rect 34756 10140 34762 10152
rect 35161 10149 35173 10152
rect 35207 10149 35219 10183
rect 35161 10143 35219 10149
rect 32815 10084 33272 10112
rect 34425 10115 34483 10121
rect 32815 10081 32827 10084
rect 32769 10075 32827 10081
rect 34425 10081 34437 10115
rect 34471 10112 34483 10115
rect 34471 10084 35388 10112
rect 34471 10081 34483 10084
rect 34425 10075 34483 10081
rect 29411 10016 29776 10044
rect 29411 10013 29423 10016
rect 29365 10007 29423 10013
rect 30650 10004 30656 10056
rect 30708 10004 30714 10056
rect 32490 10004 32496 10056
rect 32548 10044 32554 10056
rect 32861 10047 32919 10053
rect 32861 10044 32873 10047
rect 32548 10016 32873 10044
rect 32548 10004 32554 10016
rect 25332 9976 25360 10004
rect 25866 9976 25872 9988
rect 25332 9948 25872 9976
rect 25866 9936 25872 9948
rect 25924 9976 25930 9988
rect 25961 9979 26019 9985
rect 25961 9976 25973 9979
rect 25924 9948 25973 9976
rect 25924 9936 25930 9948
rect 25961 9945 25973 9948
rect 26007 9945 26019 9979
rect 30466 9976 30472 9988
rect 25961 9939 26019 9945
rect 26068 9948 30472 9976
rect 26068 9908 26096 9948
rect 30466 9936 30472 9948
rect 30524 9936 30530 9988
rect 32692 9976 32720 10016
rect 32861 10013 32873 10016
rect 32907 10013 32919 10047
rect 32861 10007 32919 10013
rect 33042 10004 33048 10056
rect 33100 10004 33106 10056
rect 33134 10004 33140 10056
rect 33192 10004 33198 10056
rect 33321 10047 33379 10053
rect 33321 10013 33333 10047
rect 33367 10044 33379 10047
rect 34333 10047 34391 10053
rect 34333 10044 34345 10047
rect 33367 10016 34345 10044
rect 33367 10013 33379 10016
rect 33321 10007 33379 10013
rect 34333 10013 34345 10016
rect 34379 10013 34391 10047
rect 34333 10007 34391 10013
rect 34517 10047 34575 10053
rect 34517 10013 34529 10047
rect 34563 10044 34575 10047
rect 34606 10044 34612 10056
rect 34563 10016 34612 10044
rect 34563 10013 34575 10016
rect 34517 10007 34575 10013
rect 33778 9976 33784 9988
rect 32692 9948 33784 9976
rect 32692 9920 32720 9948
rect 33778 9936 33784 9948
rect 33836 9936 33842 9988
rect 34348 9976 34376 10007
rect 34606 10004 34612 10016
rect 34664 10004 34670 10056
rect 34701 10047 34759 10053
rect 34701 10013 34713 10047
rect 34747 10044 34759 10047
rect 34790 10044 34796 10056
rect 34747 10016 34796 10044
rect 34747 10013 34759 10016
rect 34701 10007 34759 10013
rect 34716 9976 34744 10007
rect 34790 10004 34796 10016
rect 34848 10004 34854 10056
rect 35360 10053 35388 10084
rect 39022 10072 39028 10124
rect 39080 10112 39086 10124
rect 39080 10084 39712 10112
rect 39080 10072 39086 10084
rect 35345 10047 35403 10053
rect 35345 10013 35357 10047
rect 35391 10013 35403 10047
rect 35345 10007 35403 10013
rect 35437 10047 35495 10053
rect 35437 10013 35449 10047
rect 35483 10013 35495 10047
rect 35437 10007 35495 10013
rect 34885 9979 34943 9985
rect 34885 9976 34897 9979
rect 34348 9948 34744 9976
rect 34808 9948 34897 9976
rect 34808 9920 34836 9948
rect 34885 9945 34897 9948
rect 34931 9945 34943 9979
rect 34885 9939 34943 9945
rect 35161 9979 35219 9985
rect 35161 9945 35173 9979
rect 35207 9976 35219 9979
rect 35250 9976 35256 9988
rect 35207 9948 35256 9976
rect 35207 9945 35219 9948
rect 35161 9939 35219 9945
rect 35250 9936 35256 9948
rect 35308 9936 35314 9988
rect 35452 9976 35480 10007
rect 39206 10004 39212 10056
rect 39264 10044 39270 10056
rect 39390 10044 39396 10056
rect 39264 10016 39396 10044
rect 39264 10004 39270 10016
rect 39390 10004 39396 10016
rect 39448 10044 39454 10056
rect 39684 10053 39712 10084
rect 39758 10072 39764 10124
rect 39816 10112 39822 10124
rect 40129 10115 40187 10121
rect 40129 10112 40141 10115
rect 39816 10084 40141 10112
rect 39816 10072 39822 10084
rect 40129 10081 40141 10084
rect 40175 10081 40187 10115
rect 40129 10075 40187 10081
rect 39485 10047 39543 10053
rect 39485 10044 39497 10047
rect 39448 10016 39497 10044
rect 39448 10004 39454 10016
rect 39485 10013 39497 10016
rect 39531 10013 39543 10047
rect 39485 10007 39543 10013
rect 39669 10047 39727 10053
rect 39669 10013 39681 10047
rect 39715 10013 39727 10047
rect 39669 10007 39727 10013
rect 39850 10004 39856 10056
rect 39908 10044 39914 10056
rect 40037 10047 40095 10053
rect 40037 10044 40049 10047
rect 39908 10016 40049 10044
rect 39908 10004 39914 10016
rect 40037 10013 40049 10016
rect 40083 10013 40095 10047
rect 40037 10007 40095 10013
rect 35360 9948 35480 9976
rect 23308 9880 26096 9908
rect 27798 9868 27804 9920
rect 27856 9868 27862 9920
rect 29178 9868 29184 9920
rect 29236 9868 29242 9920
rect 32674 9868 32680 9920
rect 32732 9868 32738 9920
rect 32766 9868 32772 9920
rect 32824 9868 32830 9920
rect 34606 9868 34612 9920
rect 34664 9908 34670 9920
rect 34790 9908 34796 9920
rect 34664 9880 34796 9908
rect 34664 9868 34670 9880
rect 34790 9868 34796 9880
rect 34848 9868 34854 9920
rect 35069 9911 35127 9917
rect 35069 9877 35081 9911
rect 35115 9908 35127 9911
rect 35360 9908 35388 9948
rect 35115 9880 35388 9908
rect 35115 9877 35127 9880
rect 35069 9871 35127 9877
rect 39390 9868 39396 9920
rect 39448 9868 39454 9920
rect 39574 9868 39580 9920
rect 39632 9868 39638 9920
rect 1104 9818 41400 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 41400 9818
rect 1104 9744 41400 9766
rect 10778 9704 10784 9716
rect 3896 9676 4476 9704
rect 3896 9577 3924 9676
rect 3973 9639 4031 9645
rect 3973 9605 3985 9639
rect 4019 9636 4031 9639
rect 4448 9636 4476 9676
rect 10336 9676 10784 9704
rect 8760 9648 8812 9654
rect 4890 9636 4896 9648
rect 4019 9608 4384 9636
rect 4448 9608 4896 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 4356 9577 4384 9608
rect 4890 9596 4896 9608
rect 4948 9636 4954 9648
rect 5350 9636 5356 9648
rect 4948 9608 5356 9636
rect 4948 9596 4954 9608
rect 5350 9596 5356 9608
rect 5408 9596 5414 9648
rect 6733 9639 6791 9645
rect 6733 9605 6745 9639
rect 6779 9636 6791 9639
rect 8018 9636 8024 9648
rect 6779 9608 8024 9636
rect 6779 9605 6791 9608
rect 6733 9599 6791 9605
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 8760 9590 8812 9596
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 4614 9568 4620 9580
rect 4387 9540 4620 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 4080 9432 4108 9531
rect 4172 9500 4200 9531
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 4801 9531 4859 9537
rect 5000 9540 5457 9568
rect 4816 9500 4844 9531
rect 5000 9509 5028 9540
rect 5445 9537 5457 9540
rect 5491 9568 5503 9571
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 5491 9540 5764 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 4172 9472 4476 9500
rect 4338 9432 4344 9444
rect 4080 9404 4344 9432
rect 4338 9392 4344 9404
rect 4396 9392 4402 9444
rect 4448 9441 4476 9472
rect 4632 9472 4844 9500
rect 4985 9503 5043 9509
rect 4632 9444 4660 9472
rect 4985 9469 4997 9503
rect 5031 9469 5043 9503
rect 4985 9463 5043 9469
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5353 9503 5411 9509
rect 5353 9500 5365 9503
rect 5132 9472 5365 9500
rect 5132 9460 5138 9472
rect 5353 9469 5365 9472
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 4433 9435 4491 9441
rect 4433 9401 4445 9435
rect 4479 9401 4491 9435
rect 4433 9395 4491 9401
rect 4614 9392 4620 9444
rect 4672 9432 4678 9444
rect 5166 9432 5172 9444
rect 4672 9404 5172 9432
rect 4672 9392 4678 9404
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 5442 9364 5448 9376
rect 4203 9336 5448 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5736 9364 5764 9540
rect 5828 9540 6837 9568
rect 5828 9441 5856 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 7742 9568 7748 9580
rect 7699 9540 7748 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8110 9528 8116 9580
rect 8168 9528 8174 9580
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6512 9472 6929 9500
rect 6512 9460 6518 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 5813 9435 5871 9441
rect 5813 9401 5825 9435
rect 5859 9401 5871 9435
rect 7098 9432 7104 9444
rect 5813 9395 5871 9401
rect 5920 9404 6500 9432
rect 5920 9364 5948 9404
rect 5736 9336 5948 9364
rect 6362 9324 6368 9376
rect 6420 9324 6426 9376
rect 6472 9364 6500 9404
rect 6886 9404 7104 9432
rect 6886 9364 6914 9404
rect 7098 9392 7104 9404
rect 7156 9432 7162 9444
rect 8772 9432 8800 9590
rect 9858 9528 9864 9580
rect 9916 9528 9922 9580
rect 10336 9577 10364 9676
rect 10778 9664 10784 9676
rect 10836 9704 10842 9716
rect 11146 9704 11152 9716
rect 10836 9676 11152 9704
rect 10836 9664 10842 9676
rect 11146 9664 11152 9676
rect 11204 9704 11210 9716
rect 15381 9707 15439 9713
rect 11204 9676 12434 9704
rect 11204 9664 11210 9676
rect 10502 9596 10508 9648
rect 10560 9596 10566 9648
rect 12406 9636 12434 9676
rect 15381 9673 15393 9707
rect 15427 9704 15439 9707
rect 15470 9704 15476 9716
rect 15427 9676 15476 9704
rect 15427 9673 15439 9676
rect 15381 9667 15439 9673
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 15841 9707 15899 9713
rect 15841 9673 15853 9707
rect 15887 9704 15899 9707
rect 16298 9704 16304 9716
rect 15887 9676 16304 9704
rect 15887 9673 15899 9676
rect 15841 9667 15899 9673
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 21726 9664 21732 9716
rect 21784 9704 21790 9716
rect 21910 9704 21916 9716
rect 21784 9676 21916 9704
rect 21784 9664 21790 9676
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 25041 9707 25099 9713
rect 25041 9673 25053 9707
rect 25087 9704 25099 9707
rect 25406 9704 25412 9716
rect 25087 9676 25412 9704
rect 25087 9673 25099 9676
rect 25041 9667 25099 9673
rect 25406 9664 25412 9676
rect 25464 9664 25470 9716
rect 25792 9676 28028 9704
rect 15194 9636 15200 9648
rect 12406 9608 12558 9636
rect 15134 9608 15200 9636
rect 15194 9596 15200 9608
rect 15252 9636 15258 9648
rect 15562 9636 15568 9648
rect 15252 9608 15568 9636
rect 15252 9596 15258 9608
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 15930 9596 15936 9648
rect 15988 9596 15994 9648
rect 16853 9639 16911 9645
rect 16853 9605 16865 9639
rect 16899 9636 16911 9639
rect 19337 9639 19395 9645
rect 16899 9608 17172 9636
rect 16899 9605 16911 9608
rect 16853 9599 16911 9605
rect 17144 9580 17172 9608
rect 19337 9605 19349 9639
rect 19383 9636 19395 9639
rect 19518 9636 19524 9648
rect 19383 9608 19524 9636
rect 19383 9605 19395 9608
rect 19337 9599 19395 9605
rect 19518 9596 19524 9608
rect 19576 9636 19582 9648
rect 20070 9636 20076 9648
rect 19576 9608 20076 9636
rect 19576 9596 19582 9608
rect 20070 9596 20076 9608
rect 20128 9596 20134 9648
rect 20993 9639 21051 9645
rect 20993 9636 21005 9639
rect 20180 9608 21005 9636
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 12124 9540 12173 9568
rect 12124 9528 12130 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 13630 9528 13636 9580
rect 13688 9528 13694 9580
rect 16574 9568 16580 9580
rect 15120 9540 16580 9568
rect 13906 9460 13912 9512
rect 13964 9460 13970 9512
rect 7156 9404 8800 9432
rect 7156 9392 7162 9404
rect 6472 9336 6914 9364
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 15120 9364 15148 9540
rect 16574 9528 16580 9540
rect 16632 9568 16638 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16632 9540 16681 9568
rect 16632 9528 16638 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 16945 9571 17003 9577
rect 16945 9568 16957 9571
rect 16816 9540 16957 9568
rect 16816 9528 16822 9540
rect 16945 9537 16957 9540
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 17126 9528 17132 9580
rect 17184 9528 17190 9580
rect 20180 9568 20208 9608
rect 20993 9605 21005 9608
rect 21039 9605 21051 9639
rect 22922 9636 22928 9648
rect 20993 9599 21051 9605
rect 21192 9608 22928 9636
rect 19444 9540 20208 9568
rect 16114 9460 16120 9512
rect 16172 9460 16178 9512
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 19444 9509 19472 9540
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20772 9540 20913 9568
rect 20772 9528 20778 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 19392 9472 19441 9500
rect 19392 9460 19398 9472
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9500 19671 9503
rect 20438 9500 20444 9512
rect 19659 9472 20444 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 21192 9509 21220 9608
rect 22922 9596 22928 9608
rect 22980 9596 22986 9648
rect 23014 9596 23020 9648
rect 23072 9636 23078 9648
rect 25792 9636 25820 9676
rect 23072 9608 25820 9636
rect 26073 9639 26131 9645
rect 23072 9596 23078 9608
rect 26073 9605 26085 9639
rect 26119 9636 26131 9639
rect 26119 9608 27936 9636
rect 26119 9605 26131 9608
rect 26073 9599 26131 9605
rect 21361 9571 21419 9577
rect 21361 9537 21373 9571
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 21913 9571 21971 9577
rect 21913 9537 21925 9571
rect 21959 9568 21971 9571
rect 22002 9568 22008 9580
rect 21959 9540 22008 9568
rect 21959 9537 21971 9540
rect 21913 9531 21971 9537
rect 21177 9503 21235 9509
rect 21177 9469 21189 9503
rect 21223 9469 21235 9503
rect 21177 9463 21235 9469
rect 17221 9435 17279 9441
rect 17221 9401 17233 9435
rect 17267 9432 17279 9435
rect 17586 9432 17592 9444
rect 17267 9404 17592 9432
rect 17267 9401 17279 9404
rect 17221 9395 17279 9401
rect 17586 9392 17592 9404
rect 17644 9392 17650 9444
rect 20533 9435 20591 9441
rect 17696 9404 19334 9432
rect 7984 9336 15148 9364
rect 7984 9324 7990 9336
rect 15470 9324 15476 9376
rect 15528 9324 15534 9376
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 17696 9364 17724 9404
rect 19306 9376 19334 9404
rect 20533 9401 20545 9435
rect 20579 9432 20591 9435
rect 21376 9432 21404 9531
rect 22002 9528 22008 9540
rect 22060 9528 22066 9580
rect 25222 9528 25228 9580
rect 25280 9528 25286 9580
rect 25314 9528 25320 9580
rect 25372 9568 25378 9580
rect 25372 9540 25544 9568
rect 25372 9528 25378 9540
rect 21450 9460 21456 9512
rect 21508 9500 21514 9512
rect 25516 9509 25544 9540
rect 25682 9528 25688 9580
rect 25740 9528 25746 9580
rect 25958 9577 25964 9580
rect 25778 9571 25836 9577
rect 25778 9537 25790 9571
rect 25824 9537 25836 9571
rect 25778 9531 25836 9537
rect 25915 9571 25964 9577
rect 25915 9537 25927 9571
rect 25961 9537 25964 9571
rect 25915 9531 25964 9537
rect 25409 9503 25467 9509
rect 25409 9500 25421 9503
rect 21508 9472 25421 9500
rect 21508 9460 21514 9472
rect 25409 9469 25421 9472
rect 25455 9469 25467 9503
rect 25409 9463 25467 9469
rect 25501 9503 25559 9509
rect 25501 9469 25513 9503
rect 25547 9469 25559 9503
rect 25501 9463 25559 9469
rect 20579 9404 21404 9432
rect 25792 9432 25820 9531
rect 25958 9528 25964 9531
rect 26016 9528 26022 9580
rect 26150 9571 26208 9577
rect 26150 9537 26162 9571
rect 26196 9537 26208 9571
rect 26150 9531 26208 9537
rect 26165 9500 26193 9531
rect 26418 9528 26424 9580
rect 26476 9528 26482 9580
rect 26602 9528 26608 9580
rect 26660 9568 26666 9580
rect 27154 9568 27160 9580
rect 26660 9540 27160 9568
rect 26660 9528 26666 9540
rect 27154 9528 27160 9540
rect 27212 9568 27218 9580
rect 27341 9571 27399 9577
rect 27341 9568 27353 9571
rect 27212 9540 27353 9568
rect 27212 9528 27218 9540
rect 27341 9537 27353 9540
rect 27387 9537 27399 9571
rect 27341 9531 27399 9537
rect 27522 9528 27528 9580
rect 27580 9528 27586 9580
rect 26436 9500 26464 9528
rect 26878 9500 26884 9512
rect 26165 9472 26280 9500
rect 26436 9472 26884 9500
rect 25866 9432 25872 9444
rect 25792 9404 25872 9432
rect 20579 9401 20591 9404
rect 20533 9395 20591 9401
rect 25866 9392 25872 9404
rect 25924 9392 25930 9444
rect 26252 9432 26280 9472
rect 26878 9460 26884 9472
rect 26936 9500 26942 9512
rect 27433 9503 27491 9509
rect 27433 9500 27445 9503
rect 26936 9472 27445 9500
rect 26936 9460 26942 9472
rect 27433 9469 27445 9472
rect 27479 9469 27491 9503
rect 27540 9500 27568 9528
rect 27908 9512 27936 9608
rect 28000 9568 28028 9676
rect 30374 9664 30380 9716
rect 30432 9664 30438 9716
rect 31110 9664 31116 9716
rect 31168 9664 31174 9716
rect 32401 9707 32459 9713
rect 32401 9673 32413 9707
rect 32447 9704 32459 9707
rect 32674 9704 32680 9716
rect 32447 9676 32680 9704
rect 32447 9673 32459 9676
rect 32401 9667 32459 9673
rect 32674 9664 32680 9676
rect 32732 9664 32738 9716
rect 32858 9664 32864 9716
rect 32916 9704 32922 9716
rect 35250 9704 35256 9716
rect 32916 9676 35256 9704
rect 32916 9664 32922 9676
rect 35250 9664 35256 9676
rect 35308 9704 35314 9716
rect 38562 9704 38568 9716
rect 35308 9676 38568 9704
rect 35308 9664 35314 9676
rect 38562 9664 38568 9676
rect 38620 9664 38626 9716
rect 39206 9704 39212 9716
rect 38672 9676 39212 9704
rect 28905 9639 28963 9645
rect 28905 9605 28917 9639
rect 28951 9636 28963 9639
rect 29178 9636 29184 9648
rect 28951 9608 29184 9636
rect 28951 9605 28963 9608
rect 28905 9599 28963 9605
rect 29178 9596 29184 9608
rect 29236 9596 29242 9648
rect 29638 9596 29644 9648
rect 29696 9596 29702 9648
rect 28534 9568 28540 9580
rect 28000 9540 28540 9568
rect 28534 9528 28540 9540
rect 28592 9528 28598 9580
rect 28626 9528 28632 9580
rect 28684 9528 28690 9580
rect 30392 9568 30420 9664
rect 32217 9639 32275 9645
rect 32217 9605 32229 9639
rect 32263 9636 32275 9639
rect 32766 9636 32772 9648
rect 32263 9608 32772 9636
rect 32263 9605 32275 9608
rect 32217 9599 32275 9605
rect 32766 9596 32772 9608
rect 32824 9596 32830 9648
rect 36170 9596 36176 9648
rect 36228 9636 36234 9648
rect 37090 9636 37096 9648
rect 36228 9608 37096 9636
rect 36228 9596 36234 9608
rect 37090 9596 37096 9608
rect 37148 9596 37154 9648
rect 37182 9596 37188 9648
rect 37240 9636 37246 9648
rect 37277 9639 37335 9645
rect 37277 9636 37289 9639
rect 37240 9608 37289 9636
rect 37240 9596 37246 9608
rect 37277 9605 37289 9608
rect 37323 9636 37335 9639
rect 38672 9636 38700 9676
rect 39206 9664 39212 9676
rect 39264 9664 39270 9716
rect 39850 9664 39856 9716
rect 39908 9664 39914 9716
rect 37323 9608 38700 9636
rect 38948 9608 39804 9636
rect 37323 9605 37335 9608
rect 37277 9599 37335 9605
rect 30745 9571 30803 9577
rect 30745 9568 30757 9571
rect 30392 9540 30757 9568
rect 30745 9537 30757 9540
rect 30791 9537 30803 9571
rect 30745 9531 30803 9537
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9568 32551 9571
rect 32582 9568 32588 9580
rect 32539 9540 32588 9568
rect 32539 9537 32551 9540
rect 32493 9531 32551 9537
rect 32582 9528 32588 9540
rect 32640 9528 32646 9580
rect 37366 9568 37372 9580
rect 33152 9540 37372 9568
rect 27617 9503 27675 9509
rect 27617 9500 27629 9503
rect 27540 9472 27629 9500
rect 27433 9463 27491 9469
rect 27617 9469 27629 9472
rect 27663 9469 27675 9503
rect 27617 9463 27675 9469
rect 27890 9460 27896 9512
rect 27948 9460 27954 9512
rect 27982 9460 27988 9512
rect 28040 9460 28046 9512
rect 30650 9460 30656 9512
rect 30708 9460 30714 9512
rect 26165 9404 26280 9432
rect 26973 9435 27031 9441
rect 26165 9376 26193 9404
rect 26973 9401 26985 9435
rect 27019 9432 27031 9435
rect 28000 9432 28028 9460
rect 27019 9404 28028 9432
rect 27019 9401 27031 9404
rect 26973 9395 27031 9401
rect 33152 9376 33180 9540
rect 37366 9528 37372 9540
rect 37424 9568 37430 9580
rect 37461 9571 37519 9577
rect 37461 9568 37473 9571
rect 37424 9540 37473 9568
rect 37424 9528 37430 9540
rect 37461 9537 37473 9540
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 37737 9571 37795 9577
rect 37737 9537 37749 9571
rect 37783 9537 37795 9571
rect 37737 9531 37795 9537
rect 37752 9500 37780 9531
rect 37918 9528 37924 9580
rect 37976 9528 37982 9580
rect 38948 9577 38976 9608
rect 39408 9580 39436 9608
rect 38933 9571 38991 9577
rect 38933 9537 38945 9571
rect 38979 9537 38991 9571
rect 38933 9531 38991 9537
rect 39390 9528 39396 9580
rect 39448 9528 39454 9580
rect 39485 9571 39543 9577
rect 39485 9537 39497 9571
rect 39531 9537 39543 9571
rect 39485 9531 39543 9537
rect 38562 9500 38568 9512
rect 36464 9472 38568 9500
rect 36464 9376 36492 9472
rect 38562 9460 38568 9472
rect 38620 9500 38626 9512
rect 39117 9503 39175 9509
rect 39117 9500 39129 9503
rect 38620 9472 39129 9500
rect 38620 9460 38626 9472
rect 39117 9469 39129 9472
rect 39163 9469 39175 9503
rect 39117 9463 39175 9469
rect 37645 9435 37703 9441
rect 37645 9401 37657 9435
rect 37691 9432 37703 9435
rect 38654 9432 38660 9444
rect 37691 9404 38660 9432
rect 37691 9401 37703 9404
rect 37645 9395 37703 9401
rect 38654 9392 38660 9404
rect 38712 9392 38718 9444
rect 39500 9432 39528 9531
rect 39574 9528 39580 9580
rect 39632 9528 39638 9580
rect 39776 9577 39804 9608
rect 39761 9571 39819 9577
rect 39761 9537 39773 9571
rect 39807 9537 39819 9571
rect 39761 9531 39819 9537
rect 39945 9571 40003 9577
rect 39945 9537 39957 9571
rect 39991 9537 40003 9571
rect 39945 9531 40003 9537
rect 39592 9500 39620 9528
rect 39960 9500 39988 9531
rect 39592 9472 39988 9500
rect 39758 9432 39764 9444
rect 39500 9404 39764 9432
rect 39758 9392 39764 9404
rect 39816 9392 39822 9444
rect 15620 9336 17724 9364
rect 15620 9324 15626 9336
rect 18966 9324 18972 9376
rect 19024 9324 19030 9376
rect 19306 9336 19340 9376
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 21450 9324 21456 9376
rect 21508 9324 21514 9376
rect 22002 9324 22008 9376
rect 22060 9324 22066 9376
rect 26142 9324 26148 9376
rect 26200 9324 26206 9376
rect 26326 9324 26332 9376
rect 26384 9324 26390 9376
rect 26786 9324 26792 9376
rect 26844 9364 26850 9376
rect 28445 9367 28503 9373
rect 28445 9364 28457 9367
rect 26844 9336 28457 9364
rect 26844 9324 26850 9336
rect 28445 9333 28457 9336
rect 28491 9333 28503 9367
rect 28445 9327 28503 9333
rect 32214 9324 32220 9376
rect 32272 9324 32278 9376
rect 33134 9324 33140 9376
rect 33192 9324 33198 9376
rect 36446 9324 36452 9376
rect 36504 9324 36510 9376
rect 36906 9324 36912 9376
rect 36964 9364 36970 9376
rect 37829 9367 37887 9373
rect 37829 9364 37841 9367
rect 36964 9336 37841 9364
rect 36964 9324 36970 9336
rect 37829 9333 37841 9336
rect 37875 9333 37887 9367
rect 37829 9327 37887 9333
rect 1104 9274 41400 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 41400 9274
rect 1104 9200 41400 9222
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 4893 9163 4951 9169
rect 4893 9160 4905 9163
rect 4856 9132 4905 9160
rect 4856 9120 4862 9132
rect 4893 9129 4905 9132
rect 4939 9129 4951 9163
rect 4893 9123 4951 9129
rect 5442 9120 5448 9172
rect 5500 9120 5506 9172
rect 8570 9120 8576 9172
rect 8628 9120 8634 9172
rect 10962 9120 10968 9172
rect 11020 9120 11026 9172
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 13964 9132 14289 9160
rect 13964 9120 13970 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 15470 9120 15476 9172
rect 15528 9120 15534 9172
rect 17494 9120 17500 9172
rect 17552 9120 17558 9172
rect 19518 9120 19524 9172
rect 19576 9120 19582 9172
rect 22002 9160 22008 9172
rect 21928 9132 22008 9160
rect 4890 8984 4896 9036
rect 4948 8984 4954 9036
rect 5460 9024 5488 9120
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 9585 9095 9643 9101
rect 9585 9092 9597 9095
rect 8352 9064 9597 9092
rect 8352 9052 8358 9064
rect 9585 9061 9597 9064
rect 9631 9061 9643 9095
rect 10980 9092 11008 9120
rect 9585 9055 9643 9061
rect 10888 9064 11008 9092
rect 5460 8996 6684 9024
rect 4614 8916 4620 8968
rect 4672 8916 4678 8968
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 4908 8956 4936 8984
rect 4755 8928 4936 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 6546 8956 6552 8968
rect 6144 8928 6552 8956
rect 6144 8916 6150 8928
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6656 8965 6684 8996
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 8205 9027 8263 9033
rect 8205 9024 8217 9027
rect 7800 8996 8217 9024
rect 7800 8984 7806 8996
rect 8205 8993 8217 8996
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 9122 8984 9128 9036
rect 9180 8984 9186 9036
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 9306 9024 9312 9036
rect 9263 8996 9312 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9548 8996 10824 9024
rect 9548 8984 9554 8996
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 9140 8956 9168 8984
rect 8435 8928 9168 8956
rect 9401 8959 9459 8965
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9582 8956 9588 8968
rect 9447 8928 9588 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 10704 8888 10732 8919
rect 8536 8860 10732 8888
rect 10796 8888 10824 8996
rect 10888 8965 10916 9064
rect 10980 8996 11652 9024
rect 10980 8965 11008 8996
rect 11624 8968 11652 8996
rect 10854 8959 10916 8965
rect 10854 8925 10866 8959
rect 10900 8928 10916 8959
rect 10965 8959 11023 8965
rect 10900 8925 10912 8928
rect 10854 8919 10912 8925
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11072 8888 11100 8919
rect 11606 8916 11612 8968
rect 11664 8916 11670 8968
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8956 14519 8959
rect 15488 8956 15516 9120
rect 16853 9095 16911 9101
rect 16853 9061 16865 9095
rect 16899 9092 16911 9095
rect 19978 9092 19984 9104
rect 16899 9064 19984 9092
rect 16899 9061 16911 9064
rect 16853 9055 16911 9061
rect 19978 9052 19984 9064
rect 20036 9052 20042 9104
rect 16758 9024 16764 9036
rect 16316 8996 16764 9024
rect 14507 8928 15516 8956
rect 14507 8925 14519 8928
rect 14461 8919 14519 8925
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 16316 8965 16344 8996
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 17954 8984 17960 9036
rect 18012 9024 18018 9036
rect 20533 9027 20591 9033
rect 20533 9024 20545 9027
rect 18012 8996 20545 9024
rect 18012 8984 18018 8996
rect 20533 8993 20545 8996
rect 20579 8993 20591 9027
rect 20533 8987 20591 8993
rect 20809 9027 20867 9033
rect 20809 8993 20821 9027
rect 20855 9024 20867 9027
rect 21450 9024 21456 9036
rect 20855 8996 21456 9024
rect 20855 8993 20867 8996
rect 20809 8987 20867 8993
rect 21450 8984 21456 8996
rect 21508 8984 21514 9036
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 16264 8928 16313 8956
rect 16264 8916 16270 8928
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 16301 8919 16359 8925
rect 16482 8916 16488 8968
rect 16540 8916 16546 8968
rect 16574 8916 16580 8968
rect 16632 8916 16638 8968
rect 16669 8959 16727 8965
rect 16669 8925 16681 8959
rect 16715 8956 16727 8959
rect 16850 8956 16856 8968
rect 16715 8928 16856 8956
rect 16715 8925 16727 8928
rect 16669 8919 16727 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 16945 8959 17003 8965
rect 16945 8925 16957 8959
rect 16991 8925 17003 8959
rect 16945 8919 17003 8925
rect 16960 8888 16988 8919
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 17092 8928 17325 8956
rect 17092 8916 17098 8928
rect 17313 8925 17325 8928
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 18601 8959 18659 8965
rect 18601 8925 18613 8959
rect 18647 8956 18659 8959
rect 18966 8956 18972 8968
rect 18647 8928 18972 8956
rect 18647 8925 18659 8928
rect 18601 8919 18659 8925
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 19426 8916 19432 8968
rect 19484 8916 19490 8968
rect 21928 8956 21956 9132
rect 22002 9120 22008 9132
rect 22060 9120 22066 9172
rect 22281 9163 22339 9169
rect 22281 9129 22293 9163
rect 22327 9160 22339 9163
rect 22462 9160 22468 9172
rect 22327 9132 22468 9160
rect 22327 9129 22339 9132
rect 22281 9123 22339 9129
rect 22462 9120 22468 9132
rect 22520 9120 22526 9172
rect 23106 9120 23112 9172
rect 23164 9160 23170 9172
rect 26694 9160 26700 9172
rect 23164 9132 26700 9160
rect 23164 9120 23170 9132
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 26804 9132 27016 9160
rect 25590 9052 25596 9104
rect 25648 9092 25654 9104
rect 26804 9092 26832 9132
rect 25648 9064 26832 9092
rect 25648 9052 25654 9064
rect 26988 9036 27016 9132
rect 27614 9120 27620 9172
rect 27672 9160 27678 9172
rect 28626 9160 28632 9172
rect 27672 9132 28632 9160
rect 27672 9120 27678 9132
rect 28626 9120 28632 9132
rect 28684 9120 28690 9172
rect 34241 9163 34299 9169
rect 34241 9129 34253 9163
rect 34287 9160 34299 9163
rect 34287 9132 34468 9160
rect 34287 9129 34299 9132
rect 34241 9123 34299 9129
rect 28534 9052 28540 9104
rect 28592 9092 28598 9104
rect 28592 9064 31754 9092
rect 28592 9052 28598 9064
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 22060 8996 26740 9024
rect 22060 8984 22066 8996
rect 23750 8956 23756 8968
rect 21928 8942 23756 8956
rect 21942 8928 23756 8942
rect 23750 8916 23756 8928
rect 23808 8916 23814 8968
rect 25314 8916 25320 8968
rect 25372 8956 25378 8968
rect 26326 8956 26332 8968
rect 25372 8928 26332 8956
rect 25372 8916 25378 8928
rect 26326 8916 26332 8928
rect 26384 8916 26390 8968
rect 10796 8860 11100 8888
rect 16592 8860 16988 8888
rect 8536 8848 8542 8860
rect 16592 8832 16620 8860
rect 17126 8848 17132 8900
rect 17184 8848 17190 8900
rect 17221 8891 17279 8897
rect 17221 8857 17233 8891
rect 17267 8857 17279 8891
rect 26712 8888 26740 8996
rect 26878 8984 26884 9036
rect 26936 8984 26942 9036
rect 26970 8984 26976 9036
rect 27028 8984 27034 9036
rect 27154 8984 27160 9036
rect 27212 9024 27218 9036
rect 28997 9027 29055 9033
rect 28997 9024 29009 9027
rect 27212 8996 29009 9024
rect 27212 8984 27218 8996
rect 28997 8993 29009 8996
rect 29043 8993 29055 9027
rect 31726 9024 31754 9064
rect 32306 9052 32312 9104
rect 32364 9092 32370 9104
rect 33870 9092 33876 9104
rect 32364 9064 33876 9092
rect 32364 9052 32370 9064
rect 33870 9052 33876 9064
rect 33928 9092 33934 9104
rect 33928 9064 34376 9092
rect 33928 9052 33934 9064
rect 33134 9024 33140 9036
rect 31726 8996 33140 9024
rect 28997 8987 29055 8993
rect 33134 8984 33140 8996
rect 33192 8984 33198 9036
rect 26786 8916 26792 8968
rect 26844 8916 26850 8968
rect 27249 8959 27307 8965
rect 27249 8925 27261 8959
rect 27295 8925 27307 8959
rect 27249 8919 27307 8925
rect 27264 8888 27292 8919
rect 28626 8916 28632 8968
rect 28684 8956 28690 8968
rect 29638 8956 29644 8968
rect 28684 8928 29644 8956
rect 28684 8916 28690 8928
rect 29638 8916 29644 8928
rect 29696 8916 29702 8968
rect 30282 8916 30288 8968
rect 30340 8956 30346 8968
rect 31662 8956 31668 8968
rect 30340 8928 31668 8956
rect 30340 8916 30346 8928
rect 31662 8916 31668 8928
rect 31720 8956 31726 8968
rect 33226 8956 33232 8968
rect 31720 8928 33232 8956
rect 31720 8916 31726 8928
rect 27430 8888 27436 8900
rect 26712 8860 26832 8888
rect 27264 8860 27436 8888
rect 17221 8851 17279 8857
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8820 6331 8823
rect 7650 8820 7656 8832
rect 6319 8792 7656 8820
rect 6319 8789 6331 8792
rect 6273 8783 6331 8789
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10505 8823 10563 8829
rect 10505 8820 10517 8823
rect 10284 8792 10517 8820
rect 10284 8780 10290 8792
rect 10505 8789 10517 8792
rect 10551 8789 10563 8823
rect 10505 8783 10563 8789
rect 14090 8780 14096 8832
rect 14148 8820 14154 8832
rect 15010 8820 15016 8832
rect 14148 8792 15016 8820
rect 14148 8780 14154 8792
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 16574 8780 16580 8832
rect 16632 8780 16638 8832
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 17236 8820 17264 8851
rect 16816 8792 17264 8820
rect 16816 8780 16822 8792
rect 18414 8780 18420 8832
rect 18472 8820 18478 8832
rect 18693 8823 18751 8829
rect 18693 8820 18705 8823
rect 18472 8792 18705 8820
rect 18472 8780 18478 8792
rect 18693 8789 18705 8792
rect 18739 8789 18751 8823
rect 18693 8783 18751 8789
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 25130 8820 25136 8832
rect 23532 8792 25136 8820
rect 23532 8780 23538 8792
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 26418 8780 26424 8832
rect 26476 8780 26482 8832
rect 26804 8820 26832 8860
rect 27430 8848 27436 8860
rect 27488 8848 27494 8900
rect 27525 8891 27583 8897
rect 27525 8857 27537 8891
rect 27571 8888 27583 8891
rect 27798 8888 27804 8900
rect 27571 8860 27804 8888
rect 27571 8857 27583 8860
rect 27525 8851 27583 8857
rect 27798 8848 27804 8860
rect 27856 8848 27862 8900
rect 31754 8888 31760 8900
rect 28828 8860 31760 8888
rect 28828 8820 28856 8860
rect 31754 8848 31760 8860
rect 31812 8848 31818 8900
rect 32968 8897 32996 8928
rect 33226 8916 33232 8928
rect 33284 8956 33290 8968
rect 34348 8965 34376 9064
rect 34440 9024 34468 9132
rect 34514 9120 34520 9172
rect 34572 9160 34578 9172
rect 38749 9163 38807 9169
rect 38749 9160 38761 9163
rect 34572 9132 38761 9160
rect 34572 9120 34578 9132
rect 38749 9129 38761 9132
rect 38795 9129 38807 9163
rect 38749 9123 38807 9129
rect 39209 9095 39267 9101
rect 39209 9092 39221 9095
rect 36556 9064 37780 9092
rect 34440 8996 34744 9024
rect 34149 8959 34207 8965
rect 34149 8956 34161 8959
rect 33284 8928 33640 8956
rect 33284 8916 33290 8928
rect 33612 8900 33640 8928
rect 33704 8928 34161 8956
rect 32953 8891 33011 8897
rect 32953 8857 32965 8891
rect 32999 8857 33011 8891
rect 32953 8851 33011 8857
rect 33594 8848 33600 8900
rect 33652 8848 33658 8900
rect 26804 8792 28856 8820
rect 31110 8780 31116 8832
rect 31168 8820 31174 8832
rect 33042 8820 33048 8832
rect 31168 8792 33048 8820
rect 31168 8780 31174 8792
rect 33042 8780 33048 8792
rect 33100 8820 33106 8832
rect 33704 8820 33732 8928
rect 34149 8925 34161 8928
rect 34195 8925 34207 8959
rect 34149 8919 34207 8925
rect 34333 8959 34391 8965
rect 34333 8925 34345 8959
rect 34379 8956 34391 8959
rect 34606 8956 34612 8968
rect 34379 8928 34612 8956
rect 34379 8925 34391 8928
rect 34333 8919 34391 8925
rect 34606 8916 34612 8928
rect 34664 8916 34670 8968
rect 34716 8965 34744 8996
rect 35820 8996 36308 9024
rect 35820 8968 35848 8996
rect 34701 8959 34759 8965
rect 34701 8925 34713 8959
rect 34747 8925 34759 8959
rect 34701 8919 34759 8925
rect 34885 8959 34943 8965
rect 34885 8925 34897 8959
rect 34931 8925 34943 8959
rect 34885 8919 34943 8925
rect 34054 8848 34060 8900
rect 34112 8888 34118 8900
rect 34900 8888 34928 8919
rect 35802 8916 35808 8968
rect 35860 8916 35866 8968
rect 36078 8916 36084 8968
rect 36136 8916 36142 8968
rect 36280 8965 36308 8996
rect 36446 8984 36452 9036
rect 36504 8984 36510 9036
rect 36556 9033 36584 9064
rect 36541 9027 36599 9033
rect 36541 8993 36553 9027
rect 36587 8993 36599 9027
rect 36541 8987 36599 8993
rect 36906 8984 36912 9036
rect 36964 8984 36970 9036
rect 36265 8959 36323 8965
rect 36265 8925 36277 8959
rect 36311 8925 36323 8959
rect 36265 8919 36323 8925
rect 36633 8959 36691 8965
rect 36633 8925 36645 8959
rect 36679 8925 36691 8959
rect 36633 8919 36691 8925
rect 36726 8959 36784 8965
rect 36726 8925 36738 8959
rect 36772 8925 36784 8959
rect 36726 8919 36784 8925
rect 34112 8860 34928 8888
rect 36096 8888 36124 8916
rect 36648 8888 36676 8919
rect 36096 8860 36676 8888
rect 34112 8848 34118 8860
rect 33100 8792 33732 8820
rect 33100 8780 33106 8792
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 34793 8823 34851 8829
rect 34793 8820 34805 8823
rect 34572 8792 34805 8820
rect 34572 8780 34578 8792
rect 34793 8789 34805 8792
rect 34839 8789 34851 8823
rect 34793 8783 34851 8789
rect 36081 8823 36139 8829
rect 36081 8789 36093 8823
rect 36127 8820 36139 8823
rect 36740 8820 36768 8919
rect 36924 8897 36952 8984
rect 37090 8916 37096 8968
rect 37148 8965 37154 8968
rect 37148 8956 37156 8965
rect 37148 8928 37193 8956
rect 37148 8919 37156 8928
rect 37148 8916 37154 8919
rect 37366 8916 37372 8968
rect 37424 8916 37430 8968
rect 37752 8956 37780 9064
rect 38488 9064 39221 9092
rect 37918 8956 37924 8968
rect 37752 8928 37924 8956
rect 37918 8916 37924 8928
rect 37976 8956 37982 8968
rect 38488 8965 38516 9064
rect 39209 9061 39221 9064
rect 39255 9061 39267 9095
rect 39209 9055 39267 9061
rect 38562 8984 38568 9036
rect 38620 8984 38626 9036
rect 38654 8984 38660 9036
rect 38712 9024 38718 9036
rect 38712 8996 39068 9024
rect 38712 8984 38718 8996
rect 39040 8965 39068 8996
rect 38473 8959 38531 8965
rect 38473 8956 38485 8959
rect 37976 8928 38485 8956
rect 37976 8916 37982 8928
rect 38473 8925 38485 8928
rect 38519 8925 38531 8959
rect 38473 8919 38531 8925
rect 38841 8959 38899 8965
rect 38841 8925 38853 8959
rect 38887 8925 38899 8959
rect 38841 8919 38899 8925
rect 39025 8959 39083 8965
rect 39025 8925 39037 8959
rect 39071 8925 39083 8959
rect 39025 8919 39083 8925
rect 36909 8891 36967 8897
rect 36909 8857 36921 8891
rect 36955 8857 36967 8891
rect 36909 8851 36967 8857
rect 37001 8891 37059 8897
rect 37001 8857 37013 8891
rect 37047 8888 37059 8891
rect 38013 8891 38071 8897
rect 38013 8888 38025 8891
rect 37047 8860 38025 8888
rect 37047 8857 37059 8860
rect 37001 8851 37059 8857
rect 38013 8857 38025 8860
rect 38059 8857 38071 8891
rect 38856 8888 38884 8919
rect 38013 8851 38071 8857
rect 38120 8860 38884 8888
rect 36127 8792 36768 8820
rect 36127 8789 36139 8792
rect 36081 8783 36139 8789
rect 37274 8780 37280 8832
rect 37332 8780 37338 8832
rect 37458 8780 37464 8832
rect 37516 8820 37522 8832
rect 38120 8829 38148 8860
rect 38105 8823 38163 8829
rect 38105 8820 38117 8823
rect 37516 8792 38117 8820
rect 37516 8780 37522 8792
rect 38105 8789 38117 8792
rect 38151 8789 38163 8823
rect 38105 8783 38163 8789
rect 1104 8730 41400 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 41400 8730
rect 1104 8656 41400 8678
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 3878 8616 3884 8628
rect 3835 8588 3884 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 10042 8616 10048 8628
rect 4948 8588 10048 8616
rect 4948 8576 4954 8588
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10410 8576 10416 8628
rect 10468 8576 10474 8628
rect 10520 8588 14228 8616
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 10428 8548 10456 8576
rect 4672 8520 6776 8548
rect 4672 8508 4678 8520
rect 6748 8489 6776 8520
rect 6886 8520 10456 8548
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 4203 8452 5549 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 6886 8480 6914 8520
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 6779 8452 6914 8480
rect 7116 8452 8861 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4985 8415 5043 8421
rect 4295 8384 4936 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4614 8276 4620 8288
rect 4479 8248 4620 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 4908 8276 4936 8384
rect 4985 8381 4997 8415
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 5000 8344 5028 8375
rect 6546 8372 6552 8424
rect 6604 8412 6610 8424
rect 7116 8421 7144 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6604 8384 6653 8412
rect 6604 8372 6610 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 9048 8412 9076 8443
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 10520 8480 10548 8588
rect 13722 8548 13728 8560
rect 13570 8520 13728 8548
rect 13722 8508 13728 8520
rect 13780 8548 13786 8560
rect 14090 8548 14096 8560
rect 13780 8520 14096 8548
rect 13780 8508 13786 8520
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 14200 8548 14228 8588
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 15105 8619 15163 8625
rect 15105 8616 15117 8619
rect 14332 8588 15117 8616
rect 14332 8576 14338 8588
rect 15105 8585 15117 8588
rect 15151 8585 15163 8619
rect 15105 8579 15163 8585
rect 15286 8576 15292 8628
rect 15344 8616 15350 8628
rect 17126 8616 17132 8628
rect 15344 8588 17132 8616
rect 15344 8576 15350 8588
rect 16574 8548 16580 8560
rect 14200 8520 16580 8548
rect 16574 8508 16580 8520
rect 16632 8508 16638 8560
rect 16960 8557 16988 8588
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 18414 8616 18420 8628
rect 18248 8588 18420 8616
rect 16945 8551 17003 8557
rect 16684 8520 16896 8548
rect 9456 8452 10548 8480
rect 9456 8440 9462 8452
rect 14550 8440 14556 8492
rect 14608 8440 14614 8492
rect 14734 8440 14740 8492
rect 14792 8440 14798 8492
rect 14826 8440 14832 8492
rect 14884 8440 14890 8492
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8480 14979 8483
rect 15010 8480 15016 8492
rect 14967 8452 15016 8480
rect 14967 8449 14979 8452
rect 14921 8443 14979 8449
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 16206 8440 16212 8492
rect 16264 8440 16270 8492
rect 16684 8489 16712 8520
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 16762 8483 16820 8489
rect 16762 8449 16774 8483
rect 16808 8449 16820 8483
rect 16762 8443 16820 8449
rect 9490 8412 9496 8424
rect 8260 8384 9496 8412
rect 8260 8372 8266 8384
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10594 8412 10600 8424
rect 9732 8384 10600 8412
rect 9732 8372 9738 8384
rect 10594 8372 10600 8384
rect 10652 8412 10658 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 10652 8384 12081 8412
rect 10652 8372 10658 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8412 12403 8415
rect 12434 8412 12440 8424
rect 12391 8384 12440 8412
rect 12391 8381 12403 8384
rect 12345 8375 12403 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 16224 8412 16252 8440
rect 13872 8384 16252 8412
rect 13872 8372 13878 8384
rect 5534 8344 5540 8356
rect 5000 8316 5540 8344
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 8941 8347 8999 8353
rect 8941 8313 8953 8347
rect 8987 8344 8999 8347
rect 10042 8344 10048 8356
rect 8987 8316 10048 8344
rect 8987 8313 8999 8316
rect 8941 8307 8999 8313
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 13740 8316 13952 8344
rect 5718 8276 5724 8288
rect 4908 8248 5724 8276
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 13740 8276 13768 8316
rect 7984 8248 13768 8276
rect 13924 8276 13952 8316
rect 16776 8276 16804 8443
rect 16868 8344 16896 8520
rect 16945 8517 16957 8551
rect 16991 8517 17003 8551
rect 16945 8511 17003 8517
rect 17037 8551 17095 8557
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 17310 8548 17316 8560
rect 17083 8520 17316 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 18248 8557 18276 8588
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 20162 8576 20168 8628
rect 20220 8576 20226 8628
rect 22097 8619 22155 8625
rect 22097 8585 22109 8619
rect 22143 8585 22155 8619
rect 22097 8579 22155 8585
rect 18233 8551 18291 8557
rect 18233 8517 18245 8551
rect 18279 8517 18291 8551
rect 20180 8548 20208 8576
rect 18233 8511 18291 8517
rect 19812 8520 20208 8548
rect 22112 8548 22140 8579
rect 23290 8576 23296 8628
rect 23348 8616 23354 8628
rect 24118 8616 24124 8628
rect 23348 8588 24124 8616
rect 23348 8576 23354 8588
rect 24118 8576 24124 8588
rect 24176 8576 24182 8628
rect 26418 8576 26424 8628
rect 26476 8576 26482 8628
rect 27614 8576 27620 8628
rect 27672 8576 27678 8628
rect 27890 8576 27896 8628
rect 27948 8616 27954 8628
rect 29089 8619 29147 8625
rect 29089 8616 29101 8619
rect 27948 8588 29101 8616
rect 27948 8576 27954 8588
rect 29089 8585 29101 8588
rect 29135 8585 29147 8619
rect 29089 8579 29147 8585
rect 30561 8619 30619 8625
rect 30561 8585 30573 8619
rect 30607 8616 30619 8619
rect 30650 8616 30656 8628
rect 30607 8588 30656 8616
rect 30607 8585 30619 8588
rect 30561 8579 30619 8585
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 31386 8576 31392 8628
rect 31444 8616 31450 8628
rect 31665 8619 31723 8625
rect 31665 8616 31677 8619
rect 31444 8588 31677 8616
rect 31444 8576 31450 8588
rect 31665 8585 31677 8588
rect 31711 8585 31723 8619
rect 31665 8579 31723 8585
rect 32214 8576 32220 8628
rect 32272 8576 32278 8628
rect 32324 8588 33824 8616
rect 22649 8551 22707 8557
rect 22649 8548 22661 8551
rect 22112 8520 22661 8548
rect 17134 8483 17192 8489
rect 17134 8480 17146 8483
rect 17052 8452 17146 8480
rect 17052 8424 17080 8452
rect 17134 8449 17146 8452
rect 17180 8449 17192 8483
rect 17134 8443 17192 8449
rect 17954 8440 17960 8492
rect 18012 8440 18018 8492
rect 19334 8440 19340 8492
rect 19392 8440 19398 8492
rect 19812 8489 19840 8520
rect 22649 8517 22661 8520
rect 22695 8517 22707 8551
rect 22649 8511 22707 8517
rect 25225 8551 25283 8557
rect 25225 8517 25237 8551
rect 25271 8548 25283 8551
rect 25498 8548 25504 8560
rect 25271 8520 25504 8548
rect 25271 8517 25283 8520
rect 25225 8511 25283 8517
rect 25498 8508 25504 8520
rect 25556 8508 25562 8560
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 19945 8483 20003 8489
rect 19945 8449 19957 8483
rect 19991 8480 20003 8483
rect 19991 8449 20024 8480
rect 19945 8443 20024 8449
rect 17034 8372 17040 8424
rect 17092 8372 17098 8424
rect 18690 8412 18696 8424
rect 17328 8384 18696 8412
rect 16942 8344 16948 8356
rect 16868 8316 16948 8344
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 17328 8353 17356 8384
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 17313 8347 17371 8353
rect 17313 8313 17325 8347
rect 17359 8313 17371 8347
rect 19352 8344 19380 8440
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 19705 8415 19763 8421
rect 19705 8412 19717 8415
rect 19484 8384 19717 8412
rect 19484 8372 19490 8384
rect 19705 8381 19717 8384
rect 19751 8381 19763 8415
rect 19705 8375 19763 8381
rect 19886 8344 19892 8356
rect 19352 8316 19892 8344
rect 17313 8307 17371 8313
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 19996 8344 20024 8443
rect 20070 8440 20076 8492
rect 20128 8440 20134 8492
rect 20162 8440 20168 8492
rect 20220 8440 20226 8492
rect 20346 8489 20352 8492
rect 20303 8483 20352 8489
rect 20303 8449 20315 8483
rect 20349 8449 20352 8483
rect 20303 8443 20352 8449
rect 20346 8440 20352 8443
rect 20404 8480 20410 8492
rect 21542 8480 21548 8492
rect 20404 8452 21548 8480
rect 20404 8440 20410 8452
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 22281 8483 22339 8489
rect 22281 8480 22293 8483
rect 22244 8452 22293 8480
rect 22244 8440 22250 8452
rect 22281 8449 22293 8452
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 23750 8440 23756 8492
rect 23808 8440 23814 8492
rect 24946 8440 24952 8492
rect 25004 8440 25010 8492
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8480 25191 8483
rect 26436 8480 26464 8576
rect 27632 8548 27660 8576
rect 27356 8520 27660 8548
rect 27356 8489 27384 8520
rect 28626 8508 28632 8560
rect 28684 8508 28690 8560
rect 30098 8508 30104 8560
rect 30156 8548 30162 8560
rect 30156 8520 30972 8548
rect 30156 8508 30162 8520
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 25179 8452 25268 8480
rect 26436 8452 27169 8480
rect 25179 8449 25191 8452
rect 25133 8443 25191 8449
rect 20088 8412 20116 8440
rect 21174 8412 21180 8424
rect 20088 8384 21180 8412
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 22373 8415 22431 8421
rect 22373 8381 22385 8415
rect 22419 8381 22431 8415
rect 23768 8412 23796 8440
rect 25240 8424 25268 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 23768 8384 24532 8412
rect 22373 8375 22431 8381
rect 19996 8316 22094 8344
rect 17402 8276 17408 8288
rect 13924 8248 17408 8276
rect 7984 8236 7990 8248
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 19702 8236 19708 8288
rect 19760 8276 19766 8288
rect 20441 8279 20499 8285
rect 20441 8276 20453 8279
rect 19760 8248 20453 8276
rect 19760 8236 19766 8248
rect 20441 8245 20453 8248
rect 20487 8245 20499 8279
rect 22066 8276 22094 8316
rect 22278 8304 22284 8356
rect 22336 8344 22342 8356
rect 22388 8344 22416 8375
rect 24504 8356 24532 8384
rect 25222 8372 25228 8424
rect 25280 8372 25286 8424
rect 27617 8415 27675 8421
rect 27617 8412 27629 8415
rect 26988 8384 27629 8412
rect 22336 8316 22416 8344
rect 22336 8304 22342 8316
rect 24486 8304 24492 8356
rect 24544 8344 24550 8356
rect 26988 8353 27016 8384
rect 27617 8381 27629 8384
rect 27663 8381 27675 8415
rect 27617 8375 27675 8381
rect 26973 8347 27031 8353
rect 24544 8316 26924 8344
rect 24544 8304 24550 8316
rect 23290 8276 23296 8288
rect 22066 8248 23296 8276
rect 20441 8239 20499 8245
rect 23290 8236 23296 8248
rect 23348 8236 23354 8288
rect 26896 8276 26924 8316
rect 26973 8313 26985 8347
rect 27019 8313 27031 8347
rect 26973 8307 27031 8313
rect 28644 8276 28672 8508
rect 30282 8440 30288 8492
rect 30340 8440 30346 8492
rect 30484 8489 30512 8520
rect 30469 8483 30527 8489
rect 30469 8449 30481 8483
rect 30515 8449 30527 8483
rect 30469 8443 30527 8449
rect 30745 8483 30803 8489
rect 30745 8449 30757 8483
rect 30791 8449 30803 8483
rect 30944 8480 30972 8520
rect 31110 8508 31116 8560
rect 31168 8508 31174 8560
rect 32232 8548 32260 8576
rect 32140 8520 32260 8548
rect 31297 8483 31355 8489
rect 31297 8480 31309 8483
rect 30944 8478 31156 8480
rect 31220 8478 31309 8480
rect 30944 8452 31309 8478
rect 31128 8450 31248 8452
rect 30745 8443 30803 8449
rect 31297 8449 31309 8452
rect 31343 8480 31355 8483
rect 31573 8483 31631 8489
rect 31343 8452 31524 8480
rect 31343 8449 31355 8452
rect 31297 8443 31355 8449
rect 30377 8415 30435 8421
rect 30377 8381 30389 8415
rect 30423 8412 30435 8415
rect 30558 8412 30564 8424
rect 30423 8384 30564 8412
rect 30423 8381 30435 8384
rect 30377 8375 30435 8381
rect 30558 8372 30564 8384
rect 30616 8412 30622 8424
rect 30760 8412 30788 8443
rect 30616 8384 30788 8412
rect 31021 8415 31079 8421
rect 30616 8372 30622 8384
rect 31021 8381 31033 8415
rect 31067 8412 31079 8415
rect 31496 8412 31524 8452
rect 31573 8449 31585 8483
rect 31619 8480 31631 8483
rect 31662 8480 31668 8492
rect 31619 8452 31668 8480
rect 31619 8449 31631 8452
rect 31573 8443 31631 8449
rect 31662 8440 31668 8452
rect 31720 8440 31726 8492
rect 32140 8489 32168 8520
rect 32324 8489 32352 8588
rect 32493 8551 32551 8557
rect 32493 8517 32505 8551
rect 32539 8548 32551 8551
rect 33505 8551 33563 8557
rect 33505 8548 33517 8551
rect 32539 8520 33517 8548
rect 32539 8517 32551 8520
rect 32493 8511 32551 8517
rect 33505 8517 33517 8520
rect 33551 8517 33563 8551
rect 33505 8511 33563 8517
rect 33594 8508 33600 8560
rect 33652 8548 33658 8560
rect 33689 8551 33747 8557
rect 33689 8548 33701 8551
rect 33652 8520 33701 8548
rect 33652 8508 33658 8520
rect 33689 8517 33701 8520
rect 33735 8517 33747 8551
rect 33796 8548 33824 8588
rect 34054 8576 34060 8628
rect 34112 8576 34118 8628
rect 35802 8616 35808 8628
rect 34164 8588 35808 8616
rect 34164 8548 34192 8588
rect 34514 8548 34520 8560
rect 33796 8520 34192 8548
rect 34348 8520 34520 8548
rect 33689 8511 33747 8517
rect 31769 8483 31827 8489
rect 31769 8449 31781 8483
rect 31815 8480 31827 8483
rect 32125 8483 32183 8489
rect 31815 8452 31892 8480
rect 31815 8449 31827 8452
rect 31769 8443 31827 8449
rect 31067 8384 31248 8412
rect 31496 8384 31708 8412
rect 31067 8381 31079 8384
rect 31021 8375 31079 8381
rect 26896 8248 28672 8276
rect 30929 8279 30987 8285
rect 30929 8245 30941 8279
rect 30975 8276 30987 8279
rect 31110 8276 31116 8288
rect 30975 8248 31116 8276
rect 30975 8245 30987 8248
rect 30929 8239 30987 8245
rect 31110 8236 31116 8248
rect 31168 8236 31174 8288
rect 31220 8276 31248 8384
rect 31680 8344 31708 8384
rect 31864 8344 31892 8452
rect 32125 8449 32137 8483
rect 32171 8449 32183 8483
rect 32125 8443 32183 8449
rect 32273 8483 32352 8489
rect 32273 8449 32285 8483
rect 32319 8452 32352 8483
rect 32401 8483 32459 8489
rect 32319 8449 32331 8452
rect 32273 8443 32331 8449
rect 32401 8449 32413 8483
rect 32447 8449 32459 8483
rect 32401 8443 32459 8449
rect 32631 8483 32689 8489
rect 32631 8449 32643 8483
rect 32677 8480 32689 8483
rect 32677 8452 33824 8480
rect 32677 8449 32689 8452
rect 32631 8443 32689 8449
rect 32030 8372 32036 8424
rect 32088 8412 32094 8424
rect 32416 8412 32444 8443
rect 32088 8384 32444 8412
rect 32861 8415 32919 8421
rect 32088 8372 32094 8384
rect 32861 8381 32873 8415
rect 32907 8381 32919 8415
rect 33796 8412 33824 8452
rect 33870 8440 33876 8492
rect 33928 8440 33934 8492
rect 34348 8489 34376 8520
rect 34514 8508 34520 8520
rect 34572 8508 34578 8560
rect 34333 8483 34391 8489
rect 34333 8449 34345 8483
rect 34379 8449 34391 8483
rect 34333 8443 34391 8449
rect 34422 8440 34428 8492
rect 34480 8440 34486 8492
rect 34698 8440 34704 8492
rect 34756 8480 34762 8492
rect 34992 8489 35020 8588
rect 35802 8576 35808 8588
rect 35860 8576 35866 8628
rect 37182 8616 37188 8628
rect 36832 8588 37188 8616
rect 35161 8551 35219 8557
rect 35161 8517 35173 8551
rect 35207 8548 35219 8551
rect 36173 8551 36231 8557
rect 36173 8548 36185 8551
rect 35207 8520 36185 8548
rect 35207 8517 35219 8520
rect 35161 8511 35219 8517
rect 36173 8517 36185 8520
rect 36219 8517 36231 8551
rect 36173 8511 36231 8517
rect 36832 8489 36860 8588
rect 37182 8576 37188 8588
rect 37240 8576 37246 8628
rect 37274 8576 37280 8628
rect 37332 8616 37338 8628
rect 37332 8588 37596 8616
rect 37332 8576 37338 8588
rect 36909 8551 36967 8557
rect 36909 8517 36921 8551
rect 36955 8548 36967 8551
rect 37458 8548 37464 8560
rect 36955 8520 37464 8548
rect 36955 8517 36967 8520
rect 36909 8511 36967 8517
rect 37458 8508 37464 8520
rect 37516 8508 37522 8560
rect 37568 8557 37596 8588
rect 37660 8588 39344 8616
rect 37660 8560 37688 8588
rect 37553 8551 37611 8557
rect 37553 8517 37565 8551
rect 37599 8517 37611 8551
rect 37553 8511 37611 8517
rect 37642 8508 37648 8560
rect 37700 8508 37706 8560
rect 38838 8548 38844 8560
rect 38778 8520 38844 8548
rect 38838 8508 38844 8520
rect 38896 8508 38902 8560
rect 39316 8557 39344 8588
rect 39301 8551 39359 8557
rect 39301 8517 39313 8551
rect 39347 8517 39359 8551
rect 39301 8511 39359 8517
rect 34793 8483 34851 8489
rect 34793 8480 34805 8483
rect 34756 8452 34805 8480
rect 34756 8440 34762 8452
rect 34793 8449 34805 8452
rect 34839 8449 34851 8483
rect 34793 8443 34851 8449
rect 34941 8483 35020 8489
rect 34941 8449 34953 8483
rect 34987 8452 35020 8483
rect 35069 8483 35127 8489
rect 34987 8449 34999 8452
rect 34941 8443 34999 8449
rect 35069 8449 35081 8483
rect 35115 8449 35127 8483
rect 35299 8483 35357 8489
rect 35299 8480 35311 8483
rect 35069 8443 35127 8449
rect 35176 8452 35311 8480
rect 34241 8415 34299 8421
rect 33796 8384 33916 8412
rect 32861 8375 32919 8381
rect 32876 8344 32904 8375
rect 33686 8344 33692 8356
rect 31680 8316 33692 8344
rect 33686 8304 33692 8316
rect 33744 8304 33750 8356
rect 33888 8344 33916 8384
rect 34241 8381 34253 8415
rect 34287 8412 34299 8415
rect 34440 8412 34468 8440
rect 34287 8384 34468 8412
rect 34287 8381 34299 8384
rect 34241 8375 34299 8381
rect 34701 8347 34759 8353
rect 33888 8316 34652 8344
rect 31386 8276 31392 8288
rect 31220 8248 31392 8276
rect 31386 8236 31392 8248
rect 31444 8236 31450 8288
rect 31478 8236 31484 8288
rect 31536 8236 31542 8288
rect 32214 8236 32220 8288
rect 32272 8276 32278 8288
rect 32769 8279 32827 8285
rect 32769 8276 32781 8279
rect 32272 8248 32781 8276
rect 32272 8236 32278 8248
rect 32769 8245 32781 8248
rect 32815 8245 32827 8279
rect 34624 8276 34652 8316
rect 34701 8313 34713 8347
rect 34747 8344 34759 8347
rect 35084 8344 35112 8443
rect 34747 8316 35112 8344
rect 34747 8313 34759 8316
rect 34701 8307 34759 8313
rect 35176 8276 35204 8452
rect 35299 8449 35311 8452
rect 35345 8480 35357 8483
rect 36817 8483 36875 8489
rect 35345 8452 36216 8480
rect 35345 8449 35357 8452
rect 35299 8443 35357 8449
rect 36188 8424 36216 8452
rect 36817 8449 36829 8483
rect 36863 8449 36875 8483
rect 36817 8443 36875 8449
rect 37001 8483 37059 8489
rect 37001 8449 37013 8483
rect 37047 8480 37059 8483
rect 37182 8480 37188 8492
rect 37047 8452 37188 8480
rect 37047 8449 37059 8452
rect 37001 8443 37059 8449
rect 37182 8440 37188 8452
rect 37240 8440 37246 8492
rect 40678 8440 40684 8492
rect 40736 8440 40742 8492
rect 35526 8372 35532 8424
rect 35584 8372 35590 8424
rect 36170 8372 36176 8424
rect 36228 8372 36234 8424
rect 37274 8372 37280 8424
rect 37332 8372 37338 8424
rect 40957 8347 41015 8353
rect 40957 8313 40969 8347
rect 41003 8344 41015 8347
rect 41046 8344 41052 8356
rect 41003 8316 41052 8344
rect 41003 8313 41015 8316
rect 40957 8307 41015 8313
rect 41046 8304 41052 8316
rect 41104 8304 41110 8356
rect 34624 8248 35204 8276
rect 32769 8239 32827 8245
rect 35434 8236 35440 8288
rect 35492 8236 35498 8288
rect 1104 8186 41400 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 41400 8186
rect 1104 8112 41400 8134
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5592 8044 12388 8072
rect 5592 8032 5598 8044
rect 12360 8004 12388 8044
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12529 8075 12587 8081
rect 12529 8072 12541 8075
rect 12492 8044 12541 8072
rect 12492 8032 12498 8044
rect 12529 8041 12541 8044
rect 12575 8041 12587 8075
rect 12529 8035 12587 8041
rect 15197 8075 15255 8081
rect 15197 8041 15209 8075
rect 15243 8072 15255 8075
rect 15654 8072 15660 8084
rect 15243 8044 15660 8072
rect 15243 8041 15255 8044
rect 15197 8035 15255 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 16390 8032 16396 8084
rect 16448 8072 16454 8084
rect 16850 8072 16856 8084
rect 16448 8044 16856 8072
rect 16448 8032 16454 8044
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 20898 8032 20904 8084
rect 20956 8032 20962 8084
rect 21082 8032 21088 8084
rect 21140 8072 21146 8084
rect 21818 8072 21824 8084
rect 21140 8044 21824 8072
rect 21140 8032 21146 8044
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 22281 8075 22339 8081
rect 22281 8072 22293 8075
rect 22244 8044 22293 8072
rect 22244 8032 22250 8044
rect 22281 8041 22293 8044
rect 22327 8041 22339 8075
rect 22281 8035 22339 8041
rect 24762 8032 24768 8084
rect 24820 8072 24826 8084
rect 24857 8075 24915 8081
rect 24857 8072 24869 8075
rect 24820 8044 24869 8072
rect 24820 8032 24826 8044
rect 24857 8041 24869 8044
rect 24903 8041 24915 8075
rect 24857 8035 24915 8041
rect 25041 8075 25099 8081
rect 25041 8041 25053 8075
rect 25087 8072 25099 8075
rect 26050 8072 26056 8084
rect 25087 8044 26056 8072
rect 25087 8041 25099 8044
rect 25041 8035 25099 8041
rect 26050 8032 26056 8044
rect 26108 8032 26114 8084
rect 34241 8075 34299 8081
rect 34241 8072 34253 8075
rect 31128 8044 34253 8072
rect 14550 8004 14556 8016
rect 8220 7976 10456 8004
rect 12360 7976 14556 8004
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4614 7936 4620 7948
rect 4111 7908 4620 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 5776 7908 6285 7936
rect 5776 7896 5782 7908
rect 6273 7905 6285 7908
rect 6319 7936 6331 7939
rect 8220 7936 8248 7976
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 6319 7908 8248 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 934 7828 940 7880
rect 992 7868 998 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 992 7840 1409 7868
rect 992 7828 998 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6362 7868 6368 7880
rect 6135 7840 6368 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7769 1731 7803
rect 3804 7800 3832 7831
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 8220 7877 8248 7908
rect 8312 7908 9597 7936
rect 8312 7877 8340 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 8662 7868 8668 7880
rect 8619 7840 8668 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 4062 7800 4068 7812
rect 3804 7772 4068 7800
rect 1673 7763 1731 7769
rect 1688 7732 1716 7763
rect 4062 7760 4068 7772
rect 4120 7760 4126 7812
rect 4706 7760 4712 7812
rect 4764 7760 4770 7812
rect 7558 7800 7564 7812
rect 5368 7772 7564 7800
rect 5368 7732 5396 7772
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 8496 7800 8524 7831
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 9033 7871 9091 7877
rect 9033 7837 9045 7871
rect 9079 7868 9091 7871
rect 9079 7840 9536 7868
rect 9079 7837 9091 7840
rect 9033 7831 9091 7837
rect 7708 7772 8524 7800
rect 7708 7760 7714 7772
rect 9508 7744 9536 7840
rect 10042 7828 10048 7880
rect 10100 7828 10106 7880
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 10428 7877 10456 7976
rect 14550 7964 14556 7976
rect 14608 7964 14614 8016
rect 16666 8004 16672 8016
rect 15580 7976 16672 8004
rect 13538 7896 13544 7948
rect 13596 7896 13602 7948
rect 15580 7880 15608 7976
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 16868 8004 16896 8032
rect 17865 8007 17923 8013
rect 16868 7976 17080 8004
rect 17052 7936 17080 7976
rect 17865 7973 17877 8007
rect 17911 8004 17923 8007
rect 25409 8007 25467 8013
rect 25409 8004 25421 8007
rect 17911 7976 25421 8004
rect 17911 7973 17923 7976
rect 17865 7967 17923 7973
rect 25409 7973 25421 7976
rect 25455 7973 25467 8007
rect 28074 8004 28080 8016
rect 25409 7967 25467 7973
rect 25884 7976 28080 8004
rect 19245 7939 19303 7945
rect 16592 7908 16988 7936
rect 16592 7880 16620 7908
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7868 11023 7871
rect 11330 7868 11336 7880
rect 11011 7840 11336 7868
rect 11011 7837 11023 7840
rect 10965 7831 11023 7837
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 13265 7871 13323 7877
rect 12759 7840 12940 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 10321 7803 10379 7809
rect 10321 7769 10333 7803
rect 10367 7800 10379 7803
rect 11517 7803 11575 7809
rect 11517 7800 11529 7803
rect 10367 7772 11529 7800
rect 10367 7769 10379 7772
rect 10321 7763 10379 7769
rect 11517 7769 11529 7772
rect 11563 7769 11575 7803
rect 11517 7763 11575 7769
rect 11698 7760 11704 7812
rect 11756 7760 11762 7812
rect 1688 7704 5396 7732
rect 5718 7692 5724 7744
rect 5776 7692 5782 7744
rect 6181 7735 6239 7741
rect 6181 7701 6193 7735
rect 6227 7732 6239 7735
rect 7098 7732 7104 7744
rect 6227 7704 7104 7732
rect 6227 7701 6239 7704
rect 6181 7695 6239 7701
rect 7098 7692 7104 7704
rect 7156 7732 7162 7744
rect 7926 7732 7932 7744
rect 7156 7704 7932 7732
rect 7156 7692 7162 7704
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 8018 7692 8024 7744
rect 8076 7692 8082 7744
rect 9490 7692 9496 7744
rect 9548 7692 9554 7744
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 10192 7704 10609 7732
rect 10192 7692 10198 7704
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10597 7695 10655 7701
rect 11790 7692 11796 7744
rect 11848 7692 11854 7744
rect 12912 7741 12940 7840
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 13814 7868 13820 7880
rect 13311 7840 13820 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 13814 7828 13820 7840
rect 13872 7828 13878 7880
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 14292 7840 14657 7868
rect 14292 7744 14320 7840
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 15010 7828 15016 7880
rect 15068 7828 15074 7880
rect 15562 7828 15568 7880
rect 15620 7828 15626 7880
rect 15838 7828 15844 7880
rect 15896 7828 15902 7880
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 16390 7868 16396 7880
rect 15988 7840 16396 7868
rect 15988 7828 15994 7840
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 16482 7828 16488 7880
rect 16540 7828 16546 7880
rect 16574 7828 16580 7880
rect 16632 7828 16638 7880
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 16758 7868 16764 7880
rect 16715 7840 16764 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 16960 7877 16988 7908
rect 17052 7908 17724 7936
rect 17052 7877 17080 7908
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 17696 7877 17724 7908
rect 19245 7905 19257 7939
rect 19291 7936 19303 7939
rect 22738 7936 22744 7948
rect 19291 7908 22744 7936
rect 19291 7905 19303 7908
rect 19245 7899 19303 7905
rect 22738 7896 22744 7908
rect 22796 7896 22802 7948
rect 22922 7896 22928 7948
rect 22980 7896 22986 7948
rect 24765 7939 24823 7945
rect 24765 7905 24777 7939
rect 24811 7936 24823 7939
rect 25590 7936 25596 7948
rect 24811 7908 25596 7936
rect 24811 7905 24823 7908
rect 24765 7899 24823 7905
rect 25590 7896 25596 7908
rect 25648 7896 25654 7948
rect 17589 7871 17647 7877
rect 17589 7868 17601 7871
rect 17460 7840 17601 7868
rect 17460 7828 17466 7840
rect 17589 7837 17601 7840
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 19426 7828 19432 7880
rect 19484 7828 19490 7880
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 14734 7760 14740 7812
rect 14792 7800 14798 7812
rect 14829 7803 14887 7809
rect 14829 7800 14841 7803
rect 14792 7772 14841 7800
rect 14792 7760 14798 7772
rect 14829 7769 14841 7772
rect 14875 7769 14887 7803
rect 14829 7763 14887 7769
rect 14918 7760 14924 7812
rect 14976 7760 14982 7812
rect 15194 7760 15200 7812
rect 15252 7800 15258 7812
rect 15746 7800 15752 7812
rect 15252 7772 15752 7800
rect 15252 7760 15258 7772
rect 15746 7760 15752 7772
rect 15804 7800 15810 7812
rect 16500 7800 16528 7828
rect 16853 7803 16911 7809
rect 16853 7800 16865 7803
rect 15804 7772 16865 7800
rect 15804 7760 15810 7772
rect 16853 7769 16865 7772
rect 16899 7800 16911 7803
rect 17497 7803 17555 7809
rect 17497 7800 17509 7803
rect 16899 7772 17509 7800
rect 16899 7769 16911 7772
rect 16853 7763 16911 7769
rect 17497 7769 17509 7772
rect 17543 7769 17555 7803
rect 17497 7763 17555 7769
rect 18598 7760 18604 7812
rect 18656 7800 18662 7812
rect 19536 7800 19564 7831
rect 19702 7828 19708 7880
rect 19760 7828 19766 7880
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7868 19855 7871
rect 19978 7868 19984 7880
rect 19843 7840 19984 7868
rect 19843 7837 19855 7840
rect 19797 7831 19855 7837
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 21082 7828 21088 7880
rect 21140 7828 21146 7880
rect 21266 7828 21272 7880
rect 21324 7828 21330 7880
rect 21358 7828 21364 7880
rect 21416 7828 21422 7880
rect 21634 7828 21640 7880
rect 21692 7868 21698 7880
rect 22002 7868 22008 7880
rect 21692 7840 22008 7868
rect 21692 7828 21698 7840
rect 22002 7828 22008 7840
rect 22060 7828 22066 7880
rect 22649 7871 22707 7877
rect 22649 7837 22661 7871
rect 22695 7868 22707 7871
rect 23290 7868 23296 7880
rect 22695 7840 23296 7868
rect 22695 7837 22707 7840
rect 22649 7831 22707 7837
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7868 25007 7871
rect 25130 7868 25136 7880
rect 24995 7840 25136 7868
rect 24995 7837 25007 7840
rect 24949 7831 25007 7837
rect 24596 7800 24624 7831
rect 25130 7828 25136 7840
rect 25188 7828 25194 7880
rect 25222 7828 25228 7880
rect 25280 7828 25286 7880
rect 25314 7828 25320 7880
rect 25372 7828 25378 7880
rect 25501 7871 25559 7877
rect 25501 7837 25513 7871
rect 25547 7837 25559 7871
rect 25501 7831 25559 7837
rect 18656 7772 19564 7800
rect 19628 7772 24624 7800
rect 25148 7800 25176 7828
rect 25516 7800 25544 7831
rect 25682 7828 25688 7880
rect 25740 7828 25746 7880
rect 25884 7877 25912 7976
rect 28074 7964 28080 7976
rect 28132 7964 28138 8016
rect 31128 7948 31156 8044
rect 34241 8041 34253 8044
rect 34287 8041 34299 8075
rect 34241 8035 34299 8041
rect 34606 8032 34612 8084
rect 34664 8032 34670 8084
rect 34624 8004 34652 8032
rect 35526 8004 35532 8016
rect 34624 7976 35532 8004
rect 30558 7896 30564 7948
rect 30616 7896 30622 7948
rect 31110 7896 31116 7948
rect 31168 7896 31174 7948
rect 31665 7939 31723 7945
rect 31665 7905 31677 7939
rect 31711 7936 31723 7939
rect 34606 7936 34612 7948
rect 31711 7908 34612 7936
rect 31711 7905 31723 7908
rect 31665 7899 31723 7905
rect 34606 7896 34612 7908
rect 34664 7896 34670 7948
rect 34716 7945 34744 7976
rect 35526 7964 35532 7976
rect 35584 7964 35590 8016
rect 38105 8007 38163 8013
rect 38105 7973 38117 8007
rect 38151 8004 38163 8007
rect 38151 7976 39160 8004
rect 38151 7973 38163 7976
rect 38105 7967 38163 7973
rect 34701 7939 34759 7945
rect 34701 7905 34713 7939
rect 34747 7905 34759 7939
rect 35069 7939 35127 7945
rect 35069 7936 35081 7939
rect 34701 7899 34759 7905
rect 34808 7908 35081 7936
rect 25833 7871 25912 7877
rect 25833 7837 25845 7871
rect 25879 7840 25912 7871
rect 25879 7837 25891 7840
rect 25833 7831 25891 7837
rect 25958 7828 25964 7880
rect 26016 7828 26022 7880
rect 26142 7828 26148 7880
rect 26200 7877 26206 7880
rect 26200 7868 26208 7877
rect 30745 7871 30803 7877
rect 26200 7840 26245 7868
rect 26200 7831 26208 7840
rect 30745 7837 30757 7871
rect 30791 7837 30803 7871
rect 30745 7831 30803 7837
rect 30929 7871 30987 7877
rect 30929 7837 30941 7871
rect 30975 7868 30987 7871
rect 31205 7871 31263 7877
rect 31205 7868 31217 7871
rect 30975 7840 31217 7868
rect 30975 7837 30987 7840
rect 30929 7831 30987 7837
rect 31205 7837 31217 7840
rect 31251 7837 31263 7871
rect 31205 7831 31263 7837
rect 26200 7828 26206 7831
rect 25148 7772 25544 7800
rect 18656 7760 18662 7772
rect 12897 7735 12955 7741
rect 12897 7701 12909 7735
rect 12943 7701 12955 7735
rect 12897 7695 12955 7701
rect 13357 7735 13415 7741
rect 13357 7701 13369 7735
rect 13403 7732 13415 7735
rect 13446 7732 13452 7744
rect 13403 7704 13452 7732
rect 13403 7701 13415 7704
rect 13357 7695 13415 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 14274 7692 14280 7744
rect 14332 7692 14338 7744
rect 16114 7692 16120 7744
rect 16172 7692 16178 7744
rect 17218 7692 17224 7744
rect 17276 7692 17282 7744
rect 19058 7692 19064 7744
rect 19116 7732 19122 7744
rect 19628 7732 19656 7772
rect 19116 7704 19656 7732
rect 19116 7692 19122 7704
rect 21174 7692 21180 7744
rect 21232 7732 21238 7744
rect 22646 7732 22652 7744
rect 21232 7704 22652 7732
rect 21232 7692 21238 7704
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 22738 7692 22744 7744
rect 22796 7692 22802 7744
rect 24210 7692 24216 7744
rect 24268 7732 24274 7744
rect 25700 7732 25728 7828
rect 26050 7760 26056 7812
rect 26108 7760 26114 7812
rect 30760 7800 30788 7831
rect 31478 7828 31484 7880
rect 31536 7828 31542 7880
rect 33042 7828 33048 7880
rect 33100 7828 33106 7880
rect 33686 7828 33692 7880
rect 33744 7828 33750 7880
rect 34054 7828 34060 7880
rect 34112 7868 34118 7880
rect 34425 7871 34483 7877
rect 34425 7868 34437 7871
rect 34112 7840 34437 7868
rect 34112 7828 34118 7840
rect 34425 7837 34437 7840
rect 34471 7837 34483 7871
rect 34425 7831 34483 7837
rect 34514 7828 34520 7880
rect 34572 7828 34578 7880
rect 31496 7800 31524 7828
rect 30760 7772 31524 7800
rect 31941 7803 31999 7809
rect 31941 7769 31953 7803
rect 31987 7800 31999 7803
rect 32214 7800 32220 7812
rect 31987 7772 32220 7800
rect 31987 7769 31999 7772
rect 31941 7763 31999 7769
rect 32214 7760 32220 7772
rect 32272 7760 32278 7812
rect 34241 7803 34299 7809
rect 34241 7769 34253 7803
rect 34287 7800 34299 7803
rect 34808 7800 34836 7908
rect 35069 7905 35081 7908
rect 35115 7905 35127 7939
rect 35069 7899 35127 7905
rect 37826 7896 37832 7948
rect 37884 7936 37890 7948
rect 38657 7939 38715 7945
rect 38657 7936 38669 7939
rect 37884 7908 38669 7936
rect 37884 7896 37890 7908
rect 38657 7905 38669 7908
rect 38703 7905 38715 7939
rect 38657 7899 38715 7905
rect 34885 7871 34943 7877
rect 34885 7837 34897 7871
rect 34931 7868 34943 7871
rect 34931 7840 35020 7868
rect 34931 7837 34943 7840
rect 34885 7831 34943 7837
rect 34287 7772 34836 7800
rect 34287 7769 34299 7772
rect 34241 7763 34299 7769
rect 24268 7704 25728 7732
rect 24268 7692 24274 7704
rect 26326 7692 26332 7744
rect 26384 7692 26390 7744
rect 26970 7692 26976 7744
rect 27028 7732 27034 7744
rect 27522 7732 27528 7744
rect 27028 7704 27528 7732
rect 27028 7692 27034 7704
rect 27522 7692 27528 7704
rect 27580 7692 27586 7744
rect 31573 7735 31631 7741
rect 31573 7701 31585 7735
rect 31619 7732 31631 7735
rect 32030 7732 32036 7744
rect 31619 7704 32036 7732
rect 31619 7701 31631 7704
rect 31573 7695 31631 7701
rect 32030 7692 32036 7704
rect 32088 7692 32094 7744
rect 33594 7692 33600 7744
rect 33652 7732 33658 7744
rect 34992 7732 35020 7840
rect 38010 7828 38016 7880
rect 38068 7868 38074 7880
rect 39132 7877 39160 7976
rect 38565 7871 38623 7877
rect 38565 7868 38577 7871
rect 38068 7840 38577 7868
rect 38068 7828 38074 7840
rect 38565 7837 38577 7840
rect 38611 7837 38623 7871
rect 38565 7831 38623 7837
rect 39117 7871 39175 7877
rect 39117 7837 39129 7871
rect 39163 7837 39175 7871
rect 39117 7831 39175 7837
rect 39945 7871 40003 7877
rect 39945 7837 39957 7871
rect 39991 7868 40003 7871
rect 40678 7868 40684 7880
rect 39991 7840 40684 7868
rect 39991 7837 40003 7840
rect 39945 7831 40003 7837
rect 40678 7828 40684 7840
rect 40736 7828 40742 7880
rect 38473 7803 38531 7809
rect 38473 7769 38485 7803
rect 38519 7800 38531 7803
rect 40497 7803 40555 7809
rect 40497 7800 40509 7803
rect 38519 7772 40509 7800
rect 38519 7769 38531 7772
rect 38473 7763 38531 7769
rect 40497 7769 40509 7772
rect 40543 7769 40555 7803
rect 40497 7763 40555 7769
rect 33652 7704 35020 7732
rect 38933 7735 38991 7741
rect 33652 7692 33658 7704
rect 38933 7701 38945 7735
rect 38979 7732 38991 7735
rect 39114 7732 39120 7744
rect 38979 7704 39120 7732
rect 38979 7701 38991 7704
rect 38933 7695 38991 7701
rect 39114 7692 39120 7704
rect 39172 7692 39178 7744
rect 1104 7642 41400 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 41400 7642
rect 1104 7568 41400 7590
rect 5718 7488 5724 7540
rect 5776 7488 5782 7540
rect 9674 7528 9680 7540
rect 7760 7500 9680 7528
rect 5736 7401 5764 7488
rect 7760 7404 7788 7500
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 10134 7528 10140 7540
rect 9876 7500 10140 7528
rect 8018 7420 8024 7472
rect 8076 7420 8082 7472
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 9692 7460 9720 7488
rect 9876 7469 9904 7500
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 15286 7488 15292 7540
rect 15344 7528 15350 7540
rect 15838 7528 15844 7540
rect 15344 7500 15844 7528
rect 15344 7488 15350 7500
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16114 7488 16120 7540
rect 16172 7488 16178 7540
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 21266 7528 21272 7540
rect 17635 7500 21272 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 21637 7531 21695 7537
rect 21637 7528 21649 7531
rect 21416 7500 21649 7528
rect 21416 7488 21422 7500
rect 21637 7497 21649 7500
rect 21683 7497 21695 7531
rect 24857 7531 24915 7537
rect 21637 7491 21695 7497
rect 21744 7500 22508 7528
rect 8168 7432 8510 7460
rect 9600 7432 9720 7460
rect 9861 7463 9919 7469
rect 8168 7420 8174 7432
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 9600 7401 9628 7432
rect 9861 7429 9873 7463
rect 9907 7429 9919 7463
rect 11790 7460 11796 7472
rect 11086 7446 11796 7460
rect 9861 7423 9919 7429
rect 11072 7432 11796 7446
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 11072 7324 11100 7432
rect 11790 7420 11796 7432
rect 11848 7420 11854 7472
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 15197 7463 15255 7469
rect 15197 7460 15209 7463
rect 14608 7432 15209 7460
rect 14608 7420 14614 7432
rect 15197 7429 15209 7432
rect 15243 7429 15255 7463
rect 16132 7460 16160 7488
rect 17957 7463 18015 7469
rect 15197 7423 15255 7429
rect 15304 7432 15976 7460
rect 16132 7432 16988 7460
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 14921 7395 14979 7401
rect 14921 7392 14933 7395
rect 14884 7364 14933 7392
rect 14884 7352 14890 7364
rect 14921 7361 14933 7364
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 15010 7352 15016 7404
rect 15068 7352 15074 7404
rect 15102 7352 15108 7404
rect 15160 7352 15166 7404
rect 15304 7401 15332 7432
rect 15948 7404 15976 7432
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7361 15347 7395
rect 15289 7355 15347 7361
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 8168 7296 11100 7324
rect 15028 7324 15056 7352
rect 15580 7324 15608 7355
rect 15746 7352 15752 7404
rect 15804 7352 15810 7404
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 15028 7296 15608 7324
rect 8168 7284 8174 7296
rect 14274 7256 14280 7268
rect 11256 7228 14280 7256
rect 5534 7148 5540 7200
rect 5592 7148 5598 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 11256 7188 11284 7228
rect 14274 7216 14280 7228
rect 14332 7256 14338 7268
rect 15856 7256 15884 7355
rect 15930 7352 15936 7404
rect 15988 7352 15994 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16132 7364 16865 7392
rect 16132 7265 16160 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16960 7324 16988 7432
rect 17144 7432 17908 7460
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 17144 7401 17172 7432
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 17773 7395 17831 7401
rect 17773 7392 17785 7395
rect 17276 7364 17785 7392
rect 17276 7352 17282 7364
rect 17773 7361 17785 7364
rect 17819 7361 17831 7395
rect 17880 7392 17908 7432
rect 17957 7429 17969 7463
rect 18003 7460 18015 7463
rect 18322 7460 18328 7472
rect 18003 7432 18328 7460
rect 18003 7429 18015 7432
rect 17957 7423 18015 7429
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 21744 7460 21772 7500
rect 18524 7432 19288 7460
rect 18049 7395 18107 7401
rect 18049 7392 18061 7395
rect 17880 7364 18061 7392
rect 17773 7355 17831 7361
rect 18049 7361 18061 7364
rect 18095 7392 18107 7395
rect 18524 7392 18552 7432
rect 19260 7404 19288 7432
rect 21008 7432 21772 7460
rect 21913 7463 21971 7469
rect 18095 7364 18552 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 18598 7352 18604 7404
rect 18656 7352 18662 7404
rect 19242 7352 19248 7404
rect 19300 7352 19306 7404
rect 20254 7352 20260 7404
rect 20312 7392 20318 7404
rect 21008 7401 21036 7432
rect 21913 7429 21925 7463
rect 21959 7460 21971 7463
rect 21959 7432 22324 7460
rect 21959 7429 21971 7432
rect 21913 7423 21971 7429
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20312 7364 21005 7392
rect 20312 7352 20318 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 21082 7352 21088 7404
rect 21140 7392 21146 7404
rect 21140 7364 21185 7392
rect 21140 7352 21146 7364
rect 21266 7352 21272 7404
rect 21324 7352 21330 7404
rect 21358 7352 21364 7404
rect 21416 7352 21422 7404
rect 21542 7401 21548 7404
rect 21499 7395 21548 7401
rect 21499 7361 21511 7395
rect 21545 7361 21548 7395
rect 21499 7355 21548 7361
rect 21542 7352 21548 7355
rect 21600 7352 21606 7404
rect 21818 7352 21824 7404
rect 21876 7352 21882 7404
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 22112 7324 22140 7355
rect 16960 7296 22140 7324
rect 14332 7228 15884 7256
rect 16117 7259 16175 7265
rect 14332 7216 14338 7228
rect 16117 7225 16129 7259
rect 16163 7225 16175 7259
rect 22296 7256 22324 7432
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 22480 7324 22508 7500
rect 24857 7497 24869 7531
rect 24903 7497 24915 7531
rect 24857 7491 24915 7497
rect 22646 7420 22652 7472
rect 22704 7460 22710 7472
rect 24489 7463 24547 7469
rect 24489 7460 24501 7463
rect 22704 7432 24501 7460
rect 22704 7420 22710 7432
rect 24489 7429 24501 7432
rect 24535 7460 24547 7463
rect 24762 7460 24768 7472
rect 24535 7432 24768 7460
rect 24535 7429 24547 7432
rect 24489 7423 24547 7429
rect 24762 7420 24768 7432
rect 24820 7420 24826 7472
rect 24872 7460 24900 7491
rect 24946 7488 24952 7540
rect 25004 7488 25010 7540
rect 25222 7488 25228 7540
rect 25280 7488 25286 7540
rect 25590 7488 25596 7540
rect 25648 7528 25654 7540
rect 26421 7531 26479 7537
rect 26421 7528 26433 7531
rect 25648 7500 26433 7528
rect 25648 7488 25654 7500
rect 26421 7497 26433 7500
rect 26467 7497 26479 7531
rect 26421 7491 26479 7497
rect 26694 7488 26700 7540
rect 26752 7528 26758 7540
rect 27433 7531 27491 7537
rect 27433 7528 27445 7531
rect 26752 7500 27445 7528
rect 26752 7488 26758 7500
rect 27433 7497 27445 7500
rect 27479 7497 27491 7531
rect 27433 7491 27491 7497
rect 31754 7488 31760 7540
rect 31812 7528 31818 7540
rect 33042 7528 33048 7540
rect 31812 7500 33048 7528
rect 31812 7488 31818 7500
rect 33042 7488 33048 7500
rect 33100 7528 33106 7540
rect 40589 7531 40647 7537
rect 33100 7500 36308 7528
rect 33100 7488 33106 7500
rect 25240 7460 25268 7488
rect 26326 7460 26332 7472
rect 24872 7432 25268 7460
rect 25424 7432 26332 7460
rect 22554 7352 22560 7404
rect 22612 7352 22618 7404
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7392 22983 7395
rect 24210 7392 24216 7404
rect 22971 7364 24216 7392
rect 22971 7361 22983 7364
rect 22925 7355 22983 7361
rect 22940 7324 22968 7355
rect 24210 7352 24216 7364
rect 24268 7352 24274 7404
rect 24306 7395 24364 7401
rect 24306 7361 24318 7395
rect 24352 7361 24364 7395
rect 24306 7355 24364 7361
rect 22480 7296 22968 7324
rect 22462 7256 22468 7268
rect 16117 7219 16175 7225
rect 16592 7228 19288 7256
rect 22296 7228 22468 7256
rect 9548 7160 11284 7188
rect 9548 7148 9554 7160
rect 11330 7148 11336 7200
rect 11388 7188 11394 7200
rect 15286 7188 15292 7200
rect 11388 7160 15292 7188
rect 11388 7148 11394 7160
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15473 7191 15531 7197
rect 15473 7157 15485 7191
rect 15519 7188 15531 7191
rect 16592 7188 16620 7228
rect 15519 7160 16620 7188
rect 16669 7191 16727 7197
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 16669 7157 16681 7191
rect 16715 7188 16727 7191
rect 19058 7188 19064 7200
rect 16715 7160 19064 7188
rect 16715 7157 16727 7160
rect 16669 7151 16727 7157
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 19150 7148 19156 7200
rect 19208 7148 19214 7200
rect 19260 7188 19288 7228
rect 22462 7216 22468 7228
rect 22520 7216 22526 7268
rect 24320 7256 24348 7355
rect 24394 7352 24400 7404
rect 24452 7352 24458 7404
rect 24578 7352 24584 7404
rect 24636 7352 24642 7404
rect 24678 7395 24736 7401
rect 24678 7361 24690 7395
rect 24724 7361 24736 7395
rect 24678 7355 24736 7361
rect 25133 7395 25191 7401
rect 25133 7361 25145 7395
rect 25179 7361 25191 7395
rect 25133 7355 25191 7361
rect 24412 7324 24440 7352
rect 24688 7324 24716 7355
rect 24412 7296 24716 7324
rect 25148 7268 25176 7355
rect 25222 7352 25228 7404
rect 25280 7352 25286 7404
rect 25424 7401 25452 7432
rect 26326 7420 26332 7432
rect 26384 7420 26390 7472
rect 36280 7460 36308 7500
rect 40589 7497 40601 7531
rect 40635 7528 40647 7531
rect 40678 7528 40684 7540
rect 40635 7500 40684 7528
rect 40635 7497 40647 7500
rect 40589 7491 40647 7497
rect 40678 7488 40684 7500
rect 40736 7488 40742 7540
rect 38838 7460 38844 7472
rect 27264 7432 29132 7460
rect 36202 7432 38844 7460
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7361 25559 7395
rect 25501 7355 25559 7361
rect 24946 7256 24952 7268
rect 24320 7228 24952 7256
rect 24946 7216 24952 7228
rect 25004 7216 25010 7268
rect 25130 7216 25136 7268
rect 25188 7216 25194 7268
rect 25516 7188 25544 7355
rect 25682 7352 25688 7404
rect 25740 7392 25746 7404
rect 25777 7395 25835 7401
rect 25777 7392 25789 7395
rect 25740 7364 25789 7392
rect 25740 7352 25746 7364
rect 25777 7361 25789 7364
rect 25823 7361 25835 7395
rect 25777 7355 25835 7361
rect 25870 7395 25928 7401
rect 25870 7361 25882 7395
rect 25916 7361 25928 7395
rect 25870 7355 25928 7361
rect 25884 7256 25912 7355
rect 25958 7352 25964 7404
rect 26016 7392 26022 7404
rect 26053 7395 26111 7401
rect 26053 7392 26065 7395
rect 26016 7364 26065 7392
rect 26016 7352 26022 7364
rect 26053 7361 26065 7364
rect 26099 7361 26111 7395
rect 26053 7355 26111 7361
rect 26145 7395 26203 7401
rect 26145 7361 26157 7395
rect 26191 7361 26203 7395
rect 26145 7355 26203 7361
rect 26160 7324 26188 7355
rect 26234 7352 26240 7404
rect 26292 7401 26298 7404
rect 26292 7392 26300 7401
rect 26292 7364 26337 7392
rect 26292 7355 26300 7364
rect 26292 7352 26298 7355
rect 27264 7324 27292 7432
rect 27341 7395 27399 7401
rect 27341 7361 27353 7395
rect 27387 7392 27399 7395
rect 28445 7395 28503 7401
rect 28445 7392 28457 7395
rect 27387 7364 28457 7392
rect 27387 7361 27399 7364
rect 27341 7355 27399 7361
rect 28445 7361 28457 7364
rect 28491 7361 28503 7395
rect 28445 7355 28503 7361
rect 26160 7296 27292 7324
rect 27522 7284 27528 7336
rect 27580 7284 27586 7336
rect 27893 7327 27951 7333
rect 27893 7293 27905 7327
rect 27939 7324 27951 7327
rect 28552 7324 28580 7432
rect 28721 7395 28779 7401
rect 28721 7361 28733 7395
rect 28767 7361 28779 7395
rect 28721 7355 28779 7361
rect 27939 7296 28580 7324
rect 27939 7293 27951 7296
rect 27893 7287 27951 7293
rect 26602 7256 26608 7268
rect 25884 7228 26608 7256
rect 26602 7216 26608 7228
rect 26660 7216 26666 7268
rect 26973 7259 27031 7265
rect 26973 7225 26985 7259
rect 27019 7256 27031 7259
rect 28736 7256 28764 7355
rect 29104 7336 29132 7432
rect 38838 7420 38844 7432
rect 38896 7460 38902 7472
rect 38896 7432 39606 7460
rect 38896 7420 38902 7432
rect 34606 7352 34612 7404
rect 34664 7392 34670 7404
rect 34701 7395 34759 7401
rect 34701 7392 34713 7395
rect 34664 7364 34713 7392
rect 34664 7352 34670 7364
rect 34701 7361 34713 7364
rect 34747 7361 34759 7395
rect 34701 7355 34759 7361
rect 29086 7284 29092 7336
rect 29144 7284 29150 7336
rect 34977 7327 35035 7333
rect 34977 7293 34989 7327
rect 35023 7324 35035 7327
rect 35434 7324 35440 7336
rect 35023 7296 35440 7324
rect 35023 7293 35035 7296
rect 34977 7287 35035 7293
rect 35434 7284 35440 7296
rect 35492 7284 35498 7336
rect 35526 7284 35532 7336
rect 35584 7324 35590 7336
rect 36449 7327 36507 7333
rect 36449 7324 36461 7327
rect 35584 7296 36461 7324
rect 35584 7284 35590 7296
rect 36449 7293 36461 7296
rect 36495 7293 36507 7327
rect 36449 7287 36507 7293
rect 37274 7284 37280 7336
rect 37332 7324 37338 7336
rect 38841 7327 38899 7333
rect 38841 7324 38853 7327
rect 37332 7296 38853 7324
rect 37332 7284 37338 7296
rect 38841 7293 38853 7296
rect 38887 7293 38899 7327
rect 38841 7287 38899 7293
rect 39114 7284 39120 7336
rect 39172 7284 39178 7336
rect 27019 7228 28764 7256
rect 27019 7225 27031 7228
rect 26973 7219 27031 7225
rect 19260 7160 25544 7188
rect 28534 7148 28540 7200
rect 28592 7148 28598 7200
rect 1104 7098 41400 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 41400 7098
rect 1104 7024 41400 7046
rect 5534 6993 5540 6996
rect 5524 6987 5540 6993
rect 5524 6953 5536 6987
rect 5524 6947 5540 6953
rect 5534 6944 5540 6947
rect 5592 6944 5598 6996
rect 7009 6987 7067 6993
rect 7009 6953 7021 6987
rect 7055 6984 7067 6987
rect 7098 6984 7104 6996
rect 7055 6956 7104 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 9030 6944 9036 6996
rect 9088 6984 9094 6996
rect 13446 6984 13452 6996
rect 9088 6956 13452 6984
rect 9088 6944 9094 6956
rect 13446 6944 13452 6956
rect 13504 6984 13510 6996
rect 13504 6956 18644 6984
rect 13504 6944 13510 6956
rect 13538 6876 13544 6928
rect 13596 6916 13602 6928
rect 13596 6888 14596 6916
rect 13596 6876 13602 6888
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 5074 6848 5080 6860
rect 4120 6820 5080 6848
rect 4120 6808 4126 6820
rect 5074 6808 5080 6820
rect 5132 6848 5138 6860
rect 5261 6851 5319 6857
rect 5261 6848 5273 6851
rect 5132 6820 5273 6848
rect 5132 6808 5138 6820
rect 5261 6817 5273 6820
rect 5307 6848 5319 6851
rect 12526 6848 12532 6860
rect 5307 6820 7788 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 7760 6792 7788 6820
rect 11164 6820 12532 6848
rect 7742 6740 7748 6792
rect 7800 6740 7806 6792
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 11164 6789 11192 6820
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 13909 6851 13967 6857
rect 13909 6817 13921 6851
rect 13955 6817 13967 6851
rect 14568 6848 14596 6888
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 14568 6820 14657 6848
rect 13909 6811 13967 6817
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 14645 6811 14703 6817
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8904 6752 9137 6780
rect 8904 6740 8910 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9125 6743 9183 6749
rect 9600 6752 9873 6780
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 5994 6712 6000 6724
rect 4764 6684 6000 6712
rect 4764 6672 4770 6684
rect 5994 6672 6000 6684
rect 6052 6672 6058 6724
rect 9600 6656 9628 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 9950 6672 9956 6724
rect 10008 6712 10014 6724
rect 11440 6712 11468 6743
rect 12158 6740 12164 6792
rect 12216 6740 12222 6792
rect 13924 6780 13952 6811
rect 15378 6808 15384 6860
rect 15436 6808 15442 6860
rect 16022 6808 16028 6860
rect 16080 6808 16086 6860
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16574 6848 16580 6860
rect 16347 6820 16580 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16574 6808 16580 6820
rect 16632 6848 16638 6860
rect 17034 6848 17040 6860
rect 16632 6820 17040 6848
rect 16632 6808 16638 6820
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 18509 6851 18567 6857
rect 18509 6848 18521 6851
rect 18064 6820 18521 6848
rect 14553 6783 14611 6789
rect 13924 6752 14412 6780
rect 10008 6684 11468 6712
rect 10008 6672 10014 6684
rect 12434 6672 12440 6724
rect 12492 6672 12498 6724
rect 13814 6712 13820 6724
rect 13662 6684 13820 6712
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 9582 6604 9588 6656
rect 9640 6604 9646 6656
rect 9766 6604 9772 6656
rect 9824 6604 9830 6656
rect 10962 6604 10968 6656
rect 11020 6604 11026 6656
rect 11330 6604 11336 6656
rect 11388 6604 11394 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 14384 6644 14412 6752
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 15396 6780 15424 6808
rect 15930 6780 15936 6792
rect 14599 6752 15936 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16040 6780 16068 6808
rect 17678 6780 17684 6792
rect 16040 6752 17684 6780
rect 17678 6740 17684 6752
rect 17736 6780 17742 6792
rect 18064 6780 18092 6820
rect 18509 6817 18521 6820
rect 18555 6817 18567 6851
rect 18509 6811 18567 6817
rect 18616 6848 18644 6956
rect 19242 6944 19248 6996
rect 19300 6984 19306 6996
rect 19300 6956 21220 6984
rect 19300 6944 19306 6956
rect 20438 6916 20444 6928
rect 20088 6888 20444 6916
rect 19886 6848 19892 6860
rect 18616 6820 19892 6848
rect 17736 6752 18092 6780
rect 18417 6783 18475 6789
rect 17736 6740 17742 6752
rect 18417 6749 18429 6783
rect 18463 6780 18475 6783
rect 18616 6780 18644 6820
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 20088 6857 20116 6888
rect 20438 6876 20444 6888
rect 20496 6876 20502 6928
rect 21192 6916 21220 6956
rect 21266 6944 21272 6996
rect 21324 6984 21330 6996
rect 21634 6984 21640 6996
rect 21324 6956 21640 6984
rect 21324 6944 21330 6956
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 22005 6987 22063 6993
rect 22005 6953 22017 6987
rect 22051 6984 22063 6987
rect 22554 6984 22560 6996
rect 22051 6956 22560 6984
rect 22051 6953 22063 6956
rect 22005 6947 22063 6953
rect 22554 6944 22560 6956
rect 22612 6944 22618 6996
rect 22922 6944 22928 6996
rect 22980 6984 22986 6996
rect 22980 6956 26372 6984
rect 22980 6944 22986 6956
rect 26344 6928 26372 6956
rect 26602 6944 26608 6996
rect 26660 6984 26666 6996
rect 27430 6984 27436 6996
rect 26660 6956 27436 6984
rect 26660 6944 26666 6956
rect 27430 6944 27436 6956
rect 27488 6944 27494 6996
rect 21192 6888 21956 6916
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6817 20131 6851
rect 20073 6811 20131 6817
rect 20162 6808 20168 6860
rect 20220 6848 20226 6860
rect 20257 6851 20315 6857
rect 20257 6848 20269 6851
rect 20220 6820 20269 6848
rect 20220 6808 20226 6820
rect 20257 6817 20269 6820
rect 20303 6817 20315 6851
rect 20257 6811 20315 6817
rect 18463 6752 18644 6780
rect 19061 6783 19119 6789
rect 18463 6749 18475 6752
rect 18417 6743 18475 6749
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 19107 6752 19472 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 18325 6715 18383 6721
rect 18325 6681 18337 6715
rect 18371 6712 18383 6715
rect 19150 6712 19156 6724
rect 18371 6684 19156 6712
rect 18371 6681 18383 6684
rect 18325 6675 18383 6681
rect 19150 6672 19156 6684
rect 19208 6672 19214 6724
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 14384 6616 14473 6644
rect 14461 6613 14473 6616
rect 14507 6644 14519 6647
rect 14918 6644 14924 6656
rect 14507 6616 14924 6644
rect 14507 6613 14519 6616
rect 14461 6607 14519 6613
rect 14918 6604 14924 6616
rect 14976 6604 14982 6656
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 16853 6647 16911 6653
rect 16853 6644 16865 6647
rect 15896 6616 16865 6644
rect 15896 6604 15902 6616
rect 16853 6613 16865 6616
rect 16899 6613 16911 6647
rect 16853 6607 16911 6613
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 17957 6647 18015 6653
rect 17957 6644 17969 6647
rect 17920 6616 17969 6644
rect 17920 6604 17926 6616
rect 17957 6613 17969 6616
rect 18003 6613 18015 6647
rect 17957 6607 18015 6613
rect 18874 6604 18880 6656
rect 18932 6604 18938 6656
rect 19444 6653 19472 6752
rect 20438 6740 20444 6792
rect 20496 6780 20502 6792
rect 21192 6789 21220 6888
rect 21542 6808 21548 6860
rect 21600 6848 21606 6860
rect 21928 6848 21956 6888
rect 24394 6876 24400 6928
rect 24452 6916 24458 6928
rect 26142 6916 26148 6928
rect 24452 6888 26148 6916
rect 24452 6876 24458 6888
rect 26142 6876 26148 6888
rect 26200 6876 26206 6928
rect 26326 6876 26332 6928
rect 26384 6916 26390 6928
rect 29733 6919 29791 6925
rect 29733 6916 29745 6919
rect 26384 6888 26924 6916
rect 26384 6876 26390 6888
rect 21600 6820 21680 6848
rect 21928 6820 22094 6848
rect 21600 6808 21606 6820
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20496 6752 21005 6780
rect 20496 6740 20502 6752
rect 20993 6749 21005 6752
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21652 6780 21680 6820
rect 21821 6783 21879 6789
rect 21821 6780 21833 6783
rect 21652 6752 21833 6780
rect 21453 6743 21511 6749
rect 21821 6749 21833 6752
rect 21867 6780 21879 6783
rect 21867 6752 21956 6780
rect 21867 6749 21879 6752
rect 21821 6743 21879 6749
rect 19797 6715 19855 6721
rect 19797 6681 19809 6715
rect 19843 6712 19855 6715
rect 20901 6715 20959 6721
rect 20901 6712 20913 6715
rect 19843 6684 20913 6712
rect 19843 6681 19855 6684
rect 19797 6675 19855 6681
rect 20901 6681 20913 6684
rect 20947 6681 20959 6715
rect 20901 6675 20959 6681
rect 19429 6647 19487 6653
rect 19429 6613 19441 6647
rect 19475 6613 19487 6647
rect 19429 6607 19487 6613
rect 21358 6604 21364 6656
rect 21416 6604 21422 6656
rect 21468 6644 21496 6743
rect 21634 6672 21640 6724
rect 21692 6672 21698 6724
rect 21726 6672 21732 6724
rect 21784 6672 21790 6724
rect 21818 6644 21824 6656
rect 21468 6616 21824 6644
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 21928 6644 21956 6752
rect 22066 6712 22094 6820
rect 22186 6808 22192 6860
rect 22244 6848 22250 6860
rect 23382 6848 23388 6860
rect 22244 6820 23388 6848
rect 22244 6808 22250 6820
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 25314 6808 25320 6860
rect 25372 6808 25378 6860
rect 26694 6808 26700 6860
rect 26752 6808 26758 6860
rect 26896 6857 26924 6888
rect 29472 6888 29745 6916
rect 26881 6851 26939 6857
rect 26881 6817 26893 6851
rect 26927 6848 26939 6851
rect 27338 6848 27344 6860
rect 26927 6820 27344 6848
rect 26927 6817 26939 6820
rect 26881 6811 26939 6817
rect 27338 6808 27344 6820
rect 27396 6808 27402 6860
rect 27430 6808 27436 6860
rect 27488 6848 27494 6860
rect 28813 6851 28871 6857
rect 28813 6848 28825 6851
rect 27488 6820 28825 6848
rect 27488 6808 27494 6820
rect 28813 6817 28825 6820
rect 28859 6817 28871 6851
rect 28813 6811 28871 6817
rect 24486 6740 24492 6792
rect 24544 6740 24550 6792
rect 24854 6740 24860 6792
rect 24912 6780 24918 6792
rect 24949 6783 25007 6789
rect 24949 6780 24961 6783
rect 24912 6752 24961 6780
rect 24912 6740 24918 6752
rect 24949 6749 24961 6752
rect 24995 6749 25007 6783
rect 24949 6743 25007 6749
rect 25130 6740 25136 6792
rect 25188 6740 25194 6792
rect 26602 6740 26608 6792
rect 26660 6740 26666 6792
rect 27062 6740 27068 6792
rect 27120 6740 27126 6792
rect 28626 6740 28632 6792
rect 28684 6780 28690 6792
rect 28828 6780 28856 6811
rect 28684 6752 28856 6780
rect 29365 6783 29423 6789
rect 28684 6740 28690 6752
rect 29365 6749 29377 6783
rect 29411 6780 29423 6783
rect 29472 6780 29500 6888
rect 29733 6885 29745 6888
rect 29779 6885 29791 6919
rect 29733 6879 29791 6885
rect 29546 6808 29552 6860
rect 29604 6848 29610 6860
rect 30193 6851 30251 6857
rect 30193 6848 30205 6851
rect 29604 6820 30205 6848
rect 29604 6808 29610 6820
rect 30193 6817 30205 6820
rect 30239 6817 30251 6851
rect 30193 6811 30251 6817
rect 30285 6851 30343 6857
rect 30285 6817 30297 6851
rect 30331 6817 30343 6851
rect 30285 6811 30343 6817
rect 30300 6780 30328 6811
rect 29411 6752 29500 6780
rect 29840 6752 30328 6780
rect 30745 6783 30803 6789
rect 29411 6749 29423 6752
rect 29365 6743 29423 6749
rect 25148 6712 25176 6740
rect 22066 6684 25176 6712
rect 26142 6672 26148 6724
rect 26200 6712 26206 6724
rect 26200 6684 26832 6712
rect 26200 6672 26206 6684
rect 24394 6644 24400 6656
rect 21928 6616 24400 6644
rect 24394 6604 24400 6616
rect 24452 6604 24458 6656
rect 24670 6604 24676 6656
rect 24728 6644 24734 6656
rect 24765 6647 24823 6653
rect 24765 6644 24777 6647
rect 24728 6616 24777 6644
rect 24728 6604 24734 6616
rect 24765 6613 24777 6616
rect 24811 6613 24823 6647
rect 24765 6607 24823 6613
rect 26234 6604 26240 6656
rect 26292 6604 26298 6656
rect 26804 6644 26832 6684
rect 26970 6672 26976 6724
rect 27028 6712 27034 6724
rect 27341 6715 27399 6721
rect 27341 6712 27353 6715
rect 27028 6684 27353 6712
rect 27028 6672 27034 6684
rect 27341 6681 27353 6684
rect 27387 6681 27399 6715
rect 27341 6675 27399 6681
rect 28350 6672 28356 6724
rect 28408 6672 28414 6724
rect 29840 6712 29868 6752
rect 30745 6749 30757 6783
rect 30791 6780 30803 6783
rect 31110 6780 31116 6792
rect 30791 6752 31116 6780
rect 30791 6749 30803 6752
rect 30745 6743 30803 6749
rect 31110 6740 31116 6752
rect 31168 6740 31174 6792
rect 36630 6740 36636 6792
rect 36688 6740 36694 6792
rect 28644 6684 29868 6712
rect 30101 6715 30159 6721
rect 28644 6644 28672 6684
rect 30101 6681 30113 6715
rect 30147 6712 30159 6715
rect 31297 6715 31355 6721
rect 31297 6712 31309 6715
rect 30147 6684 31309 6712
rect 30147 6681 30159 6684
rect 30101 6675 30159 6681
rect 31297 6681 31309 6684
rect 31343 6681 31355 6715
rect 31297 6675 31355 6681
rect 37274 6672 37280 6724
rect 37332 6712 37338 6724
rect 37369 6715 37427 6721
rect 37369 6712 37381 6715
rect 37332 6684 37381 6712
rect 37332 6672 37338 6684
rect 37369 6681 37381 6684
rect 37415 6681 37427 6715
rect 37369 6675 37427 6681
rect 26804 6616 28672 6644
rect 29178 6604 29184 6656
rect 29236 6604 29242 6656
rect 1104 6554 41400 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 41400 6554
rect 1104 6480 41400 6502
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6409 4491 6443
rect 4433 6403 4491 6409
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6304 4123 6307
rect 4448 6304 4476 6403
rect 4890 6400 4896 6452
rect 4948 6400 4954 6452
rect 8110 6440 8116 6452
rect 7760 6412 8116 6440
rect 4982 6332 4988 6384
rect 5040 6372 5046 6384
rect 6454 6372 6460 6384
rect 5040 6344 6460 6372
rect 5040 6332 5046 6344
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 7760 6372 7788 6412
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9766 6440 9772 6452
rect 9355 6412 9772 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 11238 6400 11244 6452
rect 11296 6400 11302 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 11388 6412 12357 6440
rect 11388 6400 11394 6412
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12345 6403 12403 6409
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12897 6443 12955 6449
rect 12897 6440 12909 6443
rect 12492 6412 12909 6440
rect 12492 6400 12498 6412
rect 12897 6409 12909 6412
rect 12943 6409 12955 6443
rect 12897 6403 12955 6409
rect 13814 6400 13820 6452
rect 13872 6400 13878 6452
rect 14090 6400 14096 6452
rect 14148 6400 14154 6452
rect 15473 6443 15531 6449
rect 15473 6409 15485 6443
rect 15519 6409 15531 6443
rect 15473 6403 15531 6409
rect 9401 6375 9459 6381
rect 7024 6344 7866 6372
rect 4111 6276 4476 6304
rect 4801 6307 4859 6313
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 5905 6307 5963 6313
rect 5905 6304 5917 6307
rect 4847 6276 5917 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 5905 6273 5917 6276
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 7024 6304 7052 6344
rect 9401 6341 9413 6375
rect 9447 6372 9459 6375
rect 11256 6372 11284 6400
rect 14108 6372 14136 6400
rect 9447 6344 11284 6372
rect 13096 6344 14136 6372
rect 9447 6341 9459 6344
rect 9401 6335 9459 6341
rect 9582 6304 9588 6316
rect 6052 6276 7052 6304
rect 9508 6276 9588 6304
rect 6052 6264 6058 6276
rect 4982 6196 4988 6248
rect 5040 6196 5046 6248
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6205 5319 6239
rect 5261 6199 5319 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6205 7159 6239
rect 7101 6199 7159 6205
rect 5276 6168 5304 6199
rect 5000 6140 5304 6168
rect 5000 6112 5028 6140
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 4982 6060 4988 6112
rect 5040 6060 5046 6112
rect 7116 6100 7144 6199
rect 7374 6196 7380 6248
rect 7432 6196 7438 6248
rect 9508 6245 9536 6276
rect 9582 6264 9588 6276
rect 9640 6308 9646 6316
rect 13096 6313 13124 6344
rect 9640 6304 9720 6308
rect 13081 6307 13139 6313
rect 9640 6280 11836 6304
rect 9640 6264 9646 6280
rect 9692 6276 11836 6280
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 9493 6199 9551 6205
rect 11698 6196 11704 6248
rect 11756 6196 11762 6248
rect 11808 6236 11836 6276
rect 13081 6273 13093 6307
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15488 6304 15516 6403
rect 15838 6400 15844 6452
rect 15896 6400 15902 6452
rect 15930 6400 15936 6452
rect 15988 6400 15994 6452
rect 17954 6440 17960 6452
rect 16776 6412 17960 6440
rect 16776 6313 16804 6412
rect 17954 6400 17960 6412
rect 18012 6440 18018 6452
rect 18012 6412 18644 6440
rect 18012 6400 18018 6412
rect 15335 6276 15516 6304
rect 16761 6307 16819 6313
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 16761 6273 16773 6307
rect 16807 6273 16819 6307
rect 16761 6267 16819 6273
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18616 6313 18644 6412
rect 20162 6400 20168 6452
rect 20220 6440 20226 6452
rect 20349 6443 20407 6449
rect 20349 6440 20361 6443
rect 20220 6412 20361 6440
rect 20220 6400 20226 6412
rect 20349 6409 20361 6412
rect 20395 6409 20407 6443
rect 20349 6403 20407 6409
rect 21358 6400 21364 6452
rect 21416 6440 21422 6452
rect 22370 6440 22376 6452
rect 21416 6412 22376 6440
rect 21416 6400 21422 6412
rect 22370 6400 22376 6412
rect 22428 6400 22434 6452
rect 26142 6440 26148 6452
rect 22480 6412 26148 6440
rect 22480 6372 22508 6412
rect 26142 6400 26148 6412
rect 26200 6400 26206 6452
rect 26234 6400 26240 6452
rect 26292 6400 26298 6452
rect 26970 6400 26976 6452
rect 27028 6400 27034 6452
rect 28534 6440 28540 6452
rect 27632 6412 28540 6440
rect 22204 6344 22508 6372
rect 23782 6344 24716 6372
rect 18601 6307 18659 6313
rect 18104 6276 18170 6304
rect 18104 6264 18110 6276
rect 18601 6273 18613 6307
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 19978 6264 19984 6316
rect 20036 6304 20042 6316
rect 21174 6304 21180 6316
rect 20036 6276 21180 6304
rect 20036 6264 20042 6276
rect 21174 6264 21180 6276
rect 21232 6264 21238 6316
rect 11808 6208 15884 6236
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 13078 6168 13084 6180
rect 8444 6140 13084 6168
rect 8444 6128 8450 6140
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 7742 6100 7748 6112
rect 7116 6072 7748 6100
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 8846 6060 8852 6112
rect 8904 6060 8910 6112
rect 8938 6060 8944 6112
rect 8996 6060 9002 6112
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 14182 6100 14188 6112
rect 12216 6072 14188 6100
rect 12216 6060 12222 6072
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 15068 6072 15117 6100
rect 15068 6060 15074 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15856 6100 15884 6208
rect 16022 6196 16028 6248
rect 16080 6196 16086 6248
rect 17034 6196 17040 6248
rect 17092 6196 17098 6248
rect 18874 6196 18880 6248
rect 18932 6196 18938 6248
rect 18509 6171 18567 6177
rect 18509 6137 18521 6171
rect 18555 6168 18567 6171
rect 18598 6168 18604 6180
rect 18555 6140 18604 6168
rect 18555 6137 18567 6140
rect 18509 6131 18567 6137
rect 18598 6128 18604 6140
rect 18656 6128 18662 6180
rect 21818 6128 21824 6180
rect 21876 6168 21882 6180
rect 22094 6168 22100 6180
rect 21876 6140 22100 6168
rect 21876 6128 21882 6140
rect 22094 6128 22100 6140
rect 22152 6128 22158 6180
rect 22204 6100 22232 6344
rect 24688 6316 24716 6344
rect 24213 6307 24271 6313
rect 24213 6304 24225 6307
rect 24044 6276 24225 6304
rect 22278 6196 22284 6248
rect 22336 6196 22342 6248
rect 22554 6196 22560 6248
rect 22612 6196 22618 6248
rect 24044 6245 24072 6276
rect 24213 6273 24225 6276
rect 24259 6304 24271 6307
rect 24578 6304 24584 6316
rect 24259 6276 24584 6304
rect 24259 6273 24271 6276
rect 24213 6267 24271 6273
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 24670 6264 24676 6316
rect 24728 6264 24734 6316
rect 26252 6304 26280 6400
rect 27632 6381 27660 6412
rect 28534 6400 28540 6412
rect 28592 6400 28598 6452
rect 29086 6400 29092 6452
rect 29144 6400 29150 6452
rect 29178 6400 29184 6452
rect 29236 6440 29242 6452
rect 36909 6443 36967 6449
rect 29236 6412 29592 6440
rect 29236 6400 29242 6412
rect 29564 6381 29592 6412
rect 36909 6409 36921 6443
rect 36955 6440 36967 6443
rect 36955 6412 37596 6440
rect 36955 6409 36967 6412
rect 36909 6403 36967 6409
rect 37568 6381 37596 6412
rect 27617 6375 27675 6381
rect 27617 6341 27629 6375
rect 27663 6341 27675 6375
rect 27617 6335 27675 6341
rect 29549 6375 29607 6381
rect 29549 6341 29561 6375
rect 29595 6341 29607 6375
rect 29549 6335 29607 6341
rect 37553 6375 37611 6381
rect 37553 6341 37565 6375
rect 37599 6341 37611 6375
rect 38838 6372 38844 6384
rect 38778 6344 38844 6372
rect 37553 6335 37611 6341
rect 38838 6332 38844 6344
rect 38896 6332 38902 6384
rect 27157 6307 27215 6313
rect 27157 6304 27169 6307
rect 26252 6276 27169 6304
rect 27157 6273 27169 6276
rect 27203 6273 27215 6307
rect 27157 6267 27215 6273
rect 28718 6264 28724 6316
rect 28776 6264 28782 6316
rect 29270 6264 29276 6316
rect 29328 6264 29334 6316
rect 24029 6239 24087 6245
rect 24029 6205 24041 6239
rect 24075 6205 24087 6239
rect 24029 6199 24087 6205
rect 24854 6196 24860 6248
rect 24912 6196 24918 6248
rect 27341 6239 27399 6245
rect 27341 6205 27353 6239
rect 27387 6205 27399 6239
rect 27341 6199 27399 6205
rect 15856 6072 22232 6100
rect 22296 6100 22324 6196
rect 22922 6100 22928 6112
rect 22296 6072 22928 6100
rect 15105 6063 15163 6069
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 23750 6060 23756 6112
rect 23808 6100 23814 6112
rect 24765 6103 24823 6109
rect 24765 6100 24777 6103
rect 23808 6072 24777 6100
rect 23808 6060 23814 6072
rect 24765 6069 24777 6072
rect 24811 6069 24823 6103
rect 24765 6063 24823 6069
rect 25498 6060 25504 6112
rect 25556 6060 25562 6112
rect 26510 6060 26516 6112
rect 26568 6100 26574 6112
rect 27062 6100 27068 6112
rect 26568 6072 27068 6100
rect 26568 6060 26574 6072
rect 27062 6060 27068 6072
rect 27120 6100 27126 6112
rect 27356 6100 27384 6199
rect 28350 6196 28356 6248
rect 28408 6236 28414 6248
rect 30668 6236 30696 6290
rect 34606 6264 34612 6316
rect 34664 6264 34670 6316
rect 37090 6264 37096 6316
rect 37148 6264 37154 6316
rect 28408 6208 30696 6236
rect 34624 6236 34652 6264
rect 37274 6236 37280 6248
rect 34624 6208 37280 6236
rect 28408 6196 28414 6208
rect 37274 6196 37280 6208
rect 37332 6196 37338 6248
rect 39025 6239 39083 6245
rect 39025 6205 39037 6239
rect 39071 6236 39083 6239
rect 39209 6239 39267 6245
rect 39209 6236 39221 6239
rect 39071 6208 39221 6236
rect 39071 6205 39083 6208
rect 39025 6199 39083 6205
rect 39209 6205 39221 6208
rect 39255 6236 39267 6239
rect 40678 6236 40684 6248
rect 39255 6208 40684 6236
rect 39255 6205 39267 6208
rect 39209 6199 39267 6205
rect 40678 6196 40684 6208
rect 40736 6196 40742 6248
rect 29270 6128 29276 6180
rect 29328 6128 29334 6180
rect 29288 6100 29316 6128
rect 27120 6072 29316 6100
rect 31021 6103 31079 6109
rect 27120 6060 27126 6072
rect 31021 6069 31033 6103
rect 31067 6100 31079 6103
rect 31110 6100 31116 6112
rect 31067 6072 31116 6100
rect 31067 6069 31079 6072
rect 31021 6063 31079 6069
rect 31110 6060 31116 6072
rect 31168 6060 31174 6112
rect 39758 6060 39764 6112
rect 39816 6060 39822 6112
rect 1104 6010 41400 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 41400 6010
rect 1104 5936 41400 5958
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7432 5868 8033 5896
rect 7432 5856 7438 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 10492 5899 10550 5905
rect 10492 5865 10504 5899
rect 10538 5896 10550 5899
rect 10962 5896 10968 5908
rect 10538 5868 10968 5896
rect 10538 5865 10550 5868
rect 10492 5859 10550 5865
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 16393 5899 16451 5905
rect 13228 5868 15976 5896
rect 13228 5856 13234 5868
rect 7742 5720 7748 5772
rect 7800 5720 7806 5772
rect 5074 5652 5080 5704
rect 5132 5652 5138 5704
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8956 5692 8984 5856
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5760 10287 5763
rect 10594 5760 10600 5772
rect 10275 5732 10600 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 13464 5760 13492 5868
rect 15948 5828 15976 5868
rect 16393 5865 16405 5899
rect 16439 5896 16451 5899
rect 16574 5896 16580 5908
rect 16439 5868 16580 5896
rect 16439 5865 16451 5868
rect 16393 5859 16451 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 17034 5856 17040 5908
rect 17092 5896 17098 5908
rect 17589 5899 17647 5905
rect 17589 5896 17601 5899
rect 17092 5868 17601 5896
rect 17092 5856 17098 5868
rect 17589 5865 17601 5868
rect 17635 5865 17647 5899
rect 17589 5859 17647 5865
rect 17972 5868 21312 5896
rect 17972 5828 18000 5868
rect 15948 5800 18000 5828
rect 13372 5732 13492 5760
rect 8251 5664 8984 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 11790 5692 11796 5704
rect 11664 5664 11796 5692
rect 11664 5652 11670 5664
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 5353 5627 5411 5633
rect 5353 5593 5365 5627
rect 5399 5624 5411 5627
rect 5626 5624 5632 5636
rect 5399 5596 5632 5624
rect 5399 5593 5411 5596
rect 5353 5587 5411 5593
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 5994 5584 6000 5636
rect 6052 5584 6058 5636
rect 13372 5624 13400 5732
rect 13538 5720 13544 5772
rect 13596 5760 13602 5772
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 13596 5732 13645 5760
rect 13596 5720 13602 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 14182 5720 14188 5772
rect 14240 5720 14246 5772
rect 14921 5763 14979 5769
rect 14921 5729 14933 5763
rect 14967 5760 14979 5763
rect 15010 5760 15016 5772
rect 14967 5732 15016 5760
rect 14967 5729 14979 5732
rect 14921 5723 14979 5729
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 17862 5760 17868 5772
rect 17788 5732 17868 5760
rect 14200 5692 14228 5720
rect 17788 5701 17816 5732
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5760 19855 5763
rect 20070 5760 20076 5772
rect 19843 5732 20076 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 20070 5720 20076 5732
rect 20128 5720 20134 5772
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 14200 5664 14657 5692
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 21174 5652 21180 5704
rect 21232 5652 21238 5704
rect 21284 5692 21312 5868
rect 21450 5856 21456 5908
rect 21508 5896 21514 5908
rect 21545 5899 21603 5905
rect 21545 5896 21557 5899
rect 21508 5868 21557 5896
rect 21508 5856 21514 5868
rect 21545 5865 21557 5868
rect 21591 5865 21603 5899
rect 21545 5859 21603 5865
rect 21560 5760 21588 5859
rect 22554 5856 22560 5908
rect 22612 5896 22618 5908
rect 22741 5899 22799 5905
rect 22741 5896 22753 5899
rect 22612 5868 22753 5896
rect 22612 5856 22618 5868
rect 22741 5865 22753 5868
rect 22787 5865 22799 5899
rect 22741 5859 22799 5865
rect 37090 5856 37096 5908
rect 37148 5896 37154 5908
rect 37185 5899 37243 5905
rect 37185 5896 37197 5899
rect 37148 5868 37197 5896
rect 37148 5856 37154 5868
rect 37185 5865 37197 5868
rect 37231 5865 37243 5899
rect 37185 5859 37243 5865
rect 39758 5856 39764 5908
rect 39816 5856 39822 5908
rect 23017 5831 23075 5837
rect 23017 5797 23029 5831
rect 23063 5797 23075 5831
rect 23017 5791 23075 5797
rect 21637 5763 21695 5769
rect 21637 5760 21649 5763
rect 21560 5732 21649 5760
rect 21637 5729 21649 5732
rect 21683 5729 21695 5763
rect 21637 5723 21695 5729
rect 22925 5695 22983 5701
rect 21284 5664 22094 5692
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 13372 5596 13553 5624
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 13541 5587 13599 5593
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 14550 5624 14556 5636
rect 13872 5596 14556 5624
rect 13872 5584 13878 5596
rect 14550 5584 14556 5596
rect 14608 5624 14614 5636
rect 20073 5627 20131 5633
rect 14608 5596 15410 5624
rect 14608 5584 14614 5596
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 6825 5559 6883 5565
rect 6825 5556 6837 5559
rect 6788 5528 6837 5556
rect 6788 5516 6794 5528
rect 6825 5525 6837 5528
rect 6871 5525 6883 5559
rect 6825 5519 6883 5525
rect 11974 5516 11980 5568
rect 12032 5516 12038 5568
rect 13078 5516 13084 5568
rect 13136 5516 13142 5568
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 13906 5556 13912 5568
rect 13495 5528 13912 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 15304 5556 15332 5596
rect 20073 5593 20085 5627
rect 20119 5624 20131 5627
rect 20162 5624 20168 5636
rect 20119 5596 20168 5624
rect 20119 5593 20131 5596
rect 20073 5587 20131 5593
rect 20162 5584 20168 5596
rect 20220 5584 20226 5636
rect 22066 5624 22094 5664
rect 22925 5661 22937 5695
rect 22971 5692 22983 5695
rect 23032 5692 23060 5791
rect 29270 5788 29276 5840
rect 29328 5828 29334 5840
rect 29328 5800 31616 5828
rect 29328 5788 29334 5800
rect 23106 5720 23112 5772
rect 23164 5760 23170 5772
rect 23569 5763 23627 5769
rect 23569 5760 23581 5763
rect 23164 5732 23581 5760
rect 23164 5720 23170 5732
rect 23569 5729 23581 5732
rect 23615 5729 23627 5763
rect 23569 5723 23627 5729
rect 23952 5732 24532 5760
rect 22971 5664 23060 5692
rect 22971 5661 22983 5664
rect 22925 5655 22983 5661
rect 23477 5627 23535 5633
rect 23477 5624 23489 5627
rect 22066 5596 23489 5624
rect 23477 5593 23489 5596
rect 23523 5624 23535 5627
rect 23952 5624 23980 5732
rect 24029 5695 24087 5701
rect 24029 5661 24041 5695
rect 24075 5692 24087 5695
rect 24075 5664 24440 5692
rect 24075 5661 24087 5664
rect 24029 5655 24087 5661
rect 23523 5596 23980 5624
rect 23523 5593 23535 5596
rect 23477 5587 23535 5593
rect 17954 5556 17960 5568
rect 15304 5528 17960 5556
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 22278 5516 22284 5568
rect 22336 5516 22342 5568
rect 23385 5559 23443 5565
rect 23385 5525 23397 5559
rect 23431 5556 23443 5559
rect 23750 5556 23756 5568
rect 23431 5528 23756 5556
rect 23431 5525 23443 5528
rect 23385 5519 23443 5525
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 23842 5516 23848 5568
rect 23900 5516 23906 5568
rect 24412 5565 24440 5664
rect 24504 5624 24532 5732
rect 24578 5720 24584 5772
rect 24636 5760 24642 5772
rect 25041 5763 25099 5769
rect 25041 5760 25053 5763
rect 24636 5732 25053 5760
rect 24636 5720 24642 5732
rect 25041 5729 25053 5732
rect 25087 5760 25099 5763
rect 25774 5760 25780 5772
rect 25087 5732 25780 5760
rect 25087 5729 25099 5732
rect 25041 5723 25099 5729
rect 25774 5720 25780 5732
rect 25832 5720 25838 5772
rect 26510 5720 26516 5772
rect 26568 5720 26574 5772
rect 30466 5720 30472 5772
rect 30524 5760 30530 5772
rect 31205 5763 31263 5769
rect 31205 5760 31217 5763
rect 30524 5732 31217 5760
rect 30524 5720 30530 5732
rect 31205 5729 31217 5732
rect 31251 5729 31263 5763
rect 31205 5723 31263 5729
rect 31294 5720 31300 5772
rect 31352 5720 31358 5772
rect 31588 5769 31616 5800
rect 32858 5788 32864 5840
rect 32916 5828 32922 5840
rect 32916 5800 35296 5828
rect 32916 5788 32922 5800
rect 31573 5763 31631 5769
rect 31573 5729 31585 5763
rect 31619 5729 31631 5763
rect 33042 5760 33048 5772
rect 31573 5723 31631 5729
rect 32968 5732 33048 5760
rect 24765 5695 24823 5701
rect 24765 5661 24777 5695
rect 24811 5692 24823 5695
rect 25498 5692 25504 5704
rect 24811 5664 25504 5692
rect 24811 5661 24823 5664
rect 24765 5655 24823 5661
rect 25498 5652 25504 5664
rect 25556 5652 25562 5704
rect 25685 5695 25743 5701
rect 25685 5661 25697 5695
rect 25731 5692 25743 5695
rect 28810 5692 28816 5704
rect 25731 5664 28816 5692
rect 25731 5661 25743 5664
rect 25685 5655 25743 5661
rect 28810 5652 28816 5664
rect 28868 5652 28874 5704
rect 30760 5664 31524 5692
rect 32968 5678 32996 5732
rect 33042 5720 33048 5732
rect 33100 5720 33106 5772
rect 33321 5763 33379 5769
rect 33321 5729 33333 5763
rect 33367 5760 33379 5763
rect 33367 5732 34744 5760
rect 33367 5729 33379 5732
rect 33321 5723 33379 5729
rect 24857 5627 24915 5633
rect 24857 5624 24869 5627
rect 24504 5596 24869 5624
rect 24857 5593 24869 5596
rect 24903 5624 24915 5627
rect 25038 5624 25044 5636
rect 24903 5596 25044 5624
rect 24903 5593 24915 5596
rect 24857 5587 24915 5593
rect 25038 5584 25044 5596
rect 25096 5584 25102 5636
rect 30760 5565 30788 5664
rect 31496 5624 31524 5664
rect 31754 5624 31760 5636
rect 31128 5596 31432 5624
rect 31496 5596 31760 5624
rect 31128 5565 31156 5596
rect 24397 5559 24455 5565
rect 24397 5525 24409 5559
rect 24443 5525 24455 5559
rect 24397 5519 24455 5525
rect 30745 5559 30803 5565
rect 30745 5525 30757 5559
rect 30791 5525 30803 5559
rect 30745 5519 30803 5525
rect 31113 5559 31171 5565
rect 31113 5525 31125 5559
rect 31159 5525 31171 5559
rect 31404 5556 31432 5596
rect 31754 5584 31760 5596
rect 31812 5584 31818 5636
rect 31846 5584 31852 5636
rect 31904 5584 31910 5636
rect 33336 5556 33364 5723
rect 34716 5704 34744 5732
rect 34790 5720 34796 5772
rect 34848 5760 34854 5772
rect 35161 5763 35219 5769
rect 35161 5760 35173 5763
rect 34848 5732 35173 5760
rect 34848 5720 34854 5732
rect 35161 5729 35173 5732
rect 35207 5729 35219 5763
rect 35161 5723 35219 5729
rect 34698 5652 34704 5704
rect 34756 5652 34762 5704
rect 35268 5692 35296 5800
rect 35345 5763 35403 5769
rect 35345 5729 35357 5763
rect 35391 5760 35403 5763
rect 35618 5760 35624 5772
rect 35391 5732 35624 5760
rect 35391 5729 35403 5732
rect 35345 5723 35403 5729
rect 35618 5720 35624 5732
rect 35676 5760 35682 5772
rect 37737 5763 37795 5769
rect 37737 5760 37749 5763
rect 35676 5732 37749 5760
rect 35676 5720 35682 5732
rect 37737 5729 37749 5732
rect 37783 5760 37795 5763
rect 37826 5760 37832 5772
rect 37783 5732 37832 5760
rect 37783 5729 37795 5732
rect 37737 5723 37795 5729
rect 37826 5720 37832 5732
rect 37884 5720 37890 5772
rect 34992 5664 35296 5692
rect 35805 5695 35863 5701
rect 31404 5528 33364 5556
rect 31113 5519 31171 5525
rect 34514 5516 34520 5568
rect 34572 5556 34578 5568
rect 34701 5559 34759 5565
rect 34701 5556 34713 5559
rect 34572 5528 34713 5556
rect 34572 5516 34578 5528
rect 34701 5525 34713 5528
rect 34747 5525 34759 5559
rect 34992 5556 35020 5664
rect 35805 5661 35817 5695
rect 35851 5692 35863 5695
rect 36262 5692 36268 5704
rect 35851 5664 36268 5692
rect 35851 5661 35863 5664
rect 35805 5655 35863 5661
rect 36262 5652 36268 5664
rect 36320 5652 36326 5704
rect 37553 5695 37611 5701
rect 37553 5661 37565 5695
rect 37599 5692 37611 5695
rect 39776 5692 39804 5856
rect 37599 5664 39804 5692
rect 37599 5661 37611 5664
rect 37553 5655 37611 5661
rect 35069 5627 35127 5633
rect 35069 5593 35081 5627
rect 35115 5624 35127 5627
rect 36357 5627 36415 5633
rect 36357 5624 36369 5627
rect 35115 5596 36369 5624
rect 35115 5593 35127 5596
rect 35069 5587 35127 5593
rect 36357 5593 36369 5596
rect 36403 5593 36415 5627
rect 36357 5587 36415 5593
rect 37645 5559 37703 5565
rect 37645 5556 37657 5559
rect 34992 5528 37657 5556
rect 34701 5519 34759 5525
rect 37645 5525 37657 5528
rect 37691 5525 37703 5559
rect 37645 5519 37703 5525
rect 1104 5466 41400 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 41400 5466
rect 1104 5392 41400 5414
rect 3878 5352 3884 5364
rect 3528 5324 3884 5352
rect 3528 5293 3556 5324
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 5626 5312 5632 5364
rect 5684 5312 5690 5364
rect 6365 5355 6423 5361
rect 6365 5321 6377 5355
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 8386 5352 8392 5364
rect 6871 5324 8392 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 3513 5287 3571 5293
rect 3513 5253 3525 5287
rect 3559 5253 3571 5287
rect 5994 5284 6000 5296
rect 4738 5256 6000 5284
rect 3513 5247 3571 5253
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 5074 5176 5080 5228
rect 5132 5176 5138 5228
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 6380 5216 6408 5315
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 11057 5355 11115 5361
rect 11057 5321 11069 5355
rect 11103 5352 11115 5355
rect 12710 5352 12716 5364
rect 11103 5324 12716 5352
rect 11103 5321 11115 5324
rect 11057 5315 11115 5321
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 17310 5352 17316 5364
rect 13964 5324 17316 5352
rect 13964 5312 13970 5324
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 20162 5312 20168 5364
rect 20220 5352 20226 5364
rect 20257 5355 20315 5361
rect 20257 5352 20269 5355
rect 20220 5324 20269 5352
rect 20220 5312 20226 5324
rect 20257 5321 20269 5324
rect 20303 5321 20315 5355
rect 20257 5315 20315 5321
rect 20530 5312 20536 5364
rect 20588 5312 20594 5364
rect 20901 5355 20959 5361
rect 20901 5321 20913 5355
rect 20947 5352 20959 5355
rect 22278 5352 22284 5364
rect 20947 5324 22284 5352
rect 20947 5321 20959 5324
rect 20901 5315 20959 5321
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 23842 5352 23848 5364
rect 23216 5324 23848 5352
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 13814 5284 13820 5296
rect 6512 5256 11192 5284
rect 13662 5256 13820 5284
rect 6512 5244 6518 5256
rect 5859 5188 6408 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 5092 5148 5120 5176
rect 3283 5120 5120 5148
rect 6656 5148 6684 5256
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 6779 5188 7849 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10551 5188 10977 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11164 5157 11192 5256
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 20548 5284 20576 5312
rect 23106 5284 23112 5296
rect 20548 5256 23112 5284
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6656 5120 6929 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 9953 5151 10011 5157
rect 9953 5117 9965 5151
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 11149 5151 11207 5157
rect 11149 5117 11161 5151
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 4982 4972 4988 5024
rect 5040 4972 5046 5024
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 6730 5012 6736 5024
rect 5592 4984 6736 5012
rect 5592 4972 5598 4984
rect 6730 4972 6736 4984
rect 6788 5012 6794 5024
rect 7208 5012 7236 5111
rect 6788 4984 7236 5012
rect 9968 5012 9996 5111
rect 10597 5083 10655 5089
rect 10597 5049 10609 5083
rect 10643 5080 10655 5083
rect 11716 5080 11744 5179
rect 12158 5176 12164 5228
rect 12216 5176 12222 5228
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5216 20499 5219
rect 20487 5188 20576 5216
rect 20487 5185 20499 5188
rect 20441 5179 20499 5185
rect 12434 5108 12440 5160
rect 12492 5108 12498 5160
rect 20548 5089 20576 5188
rect 20898 5176 20904 5228
rect 20956 5216 20962 5228
rect 21008 5216 21036 5256
rect 23106 5244 23112 5256
rect 23164 5244 23170 5296
rect 23216 5293 23244 5324
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 24765 5355 24823 5361
rect 24765 5321 24777 5355
rect 24811 5321 24823 5355
rect 24765 5315 24823 5321
rect 23201 5287 23259 5293
rect 23201 5253 23213 5287
rect 23247 5253 23259 5287
rect 24670 5284 24676 5296
rect 24426 5256 24676 5284
rect 23201 5247 23259 5253
rect 24670 5244 24676 5256
rect 24728 5244 24734 5296
rect 24780 5284 24808 5315
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 25130 5352 25136 5364
rect 25004 5324 25136 5352
rect 25004 5312 25010 5324
rect 25130 5312 25136 5324
rect 25188 5352 25194 5364
rect 26789 5355 26847 5361
rect 26789 5352 26801 5355
rect 25188 5324 26801 5352
rect 25188 5312 25194 5324
rect 26789 5321 26801 5324
rect 26835 5352 26847 5355
rect 27706 5352 27712 5364
rect 26835 5324 27712 5352
rect 26835 5321 26847 5324
rect 26789 5315 26847 5321
rect 27706 5312 27712 5324
rect 27764 5312 27770 5364
rect 31665 5355 31723 5361
rect 31665 5321 31677 5355
rect 31711 5352 31723 5355
rect 31846 5352 31852 5364
rect 31711 5324 31852 5352
rect 31711 5321 31723 5324
rect 31665 5315 31723 5321
rect 31846 5312 31852 5324
rect 31904 5312 31910 5364
rect 34514 5352 34520 5364
rect 34440 5324 34520 5352
rect 25317 5287 25375 5293
rect 25317 5284 25329 5287
rect 24780 5256 25329 5284
rect 25317 5253 25329 5256
rect 25363 5253 25375 5287
rect 25317 5247 25375 5253
rect 20956 5188 21128 5216
rect 20956 5176 20962 5188
rect 21100 5157 21128 5188
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 24946 5176 24952 5228
rect 25004 5176 25010 5228
rect 26602 5216 26608 5228
rect 26450 5188 26608 5216
rect 26602 5176 26608 5188
rect 26660 5216 26666 5228
rect 28350 5216 28356 5228
rect 26660 5188 28356 5216
rect 26660 5176 26666 5188
rect 28350 5176 28356 5188
rect 28408 5176 28414 5228
rect 31754 5176 31760 5228
rect 31812 5216 31818 5228
rect 34440 5225 34468 5324
rect 34514 5312 34520 5324
rect 34572 5312 34578 5364
rect 34606 5312 34612 5364
rect 34664 5312 34670 5364
rect 34624 5284 34652 5312
rect 38838 5284 38844 5296
rect 34532 5256 34652 5284
rect 36018 5256 38844 5284
rect 34532 5225 34560 5256
rect 38838 5244 38844 5256
rect 38896 5244 38902 5296
rect 31849 5219 31907 5225
rect 31849 5216 31861 5219
rect 31812 5188 31861 5216
rect 31812 5176 31818 5188
rect 31849 5185 31861 5188
rect 31895 5185 31907 5219
rect 31849 5179 31907 5185
rect 34425 5219 34483 5225
rect 34425 5185 34437 5219
rect 34471 5185 34483 5219
rect 34425 5179 34483 5185
rect 34517 5219 34575 5225
rect 34517 5185 34529 5219
rect 34563 5185 34575 5219
rect 34517 5179 34575 5185
rect 20993 5151 21051 5157
rect 20993 5117 21005 5151
rect 21039 5117 21051 5151
rect 20993 5111 21051 5117
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5117 21143 5151
rect 22940 5148 22968 5176
rect 23290 5148 23296 5160
rect 22940 5120 23296 5148
rect 21085 5111 21143 5117
rect 10643 5052 11744 5080
rect 20533 5083 20591 5089
rect 10643 5049 10655 5052
rect 10597 5043 10655 5049
rect 20533 5049 20545 5083
rect 20579 5049 20591 5083
rect 21008 5080 21036 5111
rect 23290 5108 23296 5120
rect 23348 5108 23354 5160
rect 24673 5151 24731 5157
rect 24673 5117 24685 5151
rect 24719 5148 24731 5151
rect 24854 5148 24860 5160
rect 24719 5120 24860 5148
rect 24719 5117 24731 5120
rect 24673 5111 24731 5117
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 25041 5151 25099 5157
rect 25041 5117 25053 5151
rect 25087 5148 25099 5151
rect 25314 5148 25320 5160
rect 25087 5120 25320 5148
rect 25087 5117 25099 5120
rect 25041 5111 25099 5117
rect 25314 5108 25320 5120
rect 25372 5148 25378 5160
rect 26510 5148 26516 5160
rect 25372 5120 26516 5148
rect 25372 5108 25378 5120
rect 26510 5108 26516 5120
rect 26568 5108 26574 5160
rect 34793 5151 34851 5157
rect 34793 5148 34805 5151
rect 34256 5120 34805 5148
rect 21358 5080 21364 5092
rect 21008 5052 21364 5080
rect 20533 5043 20591 5049
rect 21358 5040 21364 5052
rect 21416 5080 21422 5092
rect 21910 5080 21916 5092
rect 21416 5052 21916 5080
rect 21416 5040 21422 5052
rect 21910 5040 21916 5052
rect 21968 5040 21974 5092
rect 34256 5089 34284 5120
rect 34793 5117 34805 5120
rect 34839 5117 34851 5151
rect 34793 5111 34851 5117
rect 34241 5083 34299 5089
rect 34241 5049 34253 5083
rect 34287 5049 34299 5083
rect 34241 5043 34299 5049
rect 11330 5012 11336 5024
rect 9968 4984 11336 5012
rect 6788 4972 6794 4984
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 36262 4972 36268 5024
rect 36320 4972 36326 5024
rect 1104 4922 41400 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 41400 4922
rect 1104 4848 41400 4870
rect 10308 4811 10366 4817
rect 10308 4777 10320 4811
rect 10354 4808 10366 4811
rect 11514 4808 11520 4820
rect 10354 4780 11520 4808
rect 10354 4777 10366 4780
rect 10308 4771 10366 4777
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12621 4811 12679 4817
rect 12621 4808 12633 4811
rect 12492 4780 12633 4808
rect 12492 4768 12498 4780
rect 12621 4777 12633 4780
rect 12667 4777 12679 4811
rect 12621 4771 12679 4777
rect 18322 4768 18328 4820
rect 18380 4768 18386 4820
rect 24765 4811 24823 4817
rect 24765 4777 24777 4811
rect 24811 4808 24823 4811
rect 24946 4808 24952 4820
rect 24811 4780 24952 4808
rect 24811 4777 24823 4780
rect 24765 4771 24823 4777
rect 24946 4768 24952 4780
rect 25004 4768 25010 4820
rect 26510 4768 26516 4820
rect 26568 4768 26574 4820
rect 28074 4768 28080 4820
rect 28132 4808 28138 4820
rect 28169 4811 28227 4817
rect 28169 4808 28181 4811
rect 28132 4780 28181 4808
rect 28132 4768 28138 4780
rect 28169 4777 28181 4780
rect 28215 4777 28227 4811
rect 28169 4771 28227 4777
rect 36262 4768 36268 4820
rect 36320 4808 36326 4820
rect 36320 4780 40724 4808
rect 36320 4768 36326 4780
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11790 4740 11796 4752
rect 11388 4712 11796 4740
rect 11388 4700 11394 4712
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 12158 4672 12164 4684
rect 10091 4644 12164 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 18340 4672 18368 4768
rect 25593 4743 25651 4749
rect 25593 4709 25605 4743
rect 25639 4740 25651 4743
rect 26234 4740 26240 4752
rect 25639 4712 26240 4740
rect 25639 4709 25651 4712
rect 25593 4703 25651 4709
rect 26234 4700 26240 4712
rect 26292 4700 26298 4752
rect 18417 4675 18475 4681
rect 18417 4672 18429 4675
rect 18340 4644 18429 4672
rect 18417 4641 18429 4644
rect 18463 4641 18475 4675
rect 18417 4635 18475 4641
rect 20898 4632 20904 4684
rect 20956 4632 20962 4684
rect 21266 4632 21272 4684
rect 21324 4672 21330 4684
rect 21726 4672 21732 4684
rect 21324 4644 21732 4672
rect 21324 4632 21330 4644
rect 21726 4632 21732 4644
rect 21784 4632 21790 4684
rect 22002 4632 22008 4684
rect 22060 4632 22066 4684
rect 25038 4632 25044 4684
rect 25096 4672 25102 4684
rect 25225 4675 25283 4681
rect 25225 4672 25237 4675
rect 25096 4644 25237 4672
rect 25096 4632 25102 4644
rect 25225 4641 25237 4644
rect 25271 4641 25283 4675
rect 25225 4635 25283 4641
rect 25409 4675 25467 4681
rect 25409 4641 25421 4675
rect 25455 4641 25467 4675
rect 25409 4635 25467 4641
rect 11606 4604 11612 4616
rect 11454 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4604 12863 4607
rect 13078 4604 13084 4616
rect 12851 4576 13084 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 16574 4564 16580 4616
rect 16632 4564 16638 4616
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 19058 4604 19064 4616
rect 18012 4576 19064 4604
rect 18012 4564 18018 4576
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 20809 4607 20867 4613
rect 20809 4573 20821 4607
rect 20855 4604 20867 4607
rect 20990 4604 20996 4616
rect 20855 4576 20996 4604
rect 20855 4573 20867 4576
rect 20809 4567 20867 4573
rect 20990 4564 20996 4576
rect 21048 4604 21054 4616
rect 22020 4604 22048 4632
rect 21048 4576 22048 4604
rect 21048 4564 21054 4576
rect 25130 4564 25136 4616
rect 25188 4564 25194 4616
rect 25424 4604 25452 4635
rect 25958 4632 25964 4684
rect 26016 4672 26022 4684
rect 26053 4675 26111 4681
rect 26053 4672 26065 4675
rect 26016 4644 26065 4672
rect 26016 4632 26022 4644
rect 26053 4641 26065 4644
rect 26099 4641 26111 4675
rect 26053 4635 26111 4641
rect 26145 4675 26203 4681
rect 26145 4641 26157 4675
rect 26191 4672 26203 4675
rect 26326 4672 26332 4684
rect 26191 4644 26332 4672
rect 26191 4641 26203 4644
rect 26145 4635 26203 4641
rect 26160 4604 26188 4635
rect 26326 4632 26332 4644
rect 26384 4632 26390 4684
rect 26421 4675 26479 4681
rect 26421 4641 26433 4675
rect 26467 4672 26479 4675
rect 26528 4672 26556 4768
rect 36725 4743 36783 4749
rect 36725 4709 36737 4743
rect 36771 4740 36783 4743
rect 37458 4740 37464 4752
rect 36771 4712 37464 4740
rect 36771 4709 36783 4712
rect 36725 4703 36783 4709
rect 37458 4700 37464 4712
rect 37516 4700 37522 4752
rect 37660 4712 37872 4740
rect 37660 4681 37688 4712
rect 37844 4684 37872 4712
rect 26467 4644 26556 4672
rect 37645 4675 37703 4681
rect 26467 4641 26479 4644
rect 26421 4635 26479 4641
rect 37645 4641 37657 4675
rect 37691 4641 37703 4675
rect 37645 4635 37703 4641
rect 37734 4632 37740 4684
rect 37792 4632 37798 4684
rect 37826 4632 37832 4684
rect 37884 4632 37890 4684
rect 28350 4604 28356 4616
rect 25424 4576 26188 4604
rect 27830 4576 28356 4604
rect 28350 4564 28356 4576
rect 28408 4564 28414 4616
rect 36909 4607 36967 4613
rect 36909 4573 36921 4607
rect 36955 4604 36967 4607
rect 37461 4607 37519 4613
rect 36955 4576 37044 4604
rect 36955 4573 36967 4576
rect 36909 4567 36967 4573
rect 16850 4496 16856 4548
rect 16908 4496 16914 4548
rect 20717 4539 20775 4545
rect 20717 4505 20729 4539
rect 20763 4536 20775 4539
rect 21821 4539 21879 4545
rect 21821 4536 21833 4539
rect 20763 4508 21833 4536
rect 20763 4505 20775 4508
rect 20717 4499 20775 4505
rect 21821 4505 21833 4508
rect 21867 4505 21879 4539
rect 21821 4499 21879 4505
rect 25961 4539 26019 4545
rect 25961 4505 25973 4539
rect 26007 4536 26019 4539
rect 26007 4508 26648 4536
rect 26007 4505 26019 4508
rect 25961 4499 26019 4505
rect 18414 4428 18420 4480
rect 18472 4468 18478 4480
rect 19061 4471 19119 4477
rect 19061 4468 19073 4471
rect 18472 4440 19073 4468
rect 18472 4428 18478 4440
rect 19061 4437 19073 4440
rect 19107 4437 19119 4471
rect 19061 4431 19119 4437
rect 20346 4428 20352 4480
rect 20404 4428 20410 4480
rect 26620 4468 26648 4508
rect 26694 4496 26700 4548
rect 26752 4496 26758 4548
rect 28074 4496 28080 4548
rect 28132 4496 28138 4548
rect 28092 4468 28120 4496
rect 37016 4477 37044 4576
rect 37461 4573 37473 4607
rect 37507 4604 37519 4607
rect 37752 4604 37780 4632
rect 37507 4576 37780 4604
rect 38381 4607 38439 4613
rect 37507 4573 37519 4576
rect 37461 4567 37519 4573
rect 38381 4573 38393 4607
rect 38427 4604 38439 4607
rect 39022 4604 39028 4616
rect 38427 4576 39028 4604
rect 38427 4573 38439 4576
rect 38381 4567 38439 4573
rect 39022 4564 39028 4576
rect 39080 4564 39086 4616
rect 40696 4613 40724 4780
rect 40681 4607 40739 4613
rect 40681 4573 40693 4607
rect 40727 4573 40739 4607
rect 40681 4567 40739 4573
rect 37369 4539 37427 4545
rect 37369 4505 37381 4539
rect 37415 4536 37427 4539
rect 38933 4539 38991 4545
rect 38933 4536 38945 4539
rect 37415 4508 38945 4536
rect 37415 4505 37427 4508
rect 37369 4499 37427 4505
rect 38933 4505 38945 4508
rect 38979 4505 38991 4539
rect 38933 4499 38991 4505
rect 26620 4440 28120 4468
rect 37001 4471 37059 4477
rect 37001 4437 37013 4471
rect 37047 4437 37059 4471
rect 37001 4431 37059 4437
rect 40957 4471 41015 4477
rect 40957 4437 40969 4471
rect 41003 4468 41015 4471
rect 41046 4468 41052 4480
rect 41003 4440 41052 4468
rect 41003 4437 41015 4440
rect 40957 4431 41015 4437
rect 41046 4428 41052 4440
rect 41104 4428 41110 4480
rect 1104 4378 41400 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 41400 4378
rect 1104 4304 41400 4326
rect 14182 4224 14188 4276
rect 14240 4224 14246 4276
rect 15010 4224 15016 4276
rect 15068 4264 15074 4276
rect 15562 4264 15568 4276
rect 15068 4236 15568 4264
rect 15068 4224 15074 4236
rect 15562 4224 15568 4236
rect 15620 4224 15626 4276
rect 16025 4267 16083 4273
rect 16025 4233 16037 4267
rect 16071 4264 16083 4267
rect 16482 4264 16488 4276
rect 16071 4236 16488 4264
rect 16071 4233 16083 4236
rect 16025 4227 16083 4233
rect 16482 4224 16488 4236
rect 16540 4264 16546 4276
rect 16758 4264 16764 4276
rect 16540 4236 16764 4264
rect 16540 4224 16546 4236
rect 16758 4224 16764 4236
rect 16816 4224 16822 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 17037 4267 17095 4273
rect 17037 4264 17049 4267
rect 16908 4236 17049 4264
rect 16908 4224 16914 4236
rect 17037 4233 17049 4236
rect 17083 4233 17095 4267
rect 17037 4227 17095 4233
rect 17310 4224 17316 4276
rect 17368 4224 17374 4276
rect 17681 4267 17739 4273
rect 17681 4233 17693 4267
rect 17727 4264 17739 4267
rect 18414 4264 18420 4276
rect 17727 4236 18420 4264
rect 17727 4233 17739 4236
rect 17681 4227 17739 4233
rect 18414 4224 18420 4236
rect 18472 4224 18478 4276
rect 18690 4264 18696 4276
rect 18616 4236 18696 4264
rect 14200 4196 14228 4224
rect 13832 4168 14228 4196
rect 13722 4088 13728 4140
rect 13780 4128 13786 4140
rect 13832 4137 13860 4168
rect 14550 4156 14556 4208
rect 14608 4156 14614 4208
rect 16574 4156 16580 4208
rect 16632 4196 16638 4208
rect 18616 4205 18644 4236
rect 18690 4224 18696 4236
rect 18748 4224 18754 4276
rect 21082 4224 21088 4276
rect 21140 4264 21146 4276
rect 21269 4267 21327 4273
rect 21269 4264 21281 4267
rect 21140 4236 21281 4264
rect 21140 4224 21146 4236
rect 21269 4233 21281 4236
rect 21315 4233 21327 4267
rect 21269 4227 21327 4233
rect 21358 4224 21364 4276
rect 21416 4224 21422 4276
rect 22094 4224 22100 4276
rect 22152 4264 22158 4276
rect 22189 4267 22247 4273
rect 22189 4264 22201 4267
rect 22152 4236 22201 4264
rect 22152 4224 22158 4236
rect 22189 4233 22201 4236
rect 22235 4264 22247 4267
rect 24026 4264 24032 4276
rect 22235 4236 24032 4264
rect 22235 4233 22247 4236
rect 22189 4227 22247 4233
rect 24026 4224 24032 4236
rect 24084 4224 24090 4276
rect 26234 4224 26240 4276
rect 26292 4224 26298 4276
rect 26421 4267 26479 4273
rect 26421 4233 26433 4267
rect 26467 4264 26479 4267
rect 26694 4264 26700 4276
rect 26467 4236 26700 4264
rect 26467 4233 26479 4236
rect 26421 4227 26479 4233
rect 26694 4224 26700 4236
rect 26752 4224 26758 4276
rect 18601 4199 18659 4205
rect 16632 4168 18368 4196
rect 16632 4156 16638 4168
rect 18340 4140 18368 4168
rect 18601 4165 18613 4199
rect 18647 4165 18659 4199
rect 18601 4159 18659 4165
rect 19058 4156 19064 4208
rect 19116 4156 19122 4208
rect 21376 4196 21404 4224
rect 20180 4168 21404 4196
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13780 4100 13829 4128
rect 13780 4088 13786 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4128 16175 4131
rect 16163 4100 16896 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 14090 4020 14096 4072
rect 14148 4020 14154 4072
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4029 16267 4063
rect 16868 4060 16896 4100
rect 16942 4088 16948 4140
rect 17000 4088 17006 4140
rect 17221 4131 17279 4137
rect 17221 4097 17233 4131
rect 17267 4128 17279 4131
rect 17310 4128 17316 4140
rect 17267 4100 17316 4128
rect 17267 4097 17279 4100
rect 17221 4091 17279 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 17736 4100 17908 4128
rect 17736 4088 17742 4100
rect 17880 4069 17908 4100
rect 18322 4088 18328 4140
rect 18380 4088 18386 4140
rect 20180 4128 20208 4168
rect 19812 4100 20208 4128
rect 20257 4131 20315 4137
rect 17773 4063 17831 4069
rect 17773 4060 17785 4063
rect 16868 4032 17785 4060
rect 16209 4023 16267 4029
rect 17773 4029 17785 4032
rect 17819 4029 17831 4063
rect 17773 4023 17831 4029
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4029 17923 4063
rect 19812 4060 19840 4100
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 20438 4128 20444 4140
rect 20303 4100 20444 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 17865 4023 17923 4029
rect 18156 4032 19840 4060
rect 16224 3992 16252 4023
rect 15120 3964 16252 3992
rect 17788 3992 17816 4023
rect 18156 3992 18184 4032
rect 20070 4020 20076 4072
rect 20128 4020 20134 4072
rect 20088 3992 20116 4020
rect 17788 3964 18184 3992
rect 19628 3964 20116 3992
rect 15120 3936 15148 3964
rect 15102 3884 15108 3936
rect 15160 3884 15166 3936
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 16758 3884 16764 3936
rect 16816 3884 16822 3936
rect 18414 3884 18420 3936
rect 18472 3924 18478 3936
rect 19628 3924 19656 3964
rect 18472 3896 19656 3924
rect 20073 3927 20131 3933
rect 18472 3884 18478 3896
rect 20073 3893 20085 3927
rect 20119 3924 20131 3927
rect 20272 3924 20300 4091
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 22830 4128 22836 4140
rect 21560 4100 22836 4128
rect 21560 4069 21588 4100
rect 22480 4069 22508 4100
rect 22830 4088 22836 4100
rect 22888 4088 22894 4140
rect 24118 4088 24124 4140
rect 24176 4088 24182 4140
rect 25133 4131 25191 4137
rect 25133 4097 25145 4131
rect 25179 4128 25191 4131
rect 25222 4128 25228 4140
rect 25179 4100 25228 4128
rect 25179 4097 25191 4100
rect 25133 4091 25191 4097
rect 25222 4088 25228 4100
rect 25280 4088 25286 4140
rect 25682 4088 25688 4140
rect 25740 4128 25746 4140
rect 25961 4131 26019 4137
rect 25961 4128 25973 4131
rect 25740 4100 25973 4128
rect 25740 4088 25746 4100
rect 25961 4097 25973 4100
rect 26007 4097 26019 4131
rect 26252 4128 26280 4224
rect 37458 4156 37464 4208
rect 37516 4196 37522 4208
rect 37553 4199 37611 4205
rect 37553 4196 37565 4199
rect 37516 4168 37565 4196
rect 37516 4156 37522 4168
rect 37553 4165 37565 4168
rect 37599 4165 37611 4199
rect 38838 4196 38844 4208
rect 38778 4168 38844 4196
rect 37553 4159 37611 4165
rect 38838 4156 38844 4168
rect 38896 4156 38902 4208
rect 26605 4131 26663 4137
rect 26605 4128 26617 4131
rect 26252 4100 26617 4128
rect 25961 4091 26019 4097
rect 26605 4097 26617 4100
rect 26651 4097 26663 4131
rect 26605 4091 26663 4097
rect 37274 4088 37280 4140
rect 37332 4088 37338 4140
rect 21545 4063 21603 4069
rect 21545 4029 21557 4063
rect 21591 4029 21603 4063
rect 22281 4063 22339 4069
rect 22281 4060 22293 4063
rect 21545 4023 21603 4029
rect 22066 4032 22293 4060
rect 22066 4004 22094 4032
rect 22281 4029 22293 4032
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22511 4032 22545 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 24670 4020 24676 4072
rect 24728 4060 24734 4072
rect 24728 4032 26648 4060
rect 24728 4020 24734 4032
rect 26620 4004 26648 4032
rect 22002 3952 22008 4004
rect 22060 3964 22094 4004
rect 22060 3952 22066 3964
rect 25590 3952 25596 4004
rect 25648 3992 25654 4004
rect 25777 3995 25835 4001
rect 25777 3992 25789 3995
rect 25648 3964 25789 3992
rect 25648 3952 25654 3964
rect 25777 3961 25789 3964
rect 25823 3961 25835 3995
rect 25777 3955 25835 3961
rect 26602 3952 26608 4004
rect 26660 3952 26666 4004
rect 20119 3896 20300 3924
rect 20119 3893 20131 3896
rect 20073 3887 20131 3893
rect 20806 3884 20812 3936
rect 20864 3884 20870 3936
rect 20898 3884 20904 3936
rect 20956 3884 20962 3936
rect 21818 3884 21824 3936
rect 21876 3884 21882 3936
rect 23842 3884 23848 3936
rect 23900 3924 23906 3936
rect 23937 3927 23995 3933
rect 23937 3924 23949 3927
rect 23900 3896 23949 3924
rect 23900 3884 23906 3896
rect 23937 3893 23949 3896
rect 23983 3893 23995 3927
rect 23937 3887 23995 3893
rect 24762 3884 24768 3936
rect 24820 3924 24826 3936
rect 25685 3927 25743 3933
rect 25685 3924 25697 3927
rect 24820 3896 25697 3924
rect 24820 3884 24826 3896
rect 25685 3893 25697 3896
rect 25731 3893 25743 3927
rect 25685 3887 25743 3893
rect 39022 3884 39028 3936
rect 39080 3884 39086 3936
rect 1104 3834 41400 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 41400 3834
rect 1104 3760 41400 3782
rect 13538 3680 13544 3732
rect 13596 3680 13602 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14185 3723 14243 3729
rect 14185 3720 14197 3723
rect 14148 3692 14197 3720
rect 14148 3680 14154 3692
rect 14185 3689 14197 3692
rect 14231 3689 14243 3723
rect 14185 3683 14243 3689
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 15470 3720 15476 3732
rect 14608 3692 15476 3720
rect 14608 3680 14614 3692
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15654 3680 15660 3732
rect 15712 3680 15718 3732
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 17313 3723 17371 3729
rect 17313 3720 17325 3723
rect 17000 3692 17325 3720
rect 17000 3680 17006 3692
rect 17313 3689 17325 3692
rect 17359 3689 17371 3723
rect 17313 3683 17371 3689
rect 17678 3680 17684 3732
rect 17736 3720 17742 3732
rect 17736 3692 18092 3720
rect 17736 3680 17742 3692
rect 13556 3652 13584 3680
rect 15102 3652 15108 3664
rect 13556 3624 15108 3652
rect 13556 3584 13584 3624
rect 15028 3593 15056 3624
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 13556 3556 13737 3584
rect 13725 3553 13737 3556
rect 13771 3553 13783 3587
rect 15013 3587 15071 3593
rect 13725 3547 13783 3553
rect 14292 3556 14872 3584
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 5534 3516 5540 3528
rect 1535 3488 5540 3516
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 13541 3519 13599 3525
rect 13127 3488 13216 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 934 3340 940 3392
rect 992 3380 998 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 992 3352 1593 3380
rect 992 3340 998 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 12894 3340 12900 3392
rect 12952 3340 12958 3392
rect 13188 3389 13216 3488
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 14292 3516 14320 3556
rect 14844 3528 14872 3556
rect 15013 3553 15025 3587
rect 15059 3553 15071 3587
rect 15013 3547 15071 3553
rect 13587 3488 14320 3516
rect 14369 3519 14427 3525
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14415 3488 14504 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 13173 3383 13231 3389
rect 13173 3349 13185 3383
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 14366 3380 14372 3392
rect 13679 3352 14372 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 14476 3389 14504 3488
rect 14826 3476 14832 3528
rect 14884 3476 14890 3528
rect 14921 3519 14979 3525
rect 14921 3485 14933 3519
rect 14967 3516 14979 3519
rect 15473 3519 15531 3525
rect 14967 3488 15424 3516
rect 14967 3485 14979 3488
rect 14921 3479 14979 3485
rect 15010 3448 15016 3460
rect 14844 3420 15016 3448
rect 14844 3389 14872 3420
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 15396 3448 15424 3488
rect 15473 3485 15485 3519
rect 15519 3516 15531 3519
rect 15672 3516 15700 3680
rect 17037 3655 17095 3661
rect 17037 3621 17049 3655
rect 17083 3652 17095 3655
rect 17083 3624 17816 3652
rect 17083 3621 17095 3624
rect 17037 3615 17095 3621
rect 17788 3596 17816 3624
rect 17678 3544 17684 3596
rect 17736 3544 17742 3596
rect 17770 3544 17776 3596
rect 17828 3544 17834 3596
rect 17862 3544 17868 3596
rect 17920 3544 17926 3596
rect 18064 3584 18092 3692
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 18877 3723 18935 3729
rect 18877 3720 18889 3723
rect 18748 3692 18889 3720
rect 18748 3680 18754 3692
rect 18877 3689 18889 3692
rect 18923 3689 18935 3723
rect 20806 3720 20812 3732
rect 18877 3683 18935 3689
rect 19628 3692 20812 3720
rect 19245 3655 19303 3661
rect 19245 3621 19257 3655
rect 19291 3621 19303 3655
rect 19245 3615 19303 3621
rect 18064 3556 19012 3584
rect 15519 3488 15700 3516
rect 15519 3485 15531 3488
rect 15473 3479 15531 3485
rect 15746 3476 15752 3528
rect 15804 3476 15810 3528
rect 17696 3516 17724 3544
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17696 3488 18153 3516
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 15396 3420 16528 3448
rect 14461 3383 14519 3389
rect 14461 3349 14473 3383
rect 14507 3349 14519 3383
rect 14461 3343 14519 3349
rect 14829 3383 14887 3389
rect 14829 3349 14841 3383
rect 14875 3349 14887 3383
rect 14829 3343 14887 3349
rect 15286 3340 15292 3392
rect 15344 3340 15350 3392
rect 16500 3380 16528 3420
rect 16574 3408 16580 3460
rect 16632 3408 16638 3460
rect 17681 3451 17739 3457
rect 17681 3417 17693 3451
rect 17727 3448 17739 3451
rect 18785 3451 18843 3457
rect 18785 3448 18797 3451
rect 17727 3420 18797 3448
rect 17727 3417 17739 3420
rect 17681 3411 17739 3417
rect 18785 3417 18797 3420
rect 18831 3417 18843 3451
rect 18984 3448 19012 3556
rect 19061 3519 19119 3525
rect 19061 3485 19073 3519
rect 19107 3516 19119 3519
rect 19260 3516 19288 3615
rect 19628 3525 19656 3692
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 21082 3680 21088 3732
rect 21140 3720 21146 3732
rect 22189 3723 22247 3729
rect 22189 3720 22201 3723
rect 21140 3692 22201 3720
rect 21140 3680 21146 3692
rect 22189 3689 22201 3692
rect 22235 3689 22247 3723
rect 22189 3683 22247 3689
rect 22296 3692 23612 3720
rect 22296 3652 22324 3692
rect 19812 3624 20576 3652
rect 19812 3593 19840 3624
rect 19797 3587 19855 3593
rect 19797 3584 19809 3587
rect 19720 3556 19809 3584
rect 19107 3488 19288 3516
rect 19613 3519 19671 3525
rect 19107 3485 19119 3488
rect 19061 3479 19119 3485
rect 19613 3485 19625 3519
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 19720 3448 19748 3556
rect 19797 3553 19809 3556
rect 19843 3553 19855 3587
rect 19797 3547 19855 3553
rect 20070 3544 20076 3596
rect 20128 3584 20134 3596
rect 20441 3587 20499 3593
rect 20441 3584 20453 3587
rect 20128 3556 20453 3584
rect 20128 3544 20134 3556
rect 20441 3553 20453 3556
rect 20487 3553 20499 3587
rect 20548 3584 20576 3624
rect 22066 3624 22324 3652
rect 23584 3652 23612 3692
rect 24026 3680 24032 3732
rect 24084 3680 24090 3732
rect 24118 3680 24124 3732
rect 24176 3720 24182 3732
rect 24397 3723 24455 3729
rect 24397 3720 24409 3723
rect 24176 3692 24409 3720
rect 24176 3680 24182 3692
rect 24397 3689 24409 3692
rect 24443 3689 24455 3723
rect 24397 3683 24455 3689
rect 24762 3680 24768 3732
rect 24820 3680 24826 3732
rect 25314 3680 25320 3732
rect 25372 3680 25378 3732
rect 26050 3680 26056 3732
rect 26108 3720 26114 3732
rect 26973 3723 27031 3729
rect 26973 3720 26985 3723
rect 26108 3692 26985 3720
rect 26108 3680 26114 3692
rect 26973 3689 26985 3692
rect 27019 3689 27031 3723
rect 26973 3683 27031 3689
rect 23584 3624 24624 3652
rect 22066 3584 22094 3624
rect 24596 3596 24624 3624
rect 20548 3556 22094 3584
rect 22281 3587 22339 3593
rect 20441 3547 20499 3553
rect 22281 3553 22293 3587
rect 22327 3584 22339 3587
rect 23290 3584 23296 3596
rect 22327 3556 23296 3584
rect 22327 3553 22339 3556
rect 22281 3547 22339 3553
rect 23290 3544 23296 3556
rect 23348 3544 23354 3596
rect 24578 3544 24584 3596
rect 24636 3544 24642 3596
rect 20346 3476 20352 3528
rect 20404 3476 20410 3528
rect 24670 3516 24676 3528
rect 23690 3502 24676 3516
rect 23676 3488 24676 3502
rect 18984 3420 19748 3448
rect 19812 3420 20300 3448
rect 18785 3411 18843 3417
rect 19705 3383 19763 3389
rect 19705 3380 19717 3383
rect 16500 3352 19717 3380
rect 19705 3349 19717 3352
rect 19751 3380 19763 3383
rect 19812 3380 19840 3420
rect 19751 3352 19840 3380
rect 19751 3349 19763 3352
rect 19705 3343 19763 3349
rect 20162 3340 20168 3392
rect 20220 3340 20226 3392
rect 20272 3380 20300 3420
rect 20714 3408 20720 3460
rect 20772 3408 20778 3460
rect 20990 3408 20996 3460
rect 21048 3408 21054 3460
rect 21942 3420 22094 3448
rect 21008 3380 21036 3408
rect 20272 3352 21036 3380
rect 22066 3380 22094 3420
rect 22554 3408 22560 3460
rect 22612 3408 22618 3460
rect 23676 3380 23704 3488
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 24780 3525 24808 3680
rect 24949 3587 25007 3593
rect 24949 3553 24961 3587
rect 24995 3553 25007 3587
rect 24949 3547 25007 3553
rect 25225 3587 25283 3593
rect 25225 3553 25237 3587
rect 25271 3584 25283 3587
rect 25332 3584 25360 3680
rect 25271 3556 25360 3584
rect 25501 3587 25559 3593
rect 25271 3553 25283 3556
rect 25225 3547 25283 3553
rect 25501 3553 25513 3587
rect 25547 3584 25559 3587
rect 25590 3584 25596 3596
rect 25547 3556 25596 3584
rect 25547 3553 25559 3556
rect 25501 3547 25559 3553
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 24578 3408 24584 3460
rect 24636 3448 24642 3460
rect 24964 3448 24992 3547
rect 25590 3544 25596 3556
rect 25648 3544 25654 3596
rect 26602 3476 26608 3528
rect 26660 3476 26666 3528
rect 24636 3420 24992 3448
rect 24636 3408 24642 3420
rect 22066 3352 23704 3380
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 25866 3380 25872 3392
rect 24912 3352 25872 3380
rect 24912 3340 24918 3352
rect 25866 3340 25872 3352
rect 25924 3340 25930 3392
rect 1104 3290 41400 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 41400 3290
rect 1104 3216 41400 3238
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 16574 3176 16580 3188
rect 13780 3148 16580 3176
rect 13780 3136 13786 3148
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 12989 3111 13047 3117
rect 12989 3108 13001 3111
rect 12952 3080 13001 3108
rect 12952 3068 12958 3080
rect 12989 3077 13001 3080
rect 13035 3077 13047 3111
rect 12989 3071 13047 3077
rect 14366 3068 14372 3120
rect 14424 3068 14430 3120
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2972 12771 2975
rect 13722 2972 13728 2984
rect 12759 2944 13728 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 14108 2904 14136 3026
rect 14384 2972 14412 3068
rect 14752 3049 14780 3148
rect 16574 3136 16580 3148
rect 16632 3176 16638 3188
rect 16632 3148 16712 3176
rect 16632 3136 16638 3148
rect 15013 3111 15071 3117
rect 15013 3077 15025 3111
rect 15059 3108 15071 3111
rect 15286 3108 15292 3120
rect 15059 3080 15292 3108
rect 15059 3077 15071 3080
rect 15013 3071 15071 3077
rect 15286 3068 15292 3080
rect 15344 3068 15350 3120
rect 15470 3068 15476 3120
rect 15528 3068 15534 3120
rect 16684 3049 16712 3148
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 16816 3148 16988 3176
rect 16816 3136 16822 3148
rect 16960 3117 16988 3148
rect 20070 3136 20076 3188
rect 20128 3136 20134 3188
rect 21266 3136 21272 3188
rect 21324 3136 21330 3188
rect 21818 3136 21824 3188
rect 21876 3176 21882 3188
rect 22189 3179 22247 3185
rect 21876 3148 22094 3176
rect 21876 3136 21882 3148
rect 16945 3111 17003 3117
rect 16945 3077 16957 3111
rect 16991 3077 17003 3111
rect 16945 3071 17003 3077
rect 17954 3068 17960 3120
rect 18012 3068 18018 3120
rect 20088 3108 20116 3136
rect 21174 3108 21180 3120
rect 19536 3080 20116 3108
rect 21022 3080 21180 3108
rect 19536 3049 19564 3080
rect 21174 3068 21180 3080
rect 21232 3068 21238 3120
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3009 19579 3043
rect 22066 3040 22094 3148
rect 22189 3145 22201 3179
rect 22235 3176 22247 3179
rect 22554 3176 22560 3188
rect 22235 3148 22560 3176
rect 22235 3145 22247 3148
rect 22189 3139 22247 3145
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 25222 3136 25228 3188
rect 25280 3136 25286 3188
rect 25682 3136 25688 3188
rect 25740 3136 25746 3188
rect 25958 3136 25964 3188
rect 26016 3136 26022 3188
rect 26050 3136 26056 3188
rect 26108 3136 26114 3188
rect 23753 3111 23811 3117
rect 23753 3077 23765 3111
rect 23799 3108 23811 3111
rect 23842 3108 23848 3120
rect 23799 3080 23848 3108
rect 23799 3077 23811 3080
rect 23753 3071 23811 3077
rect 23842 3068 23848 3080
rect 23900 3068 23906 3120
rect 24762 3068 24768 3120
rect 24820 3068 24826 3120
rect 25976 3108 26004 3136
rect 26145 3111 26203 3117
rect 26145 3108 26157 3111
rect 25976 3080 26157 3108
rect 26145 3077 26157 3080
rect 26191 3077 26203 3111
rect 26145 3071 26203 3077
rect 22373 3043 22431 3049
rect 22373 3040 22385 3043
rect 22066 3012 22385 3040
rect 19521 3003 19579 3009
rect 22373 3009 22385 3012
rect 22419 3009 22431 3043
rect 22373 3003 22431 3009
rect 23290 3000 23296 3052
rect 23348 3040 23354 3052
rect 23477 3043 23535 3049
rect 23477 3040 23489 3043
rect 23348 3012 23489 3040
rect 23348 3000 23354 3012
rect 23477 3009 23489 3012
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 19797 2975 19855 2981
rect 14384 2944 19656 2972
rect 14550 2904 14556 2916
rect 14108 2876 14556 2904
rect 14550 2864 14556 2876
rect 14608 2864 14614 2916
rect 16482 2864 16488 2916
rect 16540 2864 16546 2916
rect 14461 2839 14519 2845
rect 14461 2805 14473 2839
rect 14507 2836 14519 2839
rect 14826 2836 14832 2848
rect 14507 2808 14832 2836
rect 14507 2805 14519 2808
rect 14461 2799 14519 2805
rect 14826 2796 14832 2808
rect 14884 2796 14890 2848
rect 17678 2796 17684 2848
rect 17736 2836 17742 2848
rect 18417 2839 18475 2845
rect 18417 2836 18429 2839
rect 17736 2808 18429 2836
rect 17736 2796 17742 2808
rect 18417 2805 18429 2808
rect 18463 2805 18475 2839
rect 19628 2836 19656 2944
rect 19797 2941 19809 2975
rect 19843 2972 19855 2975
rect 20162 2972 20168 2984
rect 19843 2944 20168 2972
rect 19843 2941 19855 2944
rect 19797 2935 19855 2941
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 23492 2972 23520 3003
rect 25314 3000 25320 3052
rect 25372 3000 25378 3052
rect 25332 2972 25360 3000
rect 23492 2944 25360 2972
rect 26329 2975 26387 2981
rect 26329 2941 26341 2975
rect 26375 2972 26387 2975
rect 27522 2972 27528 2984
rect 26375 2944 27528 2972
rect 26375 2941 26387 2944
rect 26329 2935 26387 2941
rect 27522 2932 27528 2944
rect 27580 2932 27586 2984
rect 24854 2836 24860 2848
rect 19628 2808 24860 2836
rect 18417 2799 18475 2805
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 1104 2746 41400 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 41400 2746
rect 1104 2672 41400 2694
rect 14274 2632 14280 2644
rect 6886 2604 14280 2632
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 6886 2428 6914 2604
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 20165 2635 20223 2641
rect 20165 2601 20177 2635
rect 20211 2632 20223 2635
rect 20714 2632 20720 2644
rect 20211 2604 20720 2632
rect 20211 2601 20223 2604
rect 20165 2595 20223 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 12032 2468 23428 2496
rect 12032 2456 12038 2468
rect 1719 2400 6914 2428
rect 7929 2431 7987 2437
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8846 2428 8852 2440
rect 7975 2400 8852 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 11790 2388 11796 2440
rect 11848 2388 11854 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 17678 2428 17684 2440
rect 15703 2400 17684 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 19518 2388 19524 2440
rect 19576 2388 19582 2440
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2428 20407 2431
rect 20806 2428 20812 2440
rect 20395 2400 20812 2428
rect 20395 2397 20407 2400
rect 20349 2391 20407 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 23400 2437 23428 2468
rect 23385 2431 23443 2437
rect 23385 2397 23397 2431
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 31110 2388 31116 2440
rect 31168 2388 31174 2440
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 34977 2431 35035 2437
rect 34977 2428 34989 2431
rect 34664 2400 34989 2428
rect 34664 2388 34670 2400
rect 34977 2397 34989 2400
rect 35023 2397 35035 2431
rect 34977 2391 35035 2397
rect 38841 2431 38899 2437
rect 38841 2397 38853 2431
rect 38887 2428 38899 2431
rect 39022 2428 39028 2440
rect 38887 2400 39028 2428
rect 38887 2397 38899 2400
rect 38841 2391 38899 2397
rect 39022 2388 39028 2400
rect 39080 2388 39086 2440
rect 40678 2388 40684 2440
rect 40736 2388 40742 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 72 2332 1501 2360
rect 72 2320 78 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 4065 2363 4123 2369
rect 4065 2329 4077 2363
rect 4111 2360 4123 2363
rect 4982 2360 4988 2372
rect 4111 2332 4988 2360
rect 4111 2329 4123 2332
rect 4065 2323 4123 2329
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 27249 2363 27307 2369
rect 27249 2360 27261 2363
rect 20680 2332 27261 2360
rect 20680 2320 20686 2332
rect 27249 2329 27261 2332
rect 27295 2329 27307 2363
rect 27249 2323 27307 2329
rect 3970 2252 3976 2304
rect 4028 2292 4034 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 4028 2264 4169 2292
rect 4028 2252 4034 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15528 2264 15761 2292
rect 15528 2252 15534 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23348 2264 23489 2292
rect 23348 2252 23354 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 27062 2252 27068 2304
rect 27120 2292 27126 2304
rect 27341 2295 27399 2301
rect 27341 2292 27353 2295
rect 27120 2264 27353 2292
rect 27120 2252 27126 2264
rect 27341 2261 27353 2264
rect 27387 2261 27399 2295
rect 27341 2255 27399 2261
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30984 2264 31217 2292
rect 30984 2252 30990 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34848 2264 35081 2292
rect 34848 2252 34854 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 38654 2252 38660 2304
rect 38712 2292 38718 2304
rect 38933 2295 38991 2301
rect 38933 2292 38945 2295
rect 38712 2264 38945 2292
rect 38712 2252 38718 2264
rect 38933 2261 38945 2264
rect 38979 2261 38991 2295
rect 38933 2255 38991 2261
rect 39942 2252 39948 2304
rect 40000 2292 40006 2304
rect 40773 2295 40831 2301
rect 40773 2292 40785 2295
rect 40000 2264 40785 2292
rect 40000 2252 40006 2264
rect 40773 2261 40785 2264
rect 40819 2261 40831 2295
rect 40773 2255 40831 2261
rect 1104 2202 41400 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 41400 2202
rect 1104 2128 41400 2150
<< via1 >>
rect 10876 42508 10928 42560
rect 14556 42508 14608 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 11060 42304 11112 42356
rect 2780 42236 2832 42288
rect 7104 42236 7156 42288
rect 1492 42211 1544 42220
rect 1492 42177 1501 42211
rect 1501 42177 1535 42211
rect 1535 42177 1544 42211
rect 1492 42168 1544 42177
rect 3240 42168 3292 42220
rect 18696 42304 18748 42356
rect 29092 42304 29144 42356
rect 30380 42304 30432 42356
rect 32956 42304 33008 42356
rect 38292 42347 38344 42356
rect 38292 42313 38301 42347
rect 38301 42313 38335 42347
rect 38335 42313 38344 42347
rect 38292 42304 38344 42313
rect 41880 42304 41932 42356
rect 14648 42211 14700 42220
rect 14648 42177 14657 42211
rect 14657 42177 14691 42211
rect 14691 42177 14700 42211
rect 14648 42168 14700 42177
rect 14832 42168 14884 42220
rect 10876 42032 10928 42084
rect 16028 42168 16080 42220
rect 34520 42236 34572 42288
rect 22560 42168 22612 42220
rect 30472 42211 30524 42220
rect 30472 42177 30481 42211
rect 30481 42177 30515 42211
rect 30515 42177 30524 42211
rect 30472 42168 30524 42177
rect 38200 42211 38252 42220
rect 38200 42177 38209 42211
rect 38209 42177 38243 42211
rect 38243 42177 38252 42211
rect 38200 42168 38252 42177
rect 14004 41964 14056 42016
rect 31668 42100 31720 42152
rect 32680 42143 32732 42152
rect 32680 42109 32689 42143
rect 32689 42109 32723 42143
rect 32723 42109 32732 42143
rect 32680 42100 32732 42109
rect 16028 42032 16080 42084
rect 23480 42032 23532 42084
rect 24400 42032 24452 42084
rect 20720 41964 20772 42016
rect 33324 42007 33376 42016
rect 33324 41973 33333 42007
rect 33333 41973 33367 42007
rect 33367 41973 33376 42007
rect 33324 41964 33376 41973
rect 40868 42007 40920 42016
rect 40868 41973 40877 42007
rect 40877 41973 40911 42007
rect 40911 41973 40920 42007
rect 40868 41964 40920 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 7196 41488 7248 41540
rect 14556 41760 14608 41812
rect 14004 41692 14056 41744
rect 11060 41667 11112 41676
rect 11060 41633 11069 41667
rect 11069 41633 11103 41667
rect 11103 41633 11112 41667
rect 11060 41624 11112 41633
rect 12716 41624 12768 41676
rect 15016 41624 15068 41676
rect 11428 41599 11480 41608
rect 11428 41565 11437 41599
rect 11437 41565 11471 41599
rect 11471 41565 11480 41599
rect 11428 41556 11480 41565
rect 13452 41556 13504 41608
rect 13544 41599 13596 41608
rect 13544 41565 13553 41599
rect 13553 41565 13587 41599
rect 13587 41565 13596 41599
rect 13544 41556 13596 41565
rect 14004 41556 14056 41608
rect 17776 41760 17828 41812
rect 29000 41760 29052 41812
rect 29092 41760 29144 41812
rect 32680 41760 32732 41812
rect 19432 41692 19484 41744
rect 18696 41624 18748 41676
rect 19064 41624 19116 41676
rect 19892 41667 19944 41676
rect 19892 41633 19901 41667
rect 19901 41633 19935 41667
rect 19935 41633 19944 41667
rect 19892 41624 19944 41633
rect 20260 41692 20312 41744
rect 24492 41692 24544 41744
rect 20168 41624 20220 41676
rect 12440 41488 12492 41540
rect 10600 41463 10652 41472
rect 10600 41429 10609 41463
rect 10609 41429 10643 41463
rect 10643 41429 10652 41463
rect 10600 41420 10652 41429
rect 13268 41420 13320 41472
rect 13452 41420 13504 41472
rect 15108 41420 15160 41472
rect 23296 41624 23348 41676
rect 24308 41624 24360 41676
rect 17500 41488 17552 41540
rect 17960 41420 18012 41472
rect 18972 41488 19024 41540
rect 20076 41599 20128 41608
rect 20076 41565 20085 41599
rect 20085 41565 20119 41599
rect 20119 41565 20128 41599
rect 20076 41556 20128 41565
rect 20168 41488 20220 41540
rect 20536 41556 20588 41608
rect 22652 41556 22704 41608
rect 21456 41488 21508 41540
rect 22100 41488 22152 41540
rect 20812 41420 20864 41472
rect 22468 41488 22520 41540
rect 23480 41556 23532 41608
rect 24124 41556 24176 41608
rect 28540 41667 28592 41676
rect 28540 41633 28549 41667
rect 28549 41633 28583 41667
rect 28583 41633 28592 41667
rect 28540 41624 28592 41633
rect 32588 41667 32640 41676
rect 32588 41633 32597 41667
rect 32597 41633 32631 41667
rect 32631 41633 32640 41667
rect 32588 41624 32640 41633
rect 33324 41624 33376 41676
rect 29276 41556 29328 41608
rect 24032 41488 24084 41540
rect 25596 41488 25648 41540
rect 25872 41488 25924 41540
rect 26240 41488 26292 41540
rect 26608 41488 26660 41540
rect 22836 41420 22888 41472
rect 23204 41420 23256 41472
rect 24400 41420 24452 41472
rect 27252 41420 27304 41472
rect 27436 41488 27488 41540
rect 32404 41488 32456 41540
rect 34428 41488 34480 41540
rect 27712 41420 27764 41472
rect 31576 41420 31628 41472
rect 33876 41420 33928 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 11060 41216 11112 41268
rect 11428 41216 11480 41268
rect 13820 41216 13872 41268
rect 15016 41216 15068 41268
rect 15660 41216 15712 41268
rect 10600 41080 10652 41132
rect 10876 41080 10928 41132
rect 9496 41055 9548 41064
rect 9496 41021 9505 41055
rect 9505 41021 9539 41055
rect 9539 41021 9548 41055
rect 9496 41012 9548 41021
rect 11704 41012 11756 41064
rect 13452 41080 13504 41132
rect 12808 41055 12860 41064
rect 12808 41021 12817 41055
rect 12817 41021 12851 41055
rect 12851 41021 12860 41055
rect 12808 41012 12860 41021
rect 12992 41055 13044 41064
rect 12992 41021 13001 41055
rect 13001 41021 13035 41055
rect 13035 41021 13044 41055
rect 12992 41012 13044 41021
rect 14740 41055 14792 41064
rect 14740 41021 14749 41055
rect 14749 41021 14783 41055
rect 14783 41021 14792 41055
rect 14740 41012 14792 41021
rect 15384 41080 15436 41132
rect 15660 41123 15712 41132
rect 15660 41089 15669 41123
rect 15669 41089 15703 41123
rect 15703 41089 15712 41123
rect 15660 41080 15712 41089
rect 15752 41080 15804 41132
rect 10232 40876 10284 40928
rect 11704 40876 11756 40928
rect 15200 40919 15252 40928
rect 15200 40885 15209 40919
rect 15209 40885 15243 40919
rect 15243 40885 15252 40919
rect 15200 40876 15252 40885
rect 16212 40987 16264 40996
rect 16212 40953 16221 40987
rect 16221 40953 16255 40987
rect 16255 40953 16264 40987
rect 16212 40944 16264 40953
rect 17316 41148 17368 41200
rect 18052 41191 18104 41200
rect 18052 41157 18061 41191
rect 18061 41157 18095 41191
rect 18095 41157 18104 41191
rect 18052 41148 18104 41157
rect 16764 41123 16816 41132
rect 16764 41089 16773 41123
rect 16773 41089 16807 41123
rect 16807 41089 16816 41123
rect 16764 41080 16816 41089
rect 17132 41123 17184 41132
rect 17132 41089 17141 41123
rect 17141 41089 17175 41123
rect 17175 41089 17184 41123
rect 17132 41080 17184 41089
rect 17316 41012 17368 41064
rect 17592 41080 17644 41132
rect 17868 41123 17920 41132
rect 17868 41089 17877 41123
rect 17877 41089 17911 41123
rect 17911 41089 17920 41123
rect 17868 41080 17920 41089
rect 17960 41123 18012 41132
rect 17960 41089 17969 41123
rect 17969 41089 18003 41123
rect 18003 41089 18012 41123
rect 17960 41080 18012 41089
rect 18328 41148 18380 41200
rect 18512 41080 18564 41132
rect 18604 41123 18656 41132
rect 18604 41089 18613 41123
rect 18613 41089 18647 41123
rect 18647 41089 18656 41123
rect 18604 41080 18656 41089
rect 19156 41080 19208 41132
rect 19800 41123 19852 41132
rect 19800 41089 19809 41123
rect 19809 41089 19843 41123
rect 19843 41089 19852 41123
rect 19800 41080 19852 41089
rect 20352 41148 20404 41200
rect 21732 41216 21784 41268
rect 22008 41216 22060 41268
rect 22652 41216 22704 41268
rect 25320 41216 25372 41268
rect 26332 41216 26384 41268
rect 26608 41216 26660 41268
rect 26792 41216 26844 41268
rect 27252 41216 27304 41268
rect 20076 41123 20128 41132
rect 20076 41089 20085 41123
rect 20085 41089 20119 41123
rect 20119 41089 20128 41123
rect 20076 41080 20128 41089
rect 20168 41080 20220 41132
rect 20444 41123 20496 41132
rect 20444 41089 20453 41123
rect 20453 41089 20487 41123
rect 20487 41089 20496 41123
rect 20444 41080 20496 41089
rect 20812 41080 20864 41132
rect 21088 41080 21140 41132
rect 17500 41055 17552 41064
rect 17500 41021 17509 41055
rect 17509 41021 17543 41055
rect 17543 41021 17552 41055
rect 17500 41012 17552 41021
rect 18052 41012 18104 41064
rect 18420 41055 18472 41064
rect 18420 41021 18429 41055
rect 18429 41021 18463 41055
rect 18463 41021 18472 41055
rect 18420 41012 18472 41021
rect 19248 41055 19300 41064
rect 19248 41021 19257 41055
rect 19257 41021 19291 41055
rect 19291 41021 19300 41055
rect 19248 41012 19300 41021
rect 19340 41012 19392 41064
rect 21456 41055 21508 41064
rect 21456 41021 21465 41055
rect 21465 41021 21499 41055
rect 21499 41021 21508 41055
rect 21456 41012 21508 41021
rect 15752 40876 15804 40928
rect 16672 40876 16724 40928
rect 18144 40944 18196 40996
rect 19708 40944 19760 40996
rect 19892 40944 19944 40996
rect 23388 41080 23440 41132
rect 25688 41148 25740 41200
rect 25044 41123 25096 41132
rect 25044 41089 25053 41123
rect 25053 41089 25087 41123
rect 25087 41089 25096 41123
rect 25044 41080 25096 41089
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 25412 41123 25464 41132
rect 25412 41089 25421 41123
rect 25421 41089 25455 41123
rect 25455 41089 25464 41123
rect 25412 41080 25464 41089
rect 22376 41012 22428 41064
rect 22652 41012 22704 41064
rect 23940 41055 23992 41064
rect 23940 41021 23949 41055
rect 23949 41021 23983 41055
rect 23983 41021 23992 41055
rect 23940 41012 23992 41021
rect 24124 41012 24176 41064
rect 24400 41055 24452 41064
rect 24400 41021 24434 41055
rect 24434 41021 24452 41055
rect 24400 41012 24452 41021
rect 23020 40944 23072 40996
rect 26240 41148 26292 41200
rect 29460 41216 29512 41268
rect 26608 41123 26660 41132
rect 26608 41089 26617 41123
rect 26617 41089 26651 41123
rect 26651 41089 26660 41123
rect 26608 41080 26660 41089
rect 26884 41080 26936 41132
rect 27160 41123 27212 41132
rect 27160 41089 27169 41123
rect 27169 41089 27203 41123
rect 27203 41089 27212 41123
rect 27160 41080 27212 41089
rect 27252 41123 27304 41132
rect 27252 41089 27261 41123
rect 27261 41089 27295 41123
rect 27295 41089 27304 41123
rect 27252 41080 27304 41089
rect 26516 41055 26568 41064
rect 26516 41021 26525 41055
rect 26525 41021 26559 41055
rect 26559 41021 26568 41055
rect 26516 41012 26568 41021
rect 26792 41012 26844 41064
rect 28080 41123 28132 41132
rect 28080 41089 28090 41123
rect 28090 41089 28124 41123
rect 28124 41089 28132 41123
rect 28080 41080 28132 41089
rect 28172 41080 28224 41132
rect 28356 41123 28408 41132
rect 28356 41089 28365 41123
rect 28365 41089 28399 41123
rect 28399 41089 28408 41123
rect 28356 41080 28408 41089
rect 28448 41123 28500 41132
rect 28448 41089 28462 41123
rect 28462 41089 28496 41123
rect 28496 41089 28500 41123
rect 28448 41080 28500 41089
rect 28724 41123 28776 41132
rect 28724 41089 28733 41123
rect 28733 41089 28767 41123
rect 28767 41089 28776 41123
rect 28724 41080 28776 41089
rect 29276 41148 29328 41200
rect 28540 41012 28592 41064
rect 18696 40876 18748 40928
rect 21088 40876 21140 40928
rect 22100 40876 22152 40928
rect 22744 40876 22796 40928
rect 24768 40876 24820 40928
rect 26240 40876 26292 40928
rect 26792 40919 26844 40928
rect 26792 40885 26801 40919
rect 26801 40885 26835 40919
rect 26835 40885 26844 40919
rect 26792 40876 26844 40885
rect 26884 40876 26936 40928
rect 27160 40876 27212 40928
rect 29736 41080 29788 41132
rect 30564 41080 30616 41132
rect 30656 41055 30708 41064
rect 30656 41021 30665 41055
rect 30665 41021 30699 41055
rect 30699 41021 30708 41055
rect 30656 41012 30708 41021
rect 31668 41080 31720 41132
rect 34612 41080 34664 41132
rect 40868 41148 40920 41200
rect 41236 41080 41288 41132
rect 30840 41012 30892 41064
rect 28540 40876 28592 40928
rect 29276 40919 29328 40928
rect 29276 40885 29285 40919
rect 29285 40885 29319 40919
rect 29319 40885 29328 40919
rect 29276 40876 29328 40885
rect 30012 40944 30064 40996
rect 32404 41055 32456 41064
rect 32404 41021 32413 41055
rect 32413 41021 32447 41055
rect 32447 41021 32456 41055
rect 32404 41012 32456 41021
rect 34428 41012 34480 41064
rect 40776 41055 40828 41064
rect 40776 41021 40785 41055
rect 40785 41021 40819 41055
rect 40819 41021 40828 41055
rect 40776 41012 40828 41021
rect 30380 40876 30432 40928
rect 30472 40919 30524 40928
rect 30472 40885 30481 40919
rect 30481 40885 30515 40919
rect 30515 40885 30524 40919
rect 30472 40876 30524 40885
rect 40408 40919 40460 40928
rect 40408 40885 40417 40919
rect 40417 40885 40451 40919
rect 40451 40885 40460 40919
rect 40408 40876 40460 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 9496 40672 9548 40724
rect 14740 40672 14792 40724
rect 17316 40715 17368 40724
rect 17316 40681 17325 40715
rect 17325 40681 17359 40715
rect 17359 40681 17368 40715
rect 17316 40672 17368 40681
rect 18052 40715 18104 40724
rect 18052 40681 18061 40715
rect 18061 40681 18095 40715
rect 18095 40681 18104 40715
rect 18052 40672 18104 40681
rect 19064 40672 19116 40724
rect 20168 40672 20220 40724
rect 20536 40715 20588 40724
rect 20536 40681 20545 40715
rect 20545 40681 20579 40715
rect 20579 40681 20588 40715
rect 20536 40672 20588 40681
rect 21916 40672 21968 40724
rect 15200 40604 15252 40656
rect 11060 40579 11112 40588
rect 11060 40545 11069 40579
rect 11069 40545 11103 40579
rect 11103 40545 11112 40579
rect 11060 40536 11112 40545
rect 12624 40536 12676 40588
rect 940 40468 992 40520
rect 1676 40511 1728 40520
rect 1676 40477 1685 40511
rect 1685 40477 1719 40511
rect 1719 40477 1728 40511
rect 1676 40468 1728 40477
rect 10232 40468 10284 40520
rect 10416 40511 10468 40520
rect 10416 40477 10425 40511
rect 10425 40477 10459 40511
rect 10459 40477 10468 40511
rect 10416 40468 10468 40477
rect 12440 40468 12492 40520
rect 13452 40536 13504 40588
rect 14556 40511 14608 40520
rect 14556 40477 14565 40511
rect 14565 40477 14599 40511
rect 14599 40477 14608 40511
rect 14556 40468 14608 40477
rect 15108 40468 15160 40520
rect 10968 40400 11020 40452
rect 15476 40536 15528 40588
rect 15660 40604 15712 40656
rect 16580 40604 16632 40656
rect 16764 40604 16816 40656
rect 18328 40604 18380 40656
rect 18512 40604 18564 40656
rect 19616 40604 19668 40656
rect 16948 40536 17000 40588
rect 17132 40536 17184 40588
rect 13728 40375 13780 40384
rect 13728 40341 13737 40375
rect 13737 40341 13771 40375
rect 13771 40341 13780 40375
rect 13728 40332 13780 40341
rect 14188 40375 14240 40384
rect 14188 40341 14197 40375
rect 14197 40341 14231 40375
rect 14231 40341 14240 40375
rect 14188 40332 14240 40341
rect 14464 40332 14516 40384
rect 15936 40511 15988 40520
rect 15936 40477 15945 40511
rect 15945 40477 15979 40511
rect 15979 40477 15988 40511
rect 15936 40468 15988 40477
rect 16028 40511 16080 40520
rect 16028 40477 16037 40511
rect 16037 40477 16071 40511
rect 16071 40477 16080 40511
rect 16028 40468 16080 40477
rect 16580 40511 16632 40520
rect 16580 40477 16589 40511
rect 16589 40477 16623 40511
rect 16623 40477 16632 40511
rect 16580 40468 16632 40477
rect 17868 40536 17920 40588
rect 15568 40400 15620 40452
rect 16488 40400 16540 40452
rect 17132 40400 17184 40452
rect 17776 40468 17828 40520
rect 18144 40468 18196 40520
rect 18696 40511 18748 40520
rect 18696 40477 18705 40511
rect 18705 40477 18739 40511
rect 18739 40477 18748 40511
rect 18696 40468 18748 40477
rect 19248 40468 19300 40520
rect 19708 40468 19760 40520
rect 20444 40604 20496 40656
rect 21456 40604 21508 40656
rect 22192 40715 22244 40724
rect 22192 40681 22201 40715
rect 22201 40681 22235 40715
rect 22235 40681 22244 40715
rect 22192 40672 22244 40681
rect 23388 40672 23440 40724
rect 24124 40715 24176 40724
rect 22376 40604 22428 40656
rect 21916 40536 21968 40588
rect 22008 40536 22060 40588
rect 20076 40468 20128 40520
rect 20812 40468 20864 40520
rect 20260 40400 20312 40452
rect 15476 40332 15528 40384
rect 15844 40332 15896 40384
rect 17316 40332 17368 40384
rect 17408 40332 17460 40384
rect 17776 40375 17828 40384
rect 17776 40341 17785 40375
rect 17785 40341 17819 40375
rect 17819 40341 17828 40375
rect 17776 40332 17828 40341
rect 18328 40332 18380 40384
rect 19616 40332 19668 40384
rect 21456 40400 21508 40452
rect 24124 40681 24133 40715
rect 24133 40681 24167 40715
rect 24167 40681 24176 40715
rect 24124 40672 24176 40681
rect 23756 40647 23808 40656
rect 23756 40613 23765 40647
rect 23765 40613 23799 40647
rect 23799 40613 23808 40647
rect 23756 40604 23808 40613
rect 24032 40604 24084 40656
rect 23480 40536 23532 40588
rect 22468 40511 22520 40520
rect 22468 40477 22477 40511
rect 22477 40477 22511 40511
rect 22511 40477 22520 40511
rect 22468 40468 22520 40477
rect 23112 40468 23164 40520
rect 23204 40468 23256 40520
rect 24584 40579 24636 40588
rect 24584 40545 24593 40579
rect 24593 40545 24627 40579
rect 24627 40545 24636 40579
rect 24584 40536 24636 40545
rect 25320 40672 25372 40724
rect 26976 40672 27028 40724
rect 30012 40672 30064 40724
rect 30288 40715 30340 40724
rect 30288 40681 30297 40715
rect 30297 40681 30331 40715
rect 30331 40681 30340 40715
rect 30288 40672 30340 40681
rect 30472 40672 30524 40724
rect 24216 40511 24268 40520
rect 24216 40477 24225 40511
rect 24225 40477 24259 40511
rect 24259 40477 24268 40511
rect 24216 40468 24268 40477
rect 24676 40511 24728 40520
rect 24676 40477 24685 40511
rect 24685 40477 24719 40511
rect 24719 40477 24728 40511
rect 24676 40468 24728 40477
rect 25688 40536 25740 40588
rect 22376 40400 22428 40452
rect 20720 40332 20772 40384
rect 21088 40332 21140 40384
rect 21916 40375 21968 40384
rect 21916 40341 21925 40375
rect 21925 40341 21959 40375
rect 21959 40341 21968 40375
rect 21916 40332 21968 40341
rect 22284 40375 22336 40384
rect 22284 40341 22293 40375
rect 22293 40341 22327 40375
rect 22327 40341 22336 40375
rect 22284 40332 22336 40341
rect 22652 40443 22704 40452
rect 22652 40409 22661 40443
rect 22661 40409 22695 40443
rect 22695 40409 22704 40443
rect 22652 40400 22704 40409
rect 22928 40400 22980 40452
rect 23296 40400 23348 40452
rect 24860 40400 24912 40452
rect 25412 40468 25464 40520
rect 25780 40511 25832 40520
rect 25780 40477 25809 40511
rect 25809 40477 25832 40511
rect 25780 40468 25832 40477
rect 26056 40511 26108 40520
rect 26056 40477 26065 40511
rect 26065 40477 26099 40511
rect 26099 40477 26108 40511
rect 26056 40468 26108 40477
rect 25412 40332 25464 40384
rect 26516 40468 26568 40520
rect 26976 40511 27028 40520
rect 26976 40477 26983 40511
rect 26983 40477 27028 40511
rect 26976 40468 27028 40477
rect 27712 40604 27764 40656
rect 26700 40400 26752 40452
rect 27160 40443 27212 40452
rect 27160 40409 27169 40443
rect 27169 40409 27203 40443
rect 27203 40409 27212 40443
rect 27160 40400 27212 40409
rect 28540 40468 28592 40520
rect 29368 40468 29420 40520
rect 32588 40536 32640 40588
rect 33600 40536 33652 40588
rect 40408 40672 40460 40724
rect 27712 40400 27764 40452
rect 28080 40400 28132 40452
rect 28724 40443 28776 40452
rect 28724 40409 28733 40443
rect 28733 40409 28767 40443
rect 28767 40409 28776 40443
rect 28724 40400 28776 40409
rect 29736 40443 29788 40452
rect 29736 40409 29745 40443
rect 29745 40409 29779 40443
rect 29779 40409 29788 40443
rect 29736 40400 29788 40409
rect 29828 40443 29880 40452
rect 29828 40409 29837 40443
rect 29837 40409 29871 40443
rect 29871 40409 29880 40443
rect 29828 40400 29880 40409
rect 37648 40511 37700 40520
rect 37648 40477 37657 40511
rect 37657 40477 37691 40511
rect 37691 40477 37700 40511
rect 37648 40468 37700 40477
rect 26976 40332 27028 40384
rect 27528 40332 27580 40384
rect 29184 40332 29236 40384
rect 32220 40443 32272 40452
rect 32220 40409 32229 40443
rect 32229 40409 32263 40443
rect 32263 40409 32272 40443
rect 32220 40400 32272 40409
rect 30472 40332 30524 40384
rect 31208 40332 31260 40384
rect 31484 40332 31536 40384
rect 32772 40400 32824 40452
rect 33048 40443 33100 40452
rect 33048 40409 33057 40443
rect 33057 40409 33091 40443
rect 33091 40409 33100 40443
rect 33048 40400 33100 40409
rect 34428 40400 34480 40452
rect 38660 40400 38712 40452
rect 32588 40375 32640 40384
rect 32588 40341 32597 40375
rect 32597 40341 32631 40375
rect 32631 40341 32640 40375
rect 32588 40332 32640 40341
rect 34520 40375 34572 40384
rect 34520 40341 34529 40375
rect 34529 40341 34563 40375
rect 34563 40341 34572 40375
rect 34520 40332 34572 40341
rect 39304 40332 39356 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 12624 40128 12676 40180
rect 13728 40128 13780 40180
rect 14464 40128 14516 40180
rect 10876 40060 10928 40112
rect 10968 40060 11020 40112
rect 11060 40060 11112 40112
rect 12440 40060 12492 40112
rect 8484 40035 8536 40044
rect 8484 40001 8493 40035
rect 8493 40001 8527 40035
rect 8527 40001 8536 40035
rect 8484 39992 8536 40001
rect 9588 40035 9640 40044
rect 9588 40001 9597 40035
rect 9597 40001 9631 40035
rect 9631 40001 9640 40035
rect 9588 39992 9640 40001
rect 8300 39831 8352 39840
rect 8300 39797 8309 39831
rect 8309 39797 8343 39831
rect 8343 39797 8352 39831
rect 8300 39788 8352 39797
rect 9220 39831 9272 39840
rect 9220 39797 9229 39831
rect 9229 39797 9263 39831
rect 9263 39797 9272 39831
rect 9220 39788 9272 39797
rect 9312 39788 9364 39840
rect 10968 39924 11020 39976
rect 9864 39856 9916 39908
rect 14372 40035 14424 40044
rect 14372 40001 14381 40035
rect 14381 40001 14415 40035
rect 14415 40001 14424 40035
rect 14372 39992 14424 40001
rect 15108 40128 15160 40180
rect 15936 40128 15988 40180
rect 16120 40128 16172 40180
rect 16580 40060 16632 40112
rect 16948 40060 17000 40112
rect 17132 40128 17184 40180
rect 17316 40128 17368 40180
rect 17960 40128 18012 40180
rect 15108 40035 15160 40044
rect 15108 40001 15117 40035
rect 15117 40001 15151 40035
rect 15151 40001 15160 40035
rect 15108 39992 15160 40001
rect 15936 39992 15988 40044
rect 15568 39924 15620 39976
rect 15200 39856 15252 39908
rect 15844 39967 15896 39976
rect 15844 39933 15853 39967
rect 15853 39933 15887 39967
rect 15887 39933 15896 39967
rect 18144 40060 18196 40112
rect 19248 40128 19300 40180
rect 20076 40128 20128 40180
rect 20260 40128 20312 40180
rect 20444 40128 20496 40180
rect 22652 40128 22704 40180
rect 17592 39992 17644 40044
rect 18604 39992 18656 40044
rect 20352 40060 20404 40112
rect 20904 40060 20956 40112
rect 20812 39992 20864 40044
rect 23664 40035 23716 40044
rect 23664 40001 23673 40035
rect 23673 40001 23707 40035
rect 23707 40001 23716 40035
rect 23664 39992 23716 40001
rect 24032 40103 24084 40112
rect 24032 40069 24041 40103
rect 24041 40069 24075 40103
rect 24075 40069 24084 40103
rect 24032 40060 24084 40069
rect 27344 40171 27396 40180
rect 27344 40137 27353 40171
rect 27353 40137 27387 40171
rect 27387 40137 27396 40171
rect 27344 40128 27396 40137
rect 24124 40035 24176 40044
rect 24124 40001 24138 40035
rect 24138 40001 24172 40035
rect 24172 40001 24176 40035
rect 24124 39992 24176 40001
rect 24584 39992 24636 40044
rect 15844 39924 15896 39933
rect 25504 39924 25556 39976
rect 26056 40035 26108 40044
rect 26056 40001 26065 40035
rect 26065 40001 26099 40035
rect 26099 40001 26108 40035
rect 26056 39992 26108 40001
rect 26332 39992 26384 40044
rect 26884 39992 26936 40044
rect 28448 40060 28500 40112
rect 29092 40103 29144 40112
rect 29092 40069 29101 40103
rect 29101 40069 29135 40103
rect 29135 40069 29144 40103
rect 29092 40060 29144 40069
rect 29184 39992 29236 40044
rect 32220 40128 32272 40180
rect 32588 40128 32640 40180
rect 33048 40128 33100 40180
rect 30748 40060 30800 40112
rect 30196 39992 30248 40044
rect 27068 39967 27120 39976
rect 27068 39933 27077 39967
rect 27077 39933 27111 39967
rect 27111 39933 27120 39967
rect 27068 39924 27120 39933
rect 27896 39924 27948 39976
rect 28632 39924 28684 39976
rect 31208 39967 31260 39976
rect 31208 39933 31217 39967
rect 31217 39933 31251 39967
rect 31251 39933 31260 39967
rect 31208 39924 31260 39933
rect 31668 39924 31720 39976
rect 16028 39856 16080 39908
rect 16212 39856 16264 39908
rect 17500 39856 17552 39908
rect 19800 39856 19852 39908
rect 20168 39856 20220 39908
rect 22100 39899 22152 39908
rect 22100 39865 22109 39899
rect 22109 39865 22143 39899
rect 22143 39865 22152 39899
rect 22100 39856 22152 39865
rect 23388 39856 23440 39908
rect 12992 39788 13044 39840
rect 13636 39788 13688 39840
rect 15384 39788 15436 39840
rect 17592 39788 17644 39840
rect 19892 39788 19944 39840
rect 20536 39788 20588 39840
rect 20812 39788 20864 39840
rect 22744 39788 22796 39840
rect 25780 39788 25832 39840
rect 25964 39788 26016 39840
rect 26516 39788 26568 39840
rect 26792 39788 26844 39840
rect 27896 39788 27948 39840
rect 29276 39831 29328 39840
rect 29276 39797 29285 39831
rect 29285 39797 29319 39831
rect 29319 39797 29328 39831
rect 29276 39788 29328 39797
rect 29644 39788 29696 39840
rect 30380 39788 30432 39840
rect 32036 39788 32088 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 8484 39584 8536 39636
rect 9772 39584 9824 39636
rect 14372 39584 14424 39636
rect 15292 39584 15344 39636
rect 15660 39584 15712 39636
rect 16488 39584 16540 39636
rect 16580 39584 16632 39636
rect 18512 39584 18564 39636
rect 18696 39584 18748 39636
rect 25228 39584 25280 39636
rect 25320 39627 25372 39636
rect 25320 39593 25329 39627
rect 25329 39593 25363 39627
rect 25363 39593 25372 39627
rect 25320 39584 25372 39593
rect 9220 39559 9272 39568
rect 9220 39525 9229 39559
rect 9229 39525 9263 39559
rect 9263 39525 9272 39559
rect 9220 39516 9272 39525
rect 10968 39516 11020 39568
rect 15936 39516 15988 39568
rect 17684 39516 17736 39568
rect 11612 39448 11664 39500
rect 14556 39491 14608 39500
rect 14556 39457 14565 39491
rect 14565 39457 14599 39491
rect 14599 39457 14608 39491
rect 14556 39448 14608 39457
rect 15844 39448 15896 39500
rect 16304 39448 16356 39500
rect 16580 39448 16632 39500
rect 17592 39448 17644 39500
rect 9680 39423 9732 39432
rect 9680 39389 9689 39423
rect 9689 39389 9723 39423
rect 9723 39389 9732 39423
rect 9680 39380 9732 39389
rect 16212 39380 16264 39432
rect 16396 39380 16448 39432
rect 17960 39423 18012 39432
rect 17960 39389 17969 39423
rect 17969 39389 18003 39423
rect 18003 39389 18012 39423
rect 17960 39380 18012 39389
rect 18236 39423 18288 39432
rect 18236 39389 18245 39423
rect 18245 39389 18279 39423
rect 18279 39389 18288 39423
rect 18236 39380 18288 39389
rect 18604 39423 18656 39432
rect 18604 39389 18613 39423
rect 18613 39389 18647 39423
rect 18647 39389 18656 39423
rect 18604 39380 18656 39389
rect 18788 39423 18840 39432
rect 18788 39389 18797 39423
rect 18797 39389 18831 39423
rect 18831 39389 18840 39423
rect 18788 39380 18840 39389
rect 18972 39380 19024 39432
rect 19156 39380 19208 39432
rect 9956 39355 10008 39364
rect 9956 39321 9965 39355
rect 9965 39321 9999 39355
rect 9999 39321 10008 39355
rect 9956 39312 10008 39321
rect 10600 39312 10652 39364
rect 12164 39287 12216 39296
rect 12164 39253 12173 39287
rect 12173 39253 12207 39287
rect 12207 39253 12216 39287
rect 12164 39244 12216 39253
rect 15292 39244 15344 39296
rect 15568 39244 15620 39296
rect 16488 39244 16540 39296
rect 18328 39312 18380 39364
rect 17960 39244 18012 39296
rect 18696 39244 18748 39296
rect 18788 39244 18840 39296
rect 19432 39312 19484 39364
rect 19340 39244 19392 39296
rect 19892 39423 19944 39432
rect 19892 39389 19901 39423
rect 19901 39389 19935 39423
rect 19935 39389 19944 39423
rect 19892 39380 19944 39389
rect 20812 39516 20864 39568
rect 23204 39516 23256 39568
rect 23756 39516 23808 39568
rect 24768 39516 24820 39568
rect 23020 39448 23072 39500
rect 24308 39448 24360 39500
rect 25596 39584 25648 39636
rect 25688 39584 25740 39636
rect 26516 39584 26568 39636
rect 28356 39584 28408 39636
rect 29276 39584 29328 39636
rect 29552 39627 29604 39636
rect 29552 39593 29561 39627
rect 29561 39593 29595 39627
rect 29595 39593 29604 39627
rect 29552 39584 29604 39593
rect 30472 39584 30524 39636
rect 31852 39584 31904 39636
rect 32036 39627 32088 39636
rect 32036 39593 32045 39627
rect 32045 39593 32079 39627
rect 32079 39593 32088 39627
rect 32036 39584 32088 39593
rect 39304 39584 39356 39636
rect 20260 39380 20312 39432
rect 26240 39516 26292 39568
rect 26608 39516 26660 39568
rect 31208 39516 31260 39568
rect 29184 39448 29236 39500
rect 29644 39491 29696 39500
rect 29644 39457 29653 39491
rect 29653 39457 29687 39491
rect 29687 39457 29696 39491
rect 29644 39448 29696 39457
rect 29736 39448 29788 39500
rect 20168 39312 20220 39364
rect 24952 39312 25004 39364
rect 25872 39380 25924 39432
rect 26148 39380 26200 39432
rect 27712 39380 27764 39432
rect 28080 39380 28132 39432
rect 28264 39380 28316 39432
rect 28356 39355 28408 39364
rect 20076 39287 20128 39296
rect 20076 39253 20085 39287
rect 20085 39253 20119 39287
rect 20119 39253 20128 39287
rect 20076 39244 20128 39253
rect 23572 39244 23624 39296
rect 24032 39244 24084 39296
rect 24308 39244 24360 39296
rect 24860 39244 24912 39296
rect 25688 39287 25740 39296
rect 25688 39253 25697 39287
rect 25697 39253 25731 39287
rect 25731 39253 25740 39287
rect 25688 39244 25740 39253
rect 25780 39244 25832 39296
rect 28356 39321 28365 39355
rect 28365 39321 28399 39355
rect 28399 39321 28408 39355
rect 28356 39312 28408 39321
rect 28540 39423 28592 39432
rect 28540 39389 28549 39423
rect 28549 39389 28583 39423
rect 28583 39389 28592 39423
rect 28540 39380 28592 39389
rect 29000 39380 29052 39432
rect 30656 39380 30708 39432
rect 27620 39244 27672 39296
rect 30564 39312 30616 39364
rect 30932 39355 30984 39364
rect 30932 39321 30941 39355
rect 30941 39321 30975 39355
rect 30975 39321 30984 39355
rect 30932 39312 30984 39321
rect 28816 39244 28868 39296
rect 28908 39244 28960 39296
rect 29644 39244 29696 39296
rect 29920 39287 29972 39296
rect 29920 39253 29929 39287
rect 29929 39253 29963 39287
rect 29963 39253 29972 39287
rect 29920 39244 29972 39253
rect 31576 39423 31628 39432
rect 31576 39389 31585 39423
rect 31585 39389 31619 39423
rect 31619 39389 31628 39423
rect 31576 39380 31628 39389
rect 37648 39448 37700 39500
rect 31392 39312 31444 39364
rect 32588 39312 32640 39364
rect 33508 39423 33560 39432
rect 33508 39389 33517 39423
rect 33517 39389 33551 39423
rect 33551 39389 33560 39423
rect 33508 39380 33560 39389
rect 38660 39312 38712 39364
rect 31576 39244 31628 39296
rect 31944 39287 31996 39296
rect 31944 39253 31953 39287
rect 31953 39253 31987 39287
rect 31987 39253 31996 39287
rect 31944 39244 31996 39253
rect 32496 39287 32548 39296
rect 32496 39253 32505 39287
rect 32505 39253 32539 39287
rect 32539 39253 32548 39287
rect 32496 39244 32548 39253
rect 32680 39244 32732 39296
rect 33692 39244 33744 39296
rect 39672 39287 39724 39296
rect 39672 39253 39681 39287
rect 39681 39253 39715 39287
rect 39715 39253 39724 39287
rect 39672 39244 39724 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 8300 39040 8352 39092
rect 9588 39040 9640 39092
rect 9864 39040 9916 39092
rect 9956 39040 10008 39092
rect 12164 39040 12216 39092
rect 6920 38836 6972 38888
rect 13636 39040 13688 39092
rect 14556 39040 14608 39092
rect 16488 39040 16540 39092
rect 18880 39040 18932 39092
rect 19800 39040 19852 39092
rect 20260 39083 20312 39092
rect 20260 39049 20269 39083
rect 20269 39049 20303 39083
rect 20303 39049 20312 39083
rect 20260 39040 20312 39049
rect 20536 39040 20588 39092
rect 22376 39040 22428 39092
rect 13544 38972 13596 39024
rect 10416 38904 10468 38956
rect 10968 38904 11020 38956
rect 11428 38904 11480 38956
rect 12716 38947 12768 38956
rect 12716 38913 12725 38947
rect 12725 38913 12759 38947
rect 12759 38913 12768 38947
rect 12716 38904 12768 38913
rect 17960 38972 18012 39024
rect 18144 38972 18196 39024
rect 17776 38947 17828 38956
rect 17776 38913 17785 38947
rect 17785 38913 17819 38947
rect 17819 38913 17828 38947
rect 17776 38904 17828 38913
rect 18052 38947 18104 38956
rect 15292 38836 15344 38888
rect 18052 38913 18061 38947
rect 18061 38913 18095 38947
rect 18095 38913 18104 38947
rect 18052 38904 18104 38913
rect 19432 38904 19484 38956
rect 19984 38904 20036 38956
rect 20076 38904 20128 38956
rect 20536 38947 20588 38956
rect 20536 38913 20545 38947
rect 20545 38913 20579 38947
rect 20579 38913 20588 38947
rect 20536 38904 20588 38913
rect 9036 38768 9088 38820
rect 10600 38768 10652 38820
rect 20168 38836 20220 38888
rect 20720 38947 20772 38956
rect 20720 38913 20755 38947
rect 20755 38913 20772 38947
rect 20720 38904 20772 38913
rect 21456 38972 21508 39024
rect 23020 38972 23072 39024
rect 25504 39040 25556 39092
rect 21088 38836 21140 38888
rect 20628 38768 20680 38820
rect 21732 38904 21784 38956
rect 22192 38904 22244 38956
rect 21548 38836 21600 38888
rect 21640 38879 21692 38888
rect 21640 38845 21649 38879
rect 21649 38845 21683 38879
rect 21683 38845 21692 38879
rect 21640 38836 21692 38845
rect 22284 38836 22336 38888
rect 23020 38836 23072 38888
rect 23204 38904 23256 38956
rect 23296 38947 23348 38956
rect 23296 38913 23305 38947
rect 23305 38913 23339 38947
rect 23339 38913 23348 38947
rect 23296 38904 23348 38913
rect 23480 38947 23532 38956
rect 23480 38913 23489 38947
rect 23489 38913 23523 38947
rect 23523 38913 23532 38947
rect 23480 38904 23532 38913
rect 23848 38904 23900 38956
rect 23940 38947 23992 38956
rect 23940 38913 23949 38947
rect 23949 38913 23983 38947
rect 23983 38913 23992 38947
rect 23940 38904 23992 38913
rect 23388 38836 23440 38888
rect 24032 38836 24084 38888
rect 22008 38768 22060 38820
rect 24308 38947 24360 38956
rect 24308 38913 24317 38947
rect 24317 38913 24351 38947
rect 24351 38913 24360 38947
rect 24308 38904 24360 38913
rect 25044 38972 25096 39024
rect 27068 39040 27120 39092
rect 27620 39083 27672 39092
rect 27620 39049 27629 39083
rect 27629 39049 27663 39083
rect 27663 39049 27672 39083
rect 27620 39040 27672 39049
rect 24768 38768 24820 38820
rect 24952 38947 25004 38956
rect 24952 38913 24961 38947
rect 24961 38913 24995 38947
rect 24995 38913 25004 38947
rect 24952 38904 25004 38913
rect 25228 38947 25280 38956
rect 25228 38913 25237 38947
rect 25237 38913 25271 38947
rect 25271 38913 25280 38947
rect 25228 38904 25280 38913
rect 25504 38947 25556 38956
rect 25504 38913 25513 38947
rect 25513 38913 25547 38947
rect 25547 38913 25556 38947
rect 25504 38904 25556 38913
rect 26056 38904 26108 38956
rect 26148 38947 26200 38956
rect 26148 38913 26157 38947
rect 26157 38913 26191 38947
rect 26191 38913 26200 38947
rect 26148 38904 26200 38913
rect 25964 38836 26016 38888
rect 26516 38947 26568 38956
rect 26516 38913 26525 38947
rect 26525 38913 26559 38947
rect 26559 38913 26568 38947
rect 26516 38904 26568 38913
rect 26700 38836 26752 38888
rect 25044 38768 25096 38820
rect 26148 38768 26200 38820
rect 17592 38700 17644 38752
rect 21180 38700 21232 38752
rect 22100 38700 22152 38752
rect 22376 38700 22428 38752
rect 22560 38743 22612 38752
rect 22560 38709 22569 38743
rect 22569 38709 22603 38743
rect 22603 38709 22612 38743
rect 22560 38700 22612 38709
rect 23756 38700 23808 38752
rect 26240 38700 26292 38752
rect 26516 38768 26568 38820
rect 27712 38947 27764 38956
rect 27712 38913 27721 38947
rect 27721 38913 27755 38947
rect 27755 38913 27764 38947
rect 27712 38904 27764 38913
rect 27896 38947 27948 38956
rect 27896 38913 27905 38947
rect 27905 38913 27939 38947
rect 27939 38913 27948 38947
rect 27896 38904 27948 38913
rect 27988 38947 28040 38956
rect 27988 38913 27997 38947
rect 27997 38913 28031 38947
rect 28031 38913 28040 38947
rect 27988 38904 28040 38913
rect 28540 39040 28592 39092
rect 29552 39040 29604 39092
rect 31484 39083 31536 39092
rect 31484 39049 31493 39083
rect 31493 39049 31527 39083
rect 31527 39049 31536 39083
rect 31484 39040 31536 39049
rect 31576 39040 31628 39092
rect 28632 39015 28684 39024
rect 28632 38981 28641 39015
rect 28641 38981 28675 39015
rect 28675 38981 28684 39015
rect 28632 38972 28684 38981
rect 28816 38972 28868 39024
rect 31024 39015 31076 39024
rect 27620 38836 27672 38888
rect 28540 38700 28592 38752
rect 28724 38700 28776 38752
rect 28816 38700 28868 38752
rect 29644 38947 29696 38956
rect 29644 38913 29653 38947
rect 29653 38913 29687 38947
rect 29687 38913 29696 38947
rect 29644 38904 29696 38913
rect 31024 38981 31033 39015
rect 31033 38981 31067 39015
rect 31067 38981 31076 39015
rect 31024 38972 31076 38981
rect 32496 39040 32548 39092
rect 32588 39083 32640 39092
rect 32588 39049 32597 39083
rect 32597 39049 32631 39083
rect 32631 39049 32640 39083
rect 32588 39040 32640 39049
rect 33508 39040 33560 39092
rect 30104 38904 30156 38956
rect 31576 38947 31628 38956
rect 31576 38913 31585 38947
rect 31585 38913 31619 38947
rect 31619 38913 31628 38947
rect 31576 38904 31628 38913
rect 30472 38836 30524 38888
rect 31116 38879 31168 38888
rect 31116 38845 31125 38879
rect 31125 38845 31159 38879
rect 31159 38845 31168 38879
rect 31116 38836 31168 38845
rect 31944 38972 31996 39024
rect 31760 38947 31812 38956
rect 31760 38913 31769 38947
rect 31769 38913 31803 38947
rect 31803 38913 31812 38947
rect 31760 38904 31812 38913
rect 32128 38947 32180 38956
rect 32128 38913 32137 38947
rect 32137 38913 32171 38947
rect 32171 38913 32180 38947
rect 32128 38904 32180 38913
rect 32220 38879 32272 38888
rect 32220 38845 32229 38879
rect 32229 38845 32263 38879
rect 32263 38845 32272 38879
rect 32220 38836 32272 38845
rect 32404 38947 32456 38956
rect 32404 38913 32413 38947
rect 32413 38913 32447 38947
rect 32447 38913 32456 38947
rect 32404 38904 32456 38913
rect 32772 38947 32824 38956
rect 32772 38913 32781 38947
rect 32781 38913 32815 38947
rect 32815 38913 32824 38947
rect 32772 38904 32824 38913
rect 34612 38972 34664 39024
rect 33600 38947 33652 38956
rect 33600 38913 33609 38947
rect 33609 38913 33643 38947
rect 33643 38913 33652 38947
rect 33600 38904 33652 38913
rect 30288 38743 30340 38752
rect 30288 38709 30297 38743
rect 30297 38709 30331 38743
rect 30331 38709 30340 38743
rect 30288 38700 30340 38709
rect 30656 38743 30708 38752
rect 30656 38709 30665 38743
rect 30665 38709 30699 38743
rect 30699 38709 30708 38743
rect 30656 38700 30708 38709
rect 31024 38743 31076 38752
rect 31024 38709 31033 38743
rect 31033 38709 31067 38743
rect 31067 38709 31076 38743
rect 31024 38700 31076 38709
rect 31208 38700 31260 38752
rect 31852 38700 31904 38752
rect 32680 38743 32732 38752
rect 32680 38709 32689 38743
rect 32689 38709 32723 38743
rect 32723 38709 32732 38743
rect 32680 38700 32732 38709
rect 35348 38743 35400 38752
rect 35348 38709 35357 38743
rect 35357 38709 35391 38743
rect 35391 38709 35400 38743
rect 35348 38700 35400 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 17868 38496 17920 38548
rect 17960 38539 18012 38548
rect 17960 38505 17969 38539
rect 17969 38505 18003 38539
rect 18003 38505 18012 38539
rect 17960 38496 18012 38505
rect 18236 38496 18288 38548
rect 12992 38428 13044 38480
rect 9588 38360 9640 38412
rect 11428 38360 11480 38412
rect 12256 38360 12308 38412
rect 13452 38292 13504 38344
rect 15936 38403 15988 38412
rect 15936 38369 15945 38403
rect 15945 38369 15979 38403
rect 15979 38369 15988 38403
rect 15936 38360 15988 38369
rect 17684 38360 17736 38412
rect 17776 38360 17828 38412
rect 11796 38267 11848 38276
rect 11796 38233 11805 38267
rect 11805 38233 11839 38267
rect 11839 38233 11848 38267
rect 11796 38224 11848 38233
rect 13544 38267 13596 38276
rect 13544 38233 13553 38267
rect 13553 38233 13587 38267
rect 13587 38233 13596 38267
rect 13544 38224 13596 38233
rect 17224 38335 17276 38344
rect 17224 38301 17233 38335
rect 17233 38301 17267 38335
rect 17267 38301 17276 38335
rect 18420 38360 18472 38412
rect 19432 38360 19484 38412
rect 17224 38292 17276 38301
rect 18236 38292 18288 38344
rect 19800 38292 19852 38344
rect 20536 38428 20588 38480
rect 20904 38403 20956 38412
rect 20904 38369 20913 38403
rect 20913 38369 20947 38403
rect 20947 38369 20956 38403
rect 20904 38360 20956 38369
rect 21180 38360 21232 38412
rect 23940 38496 23992 38548
rect 25136 38496 25188 38548
rect 25780 38496 25832 38548
rect 25872 38539 25924 38548
rect 25872 38505 25881 38539
rect 25881 38505 25915 38539
rect 25915 38505 25924 38539
rect 25872 38496 25924 38505
rect 25964 38496 26016 38548
rect 22836 38428 22888 38480
rect 25596 38471 25648 38480
rect 25596 38437 25605 38471
rect 25605 38437 25639 38471
rect 25639 38437 25648 38471
rect 25596 38428 25648 38437
rect 23480 38360 23532 38412
rect 24676 38360 24728 38412
rect 24860 38360 24912 38412
rect 21548 38292 21600 38344
rect 15568 38156 15620 38208
rect 15660 38156 15712 38208
rect 15752 38156 15804 38208
rect 21180 38224 21232 38276
rect 22744 38292 22796 38344
rect 22560 38224 22612 38276
rect 23204 38292 23256 38344
rect 23296 38335 23348 38344
rect 23296 38301 23305 38335
rect 23305 38301 23339 38335
rect 23339 38301 23348 38335
rect 23296 38292 23348 38301
rect 25044 38335 25096 38344
rect 25044 38301 25053 38335
rect 25053 38301 25087 38335
rect 25087 38301 25096 38335
rect 25044 38292 25096 38301
rect 25688 38360 25740 38412
rect 26884 38428 26936 38480
rect 27068 38539 27120 38548
rect 27068 38505 27077 38539
rect 27077 38505 27111 38539
rect 27111 38505 27120 38539
rect 27068 38496 27120 38505
rect 27804 38496 27856 38548
rect 29092 38496 29144 38548
rect 27620 38428 27672 38480
rect 28080 38428 28132 38480
rect 28540 38428 28592 38480
rect 29276 38496 29328 38548
rect 29644 38496 29696 38548
rect 31024 38496 31076 38548
rect 31484 38496 31536 38548
rect 32128 38496 32180 38548
rect 29000 38360 29052 38412
rect 29276 38360 29328 38412
rect 30472 38403 30524 38412
rect 30472 38369 30481 38403
rect 30481 38369 30515 38403
rect 30515 38369 30524 38403
rect 30472 38360 30524 38369
rect 25780 38292 25832 38344
rect 26148 38335 26200 38344
rect 26148 38301 26157 38335
rect 26157 38301 26191 38335
rect 26191 38301 26200 38335
rect 26148 38292 26200 38301
rect 27252 38335 27304 38344
rect 27252 38301 27261 38335
rect 27261 38301 27295 38335
rect 27295 38301 27304 38335
rect 27252 38292 27304 38301
rect 25136 38224 25188 38276
rect 25320 38267 25372 38276
rect 25320 38233 25329 38267
rect 25329 38233 25363 38267
rect 25363 38233 25372 38267
rect 25320 38224 25372 38233
rect 25872 38267 25924 38276
rect 25872 38233 25881 38267
rect 25881 38233 25915 38267
rect 25915 38233 25924 38267
rect 25872 38224 25924 38233
rect 27620 38292 27672 38344
rect 27896 38292 27948 38344
rect 30564 38292 30616 38344
rect 27712 38224 27764 38276
rect 28724 38224 28776 38276
rect 29828 38224 29880 38276
rect 30012 38224 30064 38276
rect 30380 38267 30432 38276
rect 30380 38233 30389 38267
rect 30389 38233 30423 38267
rect 30423 38233 30432 38267
rect 30380 38224 30432 38233
rect 16488 38199 16540 38208
rect 16488 38165 16497 38199
rect 16497 38165 16531 38199
rect 16531 38165 16540 38199
rect 16488 38156 16540 38165
rect 16580 38199 16632 38208
rect 16580 38165 16589 38199
rect 16589 38165 16623 38199
rect 16623 38165 16632 38199
rect 16580 38156 16632 38165
rect 16672 38156 16724 38208
rect 16764 38199 16816 38208
rect 16764 38165 16773 38199
rect 16773 38165 16807 38199
rect 16807 38165 16816 38199
rect 16764 38156 16816 38165
rect 19340 38156 19392 38208
rect 21548 38156 21600 38208
rect 22284 38156 22336 38208
rect 23296 38156 23348 38208
rect 24952 38156 25004 38208
rect 26884 38156 26936 38208
rect 30196 38156 30248 38208
rect 30288 38156 30340 38208
rect 30840 38199 30892 38208
rect 30840 38165 30849 38199
rect 30849 38165 30883 38199
rect 30883 38165 30892 38199
rect 30840 38156 30892 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 11796 37952 11848 38004
rect 13084 37952 13136 38004
rect 9036 37884 9088 37936
rect 10600 37884 10652 37936
rect 11980 37884 12032 37936
rect 12440 37884 12492 37936
rect 14280 37884 14332 37936
rect 12992 37816 13044 37868
rect 13084 37859 13136 37868
rect 13084 37825 13093 37859
rect 13093 37825 13127 37859
rect 13127 37825 13136 37859
rect 13084 37816 13136 37825
rect 6920 37748 6972 37800
rect 7564 37791 7616 37800
rect 7564 37757 7573 37791
rect 7573 37757 7607 37791
rect 7607 37757 7616 37791
rect 7564 37748 7616 37757
rect 8576 37748 8628 37800
rect 9588 37791 9640 37800
rect 9588 37757 9597 37791
rect 9597 37757 9631 37791
rect 9631 37757 9640 37791
rect 9588 37748 9640 37757
rect 11520 37748 11572 37800
rect 12440 37748 12492 37800
rect 13636 37816 13688 37868
rect 15016 37816 15068 37868
rect 15660 37884 15712 37936
rect 15568 37859 15620 37868
rect 13544 37791 13596 37800
rect 13544 37757 13553 37791
rect 13553 37757 13587 37791
rect 13587 37757 13596 37791
rect 13544 37748 13596 37757
rect 15568 37825 15577 37859
rect 15577 37825 15611 37859
rect 15611 37825 15620 37859
rect 15568 37816 15620 37825
rect 16028 37816 16080 37868
rect 16120 37859 16172 37868
rect 16120 37825 16129 37859
rect 16129 37825 16163 37859
rect 16163 37825 16172 37859
rect 16120 37816 16172 37825
rect 15384 37748 15436 37800
rect 16396 37859 16448 37868
rect 16396 37825 16405 37859
rect 16405 37825 16439 37859
rect 16439 37825 16448 37859
rect 16396 37816 16448 37825
rect 15844 37791 15896 37800
rect 15844 37757 15853 37791
rect 15853 37757 15887 37791
rect 15887 37757 15896 37791
rect 15844 37748 15896 37757
rect 16304 37748 16356 37800
rect 16672 37748 16724 37800
rect 17224 37952 17276 38004
rect 17868 37952 17920 38004
rect 16948 37859 17000 37868
rect 16948 37825 16957 37859
rect 16957 37825 16991 37859
rect 16991 37825 17000 37859
rect 16948 37816 17000 37825
rect 18880 37816 18932 37868
rect 19432 37995 19484 38004
rect 19432 37961 19457 37995
rect 19457 37961 19484 37995
rect 19432 37952 19484 37961
rect 19984 37952 20036 38004
rect 23296 37952 23348 38004
rect 25596 37952 25648 38004
rect 26516 37952 26568 38004
rect 26884 37952 26936 38004
rect 20444 37884 20496 37936
rect 21548 37884 21600 37936
rect 21732 37884 21784 37936
rect 22652 37884 22704 37936
rect 23112 37884 23164 37936
rect 27528 37952 27580 38004
rect 27620 37995 27672 38004
rect 27620 37961 27629 37995
rect 27629 37961 27663 37995
rect 27663 37961 27672 37995
rect 27620 37952 27672 37961
rect 19340 37748 19392 37800
rect 19984 37859 20036 37868
rect 19984 37825 19993 37859
rect 19993 37825 20027 37859
rect 20027 37825 20036 37859
rect 19984 37816 20036 37825
rect 20720 37816 20772 37868
rect 22376 37816 22428 37868
rect 22836 37816 22888 37868
rect 23296 37859 23348 37868
rect 23296 37825 23305 37859
rect 23305 37825 23339 37859
rect 23339 37825 23348 37859
rect 23296 37816 23348 37825
rect 20076 37748 20128 37800
rect 21732 37748 21784 37800
rect 22192 37748 22244 37800
rect 22744 37748 22796 37800
rect 24124 37816 24176 37868
rect 24492 37816 24544 37868
rect 24676 37816 24728 37868
rect 26700 37816 26752 37868
rect 26976 37859 27028 37868
rect 26976 37825 26985 37859
rect 26985 37825 27019 37859
rect 27019 37825 27028 37859
rect 26976 37816 27028 37825
rect 24952 37748 25004 37800
rect 25136 37748 25188 37800
rect 25964 37748 26016 37800
rect 26424 37748 26476 37800
rect 27712 37816 27764 37868
rect 27804 37816 27856 37868
rect 28356 37927 28408 37936
rect 28356 37893 28361 37927
rect 28361 37893 28395 37927
rect 28395 37893 28408 37927
rect 28356 37884 28408 37893
rect 27528 37748 27580 37800
rect 18420 37680 18472 37732
rect 18512 37680 18564 37732
rect 9036 37655 9088 37664
rect 9036 37621 9045 37655
rect 9045 37621 9079 37655
rect 9079 37621 9088 37655
rect 9036 37612 9088 37621
rect 10324 37612 10376 37664
rect 12164 37612 12216 37664
rect 15476 37612 15528 37664
rect 15752 37655 15804 37664
rect 15752 37621 15761 37655
rect 15761 37621 15795 37655
rect 15795 37621 15804 37655
rect 15752 37612 15804 37621
rect 18788 37612 18840 37664
rect 18880 37655 18932 37664
rect 18880 37621 18889 37655
rect 18889 37621 18923 37655
rect 18923 37621 18932 37655
rect 18880 37612 18932 37621
rect 28632 37995 28684 38004
rect 28632 37961 28641 37995
rect 28641 37961 28675 37995
rect 28675 37961 28684 37995
rect 28632 37952 28684 37961
rect 29000 37952 29052 38004
rect 29276 37927 29328 37936
rect 29276 37893 29285 37927
rect 29285 37893 29319 37927
rect 29319 37893 29328 37927
rect 29276 37884 29328 37893
rect 30104 37952 30156 38004
rect 30840 37952 30892 38004
rect 29092 37859 29144 37868
rect 29092 37825 29102 37859
rect 29102 37825 29136 37859
rect 29136 37825 29144 37859
rect 29092 37816 29144 37825
rect 30012 37816 30064 37868
rect 28264 37748 28316 37800
rect 28632 37748 28684 37800
rect 30564 37748 30616 37800
rect 27804 37680 27856 37732
rect 30472 37680 30524 37732
rect 33600 37952 33652 38004
rect 34428 37952 34480 38004
rect 31300 37816 31352 37868
rect 31668 37816 31720 37868
rect 32220 37859 32272 37868
rect 32220 37825 32229 37859
rect 32229 37825 32263 37859
rect 32263 37825 32272 37859
rect 32220 37816 32272 37825
rect 33692 37884 33744 37936
rect 38568 37884 38620 37936
rect 31208 37748 31260 37800
rect 31944 37748 31996 37800
rect 23388 37612 23440 37664
rect 23480 37612 23532 37664
rect 31116 37612 31168 37664
rect 31484 37655 31536 37664
rect 31484 37621 31493 37655
rect 31493 37621 31527 37655
rect 31527 37621 31536 37655
rect 31484 37612 31536 37621
rect 33140 37612 33192 37664
rect 34796 37612 34848 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 7564 37408 7616 37460
rect 11520 37451 11572 37460
rect 11520 37417 11529 37451
rect 11529 37417 11563 37451
rect 11563 37417 11572 37451
rect 11520 37408 11572 37417
rect 15752 37408 15804 37460
rect 16304 37408 16356 37460
rect 18328 37408 18380 37460
rect 20720 37408 20772 37460
rect 21364 37408 21416 37460
rect 22284 37408 22336 37460
rect 23388 37408 23440 37460
rect 23480 37451 23532 37460
rect 23480 37417 23489 37451
rect 23489 37417 23523 37451
rect 23523 37417 23532 37451
rect 23480 37408 23532 37417
rect 25964 37451 26016 37460
rect 25964 37417 25973 37451
rect 25973 37417 26007 37451
rect 26007 37417 26016 37451
rect 25964 37408 26016 37417
rect 26884 37408 26936 37460
rect 29092 37408 29144 37460
rect 29828 37408 29880 37460
rect 30288 37451 30340 37460
rect 30288 37417 30297 37451
rect 30297 37417 30331 37451
rect 30331 37417 30340 37451
rect 30288 37408 30340 37417
rect 30564 37408 30616 37460
rect 8668 37247 8720 37256
rect 8668 37213 8677 37247
rect 8677 37213 8711 37247
rect 8711 37213 8720 37247
rect 8668 37204 8720 37213
rect 9036 37247 9088 37256
rect 9036 37213 9045 37247
rect 9045 37213 9079 37247
rect 9079 37213 9088 37247
rect 9036 37204 9088 37213
rect 12532 37340 12584 37392
rect 12900 37340 12952 37392
rect 18880 37340 18932 37392
rect 21548 37340 21600 37392
rect 10324 37315 10376 37324
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 10324 37272 10376 37281
rect 11336 37247 11388 37256
rect 11336 37213 11345 37247
rect 11345 37213 11379 37247
rect 11379 37213 11388 37247
rect 11336 37204 11388 37213
rect 11520 37272 11572 37324
rect 11152 37179 11204 37188
rect 11152 37145 11161 37179
rect 11161 37145 11195 37179
rect 11195 37145 11204 37179
rect 11152 37136 11204 37145
rect 11980 37136 12032 37188
rect 13084 37204 13136 37256
rect 15016 37247 15068 37256
rect 15016 37213 15025 37247
rect 15025 37213 15059 37247
rect 15059 37213 15068 37247
rect 15016 37204 15068 37213
rect 15476 37272 15528 37324
rect 16488 37272 16540 37324
rect 15292 37247 15344 37256
rect 15292 37213 15301 37247
rect 15301 37213 15335 37247
rect 15335 37213 15344 37247
rect 15292 37204 15344 37213
rect 15752 37247 15804 37256
rect 15752 37213 15761 37247
rect 15761 37213 15795 37247
rect 15795 37213 15804 37247
rect 15752 37204 15804 37213
rect 15936 37204 15988 37256
rect 16028 37204 16080 37256
rect 16580 37204 16632 37256
rect 12716 37068 12768 37120
rect 12992 37068 13044 37120
rect 13636 37136 13688 37188
rect 15660 37136 15712 37188
rect 17224 37136 17276 37188
rect 13176 37068 13228 37120
rect 14280 37068 14332 37120
rect 15016 37068 15068 37120
rect 15384 37068 15436 37120
rect 18144 37204 18196 37256
rect 19156 37272 19208 37324
rect 22192 37272 22244 37324
rect 17776 37179 17828 37188
rect 17776 37145 17785 37179
rect 17785 37145 17819 37179
rect 17819 37145 17828 37179
rect 17776 37136 17828 37145
rect 17960 37068 18012 37120
rect 19432 37204 19484 37256
rect 20536 37204 20588 37256
rect 24492 37340 24544 37392
rect 25228 37340 25280 37392
rect 25504 37340 25556 37392
rect 25964 37272 26016 37324
rect 20996 37136 21048 37188
rect 22744 37136 22796 37188
rect 23020 37247 23072 37256
rect 23020 37213 23029 37247
rect 23029 37213 23063 37247
rect 23063 37213 23072 37247
rect 23020 37204 23072 37213
rect 23112 37204 23164 37256
rect 23388 37204 23440 37256
rect 23480 37204 23532 37256
rect 23664 37136 23716 37188
rect 25044 37204 25096 37256
rect 25596 37247 25648 37256
rect 25596 37213 25605 37247
rect 25605 37213 25639 37247
rect 25639 37213 25648 37247
rect 25596 37204 25648 37213
rect 25688 37247 25740 37256
rect 25688 37213 25697 37247
rect 25697 37213 25731 37247
rect 25731 37213 25740 37247
rect 25688 37204 25740 37213
rect 25780 37247 25832 37256
rect 25780 37213 25789 37247
rect 25789 37213 25823 37247
rect 25823 37213 25832 37247
rect 25780 37204 25832 37213
rect 26332 37204 26384 37256
rect 26976 37340 27028 37392
rect 27620 37272 27672 37324
rect 28724 37272 28776 37324
rect 30104 37272 30156 37324
rect 30472 37340 30524 37392
rect 31024 37340 31076 37392
rect 26424 37179 26476 37188
rect 26424 37145 26433 37179
rect 26433 37145 26467 37179
rect 26467 37145 26476 37179
rect 26424 37136 26476 37145
rect 26516 37179 26568 37188
rect 26516 37145 26525 37179
rect 26525 37145 26559 37179
rect 26559 37145 26568 37179
rect 26516 37136 26568 37145
rect 18604 37111 18656 37120
rect 18604 37077 18613 37111
rect 18613 37077 18647 37111
rect 18647 37077 18656 37111
rect 18604 37068 18656 37077
rect 18880 37068 18932 37120
rect 20536 37111 20588 37120
rect 20536 37077 20545 37111
rect 20545 37077 20579 37111
rect 20579 37077 20588 37111
rect 20536 37068 20588 37077
rect 23388 37068 23440 37120
rect 24400 37068 24452 37120
rect 25412 37068 25464 37120
rect 26976 37247 27028 37256
rect 26976 37213 26986 37247
rect 26986 37213 27020 37247
rect 27020 37213 27028 37247
rect 26976 37204 27028 37213
rect 27528 37204 27580 37256
rect 28264 37204 28316 37256
rect 28540 37204 28592 37256
rect 28632 37204 28684 37256
rect 29368 37204 29420 37256
rect 30012 37204 30064 37256
rect 27988 37136 28040 37188
rect 28724 37136 28776 37188
rect 29000 37136 29052 37188
rect 29736 37179 29788 37188
rect 29736 37145 29745 37179
rect 29745 37145 29779 37179
rect 29779 37145 29788 37179
rect 29736 37136 29788 37145
rect 30104 37136 30156 37188
rect 30196 37179 30248 37188
rect 30196 37145 30205 37179
rect 30205 37145 30239 37179
rect 30239 37145 30248 37179
rect 30196 37136 30248 37145
rect 27344 37068 27396 37120
rect 31208 37272 31260 37324
rect 30656 37204 30708 37256
rect 30840 37247 30892 37256
rect 30840 37213 30849 37247
rect 30849 37213 30883 37247
rect 30883 37213 30892 37247
rect 30840 37204 30892 37213
rect 30932 37247 30984 37256
rect 30932 37213 30942 37247
rect 30942 37213 30976 37247
rect 30976 37213 30984 37247
rect 30932 37204 30984 37213
rect 31208 37179 31260 37188
rect 31208 37145 31217 37179
rect 31217 37145 31251 37179
rect 31251 37145 31260 37179
rect 31208 37136 31260 37145
rect 32312 37247 32364 37256
rect 32312 37213 32321 37247
rect 32321 37213 32355 37247
rect 32355 37213 32364 37247
rect 32312 37204 32364 37213
rect 32404 37247 32456 37256
rect 32404 37213 32413 37247
rect 32413 37213 32447 37247
rect 32447 37213 32456 37247
rect 32404 37204 32456 37213
rect 33140 37204 33192 37256
rect 37556 37204 37608 37256
rect 31576 37136 31628 37188
rect 32128 37179 32180 37188
rect 32128 37145 32137 37179
rect 32137 37145 32171 37179
rect 32171 37145 32180 37179
rect 32128 37136 32180 37145
rect 31484 37111 31536 37120
rect 31484 37077 31493 37111
rect 31493 37077 31527 37111
rect 31527 37077 31536 37111
rect 31484 37068 31536 37077
rect 32588 37111 32640 37120
rect 32588 37077 32597 37111
rect 32597 37077 32631 37111
rect 32631 37077 32640 37111
rect 32588 37068 32640 37077
rect 33416 37111 33468 37120
rect 33416 37077 33425 37111
rect 33425 37077 33459 37111
rect 33459 37077 33468 37111
rect 33416 37068 33468 37077
rect 40960 37111 41012 37120
rect 40960 37077 40969 37111
rect 40969 37077 41003 37111
rect 41003 37077 41012 37111
rect 40960 37068 41012 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 8668 36864 8720 36916
rect 9312 36864 9364 36916
rect 11520 36864 11572 36916
rect 8576 36796 8628 36848
rect 8760 36796 8812 36848
rect 9772 36728 9824 36780
rect 11152 36796 11204 36848
rect 12072 36907 12124 36916
rect 12072 36873 12081 36907
rect 12081 36873 12115 36907
rect 12115 36873 12124 36907
rect 12072 36864 12124 36873
rect 13360 36864 13412 36916
rect 13452 36864 13504 36916
rect 10784 36771 10836 36780
rect 10784 36737 10793 36771
rect 10793 36737 10827 36771
rect 10827 36737 10836 36771
rect 10784 36728 10836 36737
rect 11336 36728 11388 36780
rect 11428 36728 11480 36780
rect 11520 36771 11572 36780
rect 11520 36737 11529 36771
rect 11529 36737 11563 36771
rect 11563 36737 11572 36771
rect 11520 36728 11572 36737
rect 12532 36839 12584 36848
rect 12532 36805 12541 36839
rect 12541 36805 12575 36839
rect 12575 36805 12584 36839
rect 12532 36796 12584 36805
rect 11796 36771 11848 36780
rect 11796 36737 11805 36771
rect 11805 36737 11839 36771
rect 11839 36737 11848 36771
rect 11796 36728 11848 36737
rect 11980 36728 12032 36780
rect 15200 36864 15252 36916
rect 16212 36907 16264 36916
rect 16212 36873 16221 36907
rect 16221 36873 16255 36907
rect 16255 36873 16264 36907
rect 16212 36864 16264 36873
rect 18512 36864 18564 36916
rect 18604 36864 18656 36916
rect 14280 36839 14332 36848
rect 14280 36805 14289 36839
rect 14289 36805 14323 36839
rect 14323 36805 14332 36839
rect 14280 36796 14332 36805
rect 15752 36839 15804 36848
rect 15752 36805 15761 36839
rect 15761 36805 15795 36839
rect 15795 36805 15804 36839
rect 15752 36796 15804 36805
rect 15384 36771 15436 36780
rect 15384 36737 15393 36771
rect 15393 36737 15427 36771
rect 15427 36737 15436 36771
rect 15384 36728 15436 36737
rect 16396 36796 16448 36848
rect 16488 36728 16540 36780
rect 16580 36728 16632 36780
rect 16764 36728 16816 36780
rect 17684 36796 17736 36848
rect 18052 36796 18104 36848
rect 9772 36567 9824 36576
rect 9772 36533 9781 36567
rect 9781 36533 9815 36567
rect 9815 36533 9824 36567
rect 9772 36524 9824 36533
rect 16304 36660 16356 36712
rect 18144 36771 18196 36780
rect 18144 36737 18153 36771
rect 18153 36737 18187 36771
rect 18187 36737 18196 36771
rect 18144 36728 18196 36737
rect 19248 36796 19300 36848
rect 19892 36796 19944 36848
rect 10048 36635 10100 36644
rect 10048 36601 10057 36635
rect 10057 36601 10091 36635
rect 10091 36601 10100 36635
rect 10048 36592 10100 36601
rect 17960 36660 18012 36712
rect 18512 36771 18564 36780
rect 18512 36737 18521 36771
rect 18521 36737 18555 36771
rect 18555 36737 18564 36771
rect 18512 36728 18564 36737
rect 19064 36771 19116 36780
rect 19064 36737 19073 36771
rect 19073 36737 19107 36771
rect 19107 36737 19116 36771
rect 19064 36728 19116 36737
rect 19156 36728 19208 36780
rect 20812 36796 20864 36848
rect 20996 36796 21048 36848
rect 20444 36728 20496 36780
rect 21272 36728 21324 36780
rect 21364 36728 21416 36780
rect 16764 36592 16816 36644
rect 18236 36592 18288 36644
rect 18880 36592 18932 36644
rect 19064 36592 19116 36644
rect 19524 36703 19576 36712
rect 19524 36669 19533 36703
rect 19533 36669 19567 36703
rect 19567 36669 19576 36703
rect 19524 36660 19576 36669
rect 19984 36660 20036 36712
rect 11520 36524 11572 36576
rect 15016 36524 15068 36576
rect 16672 36567 16724 36576
rect 16672 36533 16681 36567
rect 16681 36533 16715 36567
rect 16715 36533 16724 36567
rect 16672 36524 16724 36533
rect 17960 36524 18012 36576
rect 18788 36524 18840 36576
rect 19156 36524 19208 36576
rect 19432 36567 19484 36576
rect 19432 36533 19441 36567
rect 19441 36533 19475 36567
rect 19475 36533 19484 36567
rect 19432 36524 19484 36533
rect 20352 36592 20404 36644
rect 20168 36524 20220 36576
rect 20628 36703 20680 36712
rect 20628 36669 20637 36703
rect 20637 36669 20671 36703
rect 20671 36669 20680 36703
rect 20628 36660 20680 36669
rect 20996 36703 21048 36712
rect 20996 36669 21005 36703
rect 21005 36669 21039 36703
rect 21039 36669 21048 36703
rect 20996 36660 21048 36669
rect 21548 36660 21600 36712
rect 22560 36864 22612 36916
rect 23204 36796 23256 36848
rect 26608 36864 26660 36916
rect 27344 36864 27396 36916
rect 24216 36796 24268 36848
rect 22744 36771 22796 36780
rect 22744 36737 22753 36771
rect 22753 36737 22787 36771
rect 22787 36737 22796 36771
rect 22744 36728 22796 36737
rect 22836 36771 22888 36780
rect 22836 36737 22845 36771
rect 22845 36737 22879 36771
rect 22879 36737 22888 36771
rect 22836 36728 22888 36737
rect 21916 36703 21968 36712
rect 21916 36669 21925 36703
rect 21925 36669 21959 36703
rect 21959 36669 21968 36703
rect 21916 36660 21968 36669
rect 22100 36703 22152 36712
rect 22100 36669 22109 36703
rect 22109 36669 22143 36703
rect 22143 36669 22152 36703
rect 22100 36660 22152 36669
rect 22192 36703 22244 36712
rect 22192 36669 22201 36703
rect 22201 36669 22235 36703
rect 22235 36669 22244 36703
rect 22192 36660 22244 36669
rect 23480 36728 23532 36780
rect 24308 36750 24360 36802
rect 24676 36796 24728 36848
rect 25596 36796 25648 36848
rect 25964 36796 26016 36848
rect 28264 36864 28316 36916
rect 28816 36864 28868 36916
rect 29828 36864 29880 36916
rect 30932 36864 30984 36916
rect 31484 36864 31536 36916
rect 24216 36703 24268 36712
rect 24216 36669 24225 36703
rect 24225 36669 24259 36703
rect 24259 36669 24268 36703
rect 24216 36660 24268 36669
rect 24952 36728 25004 36780
rect 25412 36771 25464 36780
rect 25412 36737 25421 36771
rect 25421 36737 25455 36771
rect 25455 36737 25464 36771
rect 25412 36728 25464 36737
rect 25504 36771 25556 36780
rect 25504 36737 25514 36771
rect 25514 36737 25548 36771
rect 25548 36737 25556 36771
rect 25504 36728 25556 36737
rect 25780 36771 25832 36780
rect 25780 36737 25789 36771
rect 25789 36737 25823 36771
rect 25823 36737 25832 36771
rect 25780 36728 25832 36737
rect 24676 36635 24728 36644
rect 24676 36601 24685 36635
rect 24685 36601 24719 36635
rect 24719 36601 24728 36635
rect 24676 36592 24728 36601
rect 25228 36592 25280 36644
rect 26792 36660 26844 36712
rect 28908 36796 28960 36848
rect 29000 36796 29052 36848
rect 28448 36728 28500 36780
rect 27988 36703 28040 36712
rect 27988 36669 27997 36703
rect 27997 36669 28031 36703
rect 28031 36669 28040 36703
rect 27988 36660 28040 36669
rect 28816 36771 28868 36780
rect 28816 36737 28825 36771
rect 28825 36737 28859 36771
rect 28859 36737 28868 36771
rect 28816 36728 28868 36737
rect 30932 36728 30984 36780
rect 31576 36796 31628 36848
rect 31668 36796 31720 36848
rect 32220 36864 32272 36916
rect 32404 36864 32456 36916
rect 32588 36864 32640 36916
rect 33416 36864 33468 36916
rect 32036 36796 32088 36848
rect 34612 36796 34664 36848
rect 28908 36703 28960 36712
rect 28908 36669 28917 36703
rect 28917 36669 28951 36703
rect 28951 36669 28960 36703
rect 28908 36660 28960 36669
rect 22560 36567 22612 36576
rect 22560 36533 22569 36567
rect 22569 36533 22603 36567
rect 22603 36533 22612 36567
rect 22560 36524 22612 36533
rect 25964 36524 26016 36576
rect 28264 36524 28316 36576
rect 28356 36567 28408 36576
rect 28356 36533 28365 36567
rect 28365 36533 28399 36567
rect 28399 36533 28408 36567
rect 28356 36524 28408 36533
rect 31392 36635 31444 36644
rect 31392 36601 31401 36635
rect 31401 36601 31435 36635
rect 31435 36601 31444 36635
rect 33600 36728 33652 36780
rect 31392 36592 31444 36601
rect 31484 36567 31536 36576
rect 31484 36533 31493 36567
rect 31493 36533 31527 36567
rect 31527 36533 31536 36567
rect 31484 36524 31536 36533
rect 31944 36524 31996 36576
rect 33232 36524 33284 36576
rect 35532 36567 35584 36576
rect 35532 36533 35541 36567
rect 35541 36533 35575 36567
rect 35575 36533 35584 36567
rect 35532 36524 35584 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 12072 36320 12124 36372
rect 12716 36252 12768 36304
rect 16488 36363 16540 36372
rect 16488 36329 16497 36363
rect 16497 36329 16531 36363
rect 16531 36329 16540 36363
rect 16488 36320 16540 36329
rect 16948 36320 17000 36372
rect 19156 36320 19208 36372
rect 6000 36116 6052 36168
rect 6828 36184 6880 36236
rect 11428 36227 11480 36236
rect 11428 36193 11437 36227
rect 11437 36193 11471 36227
rect 11471 36193 11480 36227
rect 11428 36184 11480 36193
rect 17592 36184 17644 36236
rect 4804 36048 4856 36100
rect 940 35980 992 36032
rect 7104 35980 7156 36032
rect 8760 36116 8812 36168
rect 9312 36116 9364 36168
rect 10048 36116 10100 36168
rect 15844 36116 15896 36168
rect 18144 36184 18196 36236
rect 18420 36184 18472 36236
rect 18880 36252 18932 36304
rect 19248 36184 19300 36236
rect 19432 36363 19484 36372
rect 19432 36329 19441 36363
rect 19441 36329 19475 36363
rect 19475 36329 19484 36363
rect 19432 36320 19484 36329
rect 19892 36320 19944 36372
rect 20168 36363 20220 36372
rect 20168 36329 20177 36363
rect 20177 36329 20211 36363
rect 20211 36329 20220 36363
rect 20168 36320 20220 36329
rect 20444 36320 20496 36372
rect 20628 36363 20680 36372
rect 20628 36329 20637 36363
rect 20637 36329 20671 36363
rect 20671 36329 20680 36363
rect 20628 36320 20680 36329
rect 22192 36320 22244 36372
rect 24400 36320 24452 36372
rect 25044 36320 25096 36372
rect 25412 36320 25464 36372
rect 26700 36320 26752 36372
rect 20352 36252 20404 36304
rect 22928 36252 22980 36304
rect 23296 36252 23348 36304
rect 23664 36252 23716 36304
rect 17776 36116 17828 36168
rect 19432 36116 19484 36168
rect 23848 36184 23900 36236
rect 24860 36184 24912 36236
rect 20444 36159 20496 36168
rect 20444 36125 20453 36159
rect 20453 36125 20487 36159
rect 20487 36125 20496 36159
rect 20444 36116 20496 36125
rect 20536 36116 20588 36168
rect 20812 36116 20864 36168
rect 22192 36116 22244 36168
rect 22560 36116 22612 36168
rect 22652 36159 22704 36168
rect 22652 36125 22661 36159
rect 22661 36125 22695 36159
rect 22695 36125 22704 36159
rect 22652 36116 22704 36125
rect 22744 36159 22796 36168
rect 22744 36125 22753 36159
rect 22753 36125 22787 36159
rect 22787 36125 22796 36159
rect 22744 36116 22796 36125
rect 23572 36159 23624 36168
rect 23572 36125 23581 36159
rect 23581 36125 23615 36159
rect 23615 36125 23624 36159
rect 23572 36116 23624 36125
rect 23664 36159 23716 36168
rect 23664 36125 23674 36159
rect 23674 36125 23708 36159
rect 23708 36125 23716 36159
rect 23664 36116 23716 36125
rect 23940 36159 23992 36168
rect 23940 36125 23949 36159
rect 23949 36125 23983 36159
rect 23983 36125 23992 36159
rect 23940 36116 23992 36125
rect 24676 36116 24728 36168
rect 25412 36116 25464 36168
rect 25596 36116 25648 36168
rect 8852 36048 8904 36100
rect 10508 36048 10560 36100
rect 10692 36091 10744 36100
rect 10692 36057 10701 36091
rect 10701 36057 10735 36091
rect 10735 36057 10744 36091
rect 10692 36048 10744 36057
rect 11336 36048 11388 36100
rect 12256 36048 12308 36100
rect 12348 36048 12400 36100
rect 14188 36048 14240 36100
rect 15016 36048 15068 36100
rect 16672 36048 16724 36100
rect 17960 36048 18012 36100
rect 19064 36048 19116 36100
rect 19248 36091 19300 36100
rect 19248 36057 19257 36091
rect 19257 36057 19291 36091
rect 19291 36057 19300 36091
rect 19248 36048 19300 36057
rect 20628 36048 20680 36100
rect 23848 36091 23900 36100
rect 23848 36057 23857 36091
rect 23857 36057 23891 36091
rect 23891 36057 23900 36091
rect 23848 36048 23900 36057
rect 9128 36023 9180 36032
rect 9128 35989 9137 36023
rect 9137 35989 9171 36023
rect 9171 35989 9180 36023
rect 9128 35980 9180 35989
rect 11796 35980 11848 36032
rect 12808 35980 12860 36032
rect 18696 35980 18748 36032
rect 24952 36048 25004 36100
rect 25136 36091 25188 36100
rect 25136 36057 25145 36091
rect 25145 36057 25179 36091
rect 25179 36057 25188 36091
rect 25136 36048 25188 36057
rect 25228 36091 25280 36100
rect 25228 36057 25237 36091
rect 25237 36057 25271 36091
rect 25271 36057 25280 36091
rect 25228 36048 25280 36057
rect 26976 36252 27028 36304
rect 25964 36159 26016 36168
rect 25964 36125 25973 36159
rect 25973 36125 26007 36159
rect 26007 36125 26016 36159
rect 25964 36116 26016 36125
rect 26700 36184 26752 36236
rect 26792 36116 26844 36168
rect 27620 36320 27672 36372
rect 28724 36320 28776 36372
rect 29368 36320 29420 36372
rect 31208 36363 31260 36372
rect 31208 36329 31217 36363
rect 31217 36329 31251 36363
rect 31251 36329 31260 36363
rect 31208 36320 31260 36329
rect 32128 36320 32180 36372
rect 27896 36252 27948 36304
rect 27712 36159 27764 36168
rect 27712 36125 27721 36159
rect 27721 36125 27755 36159
rect 27755 36125 27764 36159
rect 27712 36116 27764 36125
rect 27896 36116 27948 36168
rect 28356 36252 28408 36304
rect 28448 36252 28500 36304
rect 31944 36252 31996 36304
rect 28724 36184 28776 36236
rect 31300 36184 31352 36236
rect 31392 36227 31444 36236
rect 31392 36193 31401 36227
rect 31401 36193 31435 36227
rect 31435 36193 31444 36227
rect 31392 36184 31444 36193
rect 26976 36048 27028 36100
rect 26148 35980 26200 36032
rect 27252 35980 27304 36032
rect 28724 36048 28776 36100
rect 29920 36048 29972 36100
rect 33600 36184 33652 36236
rect 37280 36048 37332 36100
rect 32496 35980 32548 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 7104 35708 7156 35760
rect 8944 35683 8996 35692
rect 8944 35649 8953 35683
rect 8953 35649 8987 35683
rect 8987 35649 8996 35683
rect 8944 35640 8996 35649
rect 9496 35776 9548 35828
rect 6000 35572 6052 35624
rect 6736 35615 6788 35624
rect 6736 35581 6745 35615
rect 6745 35581 6779 35615
rect 6779 35581 6788 35615
rect 6736 35572 6788 35581
rect 9036 35572 9088 35624
rect 10232 35776 10284 35828
rect 12348 35776 12400 35828
rect 14004 35776 14056 35828
rect 15200 35776 15252 35828
rect 22744 35776 22796 35828
rect 23020 35819 23072 35828
rect 23020 35785 23029 35819
rect 23029 35785 23063 35819
rect 23063 35785 23072 35819
rect 23020 35776 23072 35785
rect 23572 35776 23624 35828
rect 10140 35572 10192 35624
rect 10784 35683 10836 35692
rect 10784 35649 10793 35683
rect 10793 35649 10827 35683
rect 10827 35649 10836 35683
rect 12808 35708 12860 35760
rect 12992 35708 13044 35760
rect 21548 35708 21600 35760
rect 10784 35640 10836 35649
rect 19892 35640 19944 35692
rect 21272 35640 21324 35692
rect 21732 35640 21784 35692
rect 23940 35708 23992 35760
rect 22284 35640 22336 35692
rect 22928 35640 22980 35692
rect 8024 35504 8076 35556
rect 10876 35504 10928 35556
rect 11704 35504 11756 35556
rect 11888 35504 11940 35556
rect 12992 35504 13044 35556
rect 9312 35436 9364 35488
rect 9864 35479 9916 35488
rect 9864 35445 9873 35479
rect 9873 35445 9907 35479
rect 9907 35445 9916 35479
rect 9864 35436 9916 35445
rect 10048 35479 10100 35488
rect 10048 35445 10057 35479
rect 10057 35445 10091 35479
rect 10091 35445 10100 35479
rect 10048 35436 10100 35445
rect 10232 35436 10284 35488
rect 11612 35436 11664 35488
rect 12624 35436 12676 35488
rect 12716 35436 12768 35488
rect 14740 35572 14792 35624
rect 20628 35572 20680 35624
rect 22376 35615 22428 35624
rect 22376 35581 22385 35615
rect 22385 35581 22419 35615
rect 22419 35581 22428 35615
rect 22376 35572 22428 35581
rect 23296 35683 23348 35692
rect 23296 35649 23306 35683
rect 23306 35649 23340 35683
rect 23340 35649 23348 35683
rect 23296 35640 23348 35649
rect 23388 35640 23440 35692
rect 23664 35640 23716 35692
rect 25872 35819 25924 35828
rect 25872 35785 25881 35819
rect 25881 35785 25915 35819
rect 25915 35785 25924 35819
rect 25872 35776 25924 35785
rect 25964 35776 26016 35828
rect 25596 35708 25648 35760
rect 24492 35683 24544 35692
rect 24492 35649 24501 35683
rect 24501 35649 24535 35683
rect 24535 35649 24544 35683
rect 24492 35640 24544 35649
rect 24676 35683 24728 35692
rect 24676 35649 24685 35683
rect 24685 35649 24719 35683
rect 24719 35649 24728 35683
rect 24676 35640 24728 35649
rect 23940 35572 23992 35624
rect 24584 35572 24636 35624
rect 25044 35640 25096 35692
rect 25136 35640 25188 35692
rect 13912 35504 13964 35556
rect 14832 35504 14884 35556
rect 26240 35640 26292 35692
rect 26332 35683 26384 35692
rect 26332 35649 26341 35683
rect 26341 35649 26375 35683
rect 26375 35649 26384 35683
rect 26332 35640 26384 35649
rect 27344 35776 27396 35828
rect 28724 35776 28776 35828
rect 31208 35776 31260 35828
rect 33600 35776 33652 35828
rect 26792 35640 26844 35692
rect 26884 35640 26936 35692
rect 27068 35683 27120 35692
rect 27068 35649 27077 35683
rect 27077 35649 27111 35683
rect 27111 35649 27120 35683
rect 27068 35640 27120 35649
rect 30656 35708 30708 35760
rect 27436 35683 27488 35692
rect 27436 35649 27445 35683
rect 27445 35649 27479 35683
rect 27479 35649 27488 35683
rect 27436 35640 27488 35649
rect 27528 35683 27580 35692
rect 27528 35649 27542 35683
rect 27542 35649 27576 35683
rect 27576 35649 27580 35683
rect 27528 35640 27580 35649
rect 28080 35683 28132 35692
rect 28080 35649 28089 35683
rect 28089 35649 28123 35683
rect 28123 35649 28132 35683
rect 28080 35640 28132 35649
rect 28448 35640 28500 35692
rect 29644 35683 29696 35692
rect 29644 35649 29651 35683
rect 29651 35649 29696 35683
rect 26240 35504 26292 35556
rect 26424 35504 26476 35556
rect 13360 35436 13412 35488
rect 15016 35436 15068 35488
rect 19064 35436 19116 35488
rect 19892 35479 19944 35488
rect 19892 35445 19901 35479
rect 19901 35445 19935 35479
rect 19935 35445 19944 35479
rect 19892 35436 19944 35445
rect 22744 35479 22796 35488
rect 22744 35445 22753 35479
rect 22753 35445 22787 35479
rect 22787 35445 22796 35479
rect 22744 35436 22796 35445
rect 27620 35436 27672 35488
rect 27896 35436 27948 35488
rect 28632 35572 28684 35624
rect 29644 35640 29696 35649
rect 29736 35683 29788 35692
rect 29736 35649 29745 35683
rect 29745 35649 29779 35683
rect 29779 35649 29788 35683
rect 29736 35640 29788 35649
rect 29828 35683 29880 35692
rect 29828 35649 29837 35683
rect 29837 35649 29871 35683
rect 29871 35649 29880 35683
rect 29828 35640 29880 35649
rect 30012 35640 30064 35692
rect 30748 35683 30800 35692
rect 30748 35649 30757 35683
rect 30757 35649 30791 35683
rect 30791 35649 30800 35683
rect 30748 35640 30800 35649
rect 33232 35708 33284 35760
rect 31116 35640 31168 35692
rect 32496 35683 32548 35692
rect 32496 35649 32505 35683
rect 32505 35649 32539 35683
rect 32539 35649 32548 35683
rect 32496 35640 32548 35649
rect 30288 35572 30340 35624
rect 30380 35572 30432 35624
rect 34612 35708 34664 35760
rect 33324 35683 33376 35692
rect 33324 35649 33333 35683
rect 33333 35649 33367 35683
rect 33367 35649 33376 35683
rect 33324 35640 33376 35649
rect 31484 35504 31536 35556
rect 29644 35436 29696 35488
rect 29920 35436 29972 35488
rect 30196 35436 30248 35488
rect 30840 35436 30892 35488
rect 32220 35436 32272 35488
rect 32312 35479 32364 35488
rect 32312 35445 32321 35479
rect 32321 35445 32355 35479
rect 32355 35445 32364 35479
rect 32312 35436 32364 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 6736 35275 6788 35284
rect 6736 35241 6745 35275
rect 6745 35241 6779 35275
rect 6779 35241 6788 35275
rect 6736 35232 6788 35241
rect 8024 35232 8076 35284
rect 9220 35232 9272 35284
rect 9864 35232 9916 35284
rect 10232 35232 10284 35284
rect 8668 35164 8720 35216
rect 9588 35164 9640 35216
rect 10324 35164 10376 35216
rect 9496 35096 9548 35148
rect 10508 35139 10560 35148
rect 10508 35105 10517 35139
rect 10517 35105 10551 35139
rect 10551 35105 10560 35139
rect 10508 35096 10560 35105
rect 8668 35071 8720 35080
rect 8668 35037 8677 35071
rect 8677 35037 8711 35071
rect 8711 35037 8720 35071
rect 8668 35028 8720 35037
rect 10232 35028 10284 35080
rect 13176 35232 13228 35284
rect 13268 35232 13320 35284
rect 12164 35164 12216 35216
rect 10876 35028 10928 35080
rect 11704 35096 11756 35148
rect 11796 35096 11848 35148
rect 9404 35003 9456 35012
rect 9404 34969 9413 35003
rect 9413 34969 9447 35003
rect 9447 34969 9456 35003
rect 9404 34960 9456 34969
rect 9588 34892 9640 34944
rect 10784 34960 10836 35012
rect 11520 35071 11572 35080
rect 11520 35037 11529 35071
rect 11529 35037 11563 35071
rect 11563 35037 11572 35071
rect 11520 35028 11572 35037
rect 11888 35071 11940 35080
rect 11888 35037 11897 35071
rect 11897 35037 11931 35071
rect 11931 35037 11940 35071
rect 11888 35028 11940 35037
rect 12072 35028 12124 35080
rect 14004 35096 14056 35148
rect 11060 34935 11112 34944
rect 11060 34901 11069 34935
rect 11069 34901 11103 34935
rect 11103 34901 11112 34935
rect 11060 34892 11112 34901
rect 11520 34892 11572 34944
rect 12624 35071 12676 35080
rect 12624 35037 12633 35071
rect 12633 35037 12667 35071
rect 12667 35037 12676 35071
rect 12624 35028 12676 35037
rect 13268 35028 13320 35080
rect 12808 34960 12860 35012
rect 13176 34960 13228 35012
rect 13912 35028 13964 35080
rect 14096 35071 14148 35080
rect 14096 35037 14105 35071
rect 14105 35037 14139 35071
rect 14139 35037 14148 35071
rect 14096 35028 14148 35037
rect 14280 35028 14332 35080
rect 14832 35028 14884 35080
rect 15016 35071 15068 35080
rect 15016 35037 15025 35071
rect 15025 35037 15059 35071
rect 15059 35037 15068 35071
rect 15016 35028 15068 35037
rect 15936 35207 15988 35216
rect 15936 35173 15945 35207
rect 15945 35173 15979 35207
rect 15979 35173 15988 35207
rect 15936 35164 15988 35173
rect 15384 35071 15436 35080
rect 15384 35037 15393 35071
rect 15393 35037 15427 35071
rect 15427 35037 15436 35071
rect 15384 35028 15436 35037
rect 22744 35232 22796 35284
rect 22928 35232 22980 35284
rect 23940 35232 23992 35284
rect 16488 35164 16540 35216
rect 16672 35164 16724 35216
rect 17592 35096 17644 35148
rect 18144 35164 18196 35216
rect 13636 35003 13688 35012
rect 13636 34969 13645 35003
rect 13645 34969 13679 35003
rect 13679 34969 13688 35003
rect 13636 34960 13688 34969
rect 13728 34960 13780 35012
rect 12072 34892 12124 34944
rect 14096 34892 14148 34944
rect 14556 34935 14608 34944
rect 14556 34901 14565 34935
rect 14565 34901 14599 34935
rect 14599 34901 14608 34935
rect 14556 34892 14608 34901
rect 15752 34892 15804 34944
rect 17040 35028 17092 35080
rect 20260 35028 20312 35080
rect 16028 34960 16080 35012
rect 21456 34960 21508 35012
rect 16764 34935 16816 34944
rect 16764 34901 16773 34935
rect 16773 34901 16807 34935
rect 16807 34901 16816 34935
rect 16764 34892 16816 34901
rect 18512 34892 18564 34944
rect 20904 34892 20956 34944
rect 24584 35164 24636 35216
rect 26792 35232 26844 35284
rect 27712 35232 27764 35284
rect 28816 35232 28868 35284
rect 29000 35232 29052 35284
rect 30380 35232 30432 35284
rect 26700 35164 26752 35216
rect 27620 35164 27672 35216
rect 28908 35164 28960 35216
rect 23204 35028 23256 35080
rect 24492 35028 24544 35080
rect 26884 35096 26936 35148
rect 27804 35139 27856 35148
rect 27804 35105 27813 35139
rect 27813 35105 27847 35139
rect 27847 35105 27856 35139
rect 27804 35096 27856 35105
rect 28356 35096 28408 35148
rect 25044 35028 25096 35080
rect 25412 35071 25464 35080
rect 25412 35037 25421 35071
rect 25421 35037 25455 35071
rect 25455 35037 25464 35071
rect 25412 35028 25464 35037
rect 25596 35071 25648 35080
rect 25596 35037 25605 35071
rect 25605 35037 25639 35071
rect 25639 35037 25648 35071
rect 25596 35028 25648 35037
rect 25872 35028 25924 35080
rect 26240 35028 26292 35080
rect 27528 35028 27580 35080
rect 22560 35003 22612 35012
rect 22560 34969 22569 35003
rect 22569 34969 22603 35003
rect 22603 34969 22612 35003
rect 22560 34960 22612 34969
rect 28816 35071 28868 35080
rect 28816 35037 28825 35071
rect 28825 35037 28859 35071
rect 28859 35037 28868 35071
rect 28816 35028 28868 35037
rect 29276 35071 29328 35080
rect 29276 35037 29285 35071
rect 29285 35037 29319 35071
rect 29319 35037 29328 35071
rect 29276 35028 29328 35037
rect 29368 35028 29420 35080
rect 29644 35028 29696 35080
rect 30472 35164 30524 35216
rect 31116 35232 31168 35284
rect 30932 35164 30984 35216
rect 31576 35164 31628 35216
rect 32312 35232 32364 35284
rect 30380 35071 30432 35080
rect 30380 35037 30396 35071
rect 30396 35037 30430 35071
rect 30430 35037 30432 35071
rect 30380 35028 30432 35037
rect 23296 34892 23348 34944
rect 24952 34892 25004 34944
rect 25044 34892 25096 34944
rect 27988 34960 28040 35012
rect 28356 34960 28408 35012
rect 28724 34960 28776 35012
rect 25596 34892 25648 34944
rect 28816 34892 28868 34944
rect 29092 34892 29144 34944
rect 30196 34892 30248 34944
rect 30380 34892 30432 34944
rect 30472 34892 30524 34944
rect 31116 35028 31168 35080
rect 31392 35096 31444 35148
rect 31300 35071 31352 35080
rect 31300 35037 31310 35071
rect 31310 35037 31344 35071
rect 31344 35037 31352 35071
rect 31300 35028 31352 35037
rect 31852 35028 31904 35080
rect 33324 35096 33376 35148
rect 34520 35096 34572 35148
rect 34888 35096 34940 35148
rect 32036 35028 32088 35080
rect 34612 35028 34664 35080
rect 34796 35071 34848 35080
rect 34796 35037 34805 35071
rect 34805 35037 34839 35071
rect 34839 35037 34848 35071
rect 34796 35028 34848 35037
rect 31576 35003 31628 35012
rect 31576 34969 31582 35003
rect 31582 34969 31616 35003
rect 31616 34969 31628 35003
rect 31576 34960 31628 34969
rect 30840 34892 30892 34944
rect 32036 34935 32088 34944
rect 32036 34901 32045 34935
rect 32045 34901 32079 34935
rect 32079 34901 32088 34935
rect 32036 34892 32088 34901
rect 32404 34892 32456 34944
rect 34612 34892 34664 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 9404 34688 9456 34740
rect 5540 34620 5592 34672
rect 6828 34620 6880 34672
rect 9220 34620 9272 34672
rect 11796 34620 11848 34672
rect 13176 34620 13228 34672
rect 6000 34484 6052 34536
rect 9312 34484 9364 34536
rect 10140 34552 10192 34604
rect 11888 34552 11940 34604
rect 12716 34552 12768 34604
rect 13360 34595 13412 34604
rect 11428 34484 11480 34536
rect 13360 34561 13369 34595
rect 13369 34561 13403 34595
rect 13403 34561 13412 34595
rect 13360 34552 13412 34561
rect 9036 34348 9088 34400
rect 10048 34416 10100 34468
rect 13728 34595 13780 34604
rect 13728 34561 13737 34595
rect 13737 34561 13771 34595
rect 13771 34561 13780 34595
rect 13728 34552 13780 34561
rect 14004 34688 14056 34740
rect 14096 34484 14148 34536
rect 14188 34416 14240 34468
rect 9404 34348 9456 34400
rect 9680 34348 9732 34400
rect 12624 34348 12676 34400
rect 13452 34348 13504 34400
rect 17776 34688 17828 34740
rect 16028 34620 16080 34672
rect 19156 34688 19208 34740
rect 21456 34731 21508 34740
rect 21456 34697 21465 34731
rect 21465 34697 21499 34731
rect 21499 34697 21508 34731
rect 21456 34688 21508 34697
rect 22376 34688 22428 34740
rect 26056 34731 26108 34740
rect 26056 34697 26065 34731
rect 26065 34697 26099 34731
rect 26099 34697 26108 34731
rect 26056 34688 26108 34697
rect 26884 34688 26936 34740
rect 14464 34484 14516 34536
rect 14832 34484 14884 34536
rect 16764 34552 16816 34604
rect 17132 34552 17184 34604
rect 17224 34595 17276 34604
rect 17224 34561 17233 34595
rect 17233 34561 17267 34595
rect 17267 34561 17276 34595
rect 17224 34552 17276 34561
rect 17592 34595 17644 34604
rect 17592 34561 17602 34595
rect 17602 34561 17636 34595
rect 17636 34561 17644 34595
rect 17592 34552 17644 34561
rect 17684 34484 17736 34536
rect 17868 34595 17920 34604
rect 17868 34561 17877 34595
rect 17877 34561 17911 34595
rect 17911 34561 17920 34595
rect 17868 34552 17920 34561
rect 18052 34552 18104 34604
rect 18512 34595 18564 34604
rect 18512 34561 18521 34595
rect 18521 34561 18555 34595
rect 18555 34561 18564 34595
rect 18512 34552 18564 34561
rect 18604 34595 18656 34604
rect 18604 34561 18613 34595
rect 18613 34561 18647 34595
rect 18647 34561 18656 34595
rect 18604 34552 18656 34561
rect 22560 34620 22612 34672
rect 21640 34552 21692 34604
rect 22100 34552 22152 34604
rect 22652 34552 22704 34604
rect 26056 34552 26108 34604
rect 15200 34416 15252 34468
rect 20812 34484 20864 34536
rect 25228 34484 25280 34536
rect 25596 34484 25648 34536
rect 28264 34688 28316 34740
rect 29920 34688 29972 34740
rect 27620 34663 27672 34672
rect 27620 34629 27629 34663
rect 27629 34629 27663 34663
rect 27663 34629 27672 34663
rect 27620 34620 27672 34629
rect 27712 34595 27764 34604
rect 27712 34561 27721 34595
rect 27721 34561 27755 34595
rect 27755 34561 27764 34595
rect 27712 34552 27764 34561
rect 28448 34552 28500 34604
rect 29092 34552 29144 34604
rect 29368 34552 29420 34604
rect 27068 34484 27120 34536
rect 29920 34552 29972 34604
rect 30288 34688 30340 34740
rect 30656 34688 30708 34740
rect 30840 34731 30892 34740
rect 30840 34697 30849 34731
rect 30849 34697 30883 34731
rect 30883 34697 30892 34731
rect 30840 34688 30892 34697
rect 31300 34688 31352 34740
rect 30748 34620 30800 34672
rect 30288 34595 30340 34604
rect 30288 34561 30297 34595
rect 30297 34561 30331 34595
rect 30331 34561 30340 34595
rect 30288 34552 30340 34561
rect 31852 34620 31904 34672
rect 32220 34663 32272 34672
rect 32220 34629 32229 34663
rect 32229 34629 32263 34663
rect 32263 34629 32272 34663
rect 32220 34620 32272 34629
rect 18144 34459 18196 34468
rect 18144 34425 18153 34459
rect 18153 34425 18187 34459
rect 18187 34425 18196 34459
rect 18144 34416 18196 34425
rect 21916 34416 21968 34468
rect 22284 34459 22336 34468
rect 22284 34425 22293 34459
rect 22293 34425 22327 34459
rect 22327 34425 22336 34459
rect 22284 34416 22336 34425
rect 24216 34416 24268 34468
rect 26240 34416 26292 34468
rect 29736 34484 29788 34536
rect 32036 34552 32088 34604
rect 32312 34552 32364 34604
rect 34520 34552 34572 34604
rect 34612 34552 34664 34604
rect 34704 34595 34756 34604
rect 34704 34561 34713 34595
rect 34713 34561 34747 34595
rect 34747 34561 34756 34595
rect 34704 34552 34756 34561
rect 34796 34552 34848 34604
rect 34888 34595 34940 34604
rect 34888 34561 34897 34595
rect 34897 34561 34931 34595
rect 34931 34561 34940 34595
rect 34888 34552 34940 34561
rect 31208 34416 31260 34468
rect 35532 34595 35584 34604
rect 35532 34561 35541 34595
rect 35541 34561 35575 34595
rect 35575 34561 35584 34595
rect 35532 34552 35584 34561
rect 14556 34391 14608 34400
rect 14556 34357 14565 34391
rect 14565 34357 14599 34391
rect 14599 34357 14608 34391
rect 14556 34348 14608 34357
rect 14648 34348 14700 34400
rect 16672 34391 16724 34400
rect 16672 34357 16681 34391
rect 16681 34357 16715 34391
rect 16715 34357 16724 34391
rect 16672 34348 16724 34357
rect 17040 34348 17092 34400
rect 17960 34348 18012 34400
rect 18972 34391 19024 34400
rect 18972 34357 18981 34391
rect 18981 34357 19015 34391
rect 19015 34357 19024 34391
rect 18972 34348 19024 34357
rect 19524 34348 19576 34400
rect 20076 34348 20128 34400
rect 21180 34348 21232 34400
rect 26332 34348 26384 34400
rect 26424 34348 26476 34400
rect 34428 34348 34480 34400
rect 34612 34416 34664 34468
rect 34704 34348 34756 34400
rect 35348 34391 35400 34400
rect 35348 34357 35357 34391
rect 35357 34357 35391 34391
rect 35391 34357 35400 34391
rect 35348 34348 35400 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 9680 34144 9732 34196
rect 7932 34119 7984 34128
rect 7932 34085 7941 34119
rect 7941 34085 7975 34119
rect 7975 34085 7984 34119
rect 7932 34076 7984 34085
rect 8760 34076 8812 34128
rect 9404 34076 9456 34128
rect 10232 34076 10284 34128
rect 10784 34076 10836 34128
rect 11152 34119 11204 34128
rect 11152 34085 11161 34119
rect 11161 34085 11195 34119
rect 11195 34085 11204 34119
rect 11152 34076 11204 34085
rect 9956 34008 10008 34060
rect 12072 34076 12124 34128
rect 11888 34008 11940 34060
rect 8208 33872 8260 33924
rect 9864 33983 9916 33992
rect 9864 33949 9878 33983
rect 9878 33949 9912 33983
rect 9912 33949 9916 33983
rect 9864 33940 9916 33949
rect 10508 33940 10560 33992
rect 10876 33940 10928 33992
rect 11612 33940 11664 33992
rect 12348 34076 12400 34128
rect 14096 34144 14148 34196
rect 14740 34144 14792 34196
rect 17040 34187 17092 34196
rect 17040 34153 17049 34187
rect 17049 34153 17083 34187
rect 17083 34153 17092 34187
rect 17040 34144 17092 34153
rect 18604 34144 18656 34196
rect 12992 33940 13044 33992
rect 10324 33872 10376 33924
rect 8024 33847 8076 33856
rect 8024 33813 8033 33847
rect 8033 33813 8067 33847
rect 8067 33813 8076 33847
rect 8024 33804 8076 33813
rect 9496 33804 9548 33856
rect 9956 33804 10008 33856
rect 11060 33804 11112 33856
rect 11888 33872 11940 33924
rect 15476 33940 15528 33992
rect 18972 34008 19024 34060
rect 17040 33940 17092 33992
rect 13820 33872 13872 33924
rect 14188 33872 14240 33924
rect 14372 33872 14424 33924
rect 12072 33847 12124 33856
rect 12072 33813 12081 33847
rect 12081 33813 12115 33847
rect 12115 33813 12124 33847
rect 12072 33804 12124 33813
rect 12716 33804 12768 33856
rect 13636 33804 13688 33856
rect 14004 33804 14056 33856
rect 15752 33872 15804 33924
rect 16120 33872 16172 33924
rect 16212 33872 16264 33924
rect 16764 33872 16816 33924
rect 16580 33804 16632 33856
rect 19432 34008 19484 34060
rect 19248 33983 19300 33992
rect 19248 33949 19257 33983
rect 19257 33949 19291 33983
rect 19291 33949 19300 33983
rect 19248 33940 19300 33949
rect 21640 34144 21692 34196
rect 22928 34187 22980 34196
rect 22928 34153 22937 34187
rect 22937 34153 22971 34187
rect 22971 34153 22980 34187
rect 22928 34144 22980 34153
rect 23388 34144 23440 34196
rect 24308 34144 24360 34196
rect 25044 34144 25096 34196
rect 25136 34144 25188 34196
rect 19616 33983 19668 33992
rect 19616 33949 19625 33983
rect 19625 33949 19659 33983
rect 19659 33949 19668 33983
rect 19616 33940 19668 33949
rect 20720 34008 20772 34060
rect 21456 34076 21508 34128
rect 20168 33983 20220 33992
rect 20168 33949 20178 33983
rect 20178 33949 20212 33983
rect 20212 33949 20220 33983
rect 20168 33940 20220 33949
rect 17040 33804 17092 33856
rect 17684 33847 17736 33856
rect 17684 33813 17693 33847
rect 17693 33813 17727 33847
rect 17727 33813 17736 33847
rect 17684 33804 17736 33813
rect 18512 33804 18564 33856
rect 18604 33804 18656 33856
rect 18696 33804 18748 33856
rect 19984 33804 20036 33856
rect 20168 33804 20220 33856
rect 20352 33915 20404 33924
rect 20352 33881 20361 33915
rect 20361 33881 20395 33915
rect 20395 33881 20404 33915
rect 20352 33872 20404 33881
rect 21180 33983 21232 33992
rect 21180 33949 21189 33983
rect 21189 33949 21223 33983
rect 21223 33949 21232 33983
rect 21180 33940 21232 33949
rect 23296 34008 23348 34060
rect 22100 33940 22152 33992
rect 22284 33940 22336 33992
rect 22836 33940 22888 33992
rect 22652 33872 22704 33924
rect 23388 33940 23440 33992
rect 23572 34008 23624 34060
rect 23940 33872 23992 33924
rect 24124 33872 24176 33924
rect 20720 33847 20772 33856
rect 20720 33813 20729 33847
rect 20729 33813 20763 33847
rect 20763 33813 20772 33847
rect 20720 33804 20772 33813
rect 23020 33804 23072 33856
rect 28448 34076 28500 34128
rect 30656 34144 30708 34196
rect 31576 34144 31628 34196
rect 34244 34187 34296 34196
rect 34244 34153 34253 34187
rect 34253 34153 34287 34187
rect 34287 34153 34296 34187
rect 34244 34144 34296 34153
rect 34336 34144 34388 34196
rect 35348 34144 35400 34196
rect 25504 33940 25556 33992
rect 27620 34008 27672 34060
rect 30196 34008 30248 34060
rect 34520 34076 34572 34128
rect 35532 34008 35584 34060
rect 26332 33940 26384 33992
rect 28724 33940 28776 33992
rect 30104 33940 30156 33992
rect 26240 33872 26292 33924
rect 26700 33872 26752 33924
rect 27528 33872 27580 33924
rect 28264 33872 28316 33924
rect 31852 33872 31904 33924
rect 24584 33804 24636 33856
rect 27068 33804 27120 33856
rect 32312 33940 32364 33992
rect 34612 33940 34664 33992
rect 34704 33983 34756 33992
rect 34704 33949 34713 33983
rect 34713 33949 34747 33983
rect 34747 33949 34756 33983
rect 34704 33940 34756 33949
rect 34796 33940 34848 33992
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 8024 33600 8076 33652
rect 9588 33643 9640 33652
rect 9588 33609 9597 33643
rect 9597 33609 9631 33643
rect 9631 33609 9640 33643
rect 9588 33600 9640 33609
rect 11336 33600 11388 33652
rect 11888 33600 11940 33652
rect 12624 33600 12676 33652
rect 14372 33600 14424 33652
rect 7104 33532 7156 33584
rect 8208 33507 8260 33516
rect 8208 33473 8217 33507
rect 8217 33473 8251 33507
rect 8251 33473 8260 33507
rect 8208 33464 8260 33473
rect 9496 33464 9548 33516
rect 6000 33396 6052 33448
rect 6736 33439 6788 33448
rect 6736 33405 6745 33439
rect 6745 33405 6779 33439
rect 6779 33405 6788 33439
rect 6736 33396 6788 33405
rect 9220 33396 9272 33448
rect 9864 33464 9916 33516
rect 12072 33532 12124 33584
rect 16672 33600 16724 33652
rect 17684 33600 17736 33652
rect 18420 33600 18472 33652
rect 11520 33507 11572 33516
rect 11520 33473 11529 33507
rect 11529 33473 11563 33507
rect 11563 33473 11572 33507
rect 11520 33464 11572 33473
rect 11612 33507 11664 33516
rect 11612 33473 11621 33507
rect 11621 33473 11655 33507
rect 11655 33473 11664 33507
rect 11612 33464 11664 33473
rect 13912 33464 13964 33516
rect 14188 33464 14240 33516
rect 15016 33464 15068 33516
rect 11336 33396 11388 33448
rect 9864 33328 9916 33380
rect 12532 33396 12584 33448
rect 13544 33396 13596 33448
rect 9036 33260 9088 33312
rect 11060 33260 11112 33312
rect 14556 33328 14608 33380
rect 16396 33532 16448 33584
rect 19984 33600 20036 33652
rect 19064 33532 19116 33584
rect 19248 33532 19300 33584
rect 20168 33532 20220 33584
rect 17316 33464 17368 33516
rect 18696 33507 18748 33516
rect 18696 33473 18705 33507
rect 18705 33473 18739 33507
rect 18739 33473 18748 33507
rect 18696 33464 18748 33473
rect 21364 33600 21416 33652
rect 22744 33600 22796 33652
rect 23480 33643 23532 33652
rect 23480 33609 23489 33643
rect 23489 33609 23523 33643
rect 23523 33609 23532 33643
rect 23480 33600 23532 33609
rect 24032 33600 24084 33652
rect 20352 33532 20404 33584
rect 18512 33396 18564 33448
rect 20536 33464 20588 33516
rect 20720 33464 20772 33516
rect 20904 33507 20956 33516
rect 20904 33473 20913 33507
rect 20913 33473 20947 33507
rect 20947 33473 20956 33507
rect 20904 33464 20956 33473
rect 21088 33464 21140 33516
rect 21732 33532 21784 33584
rect 23020 33575 23072 33584
rect 23020 33541 23029 33575
rect 23029 33541 23063 33575
rect 23063 33541 23072 33575
rect 23020 33532 23072 33541
rect 23204 33532 23256 33584
rect 21548 33396 21600 33448
rect 22100 33464 22152 33516
rect 22284 33396 22336 33448
rect 22560 33507 22612 33516
rect 22560 33473 22569 33507
rect 22569 33473 22603 33507
rect 22603 33473 22612 33507
rect 22560 33464 22612 33473
rect 23112 33464 23164 33516
rect 24308 33575 24360 33584
rect 24308 33541 24317 33575
rect 24317 33541 24351 33575
rect 24351 33541 24360 33575
rect 24308 33532 24360 33541
rect 23388 33396 23440 33448
rect 23940 33464 23992 33516
rect 24216 33507 24268 33516
rect 24216 33473 24225 33507
rect 24225 33473 24259 33507
rect 24259 33473 24268 33507
rect 24216 33464 24268 33473
rect 21272 33328 21324 33380
rect 21640 33328 21692 33380
rect 11704 33303 11756 33312
rect 11704 33269 11713 33303
rect 11713 33269 11747 33303
rect 11747 33269 11756 33303
rect 11704 33260 11756 33269
rect 12348 33260 12400 33312
rect 14004 33303 14056 33312
rect 14004 33269 14013 33303
rect 14013 33269 14047 33303
rect 14047 33269 14056 33303
rect 14004 33260 14056 33269
rect 14372 33303 14424 33312
rect 14372 33269 14381 33303
rect 14381 33269 14415 33303
rect 14415 33269 14424 33303
rect 14372 33260 14424 33269
rect 15292 33260 15344 33312
rect 16212 33303 16264 33312
rect 16212 33269 16221 33303
rect 16221 33269 16255 33303
rect 16255 33269 16264 33303
rect 16212 33260 16264 33269
rect 16304 33260 16356 33312
rect 18512 33303 18564 33312
rect 18512 33269 18521 33303
rect 18521 33269 18555 33303
rect 18555 33269 18564 33303
rect 18512 33260 18564 33269
rect 18972 33260 19024 33312
rect 20812 33303 20864 33312
rect 20812 33269 20821 33303
rect 20821 33269 20855 33303
rect 20855 33269 20864 33303
rect 20812 33260 20864 33269
rect 21088 33303 21140 33312
rect 21088 33269 21097 33303
rect 21097 33269 21131 33303
rect 21131 33269 21140 33303
rect 21088 33260 21140 33269
rect 23020 33328 23072 33380
rect 23296 33371 23348 33380
rect 23296 33337 23305 33371
rect 23305 33337 23339 33371
rect 23339 33337 23348 33371
rect 23296 33328 23348 33337
rect 22928 33260 22980 33312
rect 23756 33328 23808 33380
rect 24400 33507 24452 33516
rect 24400 33473 24409 33507
rect 24409 33473 24443 33507
rect 24443 33473 24452 33507
rect 24400 33464 24452 33473
rect 24860 33464 24912 33516
rect 25136 33507 25188 33516
rect 25136 33473 25145 33507
rect 25145 33473 25179 33507
rect 25179 33473 25188 33507
rect 25136 33464 25188 33473
rect 25320 33507 25372 33516
rect 25320 33473 25329 33507
rect 25329 33473 25363 33507
rect 25363 33473 25372 33507
rect 25320 33464 25372 33473
rect 24584 33439 24636 33448
rect 24584 33405 24593 33439
rect 24593 33405 24627 33439
rect 24627 33405 24636 33439
rect 24584 33396 24636 33405
rect 23940 33328 23992 33380
rect 25596 33507 25648 33516
rect 25596 33473 25605 33507
rect 25605 33473 25639 33507
rect 25639 33473 25648 33507
rect 25596 33464 25648 33473
rect 25780 33464 25832 33516
rect 26240 33575 26292 33584
rect 26240 33541 26249 33575
rect 26249 33541 26283 33575
rect 26283 33541 26292 33575
rect 26240 33532 26292 33541
rect 26608 33600 26660 33652
rect 26792 33600 26844 33652
rect 27160 33600 27212 33652
rect 28172 33643 28224 33652
rect 28172 33609 28181 33643
rect 28181 33609 28215 33643
rect 28215 33609 28224 33643
rect 28172 33600 28224 33609
rect 26884 33532 26936 33584
rect 25688 33396 25740 33448
rect 25964 33464 26016 33516
rect 26424 33464 26476 33516
rect 27068 33507 27120 33516
rect 27068 33473 27077 33507
rect 27077 33473 27111 33507
rect 27111 33473 27120 33507
rect 27068 33464 27120 33473
rect 27160 33507 27212 33516
rect 27160 33473 27169 33507
rect 27169 33473 27203 33507
rect 27203 33473 27212 33507
rect 27160 33464 27212 33473
rect 27528 33464 27580 33516
rect 27988 33464 28040 33516
rect 28264 33507 28316 33516
rect 28264 33473 28273 33507
rect 28273 33473 28307 33507
rect 28307 33473 28316 33507
rect 28264 33464 28316 33473
rect 27804 33396 27856 33448
rect 24400 33260 24452 33312
rect 24492 33303 24544 33312
rect 24492 33269 24501 33303
rect 24501 33269 24535 33303
rect 24535 33269 24544 33303
rect 24492 33260 24544 33269
rect 24860 33303 24912 33312
rect 24860 33269 24869 33303
rect 24869 33269 24903 33303
rect 24903 33269 24912 33303
rect 24860 33260 24912 33269
rect 24952 33303 25004 33312
rect 24952 33269 24961 33303
rect 24961 33269 24995 33303
rect 24995 33269 25004 33303
rect 24952 33260 25004 33269
rect 25320 33260 25372 33312
rect 27160 33328 27212 33380
rect 28540 33464 28592 33516
rect 28908 33507 28960 33516
rect 28908 33473 28917 33507
rect 28917 33473 28951 33507
rect 28951 33473 28960 33507
rect 28908 33464 28960 33473
rect 30012 33464 30064 33516
rect 30288 33464 30340 33516
rect 31484 33464 31536 33516
rect 31852 33532 31904 33584
rect 33416 33532 33468 33584
rect 35348 33532 35400 33584
rect 34244 33464 34296 33516
rect 34612 33507 34664 33516
rect 34612 33473 34621 33507
rect 34621 33473 34655 33507
rect 34655 33473 34664 33507
rect 34612 33464 34664 33473
rect 35532 33464 35584 33516
rect 30656 33396 30708 33448
rect 31576 33439 31628 33448
rect 31576 33405 31585 33439
rect 31585 33405 31619 33439
rect 31619 33405 31628 33439
rect 31576 33396 31628 33405
rect 29276 33328 29328 33380
rect 25780 33303 25832 33312
rect 25780 33269 25789 33303
rect 25789 33269 25823 33303
rect 25823 33269 25832 33303
rect 25780 33260 25832 33269
rect 26608 33260 26660 33312
rect 27436 33303 27488 33312
rect 27436 33269 27445 33303
rect 27445 33269 27479 33303
rect 27479 33269 27488 33303
rect 27436 33260 27488 33269
rect 28632 33260 28684 33312
rect 29552 33303 29604 33312
rect 29552 33269 29561 33303
rect 29561 33269 29595 33303
rect 29595 33269 29604 33303
rect 29552 33260 29604 33269
rect 34796 33260 34848 33312
rect 35624 33303 35676 33312
rect 35624 33269 35633 33303
rect 35633 33269 35667 33303
rect 35667 33269 35676 33303
rect 35624 33260 35676 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 6736 33056 6788 33108
rect 8300 33056 8352 33108
rect 13544 33056 13596 33108
rect 13636 33099 13688 33108
rect 13636 33065 13645 33099
rect 13645 33065 13679 33099
rect 13679 33065 13688 33099
rect 13636 33056 13688 33065
rect 13912 33056 13964 33108
rect 14096 33056 14148 33108
rect 15476 33056 15528 33108
rect 17408 33056 17460 33108
rect 17868 33056 17920 33108
rect 18236 33056 18288 33108
rect 18512 33056 18564 33108
rect 21180 33056 21232 33108
rect 7656 32920 7708 32972
rect 5908 32852 5960 32904
rect 6092 32895 6144 32904
rect 6092 32861 6101 32895
rect 6101 32861 6135 32895
rect 6135 32861 6144 32895
rect 6092 32852 6144 32861
rect 6276 32895 6328 32904
rect 6276 32861 6285 32895
rect 6285 32861 6319 32895
rect 6319 32861 6328 32895
rect 8484 32920 8536 32972
rect 8760 32920 8812 32972
rect 15384 32988 15436 33040
rect 20260 32988 20312 33040
rect 21640 33056 21692 33108
rect 22928 33056 22980 33108
rect 23664 33056 23716 33108
rect 24584 32988 24636 33040
rect 6276 32852 6328 32861
rect 8392 32895 8444 32904
rect 8392 32861 8401 32895
rect 8401 32861 8435 32895
rect 8435 32861 8444 32895
rect 8392 32852 8444 32861
rect 11428 32895 11480 32904
rect 11428 32861 11437 32895
rect 11437 32861 11471 32895
rect 11471 32861 11480 32895
rect 11428 32852 11480 32861
rect 6460 32784 6512 32836
rect 7840 32827 7892 32836
rect 7840 32793 7849 32827
rect 7849 32793 7883 32827
rect 7883 32793 7892 32827
rect 7840 32784 7892 32793
rect 8208 32784 8260 32836
rect 8024 32716 8076 32768
rect 8576 32784 8628 32836
rect 8852 32784 8904 32836
rect 12900 32784 12952 32836
rect 13636 32852 13688 32904
rect 14372 32895 14424 32904
rect 14372 32861 14381 32895
rect 14381 32861 14415 32895
rect 14415 32861 14424 32895
rect 14372 32852 14424 32861
rect 14556 32895 14608 32904
rect 14556 32861 14570 32895
rect 14570 32861 14604 32895
rect 14604 32861 14608 32895
rect 14556 32852 14608 32861
rect 15200 32852 15252 32904
rect 16028 32895 16080 32904
rect 16028 32861 16037 32895
rect 16037 32861 16071 32895
rect 16071 32861 16080 32895
rect 16028 32852 16080 32861
rect 16120 32895 16172 32904
rect 16120 32861 16129 32895
rect 16129 32861 16163 32895
rect 16163 32861 16172 32895
rect 16120 32852 16172 32861
rect 16212 32852 16264 32904
rect 8944 32716 8996 32768
rect 10048 32716 10100 32768
rect 11796 32716 11848 32768
rect 12164 32716 12216 32768
rect 12440 32716 12492 32768
rect 14924 32784 14976 32836
rect 15936 32784 15988 32836
rect 17040 32852 17092 32904
rect 17684 32852 17736 32904
rect 18420 32895 18472 32904
rect 18420 32861 18429 32895
rect 18429 32861 18463 32895
rect 18463 32861 18472 32895
rect 18420 32852 18472 32861
rect 18972 32852 19024 32904
rect 19524 32852 19576 32904
rect 13360 32716 13412 32768
rect 13820 32716 13872 32768
rect 14372 32716 14424 32768
rect 15660 32716 15712 32768
rect 16028 32716 16080 32768
rect 16948 32716 17000 32768
rect 17868 32716 17920 32768
rect 18696 32784 18748 32836
rect 20720 32784 20772 32836
rect 21456 32895 21508 32904
rect 21456 32861 21465 32895
rect 21465 32861 21499 32895
rect 21499 32861 21508 32895
rect 21456 32852 21508 32861
rect 21732 32852 21784 32904
rect 22008 32852 22060 32904
rect 22560 32852 22612 32904
rect 24308 32852 24360 32904
rect 21732 32759 21784 32768
rect 21732 32725 21741 32759
rect 21741 32725 21775 32759
rect 21775 32725 21784 32759
rect 21732 32716 21784 32725
rect 22836 32716 22888 32768
rect 24584 32852 24636 32904
rect 27528 33056 27580 33108
rect 28172 33056 28224 33108
rect 28540 33056 28592 33108
rect 30196 33056 30248 33108
rect 30380 33056 30432 33108
rect 31208 33056 31260 33108
rect 24952 32852 25004 32904
rect 25044 32852 25096 32904
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 27712 32988 27764 33040
rect 27252 32963 27304 32972
rect 27252 32929 27261 32963
rect 27261 32929 27295 32963
rect 27295 32929 27304 32963
rect 27252 32920 27304 32929
rect 27344 32920 27396 32972
rect 26056 32852 26108 32904
rect 26240 32852 26292 32904
rect 27620 32920 27672 32972
rect 30012 32988 30064 33040
rect 34612 33056 34664 33108
rect 35624 33056 35676 33108
rect 28172 32920 28224 32972
rect 29368 32852 29420 32904
rect 30104 32920 30156 32972
rect 34060 32963 34112 32972
rect 34060 32929 34069 32963
rect 34069 32929 34103 32963
rect 34103 32929 34112 32963
rect 34060 32920 34112 32929
rect 34520 32920 34572 32972
rect 34796 32963 34848 32972
rect 34796 32929 34805 32963
rect 34805 32929 34839 32963
rect 34839 32929 34848 32963
rect 34796 32920 34848 32929
rect 30196 32895 30248 32904
rect 30196 32861 30205 32895
rect 30205 32861 30239 32895
rect 30239 32861 30248 32895
rect 30196 32852 30248 32861
rect 31392 32852 31444 32904
rect 30380 32784 30432 32836
rect 30840 32784 30892 32836
rect 30932 32827 30984 32836
rect 30932 32793 30941 32827
rect 30941 32793 30975 32827
rect 30975 32793 30984 32827
rect 30932 32784 30984 32793
rect 31852 32852 31904 32904
rect 32404 32852 32456 32904
rect 34336 32852 34388 32904
rect 34888 32895 34940 32904
rect 25596 32716 25648 32768
rect 25964 32716 26016 32768
rect 27160 32716 27212 32768
rect 29000 32716 29052 32768
rect 29828 32716 29880 32768
rect 30104 32716 30156 32768
rect 30196 32716 30248 32768
rect 32864 32827 32916 32836
rect 32864 32793 32873 32827
rect 32873 32793 32907 32827
rect 32907 32793 32916 32827
rect 32864 32784 32916 32793
rect 32956 32784 33008 32836
rect 33784 32784 33836 32836
rect 34888 32861 34897 32895
rect 34897 32861 34931 32895
rect 34931 32861 34940 32895
rect 34888 32852 34940 32861
rect 34704 32784 34756 32836
rect 39120 32852 39172 32904
rect 34980 32716 35032 32768
rect 40960 32759 41012 32768
rect 40960 32725 40969 32759
rect 40969 32725 41003 32759
rect 41003 32725 41012 32759
rect 40960 32716 41012 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 5632 32512 5684 32564
rect 6276 32512 6328 32564
rect 6460 32555 6512 32564
rect 6460 32521 6469 32555
rect 6469 32521 6503 32555
rect 6503 32521 6512 32555
rect 6460 32512 6512 32521
rect 7104 32444 7156 32496
rect 6368 32419 6420 32428
rect 6368 32385 6377 32419
rect 6377 32385 6411 32419
rect 6411 32385 6420 32419
rect 6368 32376 6420 32385
rect 8484 32512 8536 32564
rect 8668 32512 8720 32564
rect 9312 32512 9364 32564
rect 10600 32512 10652 32564
rect 940 32172 992 32224
rect 6184 32308 6236 32360
rect 8208 32376 8260 32428
rect 8576 32419 8628 32428
rect 8576 32385 8585 32419
rect 8585 32385 8619 32419
rect 8619 32385 8628 32419
rect 8576 32376 8628 32385
rect 9036 32351 9088 32360
rect 9036 32317 9045 32351
rect 9045 32317 9079 32351
rect 9079 32317 9088 32351
rect 9036 32308 9088 32317
rect 8576 32240 8628 32292
rect 9128 32240 9180 32292
rect 10140 32308 10192 32360
rect 10600 32308 10652 32360
rect 10876 32376 10928 32428
rect 11060 32419 11112 32428
rect 11060 32385 11069 32419
rect 11069 32385 11103 32419
rect 11103 32385 11112 32419
rect 11060 32376 11112 32385
rect 11612 32376 11664 32428
rect 11888 32419 11940 32428
rect 11888 32385 11897 32419
rect 11897 32385 11931 32419
rect 11931 32385 11940 32419
rect 11888 32376 11940 32385
rect 12164 32376 12216 32428
rect 11152 32308 11204 32360
rect 12532 32512 12584 32564
rect 12900 32512 12952 32564
rect 12532 32419 12584 32428
rect 12532 32385 12541 32419
rect 12541 32385 12575 32419
rect 12575 32385 12584 32419
rect 12532 32376 12584 32385
rect 12900 32419 12952 32428
rect 12900 32385 12909 32419
rect 12909 32385 12943 32419
rect 12943 32385 12952 32419
rect 12900 32376 12952 32385
rect 13544 32444 13596 32496
rect 9312 32240 9364 32292
rect 9496 32283 9548 32292
rect 9496 32249 9505 32283
rect 9505 32249 9539 32283
rect 9539 32249 9548 32283
rect 9496 32240 9548 32249
rect 11888 32240 11940 32292
rect 13176 32240 13228 32292
rect 13820 32419 13872 32428
rect 13820 32385 13830 32419
rect 13830 32385 13864 32419
rect 13864 32385 13872 32419
rect 14556 32444 14608 32496
rect 15936 32512 15988 32564
rect 16396 32512 16448 32564
rect 17316 32555 17368 32564
rect 17316 32521 17325 32555
rect 17325 32521 17359 32555
rect 17359 32521 17368 32555
rect 17316 32512 17368 32521
rect 17960 32512 18012 32564
rect 13820 32376 13872 32385
rect 14188 32419 14240 32428
rect 14188 32385 14202 32419
rect 14202 32385 14236 32419
rect 14236 32385 14240 32419
rect 14188 32376 14240 32385
rect 13544 32308 13596 32360
rect 13820 32240 13872 32292
rect 14096 32240 14148 32292
rect 14832 32351 14884 32360
rect 14832 32317 14841 32351
rect 14841 32317 14875 32351
rect 14875 32317 14884 32351
rect 14832 32308 14884 32317
rect 15384 32376 15436 32428
rect 15568 32419 15620 32428
rect 15568 32385 15577 32419
rect 15577 32385 15611 32419
rect 15611 32385 15620 32419
rect 15568 32376 15620 32385
rect 16028 32376 16080 32428
rect 4620 32172 4672 32224
rect 6000 32172 6052 32224
rect 8116 32172 8168 32224
rect 8484 32172 8536 32224
rect 10416 32172 10468 32224
rect 10784 32172 10836 32224
rect 11060 32172 11112 32224
rect 11520 32215 11572 32224
rect 11520 32181 11529 32215
rect 11529 32181 11563 32215
rect 11563 32181 11572 32215
rect 11520 32172 11572 32181
rect 12256 32215 12308 32224
rect 12256 32181 12265 32215
rect 12265 32181 12299 32215
rect 12299 32181 12308 32215
rect 12256 32172 12308 32181
rect 15200 32215 15252 32224
rect 15200 32181 15209 32215
rect 15209 32181 15243 32215
rect 15243 32181 15252 32215
rect 15200 32172 15252 32181
rect 15292 32172 15344 32224
rect 15936 32215 15988 32224
rect 15936 32181 15945 32215
rect 15945 32181 15979 32215
rect 15979 32181 15988 32215
rect 15936 32172 15988 32181
rect 16120 32240 16172 32292
rect 16304 32376 16356 32428
rect 16396 32419 16448 32428
rect 16396 32385 16405 32419
rect 16405 32385 16439 32419
rect 16439 32385 16448 32419
rect 16396 32376 16448 32385
rect 16856 32376 16908 32428
rect 16672 32172 16724 32224
rect 17500 32351 17552 32360
rect 17500 32317 17509 32351
rect 17509 32317 17543 32351
rect 17543 32317 17552 32351
rect 17500 32308 17552 32317
rect 17592 32308 17644 32360
rect 17868 32419 17920 32428
rect 17868 32385 17877 32419
rect 17877 32385 17911 32419
rect 17911 32385 17920 32419
rect 17868 32376 17920 32385
rect 18144 32487 18196 32496
rect 18144 32453 18153 32487
rect 18153 32453 18187 32487
rect 18187 32453 18196 32487
rect 18144 32444 18196 32453
rect 18420 32444 18472 32496
rect 18604 32376 18656 32428
rect 18696 32308 18748 32360
rect 19248 32512 19300 32564
rect 22008 32512 22060 32564
rect 22100 32512 22152 32564
rect 23020 32512 23072 32564
rect 24216 32512 24268 32564
rect 19432 32376 19484 32428
rect 21548 32444 21600 32496
rect 19616 32351 19668 32360
rect 19616 32317 19625 32351
rect 19625 32317 19659 32351
rect 19659 32317 19668 32351
rect 19616 32308 19668 32317
rect 21180 32376 21232 32428
rect 21640 32376 21692 32428
rect 23572 32444 23624 32496
rect 19892 32240 19944 32292
rect 21272 32308 21324 32360
rect 25136 32444 25188 32496
rect 25412 32444 25464 32496
rect 25964 32444 26016 32496
rect 27344 32555 27396 32564
rect 27344 32521 27353 32555
rect 27353 32521 27387 32555
rect 27387 32521 27396 32555
rect 27344 32512 27396 32521
rect 28816 32512 28868 32564
rect 29092 32512 29144 32564
rect 29552 32512 29604 32564
rect 30288 32512 30340 32564
rect 27068 32444 27120 32496
rect 31208 32512 31260 32564
rect 32404 32512 32456 32564
rect 32864 32512 32916 32564
rect 34336 32512 34388 32564
rect 34888 32512 34940 32564
rect 24216 32376 24268 32428
rect 24768 32376 24820 32428
rect 20536 32240 20588 32292
rect 22100 32240 22152 32292
rect 24952 32308 25004 32360
rect 26424 32376 26476 32428
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 27712 32419 27764 32428
rect 27712 32385 27721 32419
rect 27721 32385 27755 32419
rect 27755 32385 27764 32419
rect 27712 32376 27764 32385
rect 27988 32376 28040 32428
rect 28908 32376 28960 32428
rect 30840 32444 30892 32496
rect 29092 32376 29144 32428
rect 30104 32419 30156 32428
rect 30104 32385 30113 32419
rect 30113 32385 30147 32419
rect 30147 32385 30156 32419
rect 30104 32376 30156 32385
rect 30932 32376 30984 32428
rect 31576 32376 31628 32428
rect 32680 32419 32732 32428
rect 32680 32385 32689 32419
rect 32689 32385 32723 32419
rect 32723 32385 32732 32419
rect 32680 32376 32732 32385
rect 33784 32419 33836 32428
rect 33784 32385 33793 32419
rect 33793 32385 33827 32419
rect 33827 32385 33836 32419
rect 33784 32376 33836 32385
rect 28540 32308 28592 32360
rect 28632 32308 28684 32360
rect 30196 32308 30248 32360
rect 18696 32172 18748 32224
rect 19708 32172 19760 32224
rect 20904 32172 20956 32224
rect 21916 32215 21968 32224
rect 21916 32181 21925 32215
rect 21925 32181 21959 32215
rect 21959 32181 21968 32215
rect 21916 32172 21968 32181
rect 22284 32215 22336 32224
rect 22284 32181 22293 32215
rect 22293 32181 22327 32215
rect 22327 32181 22336 32215
rect 22284 32172 22336 32181
rect 22836 32172 22888 32224
rect 23204 32172 23256 32224
rect 24308 32240 24360 32292
rect 25044 32240 25096 32292
rect 27436 32240 27488 32292
rect 31116 32308 31168 32360
rect 32864 32351 32916 32360
rect 32864 32317 32873 32351
rect 32873 32317 32907 32351
rect 32907 32317 32916 32351
rect 32864 32308 32916 32317
rect 34428 32376 34480 32428
rect 34520 32376 34572 32428
rect 34980 32419 35032 32428
rect 34980 32385 34989 32419
rect 34989 32385 35023 32419
rect 35023 32385 35032 32419
rect 34980 32376 35032 32385
rect 37280 32444 37332 32496
rect 37648 32444 37700 32496
rect 38108 32487 38160 32496
rect 38108 32453 38117 32487
rect 38117 32453 38151 32487
rect 38151 32453 38160 32487
rect 38108 32444 38160 32453
rect 30656 32283 30708 32292
rect 30656 32249 30665 32283
rect 30665 32249 30699 32283
rect 30699 32249 30708 32283
rect 30656 32240 30708 32249
rect 25320 32172 25372 32224
rect 26056 32172 26108 32224
rect 27344 32172 27396 32224
rect 27528 32215 27580 32224
rect 27528 32181 27537 32215
rect 27537 32181 27571 32215
rect 27571 32181 27580 32215
rect 27528 32172 27580 32181
rect 29184 32172 29236 32224
rect 30012 32172 30064 32224
rect 30288 32172 30340 32224
rect 30840 32215 30892 32224
rect 30840 32181 30849 32215
rect 30849 32181 30883 32215
rect 30883 32181 30892 32215
rect 30840 32172 30892 32181
rect 33508 32172 33560 32224
rect 34796 32308 34848 32360
rect 37740 32376 37792 32428
rect 35532 32308 35584 32360
rect 35624 32308 35676 32360
rect 37648 32308 37700 32360
rect 38568 32308 38620 32360
rect 34704 32240 34756 32292
rect 34888 32172 34940 32224
rect 35624 32215 35676 32224
rect 35624 32181 35633 32215
rect 35633 32181 35667 32215
rect 35667 32181 35676 32215
rect 35624 32172 35676 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 5908 31968 5960 32020
rect 6184 32011 6236 32020
rect 6184 31977 6193 32011
rect 6193 31977 6227 32011
rect 6227 31977 6236 32011
rect 6184 31968 6236 31977
rect 7932 32011 7984 32020
rect 7932 31977 7941 32011
rect 7941 31977 7975 32011
rect 7975 31977 7984 32011
rect 7932 31968 7984 31977
rect 5724 31764 5776 31816
rect 6000 31807 6052 31816
rect 6000 31773 6009 31807
rect 6009 31773 6043 31807
rect 6043 31773 6052 31807
rect 6000 31764 6052 31773
rect 8116 31807 8168 31816
rect 8116 31773 8125 31807
rect 8125 31773 8159 31807
rect 8159 31773 8168 31807
rect 8116 31764 8168 31773
rect 8484 31968 8536 32020
rect 8760 31968 8812 32020
rect 9680 31968 9732 32020
rect 9772 31968 9824 32020
rect 12256 31968 12308 32020
rect 12348 31968 12400 32020
rect 14096 31968 14148 32020
rect 9128 31900 9180 31952
rect 8944 31832 8996 31884
rect 5816 31739 5868 31748
rect 5816 31705 5825 31739
rect 5825 31705 5859 31739
rect 5859 31705 5868 31739
rect 5816 31696 5868 31705
rect 8484 31696 8536 31748
rect 9036 31696 9088 31748
rect 6368 31628 6420 31680
rect 8576 31628 8628 31680
rect 8852 31628 8904 31680
rect 9220 31628 9272 31680
rect 10232 31900 10284 31952
rect 10048 31832 10100 31884
rect 10416 31832 10468 31884
rect 10784 31943 10836 31952
rect 10784 31909 10793 31943
rect 10793 31909 10827 31943
rect 10827 31909 10836 31943
rect 10784 31900 10836 31909
rect 11888 31832 11940 31884
rect 14280 31968 14332 32020
rect 15016 31968 15068 32020
rect 15936 32011 15988 32020
rect 15936 31977 15945 32011
rect 15945 31977 15979 32011
rect 15979 31977 15988 32011
rect 15936 31968 15988 31977
rect 16672 32011 16724 32020
rect 16672 31977 16681 32011
rect 16681 31977 16715 32011
rect 16715 31977 16724 32011
rect 16672 31968 16724 31977
rect 13084 31832 13136 31884
rect 10048 31739 10100 31748
rect 10048 31705 10057 31739
rect 10057 31705 10091 31739
rect 10091 31705 10100 31739
rect 10048 31696 10100 31705
rect 9588 31628 9640 31680
rect 9772 31628 9824 31680
rect 10508 31696 10560 31748
rect 11612 31696 11664 31748
rect 12900 31807 12952 31816
rect 12900 31773 12914 31807
rect 12914 31773 12948 31807
rect 12948 31773 12952 31807
rect 12900 31764 12952 31773
rect 10968 31628 11020 31680
rect 12624 31628 12676 31680
rect 13176 31628 13228 31680
rect 13544 31832 13596 31884
rect 13912 31875 13964 31884
rect 13912 31841 13921 31875
rect 13921 31841 13955 31875
rect 13955 31841 13964 31875
rect 13912 31832 13964 31841
rect 13452 31696 13504 31748
rect 14096 31764 14148 31816
rect 17040 31943 17092 31952
rect 17040 31909 17049 31943
rect 17049 31909 17083 31943
rect 17083 31909 17092 31943
rect 17040 31900 17092 31909
rect 17868 31900 17920 31952
rect 18236 31900 18288 31952
rect 19248 31968 19300 32020
rect 20812 32011 20864 32020
rect 20812 31977 20821 32011
rect 20821 31977 20855 32011
rect 20855 31977 20864 32011
rect 20812 31968 20864 31977
rect 21088 31968 21140 32020
rect 21272 32011 21324 32020
rect 21272 31977 21281 32011
rect 21281 31977 21315 32011
rect 21315 31977 21324 32011
rect 21272 31968 21324 31977
rect 21364 31968 21416 32020
rect 19892 31900 19944 31952
rect 16580 31832 16632 31884
rect 15660 31807 15712 31816
rect 15660 31773 15669 31807
rect 15669 31773 15703 31807
rect 15703 31773 15712 31807
rect 15660 31764 15712 31773
rect 15936 31807 15988 31816
rect 15936 31773 15945 31807
rect 15945 31773 15979 31807
rect 15979 31773 15988 31807
rect 15936 31764 15988 31773
rect 16120 31764 16172 31816
rect 17408 31832 17460 31884
rect 20996 31900 21048 31952
rect 17132 31807 17184 31816
rect 17132 31773 17141 31807
rect 17141 31773 17175 31807
rect 17175 31773 17184 31807
rect 17132 31764 17184 31773
rect 17960 31807 18012 31816
rect 17960 31773 17969 31807
rect 17969 31773 18003 31807
rect 18003 31773 18012 31807
rect 17960 31764 18012 31773
rect 18328 31807 18380 31816
rect 18328 31773 18337 31807
rect 18337 31773 18371 31807
rect 18371 31773 18380 31807
rect 18328 31764 18380 31773
rect 20812 31832 20864 31884
rect 15844 31696 15896 31748
rect 16580 31696 16632 31748
rect 15016 31628 15068 31680
rect 15936 31628 15988 31680
rect 16028 31628 16080 31680
rect 18696 31807 18748 31816
rect 18696 31773 18705 31807
rect 18705 31773 18739 31807
rect 18739 31773 18748 31807
rect 18696 31764 18748 31773
rect 21272 31764 21324 31816
rect 21364 31807 21416 31816
rect 21364 31773 21373 31807
rect 21373 31773 21407 31807
rect 21407 31773 21416 31807
rect 21364 31764 21416 31773
rect 21180 31696 21232 31748
rect 21732 31875 21784 31884
rect 21732 31841 21741 31875
rect 21741 31841 21775 31875
rect 21775 31841 21784 31875
rect 21732 31832 21784 31841
rect 22468 31900 22520 31952
rect 22652 31900 22704 31952
rect 22836 31900 22888 31952
rect 24400 31900 24452 31952
rect 24584 31900 24636 31952
rect 24676 31900 24728 31952
rect 25228 31900 25280 31952
rect 25780 31900 25832 31952
rect 26240 31900 26292 31952
rect 26332 31943 26384 31952
rect 26332 31909 26341 31943
rect 26341 31909 26375 31943
rect 26375 31909 26384 31943
rect 26332 31900 26384 31909
rect 26516 31968 26568 32020
rect 28724 31968 28776 32020
rect 29736 31968 29788 32020
rect 30012 31968 30064 32020
rect 30840 31968 30892 32020
rect 30932 31968 30984 32020
rect 31300 31968 31352 32020
rect 32680 31968 32732 32020
rect 33784 32011 33836 32020
rect 33784 31977 33793 32011
rect 33793 31977 33827 32011
rect 33827 31977 33836 32011
rect 33784 31968 33836 31977
rect 35624 31968 35676 32020
rect 29000 31900 29052 31952
rect 29092 31900 29144 31952
rect 21640 31807 21692 31816
rect 21640 31773 21649 31807
rect 21649 31773 21683 31807
rect 21683 31773 21692 31807
rect 21640 31764 21692 31773
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 23020 31764 23072 31816
rect 24952 31807 25004 31816
rect 24952 31773 24961 31807
rect 24961 31773 24995 31807
rect 24995 31773 25004 31807
rect 24952 31764 25004 31773
rect 25044 31764 25096 31816
rect 22376 31739 22428 31748
rect 22376 31705 22385 31739
rect 22385 31705 22419 31739
rect 22419 31705 22428 31739
rect 25320 31764 25372 31816
rect 25964 31764 26016 31816
rect 26056 31764 26108 31816
rect 28080 31832 28132 31884
rect 28816 31832 28868 31884
rect 22376 31696 22428 31705
rect 27252 31764 27304 31816
rect 27988 31764 28040 31816
rect 26608 31696 26660 31748
rect 18788 31628 18840 31680
rect 19616 31628 19668 31680
rect 22008 31628 22060 31680
rect 23112 31628 23164 31680
rect 25596 31628 25648 31680
rect 26148 31628 26200 31680
rect 26516 31628 26568 31680
rect 26976 31628 27028 31680
rect 27252 31628 27304 31680
rect 27528 31628 27580 31680
rect 28264 31764 28316 31816
rect 28908 31807 28960 31816
rect 28908 31773 28917 31807
rect 28917 31773 28951 31807
rect 28951 31773 28960 31807
rect 28908 31764 28960 31773
rect 29092 31807 29144 31816
rect 29092 31773 29101 31807
rect 29101 31773 29135 31807
rect 29135 31773 29144 31807
rect 29092 31764 29144 31773
rect 29276 31900 29328 31952
rect 29920 31900 29972 31952
rect 29368 31807 29420 31816
rect 29368 31773 29377 31807
rect 29377 31773 29411 31807
rect 29411 31773 29420 31807
rect 29368 31764 29420 31773
rect 30288 31807 30340 31816
rect 30288 31773 30297 31807
rect 30297 31773 30331 31807
rect 30331 31773 30340 31807
rect 30288 31764 30340 31773
rect 30380 31764 30432 31816
rect 31116 31900 31168 31952
rect 33600 31832 33652 31884
rect 34428 31832 34480 31884
rect 33508 31764 33560 31816
rect 34520 31764 34572 31816
rect 28816 31628 28868 31680
rect 29184 31628 29236 31680
rect 30932 31671 30984 31680
rect 30932 31637 30941 31671
rect 30941 31637 30975 31671
rect 30975 31637 30984 31671
rect 30932 31628 30984 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 7656 31424 7708 31476
rect 7288 31356 7340 31408
rect 8024 31356 8076 31408
rect 5816 31331 5868 31340
rect 5816 31297 5825 31331
rect 5825 31297 5859 31331
rect 5859 31297 5868 31331
rect 5816 31288 5868 31297
rect 5908 31331 5960 31340
rect 5908 31297 5917 31331
rect 5917 31297 5951 31331
rect 5951 31297 5960 31331
rect 5908 31288 5960 31297
rect 6000 31331 6052 31340
rect 6000 31297 6009 31331
rect 6009 31297 6043 31331
rect 6043 31297 6052 31331
rect 6000 31288 6052 31297
rect 6092 31288 6144 31340
rect 8852 31424 8904 31476
rect 9220 31424 9272 31476
rect 9404 31356 9456 31408
rect 9588 31399 9640 31408
rect 9588 31365 9597 31399
rect 9597 31365 9631 31399
rect 9631 31365 9640 31399
rect 9588 31356 9640 31365
rect 8760 31331 8812 31340
rect 8760 31297 8769 31331
rect 8769 31297 8803 31331
rect 8803 31297 8812 31331
rect 8760 31288 8812 31297
rect 4620 31220 4672 31272
rect 8668 31152 8720 31204
rect 8944 31288 8996 31340
rect 10048 31424 10100 31476
rect 10508 31424 10560 31476
rect 13176 31424 13228 31476
rect 13360 31424 13412 31476
rect 6460 31084 6512 31136
rect 9404 31152 9456 31204
rect 9588 31220 9640 31272
rect 10968 31220 11020 31272
rect 17408 31424 17460 31476
rect 13820 31356 13872 31408
rect 12624 31331 12676 31340
rect 12624 31297 12633 31331
rect 12633 31297 12667 31331
rect 12667 31297 12676 31331
rect 12624 31288 12676 31297
rect 12716 31331 12768 31340
rect 12716 31297 12726 31331
rect 12726 31297 12760 31331
rect 12760 31297 12768 31331
rect 12716 31288 12768 31297
rect 12900 31331 12952 31340
rect 12900 31297 12909 31331
rect 12909 31297 12943 31331
rect 12943 31297 12952 31331
rect 12900 31288 12952 31297
rect 12256 31152 12308 31204
rect 12624 31152 12676 31204
rect 13636 31288 13688 31340
rect 14096 31331 14148 31340
rect 14096 31297 14105 31331
rect 14105 31297 14139 31331
rect 14139 31297 14148 31331
rect 14096 31288 14148 31297
rect 14280 31331 14332 31340
rect 14280 31297 14287 31331
rect 14287 31297 14332 31331
rect 14280 31288 14332 31297
rect 14924 31288 14976 31340
rect 15568 31356 15620 31408
rect 15936 31356 15988 31408
rect 22468 31424 22520 31476
rect 31024 31467 31076 31476
rect 16120 31288 16172 31340
rect 16304 31288 16356 31340
rect 18512 31288 18564 31340
rect 19984 31288 20036 31340
rect 16488 31220 16540 31272
rect 17408 31220 17460 31272
rect 21088 31331 21140 31340
rect 21088 31297 21097 31331
rect 21097 31297 21131 31331
rect 21131 31297 21140 31331
rect 21088 31288 21140 31297
rect 21180 31331 21232 31340
rect 21180 31297 21189 31331
rect 21189 31297 21223 31331
rect 21223 31297 21232 31331
rect 21180 31288 21232 31297
rect 21548 31331 21600 31340
rect 21548 31297 21557 31331
rect 21557 31297 21591 31331
rect 21591 31297 21600 31331
rect 21548 31288 21600 31297
rect 14556 31152 14608 31204
rect 15936 31152 15988 31204
rect 21364 31152 21416 31204
rect 22376 31288 22428 31340
rect 23480 31288 23532 31340
rect 23848 31288 23900 31340
rect 24032 31288 24084 31340
rect 24216 31288 24268 31340
rect 24676 31356 24728 31408
rect 25688 31399 25740 31408
rect 25688 31365 25697 31399
rect 25697 31365 25731 31399
rect 25731 31365 25740 31399
rect 25688 31356 25740 31365
rect 24768 31331 24820 31340
rect 24768 31297 24777 31331
rect 24777 31297 24811 31331
rect 24811 31297 24820 31331
rect 24768 31288 24820 31297
rect 25044 31331 25096 31340
rect 25044 31297 25053 31331
rect 25053 31297 25087 31331
rect 25087 31297 25096 31331
rect 25044 31288 25096 31297
rect 25136 31331 25188 31340
rect 25136 31297 25145 31331
rect 25145 31297 25179 31331
rect 25179 31297 25188 31331
rect 25136 31288 25188 31297
rect 25596 31331 25648 31340
rect 25596 31297 25605 31331
rect 25605 31297 25639 31331
rect 25639 31297 25648 31331
rect 25596 31288 25648 31297
rect 25780 31331 25832 31340
rect 25780 31297 25789 31331
rect 25789 31297 25823 31331
rect 25823 31297 25832 31331
rect 25780 31288 25832 31297
rect 25964 31356 26016 31408
rect 26056 31288 26108 31340
rect 27160 31356 27212 31408
rect 27620 31356 27672 31408
rect 28724 31356 28776 31408
rect 31024 31433 31033 31467
rect 31033 31433 31067 31467
rect 31067 31433 31076 31467
rect 31024 31424 31076 31433
rect 31208 31424 31260 31476
rect 26240 31288 26292 31340
rect 22100 31263 22152 31272
rect 22100 31229 22109 31263
rect 22109 31229 22143 31263
rect 22143 31229 22152 31263
rect 22100 31220 22152 31229
rect 22560 31220 22612 31272
rect 23112 31152 23164 31204
rect 23388 31152 23440 31204
rect 23664 31195 23716 31204
rect 23664 31161 23673 31195
rect 23673 31161 23707 31195
rect 23707 31161 23716 31195
rect 23664 31152 23716 31161
rect 24676 31220 24728 31272
rect 26516 31288 26568 31340
rect 28264 31288 28316 31340
rect 28540 31331 28592 31340
rect 28540 31297 28549 31331
rect 28549 31297 28583 31331
rect 28583 31297 28592 31331
rect 28540 31288 28592 31297
rect 29092 31288 29144 31340
rect 29368 31288 29420 31340
rect 26240 31152 26292 31204
rect 9864 31127 9916 31136
rect 9864 31093 9873 31127
rect 9873 31093 9907 31127
rect 9907 31093 9916 31127
rect 9864 31084 9916 31093
rect 10048 31084 10100 31136
rect 10416 31084 10468 31136
rect 10508 31084 10560 31136
rect 11244 31084 11296 31136
rect 11428 31084 11480 31136
rect 11796 31084 11848 31136
rect 12348 31084 12400 31136
rect 16120 31084 16172 31136
rect 19248 31084 19300 31136
rect 24492 31084 24544 31136
rect 24952 31084 25004 31136
rect 25136 31084 25188 31136
rect 25320 31127 25372 31136
rect 25320 31093 25329 31127
rect 25329 31093 25363 31127
rect 25363 31093 25372 31127
rect 25320 31084 25372 31093
rect 25596 31084 25648 31136
rect 28080 31220 28132 31272
rect 27528 31152 27580 31204
rect 28724 31220 28776 31272
rect 30196 31331 30248 31340
rect 30196 31297 30205 31331
rect 30205 31297 30239 31331
rect 30239 31297 30248 31331
rect 30196 31288 30248 31297
rect 30840 31288 30892 31340
rect 31300 31356 31352 31408
rect 33600 31356 33652 31408
rect 31208 31331 31260 31340
rect 31208 31297 31217 31331
rect 31217 31297 31251 31331
rect 31251 31297 31260 31331
rect 31208 31288 31260 31297
rect 32404 31288 32456 31340
rect 32772 31288 32824 31340
rect 29828 31220 29880 31272
rect 31944 31220 31996 31272
rect 32956 31220 33008 31272
rect 33508 31220 33560 31272
rect 26700 31084 26752 31136
rect 30104 31084 30156 31136
rect 33784 31127 33836 31136
rect 33784 31093 33793 31127
rect 33793 31093 33827 31127
rect 33827 31093 33836 31127
rect 33784 31084 33836 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7288 30923 7340 30932
rect 7288 30889 7297 30923
rect 7297 30889 7331 30923
rect 7331 30889 7340 30923
rect 7288 30880 7340 30889
rect 4528 30744 4580 30796
rect 5448 30676 5500 30728
rect 6184 30744 6236 30796
rect 6276 30719 6328 30728
rect 6276 30685 6285 30719
rect 6285 30685 6319 30719
rect 6319 30685 6328 30719
rect 6276 30676 6328 30685
rect 6460 30719 6512 30728
rect 6460 30685 6469 30719
rect 6469 30685 6503 30719
rect 6503 30685 6512 30719
rect 6460 30676 6512 30685
rect 7196 30719 7248 30728
rect 7196 30685 7205 30719
rect 7205 30685 7239 30719
rect 7239 30685 7248 30719
rect 7196 30676 7248 30685
rect 6184 30651 6236 30660
rect 6184 30617 6193 30651
rect 6193 30617 6227 30651
rect 6227 30617 6236 30651
rect 6184 30608 6236 30617
rect 9588 30880 9640 30932
rect 10968 30880 11020 30932
rect 12348 30880 12400 30932
rect 12716 30880 12768 30932
rect 15844 30880 15896 30932
rect 16396 30880 16448 30932
rect 16948 30880 17000 30932
rect 7564 30744 7616 30796
rect 9956 30744 10008 30796
rect 10692 30812 10744 30864
rect 10784 30744 10836 30796
rect 11428 30787 11480 30796
rect 11428 30753 11437 30787
rect 11437 30753 11471 30787
rect 11471 30753 11480 30787
rect 11428 30744 11480 30753
rect 9036 30608 9088 30660
rect 9588 30608 9640 30660
rect 10968 30676 11020 30728
rect 11336 30719 11388 30728
rect 11336 30685 11345 30719
rect 11345 30685 11379 30719
rect 11379 30685 11388 30719
rect 11336 30676 11388 30685
rect 15108 30812 15160 30864
rect 17224 30812 17276 30864
rect 18328 30880 18380 30932
rect 19248 30880 19300 30932
rect 22192 30880 22244 30932
rect 22468 30880 22520 30932
rect 22560 30880 22612 30932
rect 23112 30880 23164 30932
rect 24308 30880 24360 30932
rect 24952 30880 25004 30932
rect 25596 30880 25648 30932
rect 26056 30923 26108 30932
rect 26056 30889 26065 30923
rect 26065 30889 26099 30923
rect 26099 30889 26108 30923
rect 26056 30880 26108 30889
rect 26240 30923 26292 30932
rect 26240 30889 26249 30923
rect 26249 30889 26283 30923
rect 26283 30889 26292 30923
rect 26240 30880 26292 30889
rect 26608 30923 26660 30932
rect 26608 30889 26617 30923
rect 26617 30889 26651 30923
rect 26651 30889 26660 30923
rect 26608 30880 26660 30889
rect 27160 30880 27212 30932
rect 28724 30880 28776 30932
rect 29000 30880 29052 30932
rect 20260 30812 20312 30864
rect 21272 30812 21324 30864
rect 22284 30812 22336 30864
rect 14556 30744 14608 30796
rect 14924 30744 14976 30796
rect 12808 30676 12860 30728
rect 13728 30676 13780 30728
rect 14280 30676 14332 30728
rect 15568 30676 15620 30728
rect 15936 30608 15988 30660
rect 16488 30719 16540 30728
rect 16488 30685 16497 30719
rect 16497 30685 16531 30719
rect 16531 30685 16540 30719
rect 16488 30676 16540 30685
rect 17500 30676 17552 30728
rect 17684 30744 17736 30796
rect 18880 30744 18932 30796
rect 24492 30855 24544 30864
rect 24492 30821 24501 30855
rect 24501 30821 24535 30855
rect 24535 30821 24544 30855
rect 24492 30812 24544 30821
rect 27344 30812 27396 30864
rect 29368 30812 29420 30864
rect 29552 30812 29604 30864
rect 18420 30676 18472 30728
rect 18696 30676 18748 30728
rect 19432 30719 19484 30728
rect 19432 30685 19441 30719
rect 19441 30685 19475 30719
rect 19475 30685 19484 30719
rect 19432 30676 19484 30685
rect 19984 30676 20036 30728
rect 21548 30719 21600 30728
rect 21548 30685 21557 30719
rect 21557 30685 21591 30719
rect 21591 30685 21600 30719
rect 21548 30676 21600 30685
rect 21916 30676 21968 30728
rect 22744 30676 22796 30728
rect 8944 30540 8996 30592
rect 9956 30583 10008 30592
rect 9956 30549 9965 30583
rect 9965 30549 9999 30583
rect 9999 30549 10008 30583
rect 9956 30540 10008 30549
rect 10416 30540 10468 30592
rect 11336 30540 11388 30592
rect 15016 30540 15068 30592
rect 18236 30608 18288 30660
rect 19800 30651 19852 30660
rect 19800 30617 19809 30651
rect 19809 30617 19843 30651
rect 19843 30617 19852 30651
rect 19800 30608 19852 30617
rect 20260 30608 20312 30660
rect 23020 30608 23072 30660
rect 16396 30583 16448 30592
rect 16396 30549 16405 30583
rect 16405 30549 16439 30583
rect 16439 30549 16448 30583
rect 16396 30540 16448 30549
rect 17776 30540 17828 30592
rect 21364 30540 21416 30592
rect 22744 30583 22796 30592
rect 22744 30549 22753 30583
rect 22753 30549 22787 30583
rect 22787 30549 22796 30583
rect 22744 30540 22796 30549
rect 24032 30719 24084 30728
rect 24032 30685 24041 30719
rect 24041 30685 24075 30719
rect 24075 30685 24084 30719
rect 24032 30676 24084 30685
rect 25964 30744 26016 30796
rect 24952 30719 25004 30728
rect 24952 30685 24961 30719
rect 24961 30685 24995 30719
rect 24995 30685 25004 30719
rect 24952 30676 25004 30685
rect 24676 30608 24728 30660
rect 25872 30719 25924 30728
rect 25872 30685 25881 30719
rect 25881 30685 25915 30719
rect 25915 30685 25924 30719
rect 25872 30676 25924 30685
rect 27804 30787 27856 30796
rect 27804 30753 27813 30787
rect 27813 30753 27847 30787
rect 27847 30753 27856 30787
rect 27804 30744 27856 30753
rect 25596 30651 25648 30660
rect 25596 30617 25605 30651
rect 25605 30617 25639 30651
rect 25639 30617 25648 30651
rect 25596 30608 25648 30617
rect 26516 30719 26568 30728
rect 26516 30685 26525 30719
rect 26525 30685 26559 30719
rect 26559 30685 26568 30719
rect 26516 30676 26568 30685
rect 26608 30719 26660 30728
rect 26608 30685 26617 30719
rect 26617 30685 26651 30719
rect 26651 30685 26660 30719
rect 26608 30676 26660 30685
rect 26700 30676 26752 30728
rect 26884 30608 26936 30660
rect 27436 30608 27488 30660
rect 27620 30719 27672 30728
rect 27620 30685 27629 30719
rect 27629 30685 27663 30719
rect 27663 30685 27672 30719
rect 27620 30676 27672 30685
rect 27712 30676 27764 30728
rect 28172 30676 28224 30728
rect 28816 30719 28868 30728
rect 28816 30685 28825 30719
rect 28825 30685 28859 30719
rect 28859 30685 28868 30719
rect 28816 30676 28868 30685
rect 29368 30719 29420 30728
rect 29368 30685 29377 30719
rect 29377 30685 29411 30719
rect 29411 30685 29420 30719
rect 29368 30676 29420 30685
rect 29644 30744 29696 30796
rect 32680 30744 32732 30796
rect 34060 30744 34112 30796
rect 31208 30676 31260 30728
rect 33508 30676 33560 30728
rect 35440 30676 35492 30728
rect 26608 30540 26660 30592
rect 26976 30540 27028 30592
rect 27620 30540 27672 30592
rect 29092 30583 29144 30592
rect 29092 30549 29101 30583
rect 29101 30549 29135 30583
rect 29135 30549 29144 30583
rect 29092 30540 29144 30549
rect 32772 30608 32824 30660
rect 29460 30540 29512 30592
rect 31576 30540 31628 30592
rect 33232 30583 33284 30592
rect 33232 30549 33241 30583
rect 33241 30549 33275 30583
rect 33275 30549 33284 30583
rect 33232 30540 33284 30549
rect 33876 30608 33928 30660
rect 34152 30540 34204 30592
rect 34612 30540 34664 30592
rect 35900 30540 35952 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 8484 30336 8536 30388
rect 9680 30336 9732 30388
rect 11060 30336 11112 30388
rect 14004 30336 14056 30388
rect 7656 30200 7708 30252
rect 12256 30268 12308 30320
rect 13728 30268 13780 30320
rect 15660 30336 15712 30388
rect 7932 30132 7984 30184
rect 8760 30132 8812 30184
rect 10416 30200 10468 30252
rect 10692 30243 10744 30252
rect 10692 30209 10702 30243
rect 10702 30209 10736 30243
rect 10736 30209 10744 30243
rect 10692 30200 10744 30209
rect 8852 30064 8904 30116
rect 10508 30132 10560 30184
rect 11520 30175 11572 30184
rect 11520 30141 11529 30175
rect 11529 30141 11563 30175
rect 11563 30141 11572 30175
rect 11520 30132 11572 30141
rect 9588 30064 9640 30116
rect 10600 30064 10652 30116
rect 11888 30200 11940 30252
rect 12808 30200 12860 30252
rect 12992 30200 13044 30252
rect 13452 30200 13504 30252
rect 14464 30200 14516 30252
rect 15568 30268 15620 30320
rect 16396 30336 16448 30388
rect 18236 30336 18288 30388
rect 16120 30268 16172 30320
rect 12072 30132 12124 30184
rect 14004 30132 14056 30184
rect 14740 30064 14792 30116
rect 16212 30200 16264 30252
rect 16856 30243 16908 30252
rect 16856 30209 16865 30243
rect 16865 30209 16899 30243
rect 16899 30209 16908 30243
rect 16856 30200 16908 30209
rect 18788 30268 18840 30320
rect 19432 30268 19484 30320
rect 22100 30336 22152 30388
rect 22836 30336 22888 30388
rect 23020 30336 23072 30388
rect 25044 30336 25096 30388
rect 25320 30336 25372 30388
rect 25504 30336 25556 30388
rect 27988 30336 28040 30388
rect 28816 30336 28868 30388
rect 29828 30336 29880 30388
rect 35900 30379 35952 30388
rect 35900 30345 35909 30379
rect 35909 30345 35943 30379
rect 35943 30345 35952 30379
rect 35900 30336 35952 30345
rect 19340 30243 19392 30252
rect 19340 30209 19349 30243
rect 19349 30209 19383 30243
rect 19383 30209 19392 30243
rect 19340 30200 19392 30209
rect 18328 30132 18380 30184
rect 18788 30132 18840 30184
rect 19984 30243 20036 30252
rect 19984 30209 19993 30243
rect 19993 30209 20027 30243
rect 20027 30209 20036 30243
rect 19984 30200 20036 30209
rect 20168 30200 20220 30252
rect 22284 30175 22336 30184
rect 22284 30141 22293 30175
rect 22293 30141 22327 30175
rect 22327 30141 22336 30175
rect 22284 30132 22336 30141
rect 22652 30132 22704 30184
rect 23480 30243 23532 30252
rect 23480 30209 23489 30243
rect 23489 30209 23523 30243
rect 23523 30209 23532 30243
rect 23480 30200 23532 30209
rect 23572 30200 23624 30252
rect 24400 30200 24452 30252
rect 25044 30200 25096 30252
rect 25964 30200 26016 30252
rect 28172 30268 28224 30320
rect 28632 30268 28684 30320
rect 32404 30311 32456 30320
rect 32404 30277 32413 30311
rect 32413 30277 32447 30311
rect 32447 30277 32456 30311
rect 32404 30268 32456 30277
rect 24676 30132 24728 30184
rect 25504 30132 25556 30184
rect 9220 29996 9272 30048
rect 9772 29996 9824 30048
rect 10140 29996 10192 30048
rect 11060 29996 11112 30048
rect 11888 30039 11940 30048
rect 11888 30005 11897 30039
rect 11897 30005 11931 30039
rect 11931 30005 11940 30039
rect 11888 29996 11940 30005
rect 14832 29996 14884 30048
rect 14924 29996 14976 30048
rect 15384 29996 15436 30048
rect 15936 29996 15988 30048
rect 16212 30039 16264 30048
rect 16212 30005 16221 30039
rect 16221 30005 16255 30039
rect 16255 30005 16264 30039
rect 16212 29996 16264 30005
rect 16856 30039 16908 30048
rect 16856 30005 16865 30039
rect 16865 30005 16899 30039
rect 16899 30005 16908 30039
rect 16856 29996 16908 30005
rect 17040 30039 17092 30048
rect 17040 30005 17049 30039
rect 17049 30005 17083 30039
rect 17083 30005 17092 30039
rect 17040 29996 17092 30005
rect 18236 29996 18288 30048
rect 18420 29996 18472 30048
rect 19156 30064 19208 30116
rect 19800 30064 19852 30116
rect 20260 30107 20312 30116
rect 20260 30073 20269 30107
rect 20269 30073 20303 30107
rect 20303 30073 20312 30107
rect 20260 30064 20312 30073
rect 20720 30064 20772 30116
rect 26608 30200 26660 30252
rect 27804 30200 27856 30252
rect 30288 30243 30340 30252
rect 30288 30209 30297 30243
rect 30297 30209 30331 30243
rect 30331 30209 30340 30243
rect 30288 30200 30340 30209
rect 30748 30243 30800 30252
rect 30748 30209 30757 30243
rect 30757 30209 30791 30243
rect 30791 30209 30800 30243
rect 30748 30200 30800 30209
rect 27160 30132 27212 30184
rect 29920 30132 29972 30184
rect 30104 30132 30156 30184
rect 26516 30064 26568 30116
rect 31576 30243 31628 30252
rect 31576 30209 31585 30243
rect 31585 30209 31619 30243
rect 31619 30209 31628 30243
rect 31576 30200 31628 30209
rect 32680 30243 32732 30252
rect 32680 30209 32689 30243
rect 32689 30209 32723 30243
rect 32723 30209 32732 30243
rect 32680 30200 32732 30209
rect 32956 30200 33008 30252
rect 33232 30200 33284 30252
rect 33508 30200 33560 30252
rect 33600 30200 33652 30252
rect 33784 30200 33836 30252
rect 31300 30132 31352 30184
rect 32220 30132 32272 30184
rect 34152 30200 34204 30252
rect 34520 30200 34572 30252
rect 35256 30175 35308 30184
rect 35256 30141 35265 30175
rect 35265 30141 35299 30175
rect 35299 30141 35308 30175
rect 35256 30132 35308 30141
rect 20812 29996 20864 30048
rect 23480 29996 23532 30048
rect 23756 29996 23808 30048
rect 24032 29996 24084 30048
rect 26608 29996 26660 30048
rect 30104 30039 30156 30048
rect 30104 30005 30113 30039
rect 30113 30005 30147 30039
rect 30147 30005 30156 30039
rect 30104 29996 30156 30005
rect 30196 29996 30248 30048
rect 34612 30064 34664 30116
rect 34796 29996 34848 30048
rect 35532 29996 35584 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 7656 29835 7708 29844
rect 7656 29801 7665 29835
rect 7665 29801 7699 29835
rect 7699 29801 7708 29835
rect 7656 29792 7708 29801
rect 11060 29792 11112 29844
rect 11336 29792 11388 29844
rect 12256 29792 12308 29844
rect 14372 29835 14424 29844
rect 14372 29801 14381 29835
rect 14381 29801 14415 29835
rect 14415 29801 14424 29835
rect 14372 29792 14424 29801
rect 14740 29792 14792 29844
rect 16028 29792 16080 29844
rect 16396 29792 16448 29844
rect 18052 29792 18104 29844
rect 19340 29835 19392 29844
rect 19340 29801 19349 29835
rect 19349 29801 19383 29835
rect 19383 29801 19392 29835
rect 19340 29792 19392 29801
rect 20352 29792 20404 29844
rect 9496 29724 9548 29776
rect 9680 29724 9732 29776
rect 8024 29699 8076 29708
rect 8024 29665 8033 29699
rect 8033 29665 8067 29699
rect 8067 29665 8076 29699
rect 8024 29656 8076 29665
rect 5724 29631 5776 29640
rect 5724 29597 5733 29631
rect 5733 29597 5767 29631
rect 5767 29597 5776 29631
rect 5724 29588 5776 29597
rect 6092 29588 6144 29640
rect 6184 29588 6236 29640
rect 6460 29588 6512 29640
rect 5264 29520 5316 29572
rect 7932 29631 7984 29640
rect 7932 29597 7941 29631
rect 7941 29597 7975 29631
rect 7975 29597 7984 29631
rect 7932 29588 7984 29597
rect 8208 29588 8260 29640
rect 8392 29631 8444 29640
rect 8392 29597 8401 29631
rect 8401 29597 8435 29631
rect 8435 29597 8444 29631
rect 8392 29588 8444 29597
rect 8484 29631 8536 29640
rect 8484 29597 8493 29631
rect 8493 29597 8527 29631
rect 8527 29597 8536 29631
rect 8484 29588 8536 29597
rect 8944 29656 8996 29708
rect 9588 29656 9640 29708
rect 9956 29724 10008 29776
rect 9312 29631 9364 29640
rect 9312 29597 9321 29631
rect 9321 29597 9355 29631
rect 9355 29597 9364 29631
rect 9312 29588 9364 29597
rect 9680 29631 9732 29640
rect 9680 29597 9689 29631
rect 9689 29597 9723 29631
rect 9723 29597 9732 29631
rect 9680 29588 9732 29597
rect 9772 29631 9824 29640
rect 9772 29597 9782 29631
rect 9782 29597 9816 29631
rect 9816 29597 9824 29631
rect 9772 29588 9824 29597
rect 8668 29520 8720 29572
rect 8852 29520 8904 29572
rect 9588 29520 9640 29572
rect 10048 29631 10100 29640
rect 10048 29597 10057 29631
rect 10057 29597 10091 29631
rect 10091 29597 10100 29631
rect 10048 29588 10100 29597
rect 10140 29588 10192 29640
rect 10324 29588 10376 29640
rect 10508 29631 10560 29640
rect 10508 29597 10517 29631
rect 10517 29597 10551 29631
rect 10551 29597 10560 29631
rect 10508 29588 10560 29597
rect 11520 29656 11572 29708
rect 15292 29724 15344 29776
rect 16120 29724 16172 29776
rect 17868 29767 17920 29776
rect 17868 29733 17877 29767
rect 17877 29733 17911 29767
rect 17911 29733 17920 29767
rect 17868 29724 17920 29733
rect 18236 29724 18288 29776
rect 19156 29724 19208 29776
rect 19432 29724 19484 29776
rect 21548 29724 21600 29776
rect 22744 29792 22796 29844
rect 23940 29792 23992 29844
rect 27528 29792 27580 29844
rect 30196 29792 30248 29844
rect 35348 29792 35400 29844
rect 35440 29835 35492 29844
rect 35440 29801 35449 29835
rect 35449 29801 35483 29835
rect 35483 29801 35492 29835
rect 35440 29792 35492 29801
rect 37556 29835 37608 29844
rect 37556 29801 37565 29835
rect 37565 29801 37599 29835
rect 37599 29801 37608 29835
rect 37556 29792 37608 29801
rect 22284 29724 22336 29776
rect 23572 29724 23624 29776
rect 24584 29724 24636 29776
rect 26240 29724 26292 29776
rect 29828 29767 29880 29776
rect 29828 29733 29837 29767
rect 29837 29733 29871 29767
rect 29871 29733 29880 29767
rect 29828 29724 29880 29733
rect 30564 29767 30616 29776
rect 30564 29733 30573 29767
rect 30573 29733 30607 29767
rect 30607 29733 30616 29767
rect 30564 29724 30616 29733
rect 14924 29699 14976 29708
rect 12440 29588 12492 29640
rect 14924 29665 14933 29699
rect 14933 29665 14967 29699
rect 14967 29665 14976 29699
rect 14924 29656 14976 29665
rect 18696 29699 18748 29708
rect 12900 29631 12952 29640
rect 12900 29597 12909 29631
rect 12909 29597 12943 29631
rect 12943 29597 12952 29631
rect 12900 29588 12952 29597
rect 13176 29588 13228 29640
rect 13728 29588 13780 29640
rect 14372 29588 14424 29640
rect 15384 29631 15436 29640
rect 15384 29597 15393 29631
rect 15393 29597 15427 29631
rect 15427 29597 15436 29631
rect 15384 29588 15436 29597
rect 6000 29495 6052 29504
rect 6000 29461 6009 29495
rect 6009 29461 6043 29495
rect 6043 29461 6052 29495
rect 6000 29452 6052 29461
rect 8300 29452 8352 29504
rect 9036 29452 9088 29504
rect 9404 29452 9456 29504
rect 9956 29452 10008 29504
rect 11060 29520 11112 29572
rect 14924 29520 14976 29572
rect 12440 29495 12492 29504
rect 12440 29461 12449 29495
rect 12449 29461 12483 29495
rect 12483 29461 12492 29495
rect 12440 29452 12492 29461
rect 13912 29452 13964 29504
rect 16304 29631 16356 29640
rect 16304 29597 16313 29631
rect 16313 29597 16347 29631
rect 16347 29597 16356 29631
rect 16304 29588 16356 29597
rect 16396 29588 16448 29640
rect 16580 29631 16632 29640
rect 16580 29597 16589 29631
rect 16589 29597 16623 29631
rect 16623 29597 16632 29631
rect 16580 29588 16632 29597
rect 17040 29631 17092 29640
rect 17040 29597 17049 29631
rect 17049 29597 17083 29631
rect 17083 29597 17092 29631
rect 17040 29588 17092 29597
rect 17132 29588 17184 29640
rect 17592 29588 17644 29640
rect 15568 29452 15620 29504
rect 15844 29495 15896 29504
rect 15844 29461 15853 29495
rect 15853 29461 15887 29495
rect 15887 29461 15896 29495
rect 15844 29452 15896 29461
rect 16028 29452 16080 29504
rect 16120 29452 16172 29504
rect 17316 29452 17368 29504
rect 18696 29665 18705 29699
rect 18705 29665 18739 29699
rect 18739 29665 18748 29699
rect 18696 29656 18748 29665
rect 18236 29631 18288 29640
rect 18236 29597 18245 29631
rect 18245 29597 18279 29631
rect 18279 29597 18288 29631
rect 18236 29588 18288 29597
rect 18972 29588 19024 29640
rect 19340 29588 19392 29640
rect 19892 29631 19944 29640
rect 19892 29597 19901 29631
rect 19901 29597 19935 29631
rect 19935 29597 19944 29631
rect 19892 29588 19944 29597
rect 22100 29699 22152 29708
rect 22100 29665 22109 29699
rect 22109 29665 22143 29699
rect 22143 29665 22152 29699
rect 22100 29656 22152 29665
rect 22468 29699 22520 29708
rect 22468 29665 22477 29699
rect 22477 29665 22511 29699
rect 22511 29665 22520 29699
rect 22468 29656 22520 29665
rect 20720 29588 20772 29640
rect 20812 29588 20864 29640
rect 21548 29631 21600 29640
rect 21548 29597 21557 29631
rect 21557 29597 21591 29631
rect 21591 29597 21600 29631
rect 21548 29588 21600 29597
rect 18144 29452 18196 29504
rect 18236 29452 18288 29504
rect 18696 29452 18748 29504
rect 20076 29452 20128 29504
rect 21088 29520 21140 29572
rect 21916 29588 21968 29640
rect 22836 29656 22888 29708
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 22284 29520 22336 29572
rect 22836 29554 22888 29606
rect 23204 29588 23256 29640
rect 23296 29631 23348 29640
rect 23296 29597 23305 29631
rect 23305 29597 23339 29631
rect 23339 29597 23348 29631
rect 23296 29588 23348 29597
rect 24032 29656 24084 29708
rect 24308 29656 24360 29708
rect 24952 29656 25004 29708
rect 25596 29656 25648 29708
rect 27528 29656 27580 29708
rect 29000 29656 29052 29708
rect 25964 29588 26016 29640
rect 27620 29631 27672 29640
rect 27620 29597 27629 29631
rect 27629 29597 27663 29631
rect 27663 29597 27672 29631
rect 27620 29588 27672 29597
rect 27804 29588 27856 29640
rect 32220 29656 32272 29708
rect 22468 29452 22520 29504
rect 22836 29495 22888 29504
rect 22836 29461 22845 29495
rect 22845 29461 22879 29495
rect 22879 29461 22888 29495
rect 22836 29452 22888 29461
rect 23572 29520 23624 29572
rect 30104 29588 30156 29640
rect 30288 29631 30340 29640
rect 30288 29597 30297 29631
rect 30297 29597 30331 29631
rect 30331 29597 30340 29631
rect 30288 29588 30340 29597
rect 30380 29631 30432 29640
rect 30380 29597 30389 29631
rect 30389 29597 30423 29631
rect 30423 29597 30432 29631
rect 31300 29631 31352 29640
rect 30380 29588 30432 29597
rect 31300 29597 31309 29631
rect 31309 29597 31343 29631
rect 31343 29597 31352 29631
rect 31300 29588 31352 29597
rect 31484 29631 31536 29640
rect 31484 29597 31493 29631
rect 31493 29597 31527 29631
rect 31527 29597 31536 29631
rect 31484 29588 31536 29597
rect 32680 29588 32732 29640
rect 24768 29452 24820 29504
rect 25044 29452 25096 29504
rect 25596 29452 25648 29504
rect 26240 29452 26292 29504
rect 27528 29452 27580 29504
rect 30748 29520 30800 29572
rect 30932 29563 30984 29572
rect 30932 29529 30941 29563
rect 30941 29529 30975 29563
rect 30975 29529 30984 29563
rect 30932 29520 30984 29529
rect 31576 29520 31628 29572
rect 33232 29631 33284 29640
rect 33232 29597 33241 29631
rect 33241 29597 33275 29631
rect 33275 29597 33284 29631
rect 33232 29588 33284 29597
rect 33600 29631 33652 29640
rect 33600 29597 33609 29631
rect 33609 29597 33643 29631
rect 33643 29597 33652 29631
rect 33600 29588 33652 29597
rect 33784 29588 33836 29640
rect 34520 29588 34572 29640
rect 34796 29631 34848 29640
rect 34796 29597 34805 29631
rect 34805 29597 34839 29631
rect 34839 29597 34848 29631
rect 34796 29588 34848 29597
rect 35808 29699 35860 29708
rect 35808 29665 35817 29699
rect 35817 29665 35851 29699
rect 35851 29665 35860 29699
rect 35808 29656 35860 29665
rect 27988 29495 28040 29504
rect 27988 29461 27997 29495
rect 27997 29461 28031 29495
rect 28031 29461 28040 29495
rect 27988 29452 28040 29461
rect 29552 29452 29604 29504
rect 30012 29452 30064 29504
rect 30656 29452 30708 29504
rect 34612 29520 34664 29572
rect 35716 29631 35768 29640
rect 35716 29597 35725 29631
rect 35725 29597 35759 29631
rect 35759 29597 35768 29631
rect 35716 29588 35768 29597
rect 38108 29588 38160 29640
rect 31760 29452 31812 29504
rect 32956 29452 33008 29504
rect 34152 29452 34204 29504
rect 36268 29452 36320 29504
rect 37648 29520 37700 29572
rect 37924 29520 37976 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 7564 29291 7616 29300
rect 7564 29257 7573 29291
rect 7573 29257 7607 29291
rect 7607 29257 7616 29291
rect 7564 29248 7616 29257
rect 7840 29248 7892 29300
rect 8484 29248 8536 29300
rect 8760 29248 8812 29300
rect 9404 29248 9456 29300
rect 11888 29248 11940 29300
rect 12900 29291 12952 29300
rect 12900 29257 12909 29291
rect 12909 29257 12943 29291
rect 12943 29257 12952 29291
rect 12900 29248 12952 29257
rect 13544 29248 13596 29300
rect 5724 29180 5776 29232
rect 5448 29112 5500 29164
rect 3792 29044 3844 29096
rect 6000 28976 6052 29028
rect 7564 29112 7616 29164
rect 7932 29044 7984 29096
rect 8116 29044 8168 29096
rect 9588 29180 9640 29232
rect 9404 29112 9456 29164
rect 9680 29155 9732 29164
rect 9680 29121 9689 29155
rect 9689 29121 9723 29155
rect 9723 29121 9732 29155
rect 9680 29112 9732 29121
rect 9772 29155 9824 29164
rect 9772 29121 9782 29155
rect 9782 29121 9816 29155
rect 9816 29121 9824 29155
rect 10048 29155 10100 29164
rect 9772 29112 9824 29121
rect 8208 28976 8260 29028
rect 9128 28976 9180 29028
rect 9680 28976 9732 29028
rect 9772 28976 9824 29028
rect 10048 29121 10057 29155
rect 10057 29121 10091 29155
rect 10091 29121 10100 29155
rect 10048 29112 10100 29121
rect 10508 29180 10560 29232
rect 14372 29180 14424 29232
rect 14648 29180 14700 29232
rect 14924 29248 14976 29300
rect 16672 29248 16724 29300
rect 17316 29248 17368 29300
rect 18788 29248 18840 29300
rect 19248 29248 19300 29300
rect 15660 29180 15712 29232
rect 16488 29180 16540 29232
rect 19340 29180 19392 29232
rect 11060 29044 11112 29096
rect 13820 29112 13872 29164
rect 12900 29044 12952 29096
rect 13636 29044 13688 29096
rect 14740 29155 14792 29164
rect 14740 29121 14749 29155
rect 14749 29121 14783 29155
rect 14783 29121 14792 29155
rect 14740 29112 14792 29121
rect 14648 29087 14700 29096
rect 14648 29053 14657 29087
rect 14657 29053 14691 29087
rect 14691 29053 14700 29087
rect 14648 29044 14700 29053
rect 14832 29044 14884 29096
rect 15292 29044 15344 29096
rect 15476 29112 15528 29164
rect 16120 29112 16172 29164
rect 16304 29112 16356 29164
rect 16672 29112 16724 29164
rect 17040 29112 17092 29164
rect 17500 29112 17552 29164
rect 15568 29044 15620 29096
rect 16120 29019 16172 29028
rect 16120 28985 16129 29019
rect 16129 28985 16163 29019
rect 16163 28985 16172 29019
rect 16120 28976 16172 28985
rect 18604 29155 18656 29164
rect 18604 29121 18613 29155
rect 18613 29121 18647 29155
rect 18647 29121 18656 29155
rect 18604 29112 18656 29121
rect 18144 29087 18196 29096
rect 18144 29053 18153 29087
rect 18153 29053 18187 29087
rect 18187 29053 18196 29087
rect 18144 29044 18196 29053
rect 18328 29044 18380 29096
rect 19524 29112 19576 29164
rect 20628 29180 20680 29232
rect 23020 29248 23072 29300
rect 23112 29248 23164 29300
rect 19984 29112 20036 29164
rect 18880 29087 18932 29096
rect 18880 29053 18889 29087
rect 18889 29053 18923 29087
rect 18923 29053 18932 29087
rect 18880 29044 18932 29053
rect 17776 28976 17828 29028
rect 10784 28951 10836 28960
rect 10784 28917 10793 28951
rect 10793 28917 10827 28951
rect 10827 28917 10836 28951
rect 10784 28908 10836 28917
rect 13728 28908 13780 28960
rect 15660 28908 15712 28960
rect 16304 28908 16356 28960
rect 17132 28908 17184 28960
rect 17684 28908 17736 28960
rect 20168 28976 20220 29028
rect 20352 29155 20404 29164
rect 20352 29121 20361 29155
rect 20361 29121 20395 29155
rect 20395 29121 20404 29155
rect 20352 29112 20404 29121
rect 20444 29155 20496 29164
rect 20444 29121 20453 29155
rect 20453 29121 20487 29155
rect 20487 29121 20496 29155
rect 20444 29112 20496 29121
rect 21180 29223 21232 29232
rect 21180 29189 21189 29223
rect 21189 29189 21223 29223
rect 21223 29189 21232 29223
rect 21180 29180 21232 29189
rect 21272 29180 21324 29232
rect 22468 29155 22520 29164
rect 22468 29121 22477 29155
rect 22477 29121 22511 29155
rect 22511 29121 22520 29155
rect 22468 29112 22520 29121
rect 21640 29044 21692 29096
rect 22744 29155 22796 29164
rect 22744 29121 22753 29155
rect 22753 29121 22787 29155
rect 22787 29121 22796 29155
rect 22744 29112 22796 29121
rect 21364 28976 21416 29028
rect 21916 28976 21968 29028
rect 22008 29019 22060 29028
rect 22008 28985 22017 29019
rect 22017 28985 22051 29019
rect 22051 28985 22060 29019
rect 22008 28976 22060 28985
rect 22284 29019 22336 29028
rect 22284 28985 22293 29019
rect 22293 28985 22327 29019
rect 22327 28985 22336 29019
rect 22284 28976 22336 28985
rect 22560 28976 22612 29028
rect 22468 28908 22520 28960
rect 22744 28976 22796 29028
rect 23204 29044 23256 29096
rect 23940 29044 23992 29096
rect 25596 29248 25648 29300
rect 26516 29291 26568 29300
rect 26516 29257 26525 29291
rect 26525 29257 26559 29291
rect 26559 29257 26568 29291
rect 26516 29248 26568 29257
rect 26700 29248 26752 29300
rect 27344 29248 27396 29300
rect 27896 29248 27948 29300
rect 32220 29248 32272 29300
rect 32680 29248 32732 29300
rect 24308 29155 24360 29164
rect 24308 29121 24317 29155
rect 24317 29121 24351 29155
rect 24351 29121 24360 29155
rect 24308 29112 24360 29121
rect 30104 29180 30156 29232
rect 30288 29223 30340 29232
rect 30288 29189 30322 29223
rect 30322 29189 30340 29223
rect 30288 29180 30340 29189
rect 24492 29155 24544 29164
rect 24492 29121 24501 29155
rect 24501 29121 24535 29155
rect 24535 29121 24544 29155
rect 24492 29112 24544 29121
rect 24584 29044 24636 29096
rect 25228 29112 25280 29164
rect 25688 29112 25740 29164
rect 25780 29112 25832 29164
rect 25964 29112 26016 29164
rect 26424 29112 26476 29164
rect 26516 29155 26568 29164
rect 26516 29121 26525 29155
rect 26525 29121 26559 29155
rect 26559 29121 26568 29155
rect 26516 29112 26568 29121
rect 26608 29155 26660 29164
rect 26608 29121 26617 29155
rect 26617 29121 26651 29155
rect 26651 29121 26660 29155
rect 26608 29112 26660 29121
rect 27344 29112 27396 29164
rect 24952 28908 25004 28960
rect 25596 29044 25648 29096
rect 27988 29112 28040 29164
rect 28172 29155 28224 29164
rect 28172 29121 28181 29155
rect 28181 29121 28215 29155
rect 28215 29121 28224 29155
rect 28172 29112 28224 29121
rect 28448 29112 28500 29164
rect 30012 29112 30064 29164
rect 25320 28976 25372 29028
rect 27712 29044 27764 29096
rect 29000 29044 29052 29096
rect 29644 29044 29696 29096
rect 29828 29087 29880 29096
rect 29828 29053 29837 29087
rect 29837 29053 29871 29087
rect 29871 29053 29880 29087
rect 29828 29044 29880 29053
rect 25964 28976 26016 29028
rect 26240 28976 26292 29028
rect 27896 28976 27948 29028
rect 25228 28908 25280 28960
rect 25872 28951 25924 28960
rect 25872 28917 25881 28951
rect 25881 28917 25915 28951
rect 25915 28917 25924 28951
rect 25872 28908 25924 28917
rect 27620 28908 27672 28960
rect 29276 28976 29328 29028
rect 30380 29044 30432 29096
rect 31300 29155 31352 29164
rect 31300 29121 31309 29155
rect 31309 29121 31343 29155
rect 31343 29121 31352 29155
rect 31300 29112 31352 29121
rect 30748 28976 30800 29028
rect 31760 29155 31812 29164
rect 31760 29121 31794 29155
rect 31794 29121 31812 29155
rect 31760 29112 31812 29121
rect 32772 29155 32824 29164
rect 32772 29121 32781 29155
rect 32781 29121 32815 29155
rect 32815 29121 32824 29155
rect 32772 29112 32824 29121
rect 35716 29248 35768 29300
rect 37556 29248 37608 29300
rect 40960 29291 41012 29300
rect 40960 29257 40969 29291
rect 40969 29257 41003 29291
rect 41003 29257 41012 29291
rect 40960 29248 41012 29257
rect 34152 29155 34204 29164
rect 34152 29121 34161 29155
rect 34161 29121 34195 29155
rect 34195 29121 34204 29155
rect 34152 29112 34204 29121
rect 34520 29112 34572 29164
rect 36452 29087 36504 29096
rect 36452 29053 36461 29087
rect 36461 29053 36495 29087
rect 36495 29053 36504 29087
rect 36452 29044 36504 29053
rect 36544 29087 36596 29096
rect 36544 29053 36553 29087
rect 36553 29053 36587 29087
rect 36587 29053 36596 29087
rect 36544 29044 36596 29053
rect 30196 28908 30248 28960
rect 31576 28908 31628 28960
rect 41328 28976 41380 29028
rect 32772 28908 32824 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 5264 28704 5316 28756
rect 7564 28704 7616 28756
rect 10232 28704 10284 28756
rect 12256 28704 12308 28756
rect 14004 28704 14056 28756
rect 14096 28704 14148 28756
rect 15660 28704 15712 28756
rect 18604 28704 18656 28756
rect 19432 28704 19484 28756
rect 20628 28704 20680 28756
rect 22744 28704 22796 28756
rect 23204 28704 23256 28756
rect 25044 28704 25096 28756
rect 9128 28636 9180 28688
rect 6000 28568 6052 28620
rect 5540 28500 5592 28552
rect 7288 28500 7340 28552
rect 8760 28500 8812 28552
rect 9404 28500 9456 28552
rect 10416 28568 10468 28620
rect 10784 28543 10836 28552
rect 10784 28509 10793 28543
rect 10793 28509 10827 28543
rect 10827 28509 10836 28543
rect 10784 28500 10836 28509
rect 10968 28568 11020 28620
rect 6184 28432 6236 28484
rect 5908 28364 5960 28416
rect 11520 28475 11572 28484
rect 11520 28441 11529 28475
rect 11529 28441 11563 28475
rect 11563 28441 11572 28475
rect 11520 28432 11572 28441
rect 11888 28543 11940 28552
rect 11888 28509 11897 28543
rect 11897 28509 11931 28543
rect 11931 28509 11940 28543
rect 11888 28500 11940 28509
rect 12164 28543 12216 28552
rect 12164 28509 12173 28543
rect 12173 28509 12207 28543
rect 12207 28509 12216 28543
rect 12164 28500 12216 28509
rect 12072 28432 12124 28484
rect 12532 28500 12584 28552
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 13360 28568 13412 28620
rect 19340 28568 19392 28620
rect 13544 28432 13596 28484
rect 13728 28432 13780 28484
rect 16764 28432 16816 28484
rect 17224 28432 17276 28484
rect 18236 28432 18288 28484
rect 18972 28432 19024 28484
rect 19248 28475 19300 28484
rect 19248 28441 19257 28475
rect 19257 28441 19291 28475
rect 19291 28441 19300 28475
rect 19248 28432 19300 28441
rect 19984 28500 20036 28552
rect 20168 28500 20220 28552
rect 20444 28500 20496 28552
rect 20628 28500 20680 28552
rect 10876 28364 10928 28416
rect 11336 28364 11388 28416
rect 12348 28407 12400 28416
rect 12348 28373 12357 28407
rect 12357 28373 12391 28407
rect 12391 28373 12400 28407
rect 12348 28364 12400 28373
rect 12440 28364 12492 28416
rect 15108 28364 15160 28416
rect 17132 28364 17184 28416
rect 18512 28364 18564 28416
rect 18880 28364 18932 28416
rect 19156 28364 19208 28416
rect 20720 28475 20772 28484
rect 20720 28441 20729 28475
rect 20729 28441 20763 28475
rect 20763 28441 20772 28475
rect 20720 28432 20772 28441
rect 21640 28543 21692 28552
rect 21640 28509 21649 28543
rect 21649 28509 21683 28543
rect 21683 28509 21692 28543
rect 21640 28500 21692 28509
rect 21364 28432 21416 28484
rect 21548 28475 21600 28484
rect 21548 28441 21557 28475
rect 21557 28441 21591 28475
rect 21591 28441 21600 28475
rect 21548 28432 21600 28441
rect 22560 28432 22612 28484
rect 24584 28636 24636 28688
rect 25780 28636 25832 28688
rect 25872 28679 25924 28688
rect 25872 28645 25881 28679
rect 25881 28645 25915 28679
rect 25915 28645 25924 28679
rect 25872 28636 25924 28645
rect 28908 28704 28960 28756
rect 29644 28704 29696 28756
rect 39120 28747 39172 28756
rect 39120 28713 39129 28747
rect 39129 28713 39163 28747
rect 39163 28713 39172 28747
rect 39120 28704 39172 28713
rect 24308 28500 24360 28552
rect 24676 28500 24728 28552
rect 23572 28432 23624 28484
rect 21640 28364 21692 28416
rect 21916 28364 21968 28416
rect 23020 28407 23072 28416
rect 23020 28373 23029 28407
rect 23029 28373 23063 28407
rect 23063 28373 23072 28407
rect 23020 28364 23072 28373
rect 23480 28364 23532 28416
rect 26608 28543 26660 28552
rect 26608 28509 26617 28543
rect 26617 28509 26651 28543
rect 26651 28509 26660 28543
rect 26608 28500 26660 28509
rect 27160 28543 27212 28552
rect 27160 28509 27169 28543
rect 27169 28509 27203 28543
rect 27203 28509 27212 28543
rect 27160 28500 27212 28509
rect 27620 28500 27672 28552
rect 28632 28543 28684 28552
rect 28632 28509 28641 28543
rect 28641 28509 28675 28543
rect 28675 28509 28684 28543
rect 28632 28500 28684 28509
rect 28540 28432 28592 28484
rect 34244 28636 34296 28688
rect 29000 28500 29052 28552
rect 29552 28543 29604 28552
rect 29552 28509 29561 28543
rect 29561 28509 29595 28543
rect 29595 28509 29604 28543
rect 38108 28568 38160 28620
rect 29552 28500 29604 28509
rect 29828 28500 29880 28552
rect 30196 28500 30248 28552
rect 29920 28432 29972 28484
rect 34060 28500 34112 28552
rect 37280 28543 37332 28552
rect 37280 28509 37289 28543
rect 37289 28509 37323 28543
rect 37323 28509 37332 28543
rect 37280 28500 37332 28509
rect 27712 28364 27764 28416
rect 28356 28364 28408 28416
rect 28724 28407 28776 28416
rect 28724 28373 28733 28407
rect 28733 28373 28767 28407
rect 28767 28373 28776 28407
rect 28724 28364 28776 28373
rect 30288 28407 30340 28416
rect 30288 28373 30297 28407
rect 30297 28373 30331 28407
rect 30331 28373 30340 28407
rect 30288 28364 30340 28373
rect 31760 28364 31812 28416
rect 33416 28364 33468 28416
rect 37924 28432 37976 28484
rect 38108 28432 38160 28484
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 8944 28203 8996 28212
rect 8944 28169 8953 28203
rect 8953 28169 8987 28203
rect 8987 28169 8996 28203
rect 8944 28160 8996 28169
rect 8300 28135 8352 28144
rect 8300 28101 8309 28135
rect 8309 28101 8343 28135
rect 8343 28101 8352 28135
rect 8300 28092 8352 28101
rect 8576 28092 8628 28144
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 4804 28024 4856 28076
rect 5356 28024 5408 28076
rect 8024 28067 8076 28076
rect 8024 28033 8033 28067
rect 8033 28033 8067 28067
rect 8067 28033 8076 28067
rect 8024 28024 8076 28033
rect 9128 28024 9180 28076
rect 10968 28160 11020 28212
rect 11060 28203 11112 28212
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 11336 28160 11388 28212
rect 3792 27956 3844 28008
rect 5540 27956 5592 28008
rect 8300 27956 8352 28008
rect 940 27888 992 27940
rect 8944 27888 8996 27940
rect 9496 27956 9548 28008
rect 10600 27999 10652 28008
rect 10600 27965 10609 27999
rect 10609 27965 10643 27999
rect 10643 27965 10652 27999
rect 10600 27956 10652 27965
rect 12532 28135 12584 28144
rect 12532 28101 12541 28135
rect 12541 28101 12575 28135
rect 12575 28101 12584 28135
rect 12532 28092 12584 28101
rect 12440 28067 12492 28076
rect 12440 28033 12447 28067
rect 12447 28033 12492 28067
rect 10876 27931 10928 27940
rect 10876 27897 10885 27931
rect 10885 27897 10919 27931
rect 10919 27897 10928 27931
rect 10876 27888 10928 27897
rect 11152 27956 11204 28008
rect 12440 28024 12492 28033
rect 18420 28160 18472 28212
rect 12532 27956 12584 28008
rect 13636 27956 13688 28008
rect 14832 28067 14884 28076
rect 14832 28033 14841 28067
rect 14841 28033 14875 28067
rect 14875 28033 14884 28067
rect 14832 28024 14884 28033
rect 14924 28067 14976 28076
rect 14924 28033 14933 28067
rect 14933 28033 14967 28067
rect 14967 28033 14976 28067
rect 14924 28024 14976 28033
rect 15660 28092 15712 28144
rect 15200 28024 15252 28076
rect 15476 28024 15528 28076
rect 13912 27888 13964 27940
rect 14556 27888 14608 27940
rect 14648 27931 14700 27940
rect 14648 27897 14657 27931
rect 14657 27897 14691 27931
rect 14691 27897 14700 27931
rect 14648 27888 14700 27897
rect 14832 27888 14884 27940
rect 17316 28024 17368 28076
rect 16120 27956 16172 28008
rect 17960 27999 18012 28008
rect 17960 27965 17969 27999
rect 17969 27965 18003 27999
rect 18003 27965 18012 27999
rect 17960 27956 18012 27965
rect 17592 27888 17644 27940
rect 18144 27999 18196 28008
rect 18144 27965 18153 27999
rect 18153 27965 18187 27999
rect 18187 27965 18196 27999
rect 18144 27956 18196 27965
rect 18880 28160 18932 28212
rect 19064 28160 19116 28212
rect 19524 28160 19576 28212
rect 20352 28160 20404 28212
rect 27160 28203 27212 28212
rect 27160 28169 27169 28203
rect 27169 28169 27203 28203
rect 27203 28169 27212 28203
rect 27160 28160 27212 28169
rect 27344 28160 27396 28212
rect 27804 28160 27856 28212
rect 18880 28067 18932 28076
rect 18880 28033 18889 28067
rect 18889 28033 18923 28067
rect 18923 28033 18932 28067
rect 18880 28024 18932 28033
rect 19248 28135 19300 28144
rect 19248 28101 19257 28135
rect 19257 28101 19291 28135
rect 19291 28101 19300 28135
rect 19248 28092 19300 28101
rect 22744 28092 22796 28144
rect 26608 28092 26660 28144
rect 19156 28067 19208 28076
rect 19156 28033 19165 28067
rect 19165 28033 19199 28067
rect 19199 28033 19208 28067
rect 19156 28024 19208 28033
rect 20444 28024 20496 28076
rect 20720 28024 20772 28076
rect 25044 28024 25096 28076
rect 25320 28024 25372 28076
rect 26148 28024 26200 28076
rect 26516 28024 26568 28076
rect 27436 28024 27488 28076
rect 27988 28092 28040 28144
rect 31944 28160 31996 28212
rect 32680 28203 32732 28212
rect 32680 28169 32689 28203
rect 32689 28169 32723 28203
rect 32723 28169 32732 28203
rect 32680 28160 32732 28169
rect 32864 28203 32916 28212
rect 32864 28169 32873 28203
rect 32873 28169 32907 28203
rect 32907 28169 32916 28203
rect 32864 28160 32916 28169
rect 33416 28203 33468 28212
rect 33416 28169 33425 28203
rect 33425 28169 33459 28203
rect 33459 28169 33468 28203
rect 33416 28160 33468 28169
rect 34060 28160 34112 28212
rect 34244 28160 34296 28212
rect 37280 28160 37332 28212
rect 27712 28024 27764 28076
rect 30840 28135 30892 28144
rect 30840 28101 30849 28135
rect 30849 28101 30883 28135
rect 30883 28101 30892 28135
rect 30840 28092 30892 28101
rect 31024 28135 31076 28144
rect 31024 28101 31033 28135
rect 31033 28101 31067 28135
rect 31067 28101 31076 28135
rect 31024 28092 31076 28101
rect 18420 27888 18472 27940
rect 20628 27956 20680 28008
rect 20904 27956 20956 28008
rect 21456 27956 21508 28008
rect 27620 27956 27672 28008
rect 29368 27956 29420 28008
rect 31116 28024 31168 28076
rect 32404 28024 32456 28076
rect 22652 27888 22704 27940
rect 26516 27888 26568 27940
rect 26608 27888 26660 27940
rect 28632 27888 28684 27940
rect 29552 27888 29604 27940
rect 29828 27888 29880 27940
rect 5172 27820 5224 27872
rect 11520 27820 11572 27872
rect 12900 27863 12952 27872
rect 12900 27829 12909 27863
rect 12909 27829 12943 27863
rect 12943 27829 12952 27863
rect 12900 27820 12952 27829
rect 13820 27820 13872 27872
rect 15752 27820 15804 27872
rect 15936 27820 15988 27872
rect 17776 27863 17828 27872
rect 17776 27829 17785 27863
rect 17785 27829 17819 27863
rect 17819 27829 17828 27863
rect 17776 27820 17828 27829
rect 18236 27820 18288 27872
rect 19294 27820 19346 27872
rect 21640 27820 21692 27872
rect 29276 27820 29328 27872
rect 30840 27888 30892 27940
rect 31944 27999 31996 28008
rect 31944 27965 31953 27999
rect 31953 27965 31987 27999
rect 31987 27965 31996 27999
rect 31944 27956 31996 27965
rect 32036 27956 32088 28008
rect 32772 28024 32824 28076
rect 30196 27863 30248 27872
rect 30196 27829 30205 27863
rect 30205 27829 30239 27863
rect 30239 27829 30248 27863
rect 30196 27820 30248 27829
rect 30380 27820 30432 27872
rect 31760 27820 31812 27872
rect 33876 28024 33928 28076
rect 33968 28067 34020 28076
rect 33968 28033 33977 28067
rect 33977 28033 34011 28067
rect 34011 28033 34020 28067
rect 33968 28024 34020 28033
rect 34428 28092 34480 28144
rect 33600 27956 33652 28008
rect 35164 28024 35216 28076
rect 35716 28024 35768 28076
rect 35440 27956 35492 28008
rect 39120 28024 39172 28076
rect 36820 27888 36872 27940
rect 34336 27863 34388 27872
rect 34336 27829 34345 27863
rect 34345 27829 34379 27863
rect 34379 27829 34388 27863
rect 34336 27820 34388 27829
rect 35532 27863 35584 27872
rect 35532 27829 35541 27863
rect 35541 27829 35575 27863
rect 35575 27829 35584 27863
rect 35532 27820 35584 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 5632 27616 5684 27668
rect 9036 27616 9088 27668
rect 10232 27616 10284 27668
rect 11888 27616 11940 27668
rect 12256 27659 12308 27668
rect 12256 27625 12265 27659
rect 12265 27625 12299 27659
rect 12299 27625 12308 27659
rect 12256 27616 12308 27625
rect 12532 27616 12584 27668
rect 6092 27548 6144 27600
rect 6736 27548 6788 27600
rect 8944 27548 8996 27600
rect 9220 27548 9272 27600
rect 12440 27548 12492 27600
rect 13176 27616 13228 27668
rect 13268 27548 13320 27600
rect 14924 27616 14976 27668
rect 15108 27616 15160 27668
rect 14648 27548 14700 27600
rect 15384 27548 15436 27600
rect 6184 27480 6236 27532
rect 3792 27455 3844 27464
rect 3792 27421 3801 27455
rect 3801 27421 3835 27455
rect 3835 27421 3844 27455
rect 3792 27412 3844 27421
rect 5448 27412 5500 27464
rect 6276 27412 6328 27464
rect 8484 27480 8536 27532
rect 6460 27412 6512 27464
rect 6736 27455 6788 27464
rect 6736 27421 6745 27455
rect 6745 27421 6779 27455
rect 6779 27421 6788 27455
rect 6736 27412 6788 27421
rect 8852 27412 8904 27464
rect 9404 27480 9456 27532
rect 9496 27480 9548 27532
rect 9588 27412 9640 27464
rect 9772 27412 9824 27464
rect 4068 27387 4120 27396
rect 4068 27353 4077 27387
rect 4077 27353 4111 27387
rect 4111 27353 4120 27387
rect 4068 27344 4120 27353
rect 6828 27344 6880 27396
rect 10048 27412 10100 27464
rect 6276 27319 6328 27328
rect 6276 27285 6285 27319
rect 6285 27285 6319 27319
rect 6319 27285 6328 27319
rect 6276 27276 6328 27285
rect 6920 27319 6972 27328
rect 6920 27285 6929 27319
rect 6929 27285 6963 27319
rect 6963 27285 6972 27319
rect 6920 27276 6972 27285
rect 9496 27319 9548 27328
rect 9496 27285 9505 27319
rect 9505 27285 9539 27319
rect 9539 27285 9548 27319
rect 9496 27276 9548 27285
rect 10784 27344 10836 27396
rect 10600 27276 10652 27328
rect 12164 27344 12216 27396
rect 12532 27344 12584 27396
rect 13176 27344 13228 27396
rect 13268 27387 13320 27396
rect 13268 27353 13277 27387
rect 13277 27353 13311 27387
rect 13311 27353 13320 27387
rect 13268 27344 13320 27353
rect 13452 27387 13504 27396
rect 13452 27353 13461 27387
rect 13461 27353 13495 27387
rect 13495 27353 13504 27387
rect 13452 27344 13504 27353
rect 13728 27344 13780 27396
rect 14096 27480 14148 27532
rect 17132 27616 17184 27668
rect 17592 27616 17644 27668
rect 18512 27616 18564 27668
rect 18972 27616 19024 27668
rect 15752 27548 15804 27600
rect 14464 27455 14516 27464
rect 14464 27421 14473 27455
rect 14473 27421 14507 27455
rect 14507 27421 14516 27455
rect 14464 27412 14516 27421
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 14832 27412 14884 27464
rect 15200 27455 15252 27464
rect 15200 27421 15209 27455
rect 15209 27421 15243 27455
rect 15243 27421 15252 27455
rect 15200 27412 15252 27421
rect 16672 27480 16724 27532
rect 20628 27548 20680 27600
rect 13912 27276 13964 27328
rect 14556 27276 14608 27328
rect 16028 27344 16080 27396
rect 16948 27455 17000 27464
rect 16948 27421 16957 27455
rect 16957 27421 16991 27455
rect 16991 27421 17000 27455
rect 16948 27412 17000 27421
rect 17316 27412 17368 27464
rect 17960 27412 18012 27464
rect 18512 27455 18564 27464
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 20812 27480 20864 27532
rect 20996 27480 21048 27532
rect 23204 27616 23256 27668
rect 21364 27548 21416 27600
rect 21088 27455 21140 27464
rect 16764 27344 16816 27396
rect 18236 27344 18288 27396
rect 21088 27421 21097 27455
rect 21097 27421 21131 27455
rect 21131 27421 21140 27455
rect 21088 27412 21140 27421
rect 21272 27412 21324 27464
rect 21364 27455 21416 27464
rect 21364 27421 21373 27455
rect 21373 27421 21407 27455
rect 21407 27421 21416 27455
rect 21364 27412 21416 27421
rect 22928 27548 22980 27600
rect 25412 27616 25464 27668
rect 23756 27548 23808 27600
rect 18972 27344 19024 27396
rect 19432 27344 19484 27396
rect 20628 27344 20680 27396
rect 22376 27344 22428 27396
rect 22560 27455 22612 27464
rect 22560 27421 22569 27455
rect 22569 27421 22603 27455
rect 22603 27421 22612 27455
rect 22560 27412 22612 27421
rect 23296 27412 23348 27464
rect 23572 27412 23624 27464
rect 27712 27548 27764 27600
rect 27896 27616 27948 27668
rect 29000 27616 29052 27668
rect 27988 27548 28040 27600
rect 24676 27412 24728 27464
rect 15752 27276 15804 27328
rect 15844 27276 15896 27328
rect 16304 27319 16356 27328
rect 16304 27285 16313 27319
rect 16313 27285 16347 27319
rect 16347 27285 16356 27319
rect 16304 27276 16356 27285
rect 16488 27276 16540 27328
rect 17132 27319 17184 27328
rect 17132 27285 17141 27319
rect 17141 27285 17175 27319
rect 17175 27285 17184 27319
rect 17132 27276 17184 27285
rect 18144 27276 18196 27328
rect 22284 27276 22336 27328
rect 22652 27319 22704 27328
rect 22652 27285 22661 27319
rect 22661 27285 22695 27319
rect 22695 27285 22704 27319
rect 22652 27276 22704 27285
rect 23388 27344 23440 27396
rect 25412 27412 25464 27464
rect 25504 27455 25556 27464
rect 25504 27421 25513 27455
rect 25513 27421 25547 27455
rect 25547 27421 25556 27455
rect 25504 27412 25556 27421
rect 25964 27455 26016 27464
rect 25964 27421 25973 27455
rect 25973 27421 26007 27455
rect 26007 27421 26016 27455
rect 25964 27412 26016 27421
rect 26424 27412 26476 27464
rect 26608 27455 26660 27464
rect 26608 27421 26617 27455
rect 26617 27421 26651 27455
rect 26651 27421 26660 27455
rect 26608 27412 26660 27421
rect 26884 27480 26936 27532
rect 29276 27480 29328 27532
rect 29552 27480 29604 27532
rect 30380 27616 30432 27668
rect 30840 27616 30892 27668
rect 31116 27659 31168 27668
rect 31116 27625 31125 27659
rect 31125 27625 31159 27659
rect 31159 27625 31168 27659
rect 31116 27616 31168 27625
rect 32680 27616 32732 27668
rect 35532 27616 35584 27668
rect 27344 27412 27396 27464
rect 27528 27455 27580 27464
rect 27528 27421 27537 27455
rect 27537 27421 27571 27455
rect 27571 27421 27580 27455
rect 27528 27412 27580 27421
rect 28540 27412 28592 27464
rect 28816 27412 28868 27464
rect 29000 27455 29052 27464
rect 29000 27421 29009 27455
rect 29009 27421 29043 27455
rect 29043 27421 29052 27455
rect 29000 27412 29052 27421
rect 24032 27276 24084 27328
rect 24216 27276 24268 27328
rect 27896 27344 27948 27396
rect 28356 27344 28408 27396
rect 29644 27412 29696 27464
rect 31760 27480 31812 27532
rect 32404 27480 32456 27532
rect 34796 27523 34848 27532
rect 34796 27489 34805 27523
rect 34805 27489 34839 27523
rect 34839 27489 34848 27523
rect 34796 27480 34848 27489
rect 35808 27480 35860 27532
rect 36820 27523 36872 27532
rect 36820 27489 36829 27523
rect 36829 27489 36863 27523
rect 36863 27489 36872 27523
rect 36820 27480 36872 27489
rect 34336 27412 34388 27464
rect 30104 27344 30156 27396
rect 25780 27276 25832 27328
rect 26148 27276 26200 27328
rect 28724 27276 28776 27328
rect 29368 27276 29420 27328
rect 29552 27276 29604 27328
rect 30564 27319 30616 27328
rect 30564 27285 30573 27319
rect 30573 27285 30607 27319
rect 30607 27285 30616 27319
rect 30564 27276 30616 27285
rect 31300 27319 31352 27328
rect 31300 27285 31309 27319
rect 31309 27285 31343 27319
rect 31343 27285 31352 27319
rect 31300 27276 31352 27285
rect 33508 27276 33560 27328
rect 35440 27276 35492 27328
rect 38108 27276 38160 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4068 27072 4120 27124
rect 6276 27072 6328 27124
rect 6920 27072 6972 27124
rect 7288 27004 7340 27056
rect 8208 27004 8260 27056
rect 11612 27072 11664 27124
rect 11704 27072 11756 27124
rect 11888 27072 11940 27124
rect 5540 26936 5592 26988
rect 8852 27004 8904 27056
rect 9404 27004 9456 27056
rect 9496 27004 9548 27056
rect 9036 26979 9088 26988
rect 9036 26945 9045 26979
rect 9045 26945 9079 26979
rect 9079 26945 9088 26979
rect 9036 26936 9088 26945
rect 10140 27004 10192 27056
rect 10876 27004 10928 27056
rect 9772 26979 9824 26988
rect 9772 26945 9781 26979
rect 9781 26945 9815 26979
rect 9815 26945 9824 26979
rect 9772 26936 9824 26945
rect 9864 26936 9916 26988
rect 4988 26911 5040 26920
rect 4988 26877 4997 26911
rect 4997 26877 5031 26911
rect 5031 26877 5040 26911
rect 4988 26868 5040 26877
rect 5172 26911 5224 26920
rect 5172 26877 5181 26911
rect 5181 26877 5215 26911
rect 5215 26877 5224 26911
rect 5172 26868 5224 26877
rect 10140 26868 10192 26920
rect 10232 26868 10284 26920
rect 9956 26800 10008 26852
rect 8300 26732 8352 26784
rect 8852 26775 8904 26784
rect 8852 26741 8861 26775
rect 8861 26741 8895 26775
rect 8895 26741 8904 26775
rect 8852 26732 8904 26741
rect 9680 26732 9732 26784
rect 9772 26732 9824 26784
rect 12072 26979 12124 26988
rect 12072 26945 12081 26979
rect 12081 26945 12115 26979
rect 12115 26945 12124 26979
rect 12072 26936 12124 26945
rect 12440 27072 12492 27124
rect 12716 27047 12768 27056
rect 12716 27013 12725 27047
rect 12725 27013 12759 27047
rect 12759 27013 12768 27047
rect 12716 27004 12768 27013
rect 12900 27115 12952 27124
rect 12900 27081 12925 27115
rect 12925 27081 12952 27115
rect 12900 27072 12952 27081
rect 14372 27072 14424 27124
rect 16396 27072 16448 27124
rect 13084 27004 13136 27056
rect 15108 27004 15160 27056
rect 17040 27004 17092 27056
rect 18604 27072 18656 27124
rect 20628 27072 20680 27124
rect 21272 27072 21324 27124
rect 10784 26868 10836 26920
rect 13452 26868 13504 26920
rect 14004 26868 14056 26920
rect 14648 26868 14700 26920
rect 15844 26936 15896 26988
rect 16304 26979 16356 26988
rect 16304 26945 16313 26979
rect 16313 26945 16347 26979
rect 16347 26945 16356 26979
rect 16304 26936 16356 26945
rect 18144 27004 18196 27056
rect 18236 27004 18288 27056
rect 19984 27004 20036 27056
rect 12164 26800 12216 26852
rect 11244 26732 11296 26784
rect 11980 26775 12032 26784
rect 11980 26741 11989 26775
rect 11989 26741 12023 26775
rect 12023 26741 12032 26775
rect 11980 26732 12032 26741
rect 12532 26800 12584 26852
rect 15016 26868 15068 26920
rect 18788 26936 18840 26988
rect 19340 26936 19392 26988
rect 13084 26775 13136 26784
rect 13084 26741 13093 26775
rect 13093 26741 13127 26775
rect 13127 26741 13136 26775
rect 13084 26732 13136 26741
rect 13268 26732 13320 26784
rect 14280 26732 14332 26784
rect 14740 26732 14792 26784
rect 15936 26800 15988 26852
rect 17132 26800 17184 26852
rect 16764 26775 16816 26784
rect 16764 26741 16773 26775
rect 16773 26741 16807 26775
rect 16807 26741 16816 26775
rect 16764 26732 16816 26741
rect 17500 26775 17552 26784
rect 17500 26741 17509 26775
rect 17509 26741 17543 26775
rect 17543 26741 17552 26775
rect 17500 26732 17552 26741
rect 20536 26936 20588 26988
rect 20720 26936 20772 26988
rect 21272 26936 21324 26988
rect 25136 27072 25188 27124
rect 21548 26936 21600 26988
rect 22744 26936 22796 26988
rect 22928 26936 22980 26988
rect 23204 26979 23256 26988
rect 23204 26945 23213 26979
rect 23213 26945 23247 26979
rect 23247 26945 23256 26979
rect 23204 26936 23256 26945
rect 24400 26979 24452 26988
rect 24400 26945 24409 26979
rect 24409 26945 24443 26979
rect 24443 26945 24452 26979
rect 24400 26936 24452 26945
rect 24952 26979 25004 26988
rect 24952 26945 24961 26979
rect 24961 26945 24995 26979
rect 24995 26945 25004 26979
rect 24952 26936 25004 26945
rect 25136 26979 25188 26988
rect 25136 26945 25145 26979
rect 25145 26945 25179 26979
rect 25179 26945 25188 26979
rect 25136 26936 25188 26945
rect 25504 27072 25556 27124
rect 25688 27072 25740 27124
rect 26516 27072 26568 27124
rect 28264 27072 28316 27124
rect 28816 27072 28868 27124
rect 29000 27072 29052 27124
rect 30196 27072 30248 27124
rect 25688 26979 25740 26988
rect 25688 26945 25697 26979
rect 25697 26945 25731 26979
rect 25731 26945 25740 26979
rect 25688 26936 25740 26945
rect 27252 26936 27304 26988
rect 27344 26936 27396 26988
rect 18604 26800 18656 26852
rect 18788 26732 18840 26784
rect 19064 26732 19116 26784
rect 23388 26800 23440 26852
rect 23756 26911 23808 26920
rect 23756 26877 23765 26911
rect 23765 26877 23799 26911
rect 23799 26877 23808 26911
rect 23756 26868 23808 26877
rect 24124 26800 24176 26852
rect 24584 26843 24636 26852
rect 24584 26809 24593 26843
rect 24593 26809 24627 26843
rect 24627 26809 24636 26843
rect 24584 26800 24636 26809
rect 24676 26843 24728 26852
rect 24676 26809 24685 26843
rect 24685 26809 24719 26843
rect 24719 26809 24728 26843
rect 24676 26800 24728 26809
rect 24860 26911 24912 26920
rect 24860 26877 24869 26911
rect 24869 26877 24903 26911
rect 24903 26877 24912 26911
rect 25964 26911 26016 26920
rect 24860 26868 24912 26877
rect 25964 26877 25973 26911
rect 25973 26877 26007 26911
rect 26007 26877 26016 26911
rect 25964 26868 26016 26877
rect 26976 26911 27028 26920
rect 26976 26877 26985 26911
rect 26985 26877 27019 26911
rect 27019 26877 27028 26911
rect 26976 26868 27028 26877
rect 27436 26868 27488 26920
rect 27712 26979 27764 26988
rect 27712 26945 27721 26979
rect 27721 26945 27755 26979
rect 27755 26945 27764 26979
rect 27712 26936 27764 26945
rect 28172 26936 28224 26988
rect 28356 26936 28408 26988
rect 28540 26979 28592 26988
rect 28540 26945 28549 26979
rect 28549 26945 28583 26979
rect 28583 26945 28592 26979
rect 28540 26936 28592 26945
rect 28724 26936 28776 26988
rect 32864 27004 32916 27056
rect 25872 26843 25924 26852
rect 25872 26809 25881 26843
rect 25881 26809 25915 26843
rect 25915 26809 25924 26843
rect 25872 26800 25924 26809
rect 26240 26800 26292 26852
rect 29828 26936 29880 26988
rect 30564 26936 30616 26988
rect 31300 26936 31352 26988
rect 33508 27072 33560 27124
rect 33324 27047 33376 27056
rect 33324 27013 33333 27047
rect 33333 27013 33367 27047
rect 33367 27013 33376 27047
rect 33324 27004 33376 27013
rect 33600 27004 33652 27056
rect 33140 26936 33192 26988
rect 33508 26936 33560 26988
rect 34796 27072 34848 27124
rect 35440 27004 35492 27056
rect 28356 26843 28408 26852
rect 28356 26809 28365 26843
rect 28365 26809 28399 26843
rect 28399 26809 28408 26843
rect 28356 26800 28408 26809
rect 29000 26800 29052 26852
rect 19432 26732 19484 26784
rect 20168 26732 20220 26784
rect 20628 26732 20680 26784
rect 20996 26732 21048 26784
rect 21272 26775 21324 26784
rect 21272 26741 21281 26775
rect 21281 26741 21315 26775
rect 21315 26741 21324 26775
rect 21272 26732 21324 26741
rect 22008 26732 22060 26784
rect 23204 26732 23256 26784
rect 24952 26732 25004 26784
rect 25780 26732 25832 26784
rect 26148 26732 26200 26784
rect 28540 26732 28592 26784
rect 29552 26868 29604 26920
rect 30104 26800 30156 26852
rect 29644 26732 29696 26784
rect 30012 26775 30064 26784
rect 30012 26741 30021 26775
rect 30021 26741 30055 26775
rect 30055 26741 30064 26775
rect 30012 26732 30064 26741
rect 31024 26800 31076 26852
rect 34336 26868 34388 26920
rect 32588 26732 32640 26784
rect 34428 26732 34480 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 6828 26528 6880 26580
rect 13268 26528 13320 26580
rect 14096 26528 14148 26580
rect 16304 26528 16356 26580
rect 16764 26528 16816 26580
rect 1676 26324 1728 26376
rect 9496 26460 9548 26512
rect 11060 26460 11112 26512
rect 6736 26392 6788 26444
rect 8392 26392 8444 26444
rect 8208 26324 8260 26376
rect 9772 26392 9824 26444
rect 9220 26367 9272 26376
rect 9220 26333 9229 26367
rect 9229 26333 9263 26367
rect 9263 26333 9272 26367
rect 9220 26324 9272 26333
rect 9404 26367 9456 26376
rect 9404 26333 9439 26367
rect 9439 26333 9456 26367
rect 10600 26392 10652 26444
rect 9404 26324 9456 26333
rect 9956 26324 10008 26376
rect 10692 26367 10744 26376
rect 10692 26333 10701 26367
rect 10701 26333 10735 26367
rect 10735 26333 10744 26367
rect 10692 26324 10744 26333
rect 11704 26392 11756 26444
rect 15200 26392 15252 26444
rect 15384 26435 15436 26444
rect 15384 26401 15393 26435
rect 15393 26401 15427 26435
rect 15427 26401 15436 26435
rect 15384 26392 15436 26401
rect 15844 26392 15896 26444
rect 16028 26392 16080 26444
rect 6920 26256 6972 26308
rect 8668 26256 8720 26308
rect 5080 26231 5132 26240
rect 5080 26197 5089 26231
rect 5089 26197 5123 26231
rect 5123 26197 5132 26231
rect 5080 26188 5132 26197
rect 6552 26188 6604 26240
rect 8484 26188 8536 26240
rect 10232 26256 10284 26308
rect 10508 26299 10560 26308
rect 10508 26265 10517 26299
rect 10517 26265 10551 26299
rect 10551 26265 10560 26299
rect 10508 26256 10560 26265
rect 10968 26256 11020 26308
rect 14924 26324 14976 26376
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 12164 26256 12216 26308
rect 14280 26256 14332 26308
rect 16488 26324 16540 26376
rect 16948 26392 17000 26444
rect 18604 26392 18656 26444
rect 17132 26324 17184 26376
rect 17408 26324 17460 26376
rect 17960 26367 18012 26376
rect 17960 26333 17969 26367
rect 17969 26333 18003 26367
rect 18003 26333 18012 26367
rect 17960 26324 18012 26333
rect 19064 26460 19116 26512
rect 22652 26528 22704 26580
rect 23296 26528 23348 26580
rect 17868 26256 17920 26308
rect 18236 26256 18288 26308
rect 19156 26256 19208 26308
rect 15292 26188 15344 26240
rect 15476 26188 15528 26240
rect 15844 26188 15896 26240
rect 17040 26188 17092 26240
rect 18052 26188 18104 26240
rect 19064 26188 19116 26240
rect 19524 26324 19576 26376
rect 19984 26324 20036 26376
rect 20812 26392 20864 26444
rect 21364 26460 21416 26512
rect 22744 26460 22796 26512
rect 22928 26460 22980 26512
rect 20352 26256 20404 26308
rect 21180 26324 21232 26376
rect 22284 26324 22336 26376
rect 23848 26460 23900 26512
rect 24676 26460 24728 26512
rect 23572 26392 23624 26444
rect 25688 26528 25740 26580
rect 25872 26528 25924 26580
rect 27344 26528 27396 26580
rect 27436 26528 27488 26580
rect 29000 26528 29052 26580
rect 32128 26528 32180 26580
rect 33140 26571 33192 26580
rect 33140 26537 33149 26571
rect 33149 26537 33183 26571
rect 33183 26537 33192 26571
rect 33140 26528 33192 26537
rect 19340 26231 19392 26240
rect 19340 26197 19349 26231
rect 19349 26197 19383 26231
rect 19383 26197 19392 26231
rect 19340 26188 19392 26197
rect 19984 26188 20036 26240
rect 20444 26231 20496 26240
rect 20444 26197 20453 26231
rect 20453 26197 20487 26231
rect 20487 26197 20496 26231
rect 20444 26188 20496 26197
rect 25504 26392 25556 26444
rect 25964 26460 26016 26512
rect 26516 26503 26568 26512
rect 26516 26469 26525 26503
rect 26525 26469 26559 26503
rect 26559 26469 26568 26503
rect 26516 26460 26568 26469
rect 24952 26367 25004 26376
rect 24952 26333 24961 26367
rect 24961 26333 24995 26367
rect 24995 26333 25004 26367
rect 24952 26324 25004 26333
rect 25780 26367 25832 26376
rect 25780 26333 25789 26367
rect 25789 26333 25823 26367
rect 25823 26333 25832 26367
rect 25780 26324 25832 26333
rect 25872 26367 25924 26376
rect 25872 26333 25881 26367
rect 25881 26333 25915 26367
rect 25915 26333 25924 26367
rect 25872 26324 25924 26333
rect 26148 26367 26200 26376
rect 26148 26333 26157 26367
rect 26157 26333 26191 26367
rect 26191 26333 26200 26367
rect 26148 26324 26200 26333
rect 26516 26324 26568 26376
rect 26976 26324 27028 26376
rect 27068 26324 27120 26376
rect 28172 26460 28224 26512
rect 31760 26460 31812 26512
rect 30472 26392 30524 26444
rect 32496 26460 32548 26512
rect 33232 26503 33284 26512
rect 33232 26469 33241 26503
rect 33241 26469 33275 26503
rect 33275 26469 33284 26503
rect 33232 26460 33284 26469
rect 24308 26188 24360 26240
rect 24492 26231 24544 26240
rect 24492 26197 24501 26231
rect 24501 26197 24535 26231
rect 24535 26197 24544 26231
rect 24492 26188 24544 26197
rect 26424 26188 26476 26240
rect 26608 26188 26660 26240
rect 28356 26188 28408 26240
rect 32220 26324 32272 26376
rect 34612 26324 34664 26376
rect 39672 26392 39724 26444
rect 35808 26367 35860 26376
rect 35808 26333 35817 26367
rect 35817 26333 35851 26367
rect 35851 26333 35860 26367
rect 35808 26324 35860 26333
rect 31944 26256 31996 26308
rect 32404 26299 32456 26308
rect 32404 26265 32413 26299
rect 32413 26265 32447 26299
rect 32447 26265 32456 26299
rect 32404 26256 32456 26265
rect 32680 26231 32732 26240
rect 32680 26197 32689 26231
rect 32689 26197 32723 26231
rect 32723 26197 32732 26231
rect 32680 26188 32732 26197
rect 33324 26188 33376 26240
rect 34336 26188 34388 26240
rect 36084 26231 36136 26240
rect 36084 26197 36093 26231
rect 36093 26197 36127 26231
rect 36127 26197 36136 26231
rect 36084 26188 36136 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5080 25984 5132 26036
rect 6920 25984 6972 26036
rect 8484 25984 8536 26036
rect 8760 25984 8812 26036
rect 5448 25916 5500 25968
rect 8024 25916 8076 25968
rect 8576 25848 8628 25900
rect 8760 25891 8812 25900
rect 8760 25857 8769 25891
rect 8769 25857 8803 25891
rect 8803 25857 8812 25891
rect 8760 25848 8812 25857
rect 8852 25891 8904 25900
rect 8852 25857 8861 25891
rect 8861 25857 8895 25891
rect 8895 25857 8904 25891
rect 8852 25848 8904 25857
rect 3792 25780 3844 25832
rect 6552 25780 6604 25832
rect 9680 25916 9732 25968
rect 9404 25891 9456 25900
rect 9404 25857 9413 25891
rect 9413 25857 9447 25891
rect 9447 25857 9456 25891
rect 9404 25848 9456 25857
rect 10048 25959 10100 25968
rect 10048 25925 10057 25959
rect 10057 25925 10091 25959
rect 10091 25925 10100 25959
rect 10048 25916 10100 25925
rect 9956 25891 10008 25900
rect 9956 25857 9963 25891
rect 9963 25857 10008 25891
rect 9956 25848 10008 25857
rect 11060 25984 11112 26036
rect 11428 25984 11480 26036
rect 13176 25984 13228 26036
rect 14464 25984 14516 26036
rect 13084 25916 13136 25968
rect 14096 25916 14148 25968
rect 16120 25916 16172 25968
rect 9588 25780 9640 25832
rect 7288 25687 7340 25696
rect 7288 25653 7297 25687
rect 7297 25653 7331 25687
rect 7331 25653 7340 25687
rect 7288 25644 7340 25653
rect 9956 25712 10008 25764
rect 9220 25687 9272 25696
rect 9220 25653 9229 25687
rect 9229 25653 9263 25687
rect 9263 25653 9272 25687
rect 9220 25644 9272 25653
rect 9312 25644 9364 25696
rect 9588 25687 9640 25696
rect 9588 25653 9597 25687
rect 9597 25653 9631 25687
rect 9631 25653 9640 25687
rect 11152 25848 11204 25900
rect 12992 25848 13044 25900
rect 13544 25848 13596 25900
rect 14924 25848 14976 25900
rect 15568 25848 15620 25900
rect 15660 25848 15712 25900
rect 11244 25780 11296 25832
rect 12716 25780 12768 25832
rect 12900 25780 12952 25832
rect 13268 25780 13320 25832
rect 14556 25780 14608 25832
rect 15108 25780 15160 25832
rect 15844 25780 15896 25832
rect 16856 25848 16908 25900
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 17316 25916 17368 25968
rect 18880 25916 18932 25968
rect 19892 25984 19944 26036
rect 21548 25984 21600 26036
rect 17960 25848 18012 25900
rect 18328 25891 18380 25900
rect 18328 25857 18337 25891
rect 18337 25857 18371 25891
rect 18371 25857 18380 25891
rect 18328 25848 18380 25857
rect 20444 25916 20496 25968
rect 20536 25916 20588 25968
rect 17592 25780 17644 25832
rect 17868 25780 17920 25832
rect 12164 25712 12216 25764
rect 17040 25712 17092 25764
rect 17316 25712 17368 25764
rect 19340 25780 19392 25832
rect 19984 25891 20036 25900
rect 19984 25857 19993 25891
rect 19993 25857 20027 25891
rect 20027 25857 20036 25891
rect 19984 25848 20036 25857
rect 25044 25916 25096 25968
rect 20628 25848 20680 25900
rect 20720 25848 20772 25900
rect 20904 25848 20956 25900
rect 21732 25848 21784 25900
rect 24584 25848 24636 25900
rect 27344 25984 27396 26036
rect 26056 25916 26108 25968
rect 26976 25916 27028 25968
rect 21364 25780 21416 25832
rect 25320 25891 25372 25900
rect 25320 25857 25334 25891
rect 25334 25857 25368 25891
rect 25368 25857 25372 25891
rect 25320 25848 25372 25857
rect 25872 25848 25924 25900
rect 26332 25891 26384 25900
rect 26332 25857 26341 25891
rect 26341 25857 26375 25891
rect 26375 25857 26384 25891
rect 26332 25848 26384 25857
rect 26424 25891 26476 25900
rect 26424 25857 26433 25891
rect 26433 25857 26467 25891
rect 26467 25857 26476 25891
rect 26424 25848 26476 25857
rect 9588 25644 9640 25653
rect 10416 25687 10468 25696
rect 10416 25653 10425 25687
rect 10425 25653 10459 25687
rect 10459 25653 10468 25687
rect 10416 25644 10468 25653
rect 10876 25644 10928 25696
rect 12440 25644 12492 25696
rect 12900 25687 12952 25696
rect 12900 25653 12909 25687
rect 12909 25653 12943 25687
rect 12943 25653 12952 25687
rect 12900 25644 12952 25653
rect 12992 25687 13044 25696
rect 12992 25653 13001 25687
rect 13001 25653 13035 25687
rect 13035 25653 13044 25687
rect 12992 25644 13044 25653
rect 14372 25644 14424 25696
rect 14924 25644 14976 25696
rect 18052 25687 18104 25696
rect 18052 25653 18061 25687
rect 18061 25653 18095 25687
rect 18095 25653 18104 25687
rect 18052 25644 18104 25653
rect 20444 25712 20496 25764
rect 22744 25712 22796 25764
rect 25688 25823 25740 25832
rect 25688 25789 25697 25823
rect 25697 25789 25731 25823
rect 25731 25789 25740 25823
rect 25688 25780 25740 25789
rect 26148 25823 26200 25832
rect 26148 25789 26157 25823
rect 26157 25789 26191 25823
rect 26191 25789 26200 25823
rect 26148 25780 26200 25789
rect 25504 25755 25556 25764
rect 25504 25721 25513 25755
rect 25513 25721 25547 25755
rect 25547 25721 25556 25755
rect 26700 25848 26752 25900
rect 27620 25916 27672 25968
rect 27528 25891 27580 25900
rect 27528 25857 27537 25891
rect 27537 25857 27571 25891
rect 27571 25857 27580 25891
rect 27528 25848 27580 25857
rect 26976 25780 27028 25832
rect 27344 25823 27396 25832
rect 27344 25789 27353 25823
rect 27353 25789 27387 25823
rect 27387 25789 27396 25823
rect 27344 25780 27396 25789
rect 27804 25780 27856 25832
rect 30380 25848 30432 25900
rect 30564 25891 30616 25900
rect 30564 25857 30573 25891
rect 30573 25857 30607 25891
rect 30607 25857 30616 25891
rect 30564 25848 30616 25857
rect 30932 25891 30984 25900
rect 30932 25857 30941 25891
rect 30941 25857 30975 25891
rect 30975 25857 30984 25891
rect 30932 25848 30984 25857
rect 31668 25984 31720 26036
rect 31944 26027 31996 26036
rect 31944 25993 31953 26027
rect 31953 25993 31987 26027
rect 31987 25993 31996 26027
rect 31944 25984 31996 25993
rect 32496 25984 32548 26036
rect 34888 25984 34940 26036
rect 36084 25984 36136 26036
rect 36268 25916 36320 25968
rect 29552 25780 29604 25832
rect 31760 25780 31812 25832
rect 31944 25780 31996 25832
rect 33232 25848 33284 25900
rect 33508 25891 33560 25900
rect 33508 25857 33517 25891
rect 33517 25857 33551 25891
rect 33551 25857 33560 25891
rect 33508 25848 33560 25857
rect 35532 25848 35584 25900
rect 25504 25712 25556 25721
rect 20904 25644 20956 25696
rect 24584 25644 24636 25696
rect 27160 25687 27212 25696
rect 27160 25653 27169 25687
rect 27169 25653 27203 25687
rect 27203 25653 27212 25687
rect 27160 25644 27212 25653
rect 28172 25644 28224 25696
rect 28724 25687 28776 25696
rect 28724 25653 28733 25687
rect 28733 25653 28767 25687
rect 28767 25653 28776 25687
rect 28724 25644 28776 25653
rect 32404 25712 32456 25764
rect 34428 25780 34480 25832
rect 33324 25712 33376 25764
rect 34888 25712 34940 25764
rect 35808 25712 35860 25764
rect 36820 25712 36872 25764
rect 34612 25644 34664 25696
rect 36084 25687 36136 25696
rect 36084 25653 36093 25687
rect 36093 25653 36127 25687
rect 36127 25653 36136 25687
rect 36084 25644 36136 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 4712 25440 4764 25492
rect 6552 25440 6604 25492
rect 7288 25440 7340 25492
rect 3792 25347 3844 25356
rect 3792 25313 3801 25347
rect 3801 25313 3835 25347
rect 3835 25313 3844 25347
rect 3792 25304 3844 25313
rect 5448 25236 5500 25288
rect 4068 25211 4120 25220
rect 4068 25177 4077 25211
rect 4077 25177 4111 25211
rect 4111 25177 4120 25211
rect 4068 25168 4120 25177
rect 6828 25279 6880 25288
rect 6828 25245 6837 25279
rect 6837 25245 6871 25279
rect 6871 25245 6880 25279
rect 6828 25236 6880 25245
rect 8760 25440 8812 25492
rect 9772 25440 9824 25492
rect 9036 25372 9088 25424
rect 9588 25372 9640 25424
rect 8208 25304 8260 25356
rect 8024 25236 8076 25288
rect 8116 25279 8168 25288
rect 8116 25245 8125 25279
rect 8125 25245 8159 25279
rect 8159 25245 8168 25279
rect 8116 25236 8168 25245
rect 9128 25304 9180 25356
rect 9220 25304 9272 25356
rect 8484 25236 8536 25288
rect 8392 25168 8444 25220
rect 9036 25168 9088 25220
rect 6368 25143 6420 25152
rect 6368 25109 6377 25143
rect 6377 25109 6411 25143
rect 6411 25109 6420 25143
rect 6368 25100 6420 25109
rect 9404 25236 9456 25288
rect 9496 25236 9548 25288
rect 9680 25279 9732 25288
rect 9680 25245 9689 25279
rect 9689 25245 9723 25279
rect 9723 25245 9732 25279
rect 9680 25236 9732 25245
rect 11152 25279 11204 25288
rect 11152 25245 11161 25279
rect 11161 25245 11195 25279
rect 11195 25245 11204 25279
rect 11152 25236 11204 25245
rect 14924 25440 14976 25492
rect 15200 25440 15252 25492
rect 15568 25483 15620 25492
rect 15568 25449 15577 25483
rect 15577 25449 15611 25483
rect 15611 25449 15620 25483
rect 15568 25440 15620 25449
rect 15752 25440 15804 25492
rect 16580 25440 16632 25492
rect 16856 25440 16908 25492
rect 11520 25236 11572 25288
rect 11704 25236 11756 25288
rect 13360 25236 13412 25288
rect 15384 25304 15436 25356
rect 16764 25372 16816 25424
rect 20720 25440 20772 25492
rect 21180 25440 21232 25492
rect 15660 25347 15712 25356
rect 15660 25313 15669 25347
rect 15669 25313 15703 25347
rect 15703 25313 15712 25347
rect 15660 25304 15712 25313
rect 16028 25347 16080 25356
rect 16028 25313 16037 25347
rect 16037 25313 16071 25347
rect 16071 25313 16080 25347
rect 16028 25304 16080 25313
rect 16304 25304 16356 25356
rect 17040 25347 17092 25356
rect 17040 25313 17049 25347
rect 17049 25313 17083 25347
rect 17083 25313 17092 25347
rect 19248 25372 19300 25424
rect 20628 25372 20680 25424
rect 17040 25304 17092 25313
rect 17960 25347 18012 25356
rect 17960 25313 17969 25347
rect 17969 25313 18003 25347
rect 18003 25313 18012 25347
rect 17960 25304 18012 25313
rect 18052 25304 18104 25356
rect 19432 25304 19484 25356
rect 11888 25168 11940 25220
rect 14372 25168 14424 25220
rect 14832 25236 14884 25288
rect 15292 25236 15344 25288
rect 15844 25236 15896 25288
rect 15936 25236 15988 25288
rect 16764 25236 16816 25288
rect 16028 25168 16080 25220
rect 16488 25211 16540 25220
rect 16488 25177 16497 25211
rect 16497 25177 16531 25211
rect 16531 25177 16540 25211
rect 16488 25168 16540 25177
rect 16948 25279 17000 25288
rect 16948 25245 16957 25279
rect 16957 25245 16991 25279
rect 16991 25245 17000 25279
rect 16948 25236 17000 25245
rect 17408 25236 17460 25288
rect 18512 25236 18564 25288
rect 20904 25236 20956 25288
rect 21456 25304 21508 25356
rect 25504 25440 25556 25492
rect 25780 25440 25832 25492
rect 26516 25440 26568 25492
rect 27344 25440 27396 25492
rect 30656 25440 30708 25492
rect 32220 25440 32272 25492
rect 28172 25415 28224 25424
rect 28172 25381 28181 25415
rect 28181 25381 28215 25415
rect 28215 25381 28224 25415
rect 28172 25372 28224 25381
rect 9404 25100 9456 25152
rect 12256 25100 12308 25152
rect 12532 25100 12584 25152
rect 13452 25100 13504 25152
rect 13636 25100 13688 25152
rect 14280 25100 14332 25152
rect 14924 25100 14976 25152
rect 15568 25100 15620 25152
rect 15936 25143 15988 25152
rect 15936 25109 15945 25143
rect 15945 25109 15979 25143
rect 15979 25109 15988 25143
rect 15936 25100 15988 25109
rect 19432 25168 19484 25220
rect 19892 25168 19944 25220
rect 21364 25279 21416 25288
rect 21364 25245 21373 25279
rect 21373 25245 21407 25279
rect 21407 25245 21416 25279
rect 21364 25236 21416 25245
rect 22192 25236 22244 25288
rect 23020 25279 23072 25288
rect 23020 25245 23029 25279
rect 23029 25245 23063 25279
rect 23063 25245 23072 25279
rect 23020 25236 23072 25245
rect 23664 25236 23716 25288
rect 24124 25236 24176 25288
rect 25136 25279 25188 25288
rect 25136 25245 25145 25279
rect 25145 25245 25179 25279
rect 25179 25245 25188 25279
rect 25136 25236 25188 25245
rect 26332 25304 26384 25356
rect 28264 25304 28316 25356
rect 28356 25347 28408 25356
rect 28356 25313 28365 25347
rect 28365 25313 28399 25347
rect 28399 25313 28408 25347
rect 28356 25304 28408 25313
rect 25596 25236 25648 25288
rect 16948 25100 17000 25152
rect 17592 25100 17644 25152
rect 18880 25100 18932 25152
rect 26976 25168 27028 25220
rect 21548 25143 21600 25152
rect 21548 25109 21557 25143
rect 21557 25109 21591 25143
rect 21591 25109 21600 25143
rect 21548 25100 21600 25109
rect 22192 25100 22244 25152
rect 25320 25100 25372 25152
rect 25964 25100 26016 25152
rect 28724 25236 28776 25288
rect 29092 25236 29144 25288
rect 29736 25279 29788 25288
rect 29736 25245 29745 25279
rect 29745 25245 29779 25279
rect 29779 25245 29788 25279
rect 29736 25236 29788 25245
rect 30564 25304 30616 25356
rect 31944 25304 31996 25356
rect 32220 25304 32272 25356
rect 36084 25440 36136 25492
rect 30380 25236 30432 25288
rect 31116 25279 31168 25288
rect 31116 25245 31125 25279
rect 31125 25245 31159 25279
rect 31159 25245 31168 25279
rect 31116 25236 31168 25245
rect 36268 25304 36320 25356
rect 34428 25236 34480 25288
rect 34796 25279 34848 25288
rect 34796 25245 34805 25279
rect 34805 25245 34839 25279
rect 34839 25245 34848 25279
rect 34796 25236 34848 25245
rect 31668 25168 31720 25220
rect 32680 25168 32732 25220
rect 34060 25168 34112 25220
rect 28816 25143 28868 25152
rect 28816 25109 28825 25143
rect 28825 25109 28859 25143
rect 28859 25109 28868 25143
rect 28816 25100 28868 25109
rect 29000 25100 29052 25152
rect 29736 25100 29788 25152
rect 33508 25100 33560 25152
rect 35808 25100 35860 25152
rect 36820 25279 36872 25288
rect 36820 25245 36829 25279
rect 36829 25245 36863 25279
rect 36863 25245 36872 25279
rect 36820 25236 36872 25245
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4068 24896 4120 24948
rect 4712 24896 4764 24948
rect 8300 24896 8352 24948
rect 8484 24896 8536 24948
rect 8576 24896 8628 24948
rect 11520 24896 11572 24948
rect 12164 24896 12216 24948
rect 10048 24828 10100 24880
rect 12532 24828 12584 24880
rect 4712 24735 4764 24744
rect 4712 24701 4721 24735
rect 4721 24701 4755 24735
rect 4755 24701 4764 24735
rect 4712 24692 4764 24701
rect 4896 24735 4948 24744
rect 4896 24701 4905 24735
rect 4905 24701 4939 24735
rect 4939 24701 4948 24735
rect 4896 24692 4948 24701
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 8392 24760 8444 24769
rect 8668 24803 8720 24812
rect 8668 24769 8675 24803
rect 8675 24769 8720 24803
rect 8208 24692 8260 24744
rect 8668 24760 8720 24769
rect 8760 24803 8812 24812
rect 8760 24769 8769 24803
rect 8769 24769 8803 24803
rect 8803 24769 8812 24803
rect 8760 24760 8812 24769
rect 8852 24803 8904 24812
rect 8852 24769 8861 24803
rect 8861 24769 8895 24803
rect 8895 24769 8904 24803
rect 8852 24760 8904 24769
rect 9128 24760 9180 24812
rect 11428 24760 11480 24812
rect 9312 24692 9364 24744
rect 11060 24692 11112 24744
rect 9956 24624 10008 24676
rect 11612 24624 11664 24676
rect 12440 24803 12492 24812
rect 13452 24896 13504 24948
rect 13636 24871 13688 24880
rect 13636 24837 13645 24871
rect 13645 24837 13679 24871
rect 13679 24837 13688 24871
rect 13636 24828 13688 24837
rect 14832 24896 14884 24948
rect 12440 24769 12454 24803
rect 12454 24769 12488 24803
rect 12488 24769 12492 24803
rect 12440 24760 12492 24769
rect 12532 24692 12584 24744
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 13176 24803 13228 24812
rect 13176 24769 13190 24803
rect 13190 24769 13224 24803
rect 13224 24769 13228 24803
rect 13176 24760 13228 24769
rect 14004 24760 14056 24812
rect 14188 24760 14240 24812
rect 14280 24803 14332 24812
rect 14280 24769 14289 24803
rect 14289 24769 14323 24803
rect 14323 24769 14332 24803
rect 14280 24760 14332 24769
rect 15016 24760 15068 24812
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 18328 24896 18380 24948
rect 18420 24896 18472 24948
rect 15568 24871 15620 24880
rect 15568 24837 15577 24871
rect 15577 24837 15611 24871
rect 15611 24837 15620 24871
rect 15568 24828 15620 24837
rect 15660 24871 15712 24880
rect 15660 24837 15669 24871
rect 15669 24837 15703 24871
rect 15703 24837 15712 24871
rect 15660 24828 15712 24837
rect 17132 24828 17184 24880
rect 19340 24896 19392 24948
rect 16580 24760 16632 24812
rect 18236 24760 18288 24812
rect 19340 24803 19392 24812
rect 19340 24769 19349 24803
rect 19349 24769 19383 24803
rect 19383 24769 19392 24803
rect 19340 24760 19392 24769
rect 19800 24760 19852 24812
rect 20076 24760 20128 24812
rect 20168 24760 20220 24812
rect 14832 24692 14884 24744
rect 15200 24692 15252 24744
rect 15844 24692 15896 24744
rect 19524 24692 19576 24744
rect 19708 24735 19760 24744
rect 19708 24701 19717 24735
rect 19717 24701 19751 24735
rect 19751 24701 19760 24735
rect 19708 24692 19760 24701
rect 20076 24624 20128 24676
rect 20444 24760 20496 24812
rect 20720 24803 20772 24812
rect 20720 24769 20729 24803
rect 20729 24769 20763 24803
rect 20763 24769 20772 24803
rect 20720 24760 20772 24769
rect 21640 24896 21692 24948
rect 25136 24896 25188 24948
rect 27528 24896 27580 24948
rect 21272 24760 21324 24812
rect 22192 24760 22244 24812
rect 22836 24760 22888 24812
rect 23664 24760 23716 24812
rect 20904 24692 20956 24744
rect 22100 24735 22152 24744
rect 22100 24701 22109 24735
rect 22109 24701 22143 24735
rect 22143 24701 22152 24735
rect 22100 24692 22152 24701
rect 22284 24735 22336 24744
rect 22284 24701 22293 24735
rect 22293 24701 22327 24735
rect 22327 24701 22336 24735
rect 22284 24692 22336 24701
rect 22744 24692 22796 24744
rect 7840 24599 7892 24608
rect 7840 24565 7849 24599
rect 7849 24565 7883 24599
rect 7883 24565 7892 24599
rect 7840 24556 7892 24565
rect 9128 24599 9180 24608
rect 9128 24565 9137 24599
rect 9137 24565 9171 24599
rect 9171 24565 9180 24599
rect 9128 24556 9180 24565
rect 11980 24556 12032 24608
rect 13268 24556 13320 24608
rect 13360 24599 13412 24608
rect 13360 24565 13369 24599
rect 13369 24565 13403 24599
rect 13403 24565 13412 24599
rect 13360 24556 13412 24565
rect 14004 24599 14056 24608
rect 14004 24565 14013 24599
rect 14013 24565 14047 24599
rect 14047 24565 14056 24599
rect 14004 24556 14056 24565
rect 14924 24556 14976 24608
rect 15936 24599 15988 24608
rect 15936 24565 15945 24599
rect 15945 24565 15979 24599
rect 15979 24565 15988 24599
rect 15936 24556 15988 24565
rect 16948 24556 17000 24608
rect 17592 24556 17644 24608
rect 17868 24556 17920 24608
rect 18512 24556 18564 24608
rect 20352 24556 20404 24608
rect 21640 24556 21692 24608
rect 23480 24624 23532 24676
rect 24032 24760 24084 24812
rect 26884 24760 26936 24812
rect 27068 24803 27120 24812
rect 27068 24769 27077 24803
rect 27077 24769 27111 24803
rect 27111 24769 27120 24803
rect 27068 24760 27120 24769
rect 28724 24828 28776 24880
rect 28080 24760 28132 24812
rect 29276 24896 29328 24948
rect 24768 24692 24820 24744
rect 26976 24624 27028 24676
rect 30380 24760 30432 24812
rect 30748 24692 30800 24744
rect 31116 24735 31168 24744
rect 31116 24701 31125 24735
rect 31125 24701 31159 24735
rect 31159 24701 31168 24735
rect 31116 24692 31168 24701
rect 31852 24624 31904 24676
rect 41328 24624 41380 24676
rect 23756 24599 23808 24608
rect 23756 24565 23765 24599
rect 23765 24565 23799 24599
rect 23799 24565 23808 24599
rect 23756 24556 23808 24565
rect 24308 24556 24360 24608
rect 24492 24556 24544 24608
rect 24860 24556 24912 24608
rect 26792 24556 26844 24608
rect 28816 24556 28868 24608
rect 29184 24556 29236 24608
rect 31484 24599 31536 24608
rect 31484 24565 31493 24599
rect 31493 24565 31527 24599
rect 31527 24565 31536 24599
rect 31484 24556 31536 24565
rect 32404 24556 32456 24608
rect 41052 24599 41104 24608
rect 41052 24565 41061 24599
rect 41061 24565 41095 24599
rect 41095 24565 41104 24599
rect 41052 24556 41104 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 4896 24352 4948 24404
rect 11244 24352 11296 24404
rect 11704 24352 11756 24404
rect 7380 24284 7432 24336
rect 8208 24216 8260 24268
rect 11520 24284 11572 24336
rect 6092 24148 6144 24200
rect 7104 24191 7156 24200
rect 7104 24157 7113 24191
rect 7113 24157 7147 24191
rect 7147 24157 7156 24191
rect 7104 24148 7156 24157
rect 8852 24148 8904 24200
rect 9312 24191 9364 24200
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 10140 24148 10192 24200
rect 4712 24080 4764 24132
rect 9496 24080 9548 24132
rect 10968 24148 11020 24200
rect 11244 24148 11296 24200
rect 11428 24191 11480 24200
rect 11428 24157 11437 24191
rect 11437 24157 11471 24191
rect 11471 24157 11480 24191
rect 11428 24148 11480 24157
rect 11612 24191 11664 24200
rect 11612 24157 11621 24191
rect 11621 24157 11655 24191
rect 11655 24157 11664 24191
rect 11612 24148 11664 24157
rect 11796 24148 11848 24200
rect 11980 24148 12032 24200
rect 13176 24352 13228 24404
rect 13544 24352 13596 24404
rect 15200 24352 15252 24404
rect 15292 24352 15344 24404
rect 15936 24395 15988 24404
rect 15936 24361 15945 24395
rect 15945 24361 15979 24395
rect 15979 24361 15988 24395
rect 15936 24352 15988 24361
rect 12532 24284 12584 24336
rect 13728 24284 13780 24336
rect 14832 24284 14884 24336
rect 14004 24216 14056 24268
rect 12992 24191 13044 24200
rect 12992 24157 13001 24191
rect 13001 24157 13035 24191
rect 13035 24157 13044 24191
rect 12992 24148 13044 24157
rect 13268 24191 13320 24200
rect 13268 24157 13277 24191
rect 13277 24157 13311 24191
rect 13311 24157 13320 24191
rect 13268 24148 13320 24157
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 16120 24191 16172 24200
rect 16120 24157 16129 24191
rect 16129 24157 16163 24191
rect 16163 24157 16172 24191
rect 16120 24148 16172 24157
rect 14188 24123 14240 24132
rect 14188 24089 14197 24123
rect 14197 24089 14231 24123
rect 14231 24089 14240 24123
rect 14188 24080 14240 24089
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 17040 24284 17092 24336
rect 17224 24284 17276 24336
rect 17868 24352 17920 24404
rect 20352 24352 20404 24404
rect 20536 24352 20588 24404
rect 18328 24284 18380 24336
rect 19340 24284 19392 24336
rect 17408 24216 17460 24268
rect 18604 24216 18656 24268
rect 18696 24191 18748 24200
rect 940 24012 992 24064
rect 6828 24055 6880 24064
rect 6828 24021 6837 24055
rect 6837 24021 6871 24055
rect 6871 24021 6880 24055
rect 6828 24012 6880 24021
rect 7012 24012 7064 24064
rect 10048 24012 10100 24064
rect 10692 24012 10744 24064
rect 11980 24012 12032 24064
rect 14556 24012 14608 24064
rect 14832 24012 14884 24064
rect 16672 24012 16724 24064
rect 17224 24123 17276 24132
rect 17224 24089 17233 24123
rect 17233 24089 17267 24123
rect 17267 24089 17276 24123
rect 17224 24080 17276 24089
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 17776 24080 17828 24132
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 19800 24148 19852 24200
rect 21180 24284 21232 24336
rect 21732 24284 21784 24336
rect 20996 24216 21048 24268
rect 20076 24148 20128 24200
rect 21272 24148 21324 24200
rect 21456 24259 21508 24268
rect 21456 24225 21465 24259
rect 21465 24225 21499 24259
rect 21499 24225 21508 24259
rect 21456 24216 21508 24225
rect 22192 24284 22244 24336
rect 23020 24352 23072 24404
rect 23296 24352 23348 24404
rect 24308 24352 24360 24404
rect 23664 24284 23716 24336
rect 21640 24148 21692 24200
rect 22100 24148 22152 24200
rect 24676 24284 24728 24336
rect 24860 24284 24912 24336
rect 18972 24012 19024 24064
rect 19248 24055 19300 24064
rect 19248 24021 19257 24055
rect 19257 24021 19291 24055
rect 19291 24021 19300 24055
rect 19248 24012 19300 24021
rect 19340 24012 19392 24064
rect 19708 24012 19760 24064
rect 20444 24012 20496 24064
rect 20904 24123 20956 24132
rect 20904 24089 20913 24123
rect 20913 24089 20947 24123
rect 20947 24089 20956 24123
rect 20904 24080 20956 24089
rect 21456 24080 21508 24132
rect 21732 24012 21784 24064
rect 22008 24055 22060 24064
rect 22008 24021 22017 24055
rect 22017 24021 22051 24055
rect 22051 24021 22060 24055
rect 22008 24012 22060 24021
rect 22652 24191 22704 24200
rect 22652 24157 22661 24191
rect 22661 24157 22695 24191
rect 22695 24157 22704 24191
rect 22652 24148 22704 24157
rect 22744 24191 22796 24200
rect 22744 24157 22753 24191
rect 22753 24157 22787 24191
rect 22787 24157 22796 24191
rect 22744 24148 22796 24157
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 23480 24148 23532 24200
rect 22376 24080 22428 24132
rect 24032 24148 24084 24200
rect 24308 24148 24360 24200
rect 26056 24395 26108 24404
rect 26056 24361 26065 24395
rect 26065 24361 26099 24395
rect 26099 24361 26108 24395
rect 26056 24352 26108 24361
rect 38016 24395 38068 24404
rect 38016 24361 38025 24395
rect 38025 24361 38059 24395
rect 38059 24361 38068 24395
rect 38016 24352 38068 24361
rect 26884 24327 26936 24336
rect 26884 24293 26893 24327
rect 26893 24293 26927 24327
rect 26927 24293 26936 24327
rect 26884 24284 26936 24293
rect 27252 24284 27304 24336
rect 27436 24284 27488 24336
rect 28540 24284 28592 24336
rect 30196 24327 30248 24336
rect 30196 24293 30205 24327
rect 30205 24293 30239 24327
rect 30239 24293 30248 24327
rect 30196 24284 30248 24293
rect 30932 24327 30984 24336
rect 30932 24293 30941 24327
rect 30941 24293 30975 24327
rect 30975 24293 30984 24327
rect 30932 24284 30984 24293
rect 26792 24216 26844 24268
rect 27068 24148 27120 24200
rect 27436 24191 27488 24200
rect 27436 24157 27445 24191
rect 27445 24157 27479 24191
rect 27479 24157 27488 24191
rect 27436 24148 27488 24157
rect 30288 24259 30340 24268
rect 30288 24225 30297 24259
rect 30297 24225 30331 24259
rect 30331 24225 30340 24259
rect 30288 24216 30340 24225
rect 34796 24216 34848 24268
rect 25872 24012 25924 24064
rect 26424 24055 26476 24064
rect 26424 24021 26433 24055
rect 26433 24021 26467 24055
rect 26467 24021 26476 24055
rect 26424 24012 26476 24021
rect 27620 24080 27672 24132
rect 30748 24191 30800 24200
rect 30748 24157 30757 24191
rect 30757 24157 30791 24191
rect 30791 24157 30800 24191
rect 30748 24148 30800 24157
rect 30932 24191 30984 24200
rect 30932 24157 30941 24191
rect 30941 24157 30975 24191
rect 30975 24157 30984 24191
rect 30932 24148 30984 24157
rect 31484 24148 31536 24200
rect 32312 24148 32364 24200
rect 38292 24148 38344 24200
rect 27896 24080 27948 24132
rect 29276 24080 29328 24132
rect 31576 24080 31628 24132
rect 36544 24123 36596 24132
rect 36544 24089 36553 24123
rect 36553 24089 36587 24123
rect 36587 24089 36596 24123
rect 36544 24080 36596 24089
rect 27068 24055 27120 24064
rect 27068 24021 27077 24055
rect 27077 24021 27111 24055
rect 27111 24021 27120 24055
rect 27068 24012 27120 24021
rect 27528 24012 27580 24064
rect 28908 24012 28960 24064
rect 31760 24055 31812 24064
rect 31760 24021 31769 24055
rect 31769 24021 31803 24055
rect 31803 24021 31812 24055
rect 31760 24012 31812 24021
rect 35808 24012 35860 24064
rect 37004 24080 37056 24132
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 5540 23808 5592 23860
rect 4620 23783 4672 23792
rect 4620 23749 4629 23783
rect 4629 23749 4663 23783
rect 4663 23749 4672 23783
rect 4620 23740 4672 23749
rect 6092 23851 6144 23860
rect 6092 23817 6101 23851
rect 6101 23817 6135 23851
rect 6135 23817 6144 23851
rect 6092 23808 6144 23817
rect 8760 23808 8812 23860
rect 4068 23604 4120 23656
rect 7012 23604 7064 23656
rect 10416 23808 10468 23860
rect 10600 23604 10652 23656
rect 11796 23672 11848 23724
rect 11980 23715 12032 23724
rect 11980 23681 11989 23715
rect 11989 23681 12023 23715
rect 12023 23681 12032 23715
rect 11980 23672 12032 23681
rect 12624 23672 12676 23724
rect 13728 23808 13780 23860
rect 14188 23808 14240 23860
rect 15844 23808 15896 23860
rect 13360 23740 13412 23792
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 13268 23604 13320 23656
rect 11244 23536 11296 23588
rect 15108 23672 15160 23724
rect 15936 23672 15988 23724
rect 13636 23604 13688 23656
rect 16764 23740 16816 23792
rect 17040 23783 17092 23792
rect 17040 23749 17056 23783
rect 17056 23749 17090 23783
rect 17090 23749 17092 23783
rect 17040 23740 17092 23749
rect 17684 23808 17736 23860
rect 17868 23808 17920 23860
rect 18604 23808 18656 23860
rect 19248 23808 19300 23860
rect 24676 23808 24728 23860
rect 17132 23604 17184 23656
rect 8852 23511 8904 23520
rect 8852 23477 8861 23511
rect 8861 23477 8895 23511
rect 8895 23477 8904 23511
rect 8852 23468 8904 23477
rect 9128 23468 9180 23520
rect 10416 23511 10468 23520
rect 10416 23477 10425 23511
rect 10425 23477 10459 23511
rect 10459 23477 10468 23511
rect 10416 23468 10468 23477
rect 11336 23468 11388 23520
rect 12532 23511 12584 23520
rect 12532 23477 12541 23511
rect 12541 23477 12575 23511
rect 12575 23477 12584 23511
rect 12532 23468 12584 23477
rect 15844 23536 15896 23588
rect 17684 23604 17736 23656
rect 18880 23715 18932 23724
rect 18880 23681 18889 23715
rect 18889 23681 18923 23715
rect 18923 23681 18932 23715
rect 18880 23672 18932 23681
rect 20168 23672 20220 23724
rect 20444 23672 20496 23724
rect 19064 23604 19116 23656
rect 20812 23783 20864 23792
rect 20812 23749 20821 23783
rect 20821 23749 20855 23783
rect 20855 23749 20864 23783
rect 20812 23740 20864 23749
rect 20996 23715 21048 23724
rect 20996 23681 21005 23715
rect 21005 23681 21039 23715
rect 21039 23681 21048 23715
rect 20996 23672 21048 23681
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 24216 23715 24268 23724
rect 24216 23681 24225 23715
rect 24225 23681 24259 23715
rect 24259 23681 24268 23715
rect 24216 23672 24268 23681
rect 26240 23808 26292 23860
rect 26884 23808 26936 23860
rect 27252 23808 27304 23860
rect 24860 23672 24912 23724
rect 25596 23672 25648 23724
rect 30932 23808 30984 23860
rect 26148 23672 26200 23724
rect 26332 23672 26384 23724
rect 28264 23740 28316 23792
rect 33048 23808 33100 23860
rect 34704 23808 34756 23860
rect 36544 23808 36596 23860
rect 34060 23740 34112 23792
rect 15384 23468 15436 23520
rect 15568 23468 15620 23520
rect 16764 23468 16816 23520
rect 16856 23468 16908 23520
rect 18512 23536 18564 23588
rect 18972 23536 19024 23588
rect 19892 23536 19944 23588
rect 20260 23536 20312 23588
rect 21088 23647 21140 23656
rect 21088 23613 21097 23647
rect 21097 23613 21131 23647
rect 21131 23613 21140 23647
rect 21088 23604 21140 23613
rect 21180 23647 21232 23656
rect 21180 23613 21189 23647
rect 21189 23613 21223 23647
rect 21223 23613 21232 23647
rect 21180 23604 21232 23613
rect 23296 23604 23348 23656
rect 24492 23604 24544 23656
rect 17132 23468 17184 23520
rect 18420 23511 18472 23520
rect 18420 23477 18429 23511
rect 18429 23477 18463 23511
rect 18463 23477 18472 23511
rect 18420 23468 18472 23477
rect 18880 23468 18932 23520
rect 20444 23511 20496 23520
rect 20444 23477 20453 23511
rect 20453 23477 20487 23511
rect 20487 23477 20496 23511
rect 20444 23468 20496 23477
rect 24676 23536 24728 23588
rect 26700 23604 26752 23656
rect 26884 23604 26936 23656
rect 27988 23672 28040 23724
rect 31760 23672 31812 23724
rect 34796 23740 34848 23792
rect 35808 23740 35860 23792
rect 38016 23808 38068 23860
rect 37740 23783 37792 23792
rect 37740 23749 37749 23783
rect 37749 23749 37783 23783
rect 37783 23749 37792 23783
rect 37740 23740 37792 23749
rect 27528 23604 27580 23656
rect 29184 23604 29236 23656
rect 30012 23647 30064 23656
rect 30012 23613 30021 23647
rect 30021 23613 30055 23647
rect 30055 23613 30064 23647
rect 30012 23604 30064 23613
rect 30656 23604 30708 23656
rect 32680 23604 32732 23656
rect 34520 23647 34572 23656
rect 34520 23613 34529 23647
rect 34529 23613 34563 23647
rect 34563 23613 34572 23647
rect 34520 23604 34572 23613
rect 36636 23647 36688 23656
rect 36636 23613 36645 23647
rect 36645 23613 36679 23647
rect 36679 23613 36688 23647
rect 36636 23604 36688 23613
rect 36728 23647 36780 23656
rect 36728 23613 36737 23647
rect 36737 23613 36771 23647
rect 36771 23613 36780 23647
rect 36728 23604 36780 23613
rect 23112 23468 23164 23520
rect 23664 23468 23716 23520
rect 24768 23468 24820 23520
rect 25596 23536 25648 23588
rect 31852 23536 31904 23588
rect 38292 23604 38344 23656
rect 26332 23511 26384 23520
rect 26332 23477 26341 23511
rect 26341 23477 26375 23511
rect 26375 23477 26384 23511
rect 26332 23468 26384 23477
rect 26424 23468 26476 23520
rect 26792 23468 26844 23520
rect 32404 23468 32456 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1400 23264 1452 23316
rect 4620 23264 4672 23316
rect 7104 23307 7156 23316
rect 7104 23273 7113 23307
rect 7113 23273 7147 23307
rect 7147 23273 7156 23307
rect 7104 23264 7156 23273
rect 11428 23307 11480 23316
rect 11428 23273 11437 23307
rect 11437 23273 11471 23307
rect 11471 23273 11480 23307
rect 11428 23264 11480 23273
rect 11704 23264 11756 23316
rect 12900 23264 12952 23316
rect 17132 23264 17184 23316
rect 9220 23196 9272 23248
rect 10600 23196 10652 23248
rect 7840 23128 7892 23180
rect 8852 23128 8904 23180
rect 1860 23103 1912 23112
rect 1860 23069 1869 23103
rect 1869 23069 1903 23103
rect 1903 23069 1912 23103
rect 1860 23060 1912 23069
rect 6828 23060 6880 23112
rect 12440 23128 12492 23180
rect 13084 23128 13136 23180
rect 10048 23060 10100 23112
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 13912 23060 13964 23112
rect 8024 22992 8076 23044
rect 8116 22924 8168 22976
rect 9312 22992 9364 23044
rect 13084 22992 13136 23044
rect 13268 22992 13320 23044
rect 15016 23103 15068 23112
rect 15016 23069 15025 23103
rect 15025 23069 15059 23103
rect 15059 23069 15068 23103
rect 15016 23060 15068 23069
rect 15292 23060 15344 23112
rect 15568 23196 15620 23248
rect 16028 23196 16080 23248
rect 16764 23196 16816 23248
rect 27988 23264 28040 23316
rect 30012 23264 30064 23316
rect 32680 23264 32732 23316
rect 17408 23196 17460 23248
rect 20352 23196 20404 23248
rect 21180 23196 21232 23248
rect 16028 23103 16080 23112
rect 16028 23069 16037 23103
rect 16037 23069 16071 23103
rect 16071 23069 16080 23103
rect 16028 23060 16080 23069
rect 17684 23128 17736 23180
rect 16948 23060 17000 23112
rect 22744 23128 22796 23180
rect 24032 23196 24084 23248
rect 25044 23239 25096 23248
rect 25044 23205 25053 23239
rect 25053 23205 25087 23239
rect 25087 23205 25096 23239
rect 25044 23196 25096 23205
rect 25228 23239 25280 23248
rect 25228 23205 25237 23239
rect 25237 23205 25271 23239
rect 25271 23205 25280 23239
rect 25228 23196 25280 23205
rect 18604 23060 18656 23112
rect 19064 23060 19116 23112
rect 20076 23060 20128 23112
rect 11060 22924 11112 22976
rect 11888 22924 11940 22976
rect 14280 22924 14332 22976
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 15476 22924 15528 22976
rect 15568 22924 15620 22976
rect 20168 22992 20220 23044
rect 16672 22924 16724 22976
rect 17776 22924 17828 22976
rect 18144 22967 18196 22976
rect 18144 22933 18153 22967
rect 18153 22933 18187 22967
rect 18187 22933 18196 22967
rect 18144 22924 18196 22933
rect 18788 22924 18840 22976
rect 19064 22924 19116 22976
rect 20352 22924 20404 22976
rect 20628 23060 20680 23112
rect 20812 23060 20864 23112
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 20996 23060 21048 23069
rect 21088 23103 21140 23112
rect 21088 23069 21097 23103
rect 21097 23069 21131 23103
rect 21131 23069 21140 23103
rect 21088 23060 21140 23069
rect 21180 23103 21232 23112
rect 21180 23069 21189 23103
rect 21189 23069 21223 23103
rect 21223 23069 21232 23103
rect 21180 23060 21232 23069
rect 22468 23060 22520 23112
rect 23848 23128 23900 23180
rect 21364 22992 21416 23044
rect 23664 22992 23716 23044
rect 24584 22992 24636 23044
rect 25228 23060 25280 23112
rect 27528 23196 27580 23248
rect 27712 23196 27764 23248
rect 26332 23060 26384 23112
rect 27436 23171 27488 23180
rect 27436 23137 27445 23171
rect 27445 23137 27479 23171
rect 27479 23137 27488 23171
rect 27436 23128 27488 23137
rect 29000 23128 29052 23180
rect 25780 22992 25832 23044
rect 26424 23035 26476 23044
rect 26424 23001 26433 23035
rect 26433 23001 26467 23035
rect 26467 23001 26476 23035
rect 26424 22992 26476 23001
rect 23296 22924 23348 22976
rect 23572 22924 23624 22976
rect 24860 22924 24912 22976
rect 28264 23060 28316 23112
rect 28816 23103 28868 23112
rect 28816 23069 28825 23103
rect 28825 23069 28859 23103
rect 28859 23069 28868 23103
rect 28816 23060 28868 23069
rect 29092 23103 29144 23112
rect 29092 23069 29101 23103
rect 29101 23069 29135 23103
rect 29135 23069 29144 23103
rect 29092 23060 29144 23069
rect 29552 23060 29604 23112
rect 29920 23196 29972 23248
rect 30656 23239 30708 23248
rect 30656 23205 30665 23239
rect 30665 23205 30699 23239
rect 30699 23205 30708 23239
rect 30656 23196 30708 23205
rect 31576 23239 31628 23248
rect 31576 23205 31585 23239
rect 31585 23205 31619 23239
rect 31619 23205 31628 23239
rect 31576 23196 31628 23205
rect 30380 23171 30432 23180
rect 30380 23137 30389 23171
rect 30389 23137 30423 23171
rect 30423 23137 30432 23171
rect 30380 23128 30432 23137
rect 30472 23128 30524 23180
rect 35716 23128 35768 23180
rect 31668 23103 31720 23112
rect 31668 23069 31677 23103
rect 31677 23069 31711 23103
rect 31711 23069 31720 23103
rect 31668 23060 31720 23069
rect 31944 23060 31996 23112
rect 32312 23060 32364 23112
rect 32404 23103 32456 23112
rect 32404 23069 32413 23103
rect 32413 23069 32447 23103
rect 32447 23069 32456 23103
rect 32404 23060 32456 23069
rect 32680 23103 32732 23112
rect 32680 23069 32689 23103
rect 32689 23069 32723 23103
rect 32723 23069 32732 23103
rect 32680 23060 32732 23069
rect 34060 23060 34112 23112
rect 34704 23060 34756 23112
rect 28172 22967 28224 22976
rect 28172 22933 28181 22967
rect 28181 22933 28215 22967
rect 28215 22933 28224 22967
rect 28172 22924 28224 22933
rect 28448 22967 28500 22976
rect 28448 22933 28457 22967
rect 28457 22933 28491 22967
rect 28491 22933 28500 22967
rect 28448 22924 28500 22933
rect 30564 22924 30616 22976
rect 34336 22924 34388 22976
rect 34704 22967 34756 22976
rect 34704 22933 34713 22967
rect 34713 22933 34747 22967
rect 34747 22933 34756 22967
rect 34704 22924 34756 22933
rect 37372 22924 37424 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9220 22720 9272 22772
rect 11796 22763 11848 22772
rect 11796 22729 11805 22763
rect 11805 22729 11839 22763
rect 11839 22729 11848 22763
rect 11796 22720 11848 22729
rect 11888 22720 11940 22772
rect 5540 22584 5592 22636
rect 7104 22584 7156 22636
rect 10508 22627 10560 22636
rect 10508 22593 10517 22627
rect 10517 22593 10551 22627
rect 10551 22593 10560 22627
rect 10508 22584 10560 22593
rect 4896 22516 4948 22568
rect 6552 22516 6604 22568
rect 9128 22516 9180 22568
rect 10784 22559 10836 22568
rect 10784 22525 10793 22559
rect 10793 22525 10827 22559
rect 10827 22525 10836 22559
rect 10784 22516 10836 22525
rect 12440 22720 12492 22772
rect 12992 22695 13044 22704
rect 12992 22661 13001 22695
rect 13001 22661 13035 22695
rect 13035 22661 13044 22695
rect 12992 22652 13044 22661
rect 13728 22652 13780 22704
rect 14832 22695 14884 22704
rect 14832 22661 14841 22695
rect 14841 22661 14875 22695
rect 14875 22661 14884 22695
rect 14832 22652 14884 22661
rect 13084 22584 13136 22636
rect 13176 22627 13228 22636
rect 13176 22593 13185 22627
rect 13185 22593 13219 22627
rect 13219 22593 13228 22627
rect 13176 22584 13228 22593
rect 5724 22423 5776 22432
rect 5724 22389 5733 22423
rect 5733 22389 5767 22423
rect 5767 22389 5776 22423
rect 5724 22380 5776 22389
rect 10140 22380 10192 22432
rect 12624 22448 12676 22500
rect 14004 22584 14056 22636
rect 14648 22584 14700 22636
rect 14924 22584 14976 22636
rect 15568 22652 15620 22704
rect 18328 22720 18380 22772
rect 16396 22652 16448 22704
rect 16580 22652 16632 22704
rect 19340 22652 19392 22704
rect 15660 22584 15712 22636
rect 16580 22448 16632 22500
rect 16856 22584 16908 22636
rect 16948 22627 17000 22636
rect 16948 22593 16957 22627
rect 16957 22593 16991 22627
rect 16991 22593 17000 22627
rect 16948 22584 17000 22593
rect 18144 22584 18196 22636
rect 18512 22584 18564 22636
rect 18604 22584 18656 22636
rect 18788 22584 18840 22636
rect 18328 22559 18380 22568
rect 18328 22525 18337 22559
rect 18337 22525 18371 22559
rect 18371 22525 18380 22559
rect 18328 22516 18380 22525
rect 18972 22584 19024 22636
rect 19892 22516 19944 22568
rect 22008 22720 22060 22772
rect 28448 22720 28500 22772
rect 30472 22720 30524 22772
rect 34520 22720 34572 22772
rect 34704 22720 34756 22772
rect 20168 22652 20220 22704
rect 20352 22584 20404 22636
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 20720 22584 20772 22593
rect 21824 22695 21876 22704
rect 21824 22661 21833 22695
rect 21833 22661 21867 22695
rect 21867 22661 21876 22695
rect 21824 22652 21876 22661
rect 23664 22695 23716 22704
rect 23664 22661 23673 22695
rect 23673 22661 23707 22695
rect 23707 22661 23716 22695
rect 23664 22652 23716 22661
rect 24032 22652 24084 22704
rect 22284 22584 22336 22636
rect 24308 22627 24360 22636
rect 24308 22593 24317 22627
rect 24317 22593 24351 22627
rect 24351 22593 24360 22627
rect 24308 22584 24360 22593
rect 24492 22627 24544 22636
rect 24492 22593 24501 22627
rect 24501 22593 24535 22627
rect 24535 22593 24544 22627
rect 24492 22584 24544 22593
rect 26608 22584 26660 22636
rect 29000 22584 29052 22636
rect 29184 22516 29236 22568
rect 29736 22627 29788 22636
rect 29736 22593 29745 22627
rect 29745 22593 29779 22627
rect 29779 22593 29788 22627
rect 29736 22584 29788 22593
rect 30380 22652 30432 22704
rect 31116 22652 31168 22704
rect 29920 22584 29972 22636
rect 37004 22652 37056 22704
rect 14280 22380 14332 22432
rect 14556 22380 14608 22432
rect 15108 22423 15160 22432
rect 15108 22389 15117 22423
rect 15117 22389 15151 22423
rect 15151 22389 15160 22423
rect 15108 22380 15160 22389
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 15476 22423 15528 22432
rect 15476 22389 15485 22423
rect 15485 22389 15519 22423
rect 15519 22389 15528 22423
rect 15476 22380 15528 22389
rect 15936 22423 15988 22432
rect 15936 22389 15945 22423
rect 15945 22389 15979 22423
rect 15979 22389 15988 22423
rect 15936 22380 15988 22389
rect 16672 22423 16724 22432
rect 16672 22389 16681 22423
rect 16681 22389 16715 22423
rect 16715 22389 16724 22423
rect 16672 22380 16724 22389
rect 18236 22423 18288 22432
rect 18236 22389 18245 22423
rect 18245 22389 18279 22423
rect 18279 22389 18288 22423
rect 18236 22380 18288 22389
rect 18604 22423 18656 22432
rect 18604 22389 18613 22423
rect 18613 22389 18647 22423
rect 18647 22389 18656 22423
rect 18604 22380 18656 22389
rect 19432 22380 19484 22432
rect 20076 22380 20128 22432
rect 22100 22448 22152 22500
rect 23296 22491 23348 22500
rect 23296 22457 23305 22491
rect 23305 22457 23339 22491
rect 23339 22457 23348 22491
rect 23296 22448 23348 22457
rect 32312 22448 32364 22500
rect 35808 22448 35860 22500
rect 24032 22380 24084 22432
rect 24584 22380 24636 22432
rect 29552 22380 29604 22432
rect 37556 22559 37608 22568
rect 37556 22525 37565 22559
rect 37565 22525 37599 22559
rect 37599 22525 37608 22559
rect 37556 22516 37608 22525
rect 39304 22559 39356 22568
rect 39304 22525 39313 22559
rect 39313 22525 39347 22559
rect 39347 22525 39356 22559
rect 39304 22516 39356 22525
rect 38292 22380 38344 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1860 22176 1912 22228
rect 5540 22219 5592 22228
rect 5540 22185 5549 22219
rect 5549 22185 5583 22219
rect 5583 22185 5592 22219
rect 5540 22176 5592 22185
rect 7380 22176 7432 22228
rect 12992 22176 13044 22228
rect 4068 22040 4120 22092
rect 5356 22040 5408 22092
rect 8116 22040 8168 22092
rect 2228 22015 2280 22024
rect 2228 21981 2237 22015
rect 2237 21981 2271 22015
rect 2271 21981 2280 22015
rect 2228 21972 2280 21981
rect 8576 22083 8628 22092
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 8576 22040 8628 22049
rect 4528 21904 4580 21956
rect 8208 21947 8260 21956
rect 8208 21913 8217 21947
rect 8217 21913 8251 21947
rect 8251 21913 8260 21947
rect 8208 21904 8260 21913
rect 9772 21972 9824 22024
rect 10968 22108 11020 22160
rect 10140 22015 10192 22024
rect 10140 21981 10149 22015
rect 10149 21981 10183 22015
rect 10183 21981 10192 22015
rect 10140 21972 10192 21981
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 11520 21972 11572 22024
rect 12624 22040 12676 22092
rect 13452 22176 13504 22228
rect 14004 22176 14056 22228
rect 15844 22176 15896 22228
rect 18144 22176 18196 22228
rect 20076 22176 20128 22228
rect 20628 22176 20680 22228
rect 21456 22176 21508 22228
rect 23112 22219 23164 22228
rect 23112 22185 23121 22219
rect 23121 22185 23155 22219
rect 23155 22185 23164 22219
rect 23112 22176 23164 22185
rect 25228 22176 25280 22228
rect 25872 22176 25924 22228
rect 26148 22176 26200 22228
rect 29000 22176 29052 22228
rect 37556 22176 37608 22228
rect 13360 22108 13412 22160
rect 16028 22108 16080 22160
rect 10876 21904 10928 21956
rect 2964 21836 3016 21888
rect 4436 21836 4488 21888
rect 5540 21836 5592 21888
rect 5816 21836 5868 21888
rect 7932 21879 7984 21888
rect 7932 21845 7941 21879
rect 7941 21845 7975 21879
rect 7975 21845 7984 21879
rect 7932 21836 7984 21845
rect 9128 21836 9180 21888
rect 10508 21836 10560 21888
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 14464 22083 14516 22092
rect 14464 22049 14473 22083
rect 14473 22049 14507 22083
rect 14507 22049 14516 22083
rect 14464 22040 14516 22049
rect 11244 21879 11296 21888
rect 11244 21845 11253 21879
rect 11253 21845 11287 21879
rect 11287 21845 11296 21879
rect 11244 21836 11296 21845
rect 12348 21904 12400 21956
rect 11428 21836 11480 21888
rect 11520 21879 11572 21888
rect 11520 21845 11529 21879
rect 11529 21845 11563 21879
rect 11563 21845 11572 21879
rect 11520 21836 11572 21845
rect 12072 21879 12124 21888
rect 12072 21845 12081 21879
rect 12081 21845 12115 21879
rect 12115 21845 12124 21879
rect 12072 21836 12124 21845
rect 12716 21836 12768 21888
rect 12808 21836 12860 21888
rect 13176 22015 13228 22024
rect 13176 21981 13185 22015
rect 13185 21981 13219 22015
rect 13219 21981 13228 22015
rect 13176 21972 13228 21981
rect 13268 21972 13320 22024
rect 13820 21972 13872 22024
rect 14556 22015 14608 22024
rect 14556 21981 14565 22015
rect 14565 21981 14599 22015
rect 14599 21981 14608 22015
rect 14556 21972 14608 21981
rect 13452 21904 13504 21956
rect 14280 21904 14332 21956
rect 15660 21904 15712 21956
rect 17224 21904 17276 21956
rect 17776 21972 17828 22024
rect 18328 21972 18380 22024
rect 15292 21836 15344 21888
rect 17776 21836 17828 21888
rect 18512 22083 18564 22092
rect 18512 22049 18521 22083
rect 18521 22049 18555 22083
rect 18555 22049 18564 22083
rect 18512 22040 18564 22049
rect 18788 22151 18840 22160
rect 18788 22117 18797 22151
rect 18797 22117 18831 22151
rect 18831 22117 18840 22151
rect 18788 22108 18840 22117
rect 19064 22015 19116 22024
rect 19064 21981 19073 22015
rect 19073 21981 19107 22015
rect 19107 21981 19116 22015
rect 19064 21972 19116 21981
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 19340 21972 19392 22024
rect 19524 22040 19576 22092
rect 20720 22108 20772 22160
rect 21088 22151 21140 22160
rect 21088 22117 21097 22151
rect 21097 22117 21131 22151
rect 21131 22117 21140 22151
rect 21088 22108 21140 22117
rect 22284 22108 22336 22160
rect 24952 22151 25004 22160
rect 19616 21972 19668 22024
rect 20076 21972 20128 22024
rect 20628 22015 20680 22024
rect 20628 21981 20637 22015
rect 20637 21981 20671 22015
rect 20671 21981 20680 22015
rect 20628 21972 20680 21981
rect 21916 22040 21968 22092
rect 24952 22117 24961 22151
rect 24961 22117 24995 22151
rect 24995 22117 25004 22151
rect 24952 22108 25004 22117
rect 20168 21904 20220 21956
rect 19340 21879 19392 21888
rect 19340 21845 19349 21879
rect 19349 21845 19383 21879
rect 19383 21845 19392 21879
rect 19340 21836 19392 21845
rect 19892 21836 19944 21888
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 23020 22015 23072 22024
rect 23020 21981 23029 22015
rect 23029 21981 23063 22015
rect 23063 21981 23072 22015
rect 23020 21972 23072 21981
rect 23388 22040 23440 22092
rect 23756 22040 23808 22092
rect 24124 22083 24176 22092
rect 24124 22049 24133 22083
rect 24133 22049 24167 22083
rect 24167 22049 24176 22083
rect 24124 22040 24176 22049
rect 24400 22040 24452 22092
rect 24860 22083 24912 22092
rect 24860 22049 24869 22083
rect 24869 22049 24903 22083
rect 24903 22049 24912 22083
rect 24860 22040 24912 22049
rect 28908 22108 28960 22160
rect 29552 22108 29604 22160
rect 37740 22108 37792 22160
rect 23664 21972 23716 22024
rect 23848 22015 23900 22024
rect 23848 21981 23857 22015
rect 23857 21981 23891 22015
rect 23891 21981 23900 22015
rect 23848 21972 23900 21981
rect 21364 21947 21416 21956
rect 21364 21913 21373 21947
rect 21373 21913 21407 21947
rect 21407 21913 21416 21947
rect 21364 21904 21416 21913
rect 22100 21904 22152 21956
rect 24216 21972 24268 22024
rect 24308 21972 24360 22024
rect 27528 21947 27580 21956
rect 27528 21913 27537 21947
rect 27537 21913 27571 21947
rect 27571 21913 27580 21947
rect 27528 21904 27580 21913
rect 24400 21879 24452 21888
rect 24400 21845 24409 21879
rect 24409 21845 24443 21879
rect 24443 21845 24452 21879
rect 24400 21836 24452 21845
rect 25596 21836 25648 21888
rect 26332 21836 26384 21888
rect 27436 21836 27488 21888
rect 28632 21972 28684 22024
rect 35440 22040 35492 22092
rect 35348 21972 35400 22024
rect 36636 21972 36688 22024
rect 30012 21904 30064 21956
rect 37648 22083 37700 22092
rect 37648 22049 37657 22083
rect 37657 22049 37691 22083
rect 37691 22049 37700 22083
rect 37648 22040 37700 22049
rect 37556 22015 37608 22024
rect 37556 21981 37565 22015
rect 37565 21981 37599 22015
rect 37599 21981 37608 22015
rect 39304 22040 39356 22092
rect 37556 21972 37608 21981
rect 28264 21836 28316 21888
rect 36820 21836 36872 21888
rect 37464 21879 37516 21888
rect 37464 21845 37473 21879
rect 37473 21845 37507 21879
rect 37507 21845 37516 21879
rect 37464 21836 37516 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 5356 21607 5408 21616
rect 5356 21573 5365 21607
rect 5365 21573 5399 21607
rect 5399 21573 5408 21607
rect 5356 21564 5408 21573
rect 4068 21496 4120 21548
rect 4528 21496 4580 21548
rect 4804 21496 4856 21548
rect 5172 21496 5224 21548
rect 1400 21428 1452 21480
rect 2228 21428 2280 21480
rect 2964 21471 3016 21480
rect 2964 21437 2973 21471
rect 2973 21437 3007 21471
rect 3007 21437 3016 21471
rect 2964 21428 3016 21437
rect 4896 21428 4948 21480
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 6552 21564 6604 21616
rect 7104 21564 7156 21616
rect 9772 21632 9824 21684
rect 9220 21564 9272 21616
rect 6644 21471 6696 21480
rect 6644 21437 6653 21471
rect 6653 21437 6687 21471
rect 6687 21437 6696 21471
rect 6644 21428 6696 21437
rect 7012 21428 7064 21480
rect 8116 21428 8168 21480
rect 8392 21539 8444 21548
rect 8392 21505 8401 21539
rect 8401 21505 8435 21539
rect 8435 21505 8444 21539
rect 8392 21496 8444 21505
rect 10600 21632 10652 21684
rect 10600 21539 10652 21548
rect 10600 21505 10609 21539
rect 10609 21505 10643 21539
rect 10643 21505 10652 21539
rect 10600 21496 10652 21505
rect 10692 21539 10744 21548
rect 10692 21505 10701 21539
rect 10701 21505 10735 21539
rect 10735 21505 10744 21539
rect 10692 21496 10744 21505
rect 11244 21632 11296 21684
rect 10876 21496 10928 21548
rect 12072 21564 12124 21616
rect 14740 21632 14792 21684
rect 16396 21632 16448 21684
rect 17224 21675 17276 21684
rect 17224 21641 17233 21675
rect 17233 21641 17267 21675
rect 17267 21641 17276 21675
rect 17224 21632 17276 21641
rect 13820 21564 13872 21616
rect 13452 21539 13504 21548
rect 13452 21505 13461 21539
rect 13461 21505 13495 21539
rect 13495 21505 13504 21539
rect 13452 21496 13504 21505
rect 13636 21496 13688 21548
rect 15936 21496 15988 21548
rect 20076 21632 20128 21684
rect 20444 21632 20496 21684
rect 21640 21632 21692 21684
rect 23020 21632 23072 21684
rect 24400 21632 24452 21684
rect 25504 21632 25556 21684
rect 14280 21428 14332 21480
rect 18144 21564 18196 21616
rect 17776 21496 17828 21548
rect 17868 21539 17920 21548
rect 17868 21505 17877 21539
rect 17877 21505 17911 21539
rect 17911 21505 17920 21539
rect 17868 21496 17920 21505
rect 5816 21292 5868 21344
rect 5908 21335 5960 21344
rect 5908 21301 5917 21335
rect 5917 21301 5951 21335
rect 5951 21301 5960 21335
rect 13820 21360 13872 21412
rect 14096 21360 14148 21412
rect 17776 21403 17828 21412
rect 17776 21369 17785 21403
rect 17785 21369 17819 21403
rect 17819 21369 17828 21403
rect 17776 21360 17828 21369
rect 18144 21428 18196 21480
rect 18420 21539 18472 21548
rect 18420 21505 18429 21539
rect 18429 21505 18463 21539
rect 18463 21505 18472 21539
rect 18420 21496 18472 21505
rect 18604 21496 18656 21548
rect 20628 21564 20680 21616
rect 19064 21539 19116 21548
rect 19064 21505 19073 21539
rect 19073 21505 19107 21539
rect 19107 21505 19116 21539
rect 19064 21496 19116 21505
rect 20352 21496 20404 21548
rect 21548 21496 21600 21548
rect 21916 21496 21968 21548
rect 23480 21607 23532 21616
rect 23480 21573 23489 21607
rect 23489 21573 23523 21607
rect 23523 21573 23532 21607
rect 23480 21564 23532 21573
rect 20168 21428 20220 21480
rect 21640 21428 21692 21480
rect 25228 21564 25280 21616
rect 23756 21496 23808 21548
rect 25596 21539 25648 21548
rect 25596 21505 25605 21539
rect 25605 21505 25639 21539
rect 25639 21505 25648 21539
rect 25596 21496 25648 21505
rect 25688 21539 25740 21548
rect 25688 21505 25698 21539
rect 25698 21505 25732 21539
rect 25732 21505 25740 21539
rect 25688 21496 25740 21505
rect 25872 21539 25924 21548
rect 25872 21505 25881 21539
rect 25881 21505 25915 21539
rect 25915 21505 25924 21539
rect 25872 21496 25924 21505
rect 26148 21496 26200 21548
rect 26332 21539 26384 21548
rect 26332 21505 26341 21539
rect 26341 21505 26375 21539
rect 26375 21505 26384 21539
rect 26332 21496 26384 21505
rect 26608 21471 26660 21480
rect 26608 21437 26617 21471
rect 26617 21437 26651 21471
rect 26651 21437 26660 21471
rect 26608 21428 26660 21437
rect 26792 21428 26844 21480
rect 30012 21632 30064 21684
rect 28632 21564 28684 21616
rect 30564 21564 30616 21616
rect 31484 21632 31536 21684
rect 31576 21675 31628 21684
rect 31576 21641 31585 21675
rect 31585 21641 31619 21675
rect 31619 21641 31628 21675
rect 31576 21632 31628 21641
rect 32220 21632 32272 21684
rect 19248 21360 19300 21412
rect 22652 21403 22704 21412
rect 22652 21369 22661 21403
rect 22661 21369 22695 21403
rect 22695 21369 22704 21403
rect 22652 21360 22704 21369
rect 23848 21360 23900 21412
rect 28540 21428 28592 21480
rect 5908 21292 5960 21301
rect 12072 21292 12124 21344
rect 12532 21292 12584 21344
rect 17960 21292 18012 21344
rect 18512 21292 18564 21344
rect 18604 21335 18656 21344
rect 18604 21301 18613 21335
rect 18613 21301 18647 21335
rect 18647 21301 18656 21335
rect 18604 21292 18656 21301
rect 22008 21292 22060 21344
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 29368 21471 29420 21480
rect 29368 21437 29377 21471
rect 29377 21437 29411 21471
rect 29411 21437 29420 21471
rect 29368 21428 29420 21437
rect 29460 21471 29512 21480
rect 29460 21437 29469 21471
rect 29469 21437 29503 21471
rect 29503 21437 29512 21471
rect 29460 21428 29512 21437
rect 28632 21360 28684 21412
rect 31484 21496 31536 21548
rect 31576 21428 31628 21480
rect 28908 21335 28960 21344
rect 28908 21301 28917 21335
rect 28917 21301 28951 21335
rect 28951 21301 28960 21335
rect 28908 21292 28960 21301
rect 31024 21292 31076 21344
rect 31208 21292 31260 21344
rect 31392 21335 31444 21344
rect 31392 21301 31401 21335
rect 31401 21301 31435 21335
rect 31435 21301 31444 21335
rect 31392 21292 31444 21301
rect 32496 21428 32548 21480
rect 33140 21428 33192 21480
rect 33692 21496 33744 21548
rect 37464 21632 37516 21684
rect 32220 21292 32272 21344
rect 36084 21428 36136 21480
rect 36820 21539 36872 21548
rect 36820 21505 36829 21539
rect 36829 21505 36863 21539
rect 36863 21505 36872 21539
rect 36820 21496 36872 21505
rect 37280 21496 37332 21548
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4620 21088 4672 21140
rect 5908 21088 5960 21140
rect 6644 21088 6696 21140
rect 6736 21088 6788 21140
rect 7932 21088 7984 21140
rect 5632 20884 5684 20936
rect 6920 21020 6972 21072
rect 6460 20995 6512 21004
rect 6460 20961 6469 20995
rect 6469 20961 6503 20995
rect 6503 20961 6512 20995
rect 6460 20952 6512 20961
rect 6644 20884 6696 20936
rect 6920 20927 6972 20936
rect 6920 20893 6929 20927
rect 6929 20893 6963 20927
rect 6963 20893 6972 20927
rect 6920 20884 6972 20893
rect 7564 20952 7616 21004
rect 9220 21020 9272 21072
rect 10692 21088 10744 21140
rect 11520 21088 11572 21140
rect 13544 21088 13596 21140
rect 13820 21088 13872 21140
rect 16120 21088 16172 21140
rect 17500 21088 17552 21140
rect 17776 21088 17828 21140
rect 18236 21088 18288 21140
rect 18420 21088 18472 21140
rect 18604 21088 18656 21140
rect 10232 20952 10284 21004
rect 13912 21020 13964 21072
rect 18788 21020 18840 21072
rect 23480 21088 23532 21140
rect 23388 21020 23440 21072
rect 12164 20995 12216 21004
rect 12164 20961 12173 20995
rect 12173 20961 12207 20995
rect 12207 20961 12216 20995
rect 12164 20952 12216 20961
rect 12256 20995 12308 21004
rect 12256 20961 12265 20995
rect 12265 20961 12299 20995
rect 12299 20961 12308 20995
rect 12256 20952 12308 20961
rect 12532 20995 12584 21004
rect 12532 20961 12541 20995
rect 12541 20961 12575 20995
rect 12575 20961 12584 20995
rect 12532 20952 12584 20961
rect 13820 20952 13872 21004
rect 16028 20995 16080 21004
rect 16028 20961 16037 20995
rect 16037 20961 16071 20995
rect 16071 20961 16080 20995
rect 16028 20952 16080 20961
rect 16304 20952 16356 21004
rect 24768 21020 24820 21072
rect 25872 21020 25924 21072
rect 28264 21131 28316 21140
rect 28264 21097 28273 21131
rect 28273 21097 28307 21131
rect 28307 21097 28316 21131
rect 28264 21088 28316 21097
rect 28448 21088 28500 21140
rect 5816 20859 5868 20868
rect 5816 20825 5825 20859
rect 5825 20825 5859 20859
rect 5859 20825 5868 20859
rect 10508 20927 10560 20936
rect 10508 20893 10517 20927
rect 10517 20893 10551 20927
rect 10551 20893 10560 20927
rect 10508 20884 10560 20893
rect 11152 20884 11204 20936
rect 12072 20884 12124 20936
rect 12624 20884 12676 20936
rect 15936 20884 15988 20936
rect 16396 20927 16448 20936
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 16396 20884 16448 20893
rect 16488 20884 16540 20936
rect 5816 20816 5868 20825
rect 6920 20748 6972 20800
rect 12900 20748 12952 20800
rect 14188 20816 14240 20868
rect 15844 20859 15896 20868
rect 15844 20825 15853 20859
rect 15853 20825 15887 20859
rect 15887 20825 15896 20859
rect 15844 20816 15896 20825
rect 16856 20816 16908 20868
rect 16212 20748 16264 20800
rect 17132 20884 17184 20936
rect 17960 20884 18012 20936
rect 18972 20884 19024 20936
rect 23940 20952 23992 21004
rect 20260 20884 20312 20936
rect 21640 20884 21692 20936
rect 27160 20952 27212 21004
rect 24860 20927 24912 20936
rect 24860 20893 24869 20927
rect 24869 20893 24903 20927
rect 24903 20893 24912 20927
rect 24860 20884 24912 20893
rect 27528 20952 27580 21004
rect 29276 21088 29328 21140
rect 29368 21088 29420 21140
rect 39120 21088 39172 21140
rect 27436 20884 27488 20936
rect 35808 21020 35860 21072
rect 29552 20995 29604 21004
rect 29552 20961 29561 20995
rect 29561 20961 29595 20995
rect 29595 20961 29604 20995
rect 29552 20952 29604 20961
rect 30288 20952 30340 21004
rect 28908 20884 28960 20936
rect 29000 20927 29052 20936
rect 29000 20893 29009 20927
rect 29009 20893 29043 20927
rect 29043 20893 29052 20927
rect 29000 20884 29052 20893
rect 31300 20952 31352 21004
rect 28172 20816 28224 20868
rect 31208 20884 31260 20936
rect 31484 20884 31536 20936
rect 31300 20859 31352 20868
rect 31300 20825 31309 20859
rect 31309 20825 31343 20859
rect 31343 20825 31352 20859
rect 31300 20816 31352 20825
rect 17040 20748 17092 20800
rect 17868 20748 17920 20800
rect 18328 20748 18380 20800
rect 19892 20791 19944 20800
rect 19892 20757 19901 20791
rect 19901 20757 19935 20791
rect 19935 20757 19944 20791
rect 19892 20748 19944 20757
rect 19984 20748 20036 20800
rect 25044 20791 25096 20800
rect 25044 20757 25053 20791
rect 25053 20757 25087 20791
rect 25087 20757 25096 20791
rect 25044 20748 25096 20757
rect 25872 20748 25924 20800
rect 26424 20748 26476 20800
rect 27160 20791 27212 20800
rect 27160 20757 27169 20791
rect 27169 20757 27203 20791
rect 27203 20757 27212 20791
rect 27160 20748 27212 20757
rect 28540 20791 28592 20800
rect 28540 20757 28549 20791
rect 28549 20757 28583 20791
rect 28583 20757 28592 20791
rect 28540 20748 28592 20757
rect 28908 20791 28960 20800
rect 28908 20757 28917 20791
rect 28917 20757 28951 20791
rect 28951 20757 28960 20791
rect 28908 20748 28960 20757
rect 34520 20952 34572 21004
rect 35256 20884 35308 20936
rect 35900 20893 35903 20902
rect 35903 20893 35937 20902
rect 35937 20893 35952 20902
rect 35532 20816 35584 20868
rect 35900 20850 35952 20893
rect 35992 20927 36044 20936
rect 35992 20893 36001 20927
rect 36001 20893 36035 20927
rect 36035 20893 36044 20927
rect 35992 20884 36044 20893
rect 37648 20816 37700 20868
rect 38568 20816 38620 20868
rect 38844 20859 38896 20868
rect 38844 20825 38853 20859
rect 38853 20825 38887 20859
rect 38887 20825 38896 20859
rect 38844 20816 38896 20825
rect 39028 20859 39080 20868
rect 39028 20825 39037 20859
rect 39037 20825 39071 20859
rect 39071 20825 39080 20859
rect 39028 20816 39080 20825
rect 32404 20791 32456 20800
rect 32404 20757 32413 20791
rect 32413 20757 32447 20791
rect 32447 20757 32456 20791
rect 32404 20748 32456 20757
rect 34704 20748 34756 20800
rect 34796 20748 34848 20800
rect 35808 20791 35860 20800
rect 35808 20757 35817 20791
rect 35817 20757 35851 20791
rect 35851 20757 35860 20791
rect 35808 20748 35860 20757
rect 36084 20791 36136 20800
rect 36084 20757 36093 20791
rect 36093 20757 36127 20791
rect 36127 20757 36136 20791
rect 36084 20748 36136 20757
rect 36176 20748 36228 20800
rect 36452 20748 36504 20800
rect 37096 20748 37148 20800
rect 39212 20791 39264 20800
rect 39212 20757 39221 20791
rect 39221 20757 39255 20791
rect 39255 20757 39264 20791
rect 39212 20748 39264 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 41512 20680 41564 20732
rect 12716 20544 12768 20596
rect 8576 20408 8628 20460
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 12164 20408 12216 20417
rect 12256 20451 12308 20460
rect 12256 20417 12265 20451
rect 12265 20417 12299 20451
rect 12299 20417 12308 20451
rect 12256 20408 12308 20417
rect 12532 20408 12584 20460
rect 12624 20408 12676 20460
rect 12992 20519 13044 20528
rect 12992 20485 13001 20519
rect 13001 20485 13035 20519
rect 13035 20485 13044 20519
rect 12992 20476 13044 20485
rect 12900 20408 12952 20460
rect 15016 20587 15068 20596
rect 15016 20553 15025 20587
rect 15025 20553 15059 20587
rect 15059 20553 15068 20587
rect 15016 20544 15068 20553
rect 15936 20544 15988 20596
rect 13544 20408 13596 20460
rect 14832 20451 14884 20460
rect 14832 20417 14841 20451
rect 14841 20417 14875 20451
rect 14875 20417 14884 20451
rect 14832 20408 14884 20417
rect 15752 20408 15804 20460
rect 15844 20408 15896 20460
rect 16488 20408 16540 20460
rect 4896 20272 4948 20324
rect 14188 20272 14240 20324
rect 16212 20383 16264 20392
rect 16212 20349 16221 20383
rect 16221 20349 16255 20383
rect 16255 20349 16264 20383
rect 16212 20340 16264 20349
rect 16304 20383 16356 20392
rect 16304 20349 16313 20383
rect 16313 20349 16347 20383
rect 16347 20349 16356 20383
rect 16304 20340 16356 20349
rect 17408 20519 17460 20528
rect 17408 20485 17417 20519
rect 17417 20485 17451 20519
rect 17451 20485 17460 20519
rect 17408 20476 17460 20485
rect 20444 20544 20496 20596
rect 20720 20544 20772 20596
rect 21916 20544 21968 20596
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 17316 20451 17368 20460
rect 17316 20417 17325 20451
rect 17325 20417 17359 20451
rect 17359 20417 17368 20451
rect 17316 20408 17368 20417
rect 17776 20408 17828 20460
rect 18972 20408 19024 20460
rect 19064 20451 19116 20460
rect 19064 20417 19073 20451
rect 19073 20417 19107 20451
rect 19107 20417 19116 20451
rect 19064 20408 19116 20417
rect 17960 20383 18012 20392
rect 17960 20349 17969 20383
rect 17969 20349 18003 20383
rect 18003 20349 18012 20383
rect 17960 20340 18012 20349
rect 19524 20451 19576 20460
rect 19524 20417 19533 20451
rect 19533 20417 19567 20451
rect 19567 20417 19576 20451
rect 19524 20408 19576 20417
rect 20996 20519 21048 20528
rect 20996 20485 21005 20519
rect 21005 20485 21039 20519
rect 21039 20485 21048 20519
rect 21824 20519 21876 20528
rect 20996 20476 21048 20485
rect 21824 20485 21833 20519
rect 21833 20485 21867 20519
rect 21867 20485 21876 20519
rect 21824 20476 21876 20485
rect 19984 20340 20036 20392
rect 20628 20408 20680 20460
rect 21364 20451 21416 20460
rect 21364 20417 21373 20451
rect 21373 20417 21407 20451
rect 21407 20417 21416 20451
rect 21364 20408 21416 20417
rect 21732 20408 21784 20460
rect 25228 20544 25280 20596
rect 26148 20587 26200 20596
rect 26148 20553 26157 20587
rect 26157 20553 26191 20587
rect 26191 20553 26200 20587
rect 26148 20544 26200 20553
rect 32404 20544 32456 20596
rect 32496 20544 32548 20596
rect 35348 20544 35400 20596
rect 35624 20544 35676 20596
rect 38844 20544 38896 20596
rect 22560 20476 22612 20528
rect 25044 20476 25096 20528
rect 27160 20476 27212 20528
rect 28540 20519 28592 20528
rect 28540 20485 28549 20519
rect 28549 20485 28583 20519
rect 28583 20485 28592 20519
rect 28540 20476 28592 20485
rect 30288 20519 30340 20528
rect 30288 20485 30297 20519
rect 30297 20485 30331 20519
rect 30331 20485 30340 20519
rect 30288 20476 30340 20485
rect 26792 20408 26844 20460
rect 22100 20340 22152 20392
rect 22652 20340 22704 20392
rect 25136 20340 25188 20392
rect 17684 20272 17736 20324
rect 19616 20272 19668 20324
rect 5264 20247 5316 20256
rect 5264 20213 5273 20247
rect 5273 20213 5307 20247
rect 5307 20213 5316 20247
rect 5264 20204 5316 20213
rect 13268 20247 13320 20256
rect 13268 20213 13277 20247
rect 13277 20213 13311 20247
rect 13311 20213 13320 20247
rect 13268 20204 13320 20213
rect 14280 20247 14332 20256
rect 14280 20213 14289 20247
rect 14289 20213 14323 20247
rect 14323 20213 14332 20247
rect 14280 20204 14332 20213
rect 15936 20247 15988 20256
rect 15936 20213 15945 20247
rect 15945 20213 15979 20247
rect 15979 20213 15988 20247
rect 15936 20204 15988 20213
rect 16856 20204 16908 20256
rect 19156 20204 19208 20256
rect 19340 20204 19392 20256
rect 19800 20204 19852 20256
rect 20996 20204 21048 20256
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 22836 20247 22888 20256
rect 22836 20213 22845 20247
rect 22845 20213 22879 20247
rect 22879 20213 22888 20247
rect 22836 20204 22888 20213
rect 23756 20204 23808 20256
rect 24952 20204 25004 20256
rect 28540 20340 28592 20392
rect 32128 20451 32180 20460
rect 32128 20417 32137 20451
rect 32137 20417 32171 20451
rect 32171 20417 32180 20451
rect 32128 20408 32180 20417
rect 32220 20451 32272 20460
rect 32220 20417 32230 20451
rect 32230 20417 32264 20451
rect 32264 20417 32272 20451
rect 32220 20408 32272 20417
rect 25412 20247 25464 20256
rect 25412 20213 25421 20247
rect 25421 20213 25455 20247
rect 25455 20213 25464 20247
rect 25412 20204 25464 20213
rect 26608 20204 26660 20256
rect 27160 20204 27212 20256
rect 30840 20204 30892 20256
rect 31760 20204 31812 20256
rect 32496 20451 32548 20460
rect 32496 20417 32505 20451
rect 32505 20417 32539 20451
rect 32539 20417 32548 20451
rect 32496 20408 32548 20417
rect 33140 20476 33192 20528
rect 32772 20408 32824 20460
rect 35900 20408 35952 20460
rect 36176 20408 36228 20460
rect 33600 20383 33652 20392
rect 33600 20349 33609 20383
rect 33609 20349 33643 20383
rect 33643 20349 33652 20383
rect 33600 20340 33652 20349
rect 35348 20383 35400 20392
rect 35348 20349 35357 20383
rect 35357 20349 35391 20383
rect 35391 20349 35400 20383
rect 35348 20340 35400 20349
rect 35532 20340 35584 20392
rect 36544 20451 36596 20460
rect 36544 20417 36553 20451
rect 36553 20417 36587 20451
rect 36587 20417 36596 20451
rect 36544 20408 36596 20417
rect 36728 20451 36780 20460
rect 36728 20417 36737 20451
rect 36737 20417 36771 20451
rect 36771 20417 36780 20451
rect 36728 20408 36780 20417
rect 37372 20408 37424 20460
rect 39120 20476 39172 20528
rect 34704 20272 34756 20324
rect 33968 20204 34020 20256
rect 34612 20204 34664 20256
rect 37280 20315 37332 20324
rect 37280 20281 37289 20315
rect 37289 20281 37323 20315
rect 37323 20281 37332 20315
rect 37280 20272 37332 20281
rect 37832 20383 37884 20392
rect 37832 20349 37841 20383
rect 37841 20349 37875 20383
rect 37875 20349 37884 20383
rect 37832 20340 37884 20349
rect 38384 20383 38436 20392
rect 38384 20349 38393 20383
rect 38393 20349 38427 20383
rect 38427 20349 38436 20383
rect 38384 20340 38436 20349
rect 38660 20383 38712 20392
rect 38660 20349 38669 20383
rect 38669 20349 38703 20383
rect 38703 20349 38712 20383
rect 38660 20340 38712 20349
rect 39028 20204 39080 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6644 20043 6696 20052
rect 6644 20009 6653 20043
rect 6653 20009 6687 20043
rect 6687 20009 6696 20043
rect 6644 20000 6696 20009
rect 13084 20000 13136 20052
rect 13268 20000 13320 20052
rect 13544 20000 13596 20052
rect 7196 19932 7248 19984
rect 9588 19932 9640 19984
rect 10048 19932 10100 19984
rect 10324 19932 10376 19984
rect 11612 19932 11664 19984
rect 6920 19864 6972 19916
rect 10600 19864 10652 19916
rect 4804 19796 4856 19848
rect 5172 19796 5224 19848
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 940 19728 992 19780
rect 1676 19771 1728 19780
rect 1676 19737 1685 19771
rect 1685 19737 1719 19771
rect 1719 19737 1728 19771
rect 1676 19728 1728 19737
rect 6828 19796 6880 19848
rect 7196 19839 7248 19848
rect 7196 19805 7205 19839
rect 7205 19805 7239 19839
rect 7239 19805 7248 19839
rect 7196 19796 7248 19805
rect 7380 19796 7432 19848
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 4712 19703 4764 19712
rect 4712 19669 4721 19703
rect 4721 19669 4755 19703
rect 4755 19669 4764 19703
rect 4712 19660 4764 19669
rect 4988 19660 5040 19712
rect 6828 19703 6880 19712
rect 6828 19669 6837 19703
rect 6837 19669 6871 19703
rect 6871 19669 6880 19703
rect 6828 19660 6880 19669
rect 7196 19660 7248 19712
rect 8208 19728 8260 19780
rect 8944 19728 8996 19780
rect 9404 19660 9456 19712
rect 11244 19728 11296 19780
rect 12624 19796 12676 19848
rect 12808 19839 12860 19848
rect 12808 19805 12817 19839
rect 12817 19805 12851 19839
rect 12851 19805 12860 19839
rect 12808 19796 12860 19805
rect 12900 19796 12952 19848
rect 13912 19932 13964 19984
rect 16120 20000 16172 20052
rect 16672 20000 16724 20052
rect 16856 20000 16908 20052
rect 14280 19907 14332 19916
rect 14280 19873 14289 19907
rect 14289 19873 14323 19907
rect 14323 19873 14332 19907
rect 14280 19864 14332 19873
rect 13820 19839 13872 19848
rect 13820 19805 13829 19839
rect 13829 19805 13863 19839
rect 13863 19805 13872 19839
rect 13820 19796 13872 19805
rect 14004 19796 14056 19848
rect 16120 19864 16172 19916
rect 16948 19864 17000 19916
rect 11428 19728 11480 19780
rect 11796 19771 11848 19780
rect 11796 19737 11805 19771
rect 11805 19737 11839 19771
rect 11839 19737 11848 19771
rect 11796 19728 11848 19737
rect 16580 19839 16632 19848
rect 16580 19805 16589 19839
rect 16589 19805 16623 19839
rect 16623 19805 16632 19839
rect 16580 19796 16632 19805
rect 17224 19864 17276 19916
rect 16212 19771 16264 19780
rect 16212 19737 16221 19771
rect 16221 19737 16255 19771
rect 16255 19737 16264 19771
rect 16212 19728 16264 19737
rect 17408 19796 17460 19848
rect 19064 20000 19116 20052
rect 19156 20000 19208 20052
rect 22284 20000 22336 20052
rect 23848 20000 23900 20052
rect 25504 20000 25556 20052
rect 27252 20000 27304 20052
rect 27528 20043 27580 20052
rect 27528 20009 27537 20043
rect 27537 20009 27571 20043
rect 27571 20009 27580 20043
rect 27528 20000 27580 20009
rect 31484 20043 31536 20052
rect 31484 20009 31493 20043
rect 31493 20009 31527 20043
rect 31527 20009 31536 20043
rect 31484 20000 31536 20009
rect 31760 20000 31812 20052
rect 33140 20000 33192 20052
rect 33600 20000 33652 20052
rect 34704 20000 34756 20052
rect 34980 20000 35032 20052
rect 35900 20000 35952 20052
rect 36176 20043 36228 20052
rect 36176 20009 36185 20043
rect 36185 20009 36219 20043
rect 36219 20009 36228 20043
rect 36176 20000 36228 20009
rect 36728 20000 36780 20052
rect 38660 20000 38712 20052
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 18328 19864 18380 19916
rect 18972 19864 19024 19916
rect 17684 19728 17736 19780
rect 19432 19864 19484 19916
rect 20168 19864 20220 19916
rect 20536 19864 20588 19916
rect 19800 19839 19852 19848
rect 19800 19805 19809 19839
rect 19809 19805 19843 19839
rect 19843 19805 19852 19839
rect 19800 19796 19852 19805
rect 19984 19796 20036 19848
rect 20076 19839 20128 19848
rect 20076 19805 20085 19839
rect 20085 19805 20119 19839
rect 20119 19805 20128 19839
rect 20076 19796 20128 19805
rect 20260 19728 20312 19780
rect 21732 19907 21784 19916
rect 21732 19873 21741 19907
rect 21741 19873 21775 19907
rect 21775 19873 21784 19907
rect 21732 19864 21784 19873
rect 23756 19975 23808 19984
rect 23756 19941 23765 19975
rect 23765 19941 23799 19975
rect 23799 19941 23808 19975
rect 23756 19932 23808 19941
rect 24492 19932 24544 19984
rect 21916 19796 21968 19848
rect 22100 19839 22152 19848
rect 22100 19805 22109 19839
rect 22109 19805 22143 19839
rect 22143 19805 22152 19839
rect 22100 19796 22152 19805
rect 22560 19839 22612 19848
rect 22560 19805 22569 19839
rect 22569 19805 22603 19839
rect 22603 19805 22612 19839
rect 22560 19796 22612 19805
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 23480 19796 23532 19805
rect 14188 19660 14240 19712
rect 14372 19703 14424 19712
rect 14372 19669 14381 19703
rect 14381 19669 14415 19703
rect 14415 19669 14424 19703
rect 14372 19660 14424 19669
rect 17776 19660 17828 19712
rect 17960 19703 18012 19712
rect 17960 19669 17969 19703
rect 17969 19669 18003 19703
rect 18003 19669 18012 19703
rect 17960 19660 18012 19669
rect 19340 19660 19392 19712
rect 20628 19660 20680 19712
rect 21364 19703 21416 19712
rect 21364 19669 21373 19703
rect 21373 19669 21407 19703
rect 21407 19669 21416 19703
rect 21364 19660 21416 19669
rect 22560 19660 22612 19712
rect 23664 19728 23716 19780
rect 25228 19932 25280 19984
rect 23940 19728 23992 19780
rect 23572 19703 23624 19712
rect 23572 19669 23581 19703
rect 23581 19669 23615 19703
rect 23615 19669 23624 19703
rect 23572 19660 23624 19669
rect 23756 19660 23808 19712
rect 24676 19771 24728 19780
rect 24676 19737 24685 19771
rect 24685 19737 24719 19771
rect 24719 19737 24728 19771
rect 24676 19728 24728 19737
rect 24768 19771 24820 19780
rect 24768 19737 24777 19771
rect 24777 19737 24811 19771
rect 24811 19737 24820 19771
rect 24768 19728 24820 19737
rect 25136 19796 25188 19848
rect 25504 19839 25556 19848
rect 25504 19805 25513 19839
rect 25513 19805 25547 19839
rect 25547 19805 25556 19839
rect 25504 19796 25556 19805
rect 26792 19864 26844 19916
rect 27160 19796 27212 19848
rect 28540 19728 28592 19780
rect 31392 19660 31444 19712
rect 32496 19932 32548 19984
rect 34520 19932 34572 19984
rect 32036 19796 32088 19848
rect 35808 19864 35860 19916
rect 33692 19839 33744 19848
rect 33692 19805 33699 19839
rect 33699 19805 33744 19839
rect 33692 19796 33744 19805
rect 33968 19839 34020 19848
rect 33968 19805 33982 19839
rect 33982 19805 34016 19839
rect 34016 19805 34020 19839
rect 33968 19796 34020 19805
rect 34612 19796 34664 19848
rect 34796 19796 34848 19848
rect 34980 19796 35032 19848
rect 35348 19839 35400 19848
rect 35348 19805 35357 19839
rect 35357 19805 35391 19839
rect 35391 19805 35400 19839
rect 35348 19796 35400 19805
rect 36084 19864 36136 19916
rect 37556 19864 37608 19916
rect 38936 19932 38988 19984
rect 33232 19660 33284 19712
rect 33324 19660 33376 19712
rect 33784 19771 33836 19780
rect 33784 19737 33793 19771
rect 33793 19737 33827 19771
rect 33827 19737 33836 19771
rect 33784 19728 33836 19737
rect 36360 19796 36412 19848
rect 37280 19796 37332 19848
rect 37832 19796 37884 19848
rect 39212 19864 39264 19916
rect 34244 19660 34296 19712
rect 37648 19728 37700 19780
rect 38844 19796 38896 19848
rect 39028 19796 39080 19848
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4896 19456 4948 19508
rect 4988 19456 5040 19508
rect 6828 19456 6880 19508
rect 10140 19456 10192 19508
rect 10416 19456 10468 19508
rect 10600 19456 10652 19508
rect 4804 19388 4856 19440
rect 4344 19252 4396 19304
rect 4620 19363 4672 19372
rect 4620 19329 4629 19363
rect 4629 19329 4663 19363
rect 4663 19329 4672 19363
rect 4620 19320 4672 19329
rect 4712 19320 4764 19372
rect 5448 19320 5500 19372
rect 4528 19252 4580 19304
rect 6644 19363 6696 19372
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 7288 19320 7340 19372
rect 6000 19252 6052 19304
rect 5816 19184 5868 19236
rect 3884 19159 3936 19168
rect 3884 19125 3893 19159
rect 3893 19125 3927 19159
rect 3927 19125 3936 19159
rect 3884 19116 3936 19125
rect 4620 19116 4672 19168
rect 4804 19116 4856 19168
rect 5172 19116 5224 19168
rect 6368 19116 6420 19168
rect 7012 19116 7064 19168
rect 7748 19116 7800 19168
rect 8576 19295 8628 19304
rect 8576 19261 8585 19295
rect 8585 19261 8619 19295
rect 8619 19261 8628 19295
rect 8576 19252 8628 19261
rect 8668 19252 8720 19304
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 9312 19363 9364 19372
rect 9312 19329 9321 19363
rect 9321 19329 9355 19363
rect 9355 19329 9364 19363
rect 9312 19320 9364 19329
rect 9404 19320 9456 19372
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 9956 19388 10008 19440
rect 10324 19320 10376 19372
rect 12532 19456 12584 19508
rect 11336 19388 11388 19440
rect 12348 19388 12400 19440
rect 16488 19456 16540 19508
rect 17408 19456 17460 19508
rect 13820 19388 13872 19440
rect 14188 19388 14240 19440
rect 14832 19388 14884 19440
rect 15016 19388 15068 19440
rect 10968 19252 11020 19304
rect 12716 19320 12768 19372
rect 12992 19363 13044 19372
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 14004 19320 14056 19372
rect 9220 19116 9272 19168
rect 9588 19116 9640 19168
rect 10416 19116 10468 19168
rect 11336 19159 11388 19168
rect 11336 19125 11345 19159
rect 11345 19125 11379 19159
rect 11379 19125 11388 19159
rect 11336 19116 11388 19125
rect 11796 19184 11848 19236
rect 14280 19184 14332 19236
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 16948 19320 17000 19329
rect 17684 19320 17736 19372
rect 20628 19456 20680 19508
rect 24952 19456 25004 19508
rect 25504 19456 25556 19508
rect 31668 19456 31720 19508
rect 17868 19388 17920 19440
rect 20076 19388 20128 19440
rect 18328 19320 18380 19372
rect 19156 19320 19208 19372
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 19432 19320 19484 19372
rect 20168 19363 20220 19372
rect 20168 19329 20177 19363
rect 20177 19329 20211 19363
rect 20211 19329 20220 19363
rect 20168 19320 20220 19329
rect 20260 19363 20312 19372
rect 20260 19329 20269 19363
rect 20269 19329 20303 19363
rect 20303 19329 20312 19363
rect 20260 19320 20312 19329
rect 21640 19320 21692 19372
rect 21732 19320 21784 19372
rect 21824 19363 21876 19372
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 21916 19320 21968 19372
rect 22192 19320 22244 19372
rect 22284 19363 22336 19372
rect 22284 19329 22293 19363
rect 22293 19329 22327 19363
rect 22327 19329 22336 19363
rect 22284 19320 22336 19329
rect 22652 19320 22704 19372
rect 27436 19431 27488 19440
rect 20720 19252 20772 19304
rect 22376 19252 22428 19304
rect 16396 19184 16448 19236
rect 21732 19184 21784 19236
rect 22284 19184 22336 19236
rect 22836 19252 22888 19304
rect 23480 19252 23532 19304
rect 24032 19252 24084 19304
rect 24952 19320 25004 19372
rect 27436 19397 27445 19431
rect 27445 19397 27479 19431
rect 27479 19397 27488 19431
rect 27436 19388 27488 19397
rect 31760 19388 31812 19440
rect 33232 19388 33284 19440
rect 34244 19456 34296 19508
rect 25044 19252 25096 19304
rect 26516 19320 26568 19372
rect 27712 19320 27764 19372
rect 25964 19252 26016 19304
rect 26700 19184 26752 19236
rect 28632 19320 28684 19372
rect 29184 19320 29236 19372
rect 31484 19320 31536 19372
rect 37372 19320 37424 19372
rect 39120 19320 39172 19372
rect 40040 19320 40092 19372
rect 29276 19252 29328 19304
rect 29552 19252 29604 19304
rect 30196 19295 30248 19304
rect 30196 19261 30205 19295
rect 30205 19261 30239 19295
rect 30239 19261 30248 19295
rect 30196 19252 30248 19261
rect 30288 19252 30340 19304
rect 35992 19252 36044 19304
rect 37280 19252 37332 19304
rect 36084 19184 36136 19236
rect 11888 19159 11940 19168
rect 11888 19125 11897 19159
rect 11897 19125 11931 19159
rect 11931 19125 11940 19159
rect 11888 19116 11940 19125
rect 12624 19116 12676 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 15568 19116 15620 19168
rect 16856 19116 16908 19168
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 18052 19116 18104 19168
rect 18788 19116 18840 19168
rect 24676 19116 24728 19168
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 26976 19159 27028 19168
rect 26976 19125 26985 19159
rect 26985 19125 27019 19159
rect 27019 19125 27028 19159
rect 26976 19116 27028 19125
rect 29000 19116 29052 19168
rect 30288 19116 30340 19168
rect 30380 19116 30432 19168
rect 31392 19116 31444 19168
rect 32220 19159 32272 19168
rect 32220 19125 32229 19159
rect 32229 19125 32263 19159
rect 32263 19125 32272 19159
rect 32220 19116 32272 19125
rect 32864 19116 32916 19168
rect 33968 19116 34020 19168
rect 34152 19159 34204 19168
rect 34152 19125 34161 19159
rect 34161 19125 34195 19159
rect 34195 19125 34204 19159
rect 34152 19116 34204 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4528 18912 4580 18964
rect 6920 18912 6972 18964
rect 11520 18912 11572 18964
rect 15200 18912 15252 18964
rect 16028 18912 16080 18964
rect 3884 18776 3936 18828
rect 4528 18819 4580 18828
rect 4528 18785 4537 18819
rect 4537 18785 4571 18819
rect 4571 18785 4580 18819
rect 4528 18776 4580 18785
rect 4896 18819 4948 18828
rect 4896 18785 4905 18819
rect 4905 18785 4939 18819
rect 4939 18785 4948 18819
rect 4896 18776 4948 18785
rect 5356 18819 5408 18828
rect 5356 18785 5365 18819
rect 5365 18785 5399 18819
rect 5399 18785 5408 18819
rect 5356 18776 5408 18785
rect 4344 18751 4396 18760
rect 4344 18717 4353 18751
rect 4353 18717 4387 18751
rect 4387 18717 4396 18751
rect 4344 18708 4396 18717
rect 5448 18708 5500 18760
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 5816 18844 5868 18896
rect 6828 18844 6880 18896
rect 8208 18844 8260 18896
rect 6368 18776 6420 18828
rect 3884 18615 3936 18624
rect 3884 18581 3893 18615
rect 3893 18581 3927 18615
rect 3927 18581 3936 18615
rect 3884 18572 3936 18581
rect 6368 18640 6420 18692
rect 6552 18683 6604 18692
rect 6552 18649 6571 18683
rect 6571 18649 6604 18683
rect 6552 18640 6604 18649
rect 6828 18683 6880 18692
rect 6828 18649 6837 18683
rect 6837 18649 6871 18683
rect 6871 18649 6880 18683
rect 6828 18640 6880 18649
rect 7288 18708 7340 18760
rect 7380 18751 7432 18760
rect 7380 18717 7389 18751
rect 7389 18717 7423 18751
rect 7423 18717 7432 18751
rect 7380 18708 7432 18717
rect 7472 18683 7524 18692
rect 7472 18649 7481 18683
rect 7481 18649 7515 18683
rect 7515 18649 7524 18683
rect 7472 18640 7524 18649
rect 7748 18708 7800 18760
rect 7932 18751 7984 18760
rect 7932 18717 7941 18751
rect 7941 18717 7975 18751
rect 7975 18717 7984 18751
rect 7932 18708 7984 18717
rect 8668 18844 8720 18896
rect 9220 18844 9272 18896
rect 9864 18844 9916 18896
rect 17684 18912 17736 18964
rect 18144 18912 18196 18964
rect 18696 18955 18748 18964
rect 18696 18921 18705 18955
rect 18705 18921 18739 18955
rect 18739 18921 18748 18955
rect 18696 18912 18748 18921
rect 19892 18955 19944 18964
rect 19892 18921 19901 18955
rect 19901 18921 19935 18955
rect 19935 18921 19944 18955
rect 19892 18912 19944 18921
rect 20260 18912 20312 18964
rect 9312 18683 9364 18692
rect 9312 18649 9321 18683
rect 9321 18649 9355 18683
rect 9355 18649 9364 18683
rect 9312 18640 9364 18649
rect 9496 18640 9548 18692
rect 10416 18640 10468 18692
rect 4988 18572 5040 18624
rect 6736 18572 6788 18624
rect 7196 18572 7248 18624
rect 8576 18572 8628 18624
rect 10968 18572 11020 18624
rect 11980 18572 12032 18624
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12440 18708 12492 18717
rect 12624 18751 12676 18760
rect 12624 18717 12633 18751
rect 12633 18717 12667 18751
rect 12667 18717 12676 18751
rect 16396 18819 16448 18828
rect 16396 18785 16405 18819
rect 16405 18785 16439 18819
rect 16439 18785 16448 18819
rect 16396 18776 16448 18785
rect 16580 18819 16632 18828
rect 16580 18785 16589 18819
rect 16589 18785 16623 18819
rect 16623 18785 16632 18819
rect 16580 18776 16632 18785
rect 16672 18819 16724 18828
rect 16672 18785 16681 18819
rect 16681 18785 16715 18819
rect 16715 18785 16724 18819
rect 16672 18776 16724 18785
rect 17868 18844 17920 18896
rect 22376 18912 22428 18964
rect 22468 18912 22520 18964
rect 23296 18912 23348 18964
rect 21548 18844 21600 18896
rect 22928 18844 22980 18896
rect 12624 18708 12676 18717
rect 13912 18708 13964 18760
rect 12256 18640 12308 18692
rect 13084 18572 13136 18624
rect 14832 18708 14884 18760
rect 15016 18708 15068 18760
rect 16212 18708 16264 18760
rect 15292 18640 15344 18692
rect 17500 18708 17552 18760
rect 18880 18776 18932 18828
rect 21916 18776 21968 18828
rect 23664 18844 23716 18896
rect 24400 18844 24452 18896
rect 23388 18776 23440 18828
rect 23480 18776 23532 18828
rect 19432 18708 19484 18760
rect 20168 18708 20220 18760
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 23572 18708 23624 18760
rect 23664 18708 23716 18760
rect 24216 18751 24268 18760
rect 24216 18717 24225 18751
rect 24225 18717 24259 18751
rect 24259 18717 24268 18751
rect 24216 18708 24268 18717
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 25044 18751 25096 18760
rect 25044 18717 25053 18751
rect 25053 18717 25087 18751
rect 25087 18717 25096 18751
rect 25044 18708 25096 18717
rect 27252 18844 27304 18896
rect 29552 18912 29604 18964
rect 33784 18912 33836 18964
rect 33876 18912 33928 18964
rect 15476 18572 15528 18624
rect 17500 18572 17552 18624
rect 17776 18615 17828 18624
rect 17776 18581 17785 18615
rect 17785 18581 17819 18615
rect 17819 18581 17828 18615
rect 17776 18572 17828 18581
rect 18052 18572 18104 18624
rect 19064 18572 19116 18624
rect 21364 18572 21416 18624
rect 24492 18640 24544 18692
rect 22652 18572 22704 18624
rect 23296 18615 23348 18624
rect 23296 18581 23305 18615
rect 23305 18581 23339 18615
rect 23339 18581 23348 18615
rect 23296 18572 23348 18581
rect 23572 18615 23624 18624
rect 23572 18581 23581 18615
rect 23581 18581 23615 18615
rect 23615 18581 23624 18615
rect 23572 18572 23624 18581
rect 24308 18572 24360 18624
rect 25228 18640 25280 18692
rect 29276 18776 29328 18828
rect 26976 18708 27028 18760
rect 30288 18776 30340 18828
rect 33232 18819 33284 18828
rect 33232 18785 33241 18819
rect 33241 18785 33275 18819
rect 33275 18785 33284 18819
rect 33232 18776 33284 18785
rect 30380 18708 30432 18760
rect 31484 18708 31536 18760
rect 27160 18572 27212 18624
rect 28540 18640 28592 18692
rect 32220 18751 32272 18760
rect 32220 18717 32229 18751
rect 32229 18717 32263 18751
rect 32263 18717 32272 18751
rect 32220 18708 32272 18717
rect 33140 18751 33192 18760
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 33140 18708 33192 18717
rect 33784 18751 33836 18760
rect 33784 18717 33793 18751
rect 33793 18717 33827 18751
rect 33827 18717 33836 18751
rect 33784 18708 33836 18717
rect 33968 18751 34020 18760
rect 33968 18717 33977 18751
rect 33977 18717 34011 18751
rect 34011 18717 34020 18751
rect 33968 18708 34020 18717
rect 34336 18708 34388 18760
rect 35808 18912 35860 18964
rect 37648 18912 37700 18964
rect 38568 18912 38620 18964
rect 37372 18776 37424 18828
rect 36084 18708 36136 18760
rect 36820 18751 36872 18760
rect 36820 18717 36829 18751
rect 36829 18717 36863 18751
rect 36863 18717 36872 18751
rect 36820 18708 36872 18717
rect 39672 18776 39724 18828
rect 29552 18615 29604 18624
rect 29552 18581 29561 18615
rect 29561 18581 29595 18615
rect 29595 18581 29604 18615
rect 29552 18572 29604 18581
rect 29644 18572 29696 18624
rect 30656 18572 30708 18624
rect 31944 18572 31996 18624
rect 32036 18615 32088 18624
rect 32036 18581 32045 18615
rect 32045 18581 32079 18615
rect 32079 18581 32088 18615
rect 32036 18572 32088 18581
rect 33324 18572 33376 18624
rect 34152 18572 34204 18624
rect 35992 18572 36044 18624
rect 36728 18640 36780 18692
rect 37096 18683 37148 18692
rect 37096 18649 37131 18683
rect 37131 18649 37148 18683
rect 37096 18640 37148 18649
rect 39304 18683 39356 18692
rect 39304 18649 39313 18683
rect 39313 18649 39347 18683
rect 39347 18649 39356 18683
rect 39304 18640 39356 18649
rect 38752 18572 38804 18624
rect 39856 18615 39908 18624
rect 39856 18581 39865 18615
rect 39865 18581 39899 18615
rect 39899 18581 39908 18615
rect 39856 18572 39908 18581
rect 40960 18572 41012 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1492 18368 1544 18420
rect 4068 18368 4120 18420
rect 4988 18368 5040 18420
rect 5172 18368 5224 18420
rect 3056 18300 3108 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 5540 18368 5592 18420
rect 5448 18343 5500 18352
rect 5448 18309 5457 18343
rect 5457 18309 5491 18343
rect 5491 18309 5500 18343
rect 5448 18300 5500 18309
rect 4988 18232 5040 18241
rect 6000 18368 6052 18420
rect 7932 18368 7984 18420
rect 8024 18368 8076 18420
rect 11244 18368 11296 18420
rect 11980 18411 12032 18420
rect 11980 18377 11989 18411
rect 11989 18377 12023 18411
rect 12023 18377 12032 18411
rect 11980 18368 12032 18377
rect 7380 18300 7432 18352
rect 11060 18300 11112 18352
rect 7196 18232 7248 18284
rect 8392 18232 8444 18284
rect 9128 18232 9180 18284
rect 9588 18232 9640 18284
rect 10508 18275 10560 18284
rect 10508 18241 10517 18275
rect 10517 18241 10551 18275
rect 10551 18241 10560 18275
rect 10508 18232 10560 18241
rect 11336 18232 11388 18284
rect 14648 18368 14700 18420
rect 15476 18368 15528 18420
rect 12256 18232 12308 18284
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 5540 18164 5592 18216
rect 7932 18096 7984 18148
rect 10600 18207 10652 18216
rect 10600 18173 10609 18207
rect 10609 18173 10643 18207
rect 10643 18173 10652 18207
rect 10600 18164 10652 18173
rect 4528 18028 4580 18080
rect 4804 18028 4856 18080
rect 5356 18028 5408 18080
rect 7288 18028 7340 18080
rect 8300 18028 8352 18080
rect 12164 18096 12216 18148
rect 11336 18028 11388 18080
rect 14372 18232 14424 18284
rect 15384 18300 15436 18352
rect 15292 18275 15344 18284
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 15568 18275 15620 18284
rect 15568 18241 15577 18275
rect 15577 18241 15611 18275
rect 15611 18241 15620 18275
rect 15568 18232 15620 18241
rect 16580 18232 16632 18284
rect 16764 18232 16816 18284
rect 17684 18275 17736 18284
rect 17684 18241 17693 18275
rect 17693 18241 17727 18275
rect 17727 18241 17736 18275
rect 17684 18232 17736 18241
rect 17776 18275 17828 18284
rect 17776 18241 17785 18275
rect 17785 18241 17819 18275
rect 17819 18241 17828 18275
rect 17776 18232 17828 18241
rect 18236 18275 18288 18284
rect 18236 18241 18245 18275
rect 18245 18241 18279 18275
rect 18279 18241 18288 18275
rect 18236 18232 18288 18241
rect 23388 18368 23440 18420
rect 24032 18411 24084 18420
rect 24032 18377 24041 18411
rect 24041 18377 24075 18411
rect 24075 18377 24084 18411
rect 24032 18368 24084 18377
rect 24584 18368 24636 18420
rect 15108 18139 15160 18148
rect 15108 18105 15117 18139
rect 15117 18105 15151 18139
rect 15151 18105 15160 18139
rect 15108 18096 15160 18105
rect 15752 18096 15804 18148
rect 17132 18096 17184 18148
rect 18328 18096 18380 18148
rect 23112 18300 23164 18352
rect 18880 18232 18932 18284
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 19248 18275 19300 18284
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 19432 18232 19484 18284
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 20076 18232 20128 18284
rect 20260 18275 20312 18284
rect 20260 18241 20269 18275
rect 20269 18241 20303 18275
rect 20303 18241 20312 18275
rect 20260 18232 20312 18241
rect 20352 18232 20404 18284
rect 21548 18232 21600 18284
rect 22284 18232 22336 18284
rect 23020 18275 23072 18284
rect 23020 18241 23029 18275
rect 23029 18241 23063 18275
rect 23063 18241 23072 18275
rect 23020 18232 23072 18241
rect 21456 18164 21508 18216
rect 22744 18164 22796 18216
rect 23296 18232 23348 18284
rect 23572 18232 23624 18284
rect 24032 18232 24084 18284
rect 24308 18232 24360 18284
rect 24400 18275 24452 18284
rect 24400 18241 24409 18275
rect 24409 18241 24443 18275
rect 24443 18241 24452 18275
rect 24400 18232 24452 18241
rect 24584 18232 24636 18284
rect 26884 18232 26936 18284
rect 27160 18368 27212 18420
rect 27804 18368 27856 18420
rect 22468 18096 22520 18148
rect 23572 18096 23624 18148
rect 15660 18028 15712 18080
rect 15936 18071 15988 18080
rect 15936 18037 15945 18071
rect 15945 18037 15979 18071
rect 15979 18037 15988 18071
rect 15936 18028 15988 18037
rect 17040 18028 17092 18080
rect 17408 18028 17460 18080
rect 18788 18071 18840 18080
rect 18788 18037 18797 18071
rect 18797 18037 18831 18071
rect 18831 18037 18840 18071
rect 18788 18028 18840 18037
rect 18972 18028 19024 18080
rect 19984 18028 20036 18080
rect 20168 18028 20220 18080
rect 20352 18028 20404 18080
rect 22192 18028 22244 18080
rect 22284 18071 22336 18080
rect 22284 18037 22293 18071
rect 22293 18037 22327 18071
rect 22327 18037 22336 18071
rect 22284 18028 22336 18037
rect 22744 18071 22796 18080
rect 22744 18037 22753 18071
rect 22753 18037 22787 18071
rect 22787 18037 22796 18071
rect 22744 18028 22796 18037
rect 23204 18028 23256 18080
rect 24860 18096 24912 18148
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 27528 18232 27580 18284
rect 27712 18275 27764 18284
rect 27712 18241 27721 18275
rect 27721 18241 27755 18275
rect 27755 18241 27764 18275
rect 27712 18232 27764 18241
rect 27988 18275 28040 18284
rect 27988 18241 27997 18275
rect 27997 18241 28031 18275
rect 28031 18241 28040 18275
rect 27988 18232 28040 18241
rect 28080 18275 28132 18284
rect 28080 18241 28089 18275
rect 28089 18241 28123 18275
rect 28123 18241 28132 18275
rect 28080 18232 28132 18241
rect 28356 18164 28408 18216
rect 29092 18164 29144 18216
rect 29552 18368 29604 18420
rect 30196 18368 30248 18420
rect 32128 18368 32180 18420
rect 33232 18368 33284 18420
rect 34704 18368 34756 18420
rect 35440 18368 35492 18420
rect 36728 18368 36780 18420
rect 36820 18368 36872 18420
rect 32220 18343 32272 18352
rect 32220 18309 32229 18343
rect 32229 18309 32263 18343
rect 32263 18309 32272 18343
rect 32220 18300 32272 18309
rect 30656 18232 30708 18284
rect 31484 18275 31536 18284
rect 31484 18241 31493 18275
rect 31493 18241 31527 18275
rect 31527 18241 31536 18275
rect 31484 18232 31536 18241
rect 31944 18232 31996 18284
rect 34612 18300 34664 18352
rect 33600 18275 33652 18284
rect 33600 18241 33609 18275
rect 33609 18241 33643 18275
rect 33643 18241 33652 18275
rect 33600 18232 33652 18241
rect 33784 18275 33836 18284
rect 33784 18241 33793 18275
rect 33793 18241 33827 18275
rect 33827 18241 33836 18275
rect 33784 18232 33836 18241
rect 33140 18164 33192 18216
rect 34152 18207 34204 18216
rect 34152 18173 34161 18207
rect 34161 18173 34195 18207
rect 34195 18173 34204 18207
rect 34152 18164 34204 18173
rect 35900 18164 35952 18216
rect 36544 18232 36596 18284
rect 38384 18300 38436 18352
rect 39856 18368 39908 18420
rect 40960 18411 41012 18420
rect 40960 18377 40969 18411
rect 40969 18377 41003 18411
rect 41003 18377 41012 18411
rect 40960 18368 41012 18377
rect 37096 18232 37148 18284
rect 37464 18275 37516 18284
rect 37464 18241 37473 18275
rect 37473 18241 37507 18275
rect 37507 18241 37516 18275
rect 37464 18232 37516 18241
rect 38752 18232 38804 18284
rect 40040 18300 40092 18352
rect 37832 18164 37884 18216
rect 38844 18207 38896 18216
rect 38844 18173 38853 18207
rect 38853 18173 38887 18207
rect 38887 18173 38896 18207
rect 38844 18164 38896 18173
rect 39120 18164 39172 18216
rect 26884 18028 26936 18080
rect 27252 18028 27304 18080
rect 27712 18028 27764 18080
rect 30012 18028 30064 18080
rect 30288 18028 30340 18080
rect 33232 18028 33284 18080
rect 33324 18071 33376 18080
rect 33324 18037 33333 18071
rect 33333 18037 33367 18071
rect 33367 18037 33376 18071
rect 33324 18028 33376 18037
rect 33508 18028 33560 18080
rect 33784 18028 33836 18080
rect 34520 18028 34572 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1676 17824 1728 17876
rect 9496 17824 9548 17876
rect 10140 17867 10192 17876
rect 10140 17833 10149 17867
rect 10149 17833 10183 17867
rect 10183 17833 10192 17867
rect 10140 17824 10192 17833
rect 12440 17824 12492 17876
rect 15660 17824 15712 17876
rect 4068 17756 4120 17808
rect 1492 17688 1544 17740
rect 11520 17756 11572 17808
rect 12072 17756 12124 17808
rect 13360 17756 13412 17808
rect 22744 17824 22796 17876
rect 23020 17824 23072 17876
rect 24032 17824 24084 17876
rect 26056 17824 26108 17876
rect 27436 17824 27488 17876
rect 31484 17824 31536 17876
rect 33876 17824 33928 17876
rect 35900 17824 35952 17876
rect 5448 17688 5500 17740
rect 9588 17688 9640 17740
rect 2964 17620 3016 17672
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 9312 17620 9364 17629
rect 10048 17663 10100 17672
rect 10048 17629 10057 17663
rect 10057 17629 10091 17663
rect 10091 17629 10100 17663
rect 10048 17620 10100 17629
rect 11796 17688 11848 17740
rect 12992 17688 13044 17740
rect 10140 17552 10192 17604
rect 11612 17663 11664 17672
rect 11612 17629 11621 17663
rect 11621 17629 11655 17663
rect 11655 17629 11664 17663
rect 11612 17620 11664 17629
rect 11704 17663 11756 17672
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 5540 17484 5592 17536
rect 9036 17484 9088 17536
rect 12256 17620 12308 17672
rect 13820 17620 13872 17672
rect 14556 17688 14608 17740
rect 15568 17688 15620 17740
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 15292 17620 15344 17672
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 18788 17688 18840 17740
rect 19984 17688 20036 17740
rect 13176 17595 13228 17604
rect 13176 17561 13185 17595
rect 13185 17561 13219 17595
rect 13219 17561 13228 17595
rect 13176 17552 13228 17561
rect 14832 17552 14884 17604
rect 16304 17552 16356 17604
rect 17960 17552 18012 17604
rect 18972 17620 19024 17672
rect 18788 17552 18840 17604
rect 19156 17552 19208 17604
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 15200 17484 15252 17536
rect 18420 17484 18472 17536
rect 18972 17484 19024 17536
rect 20076 17552 20128 17604
rect 22376 17688 22428 17740
rect 22560 17663 22612 17672
rect 22560 17629 22569 17663
rect 22569 17629 22603 17663
rect 22603 17629 22612 17663
rect 22560 17620 22612 17629
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 23296 17688 23348 17740
rect 22836 17663 22888 17672
rect 22836 17629 22871 17663
rect 22871 17629 22888 17663
rect 22836 17620 22888 17629
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 24032 17620 24084 17672
rect 26976 17663 27028 17672
rect 26976 17629 26985 17663
rect 26985 17629 27019 17663
rect 27019 17629 27028 17663
rect 26976 17620 27028 17629
rect 27252 17663 27304 17672
rect 27252 17629 27261 17663
rect 27261 17629 27295 17663
rect 27295 17629 27304 17663
rect 27252 17620 27304 17629
rect 27712 17620 27764 17672
rect 29000 17620 29052 17672
rect 26056 17552 26108 17604
rect 30748 17731 30800 17740
rect 30748 17697 30757 17731
rect 30757 17697 30791 17731
rect 30791 17697 30800 17731
rect 30748 17688 30800 17697
rect 31300 17663 31352 17672
rect 31300 17629 31309 17663
rect 31309 17629 31343 17663
rect 31343 17629 31352 17663
rect 31300 17620 31352 17629
rect 33692 17620 33744 17672
rect 34704 17620 34756 17672
rect 35900 17731 35952 17740
rect 35900 17697 35909 17731
rect 35909 17697 35943 17731
rect 35943 17697 35952 17731
rect 35900 17688 35952 17697
rect 36544 17731 36596 17740
rect 36544 17697 36553 17731
rect 36553 17697 36587 17731
rect 36587 17697 36596 17731
rect 36544 17688 36596 17697
rect 20168 17484 20220 17536
rect 21088 17484 21140 17536
rect 23848 17484 23900 17536
rect 24124 17484 24176 17536
rect 26332 17484 26384 17536
rect 26700 17527 26752 17536
rect 26700 17493 26709 17527
rect 26709 17493 26743 17527
rect 26743 17493 26752 17527
rect 26700 17484 26752 17493
rect 34612 17552 34664 17604
rect 35532 17620 35584 17672
rect 38844 17824 38896 17876
rect 28540 17484 28592 17536
rect 29644 17484 29696 17536
rect 34520 17484 34572 17536
rect 36360 17552 36412 17604
rect 40592 17620 40644 17672
rect 37832 17484 37884 17536
rect 39396 17595 39448 17604
rect 39396 17561 39405 17595
rect 39405 17561 39439 17595
rect 39439 17561 39448 17595
rect 39396 17552 39448 17561
rect 40500 17552 40552 17604
rect 39488 17484 39540 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 41512 17416 41564 17468
rect 4896 17280 4948 17332
rect 7196 17280 7248 17332
rect 10140 17280 10192 17332
rect 11612 17280 11664 17332
rect 13176 17280 13228 17332
rect 13268 17280 13320 17332
rect 15384 17280 15436 17332
rect 15568 17280 15620 17332
rect 15660 17323 15712 17332
rect 15660 17289 15669 17323
rect 15669 17289 15703 17323
rect 15703 17289 15712 17323
rect 15660 17280 15712 17289
rect 17592 17280 17644 17332
rect 18420 17280 18472 17332
rect 26976 17280 27028 17332
rect 29644 17280 29696 17332
rect 30656 17323 30708 17332
rect 30656 17289 30665 17323
rect 30665 17289 30699 17323
rect 30699 17289 30708 17323
rect 30656 17280 30708 17289
rect 30748 17280 30800 17332
rect 33324 17280 33376 17332
rect 37372 17280 37424 17332
rect 5816 17212 5868 17264
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 5080 17187 5132 17196
rect 5080 17153 5089 17187
rect 5089 17153 5123 17187
rect 5123 17153 5132 17187
rect 5080 17144 5132 17153
rect 5356 17144 5408 17196
rect 6000 17144 6052 17196
rect 6736 17144 6788 17196
rect 7932 17144 7984 17196
rect 8484 17255 8536 17264
rect 8484 17221 8493 17255
rect 8493 17221 8527 17255
rect 8527 17221 8536 17255
rect 8484 17212 8536 17221
rect 9312 17212 9364 17264
rect 9404 17255 9456 17264
rect 9404 17221 9413 17255
rect 9413 17221 9447 17255
rect 9447 17221 9456 17255
rect 9404 17212 9456 17221
rect 11520 17255 11572 17264
rect 11520 17221 11529 17255
rect 11529 17221 11563 17255
rect 11563 17221 11572 17255
rect 11520 17212 11572 17221
rect 11888 17212 11940 17264
rect 5540 17076 5592 17128
rect 8760 17144 8812 17196
rect 8852 17187 8904 17196
rect 8852 17153 8861 17187
rect 8861 17153 8895 17187
rect 8895 17153 8904 17187
rect 8852 17144 8904 17153
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9036 17144 9088 17153
rect 9128 17187 9180 17196
rect 9128 17153 9163 17187
rect 9163 17153 9180 17187
rect 9128 17144 9180 17153
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 12256 17144 12308 17196
rect 14188 17212 14240 17264
rect 14832 17187 14884 17196
rect 14832 17153 14841 17187
rect 14841 17153 14875 17187
rect 14875 17153 14884 17187
rect 14832 17144 14884 17153
rect 9312 17119 9364 17128
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 13176 17119 13228 17128
rect 13176 17085 13185 17119
rect 13185 17085 13219 17119
rect 13219 17085 13228 17119
rect 13176 17076 13228 17085
rect 7380 17008 7432 17060
rect 8484 17008 8536 17060
rect 8852 17008 8904 17060
rect 10048 17008 10100 17060
rect 12164 17008 12216 17060
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 15292 17187 15344 17196
rect 15292 17153 15306 17187
rect 15306 17153 15340 17187
rect 15340 17153 15344 17187
rect 15292 17144 15344 17153
rect 3424 16940 3476 16992
rect 7472 16940 7524 16992
rect 8116 16940 8168 16992
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 11704 16940 11756 16992
rect 14280 16940 14332 16992
rect 17224 17144 17276 17196
rect 18052 17187 18104 17196
rect 18052 17153 18061 17187
rect 18061 17153 18095 17187
rect 18095 17153 18104 17187
rect 18052 17144 18104 17153
rect 18696 17144 18748 17196
rect 18972 17212 19024 17264
rect 20536 17212 20588 17264
rect 15568 17076 15620 17128
rect 16764 17076 16816 17128
rect 17592 17076 17644 17128
rect 19984 17076 20036 17128
rect 16120 17008 16172 17060
rect 18144 17008 18196 17060
rect 19432 17008 19484 17060
rect 20168 17144 20220 17196
rect 20444 17187 20496 17196
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20996 17212 21048 17264
rect 21272 17212 21324 17264
rect 21732 17212 21784 17264
rect 20444 17144 20496 17153
rect 21824 17144 21876 17196
rect 22100 17212 22152 17264
rect 23112 17187 23164 17196
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 23940 17144 23992 17196
rect 24032 17187 24084 17196
rect 24032 17153 24041 17187
rect 24041 17153 24075 17187
rect 24075 17153 24084 17187
rect 24032 17144 24084 17153
rect 20168 17008 20220 17060
rect 20720 17008 20772 17060
rect 20812 17008 20864 17060
rect 21640 17008 21692 17060
rect 23664 17008 23716 17060
rect 17316 16940 17368 16992
rect 20076 16940 20128 16992
rect 20260 16940 20312 16992
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 21732 16940 21784 16992
rect 22468 16940 22520 16992
rect 23020 16940 23072 16992
rect 23480 16983 23532 16992
rect 23480 16949 23489 16983
rect 23489 16949 23523 16983
rect 23523 16949 23532 16983
rect 23480 16940 23532 16949
rect 24400 17008 24452 17060
rect 25044 17187 25096 17196
rect 25044 17153 25053 17187
rect 25053 17153 25087 17187
rect 25087 17153 25096 17187
rect 25044 17144 25096 17153
rect 27436 17144 27488 17196
rect 29736 17144 29788 17196
rect 30104 17144 30156 17196
rect 30656 17187 30708 17196
rect 30656 17153 30665 17187
rect 30665 17153 30699 17187
rect 30699 17153 30708 17187
rect 30656 17144 30708 17153
rect 30932 17144 30984 17196
rect 25504 16983 25556 16992
rect 25504 16949 25513 16983
rect 25513 16949 25547 16983
rect 25547 16949 25556 16983
rect 25504 16940 25556 16949
rect 26608 16940 26660 16992
rect 26976 16940 27028 16992
rect 29460 16940 29512 16992
rect 29920 16983 29972 16992
rect 29920 16949 29929 16983
rect 29929 16949 29963 16983
rect 29963 16949 29972 16983
rect 31300 17008 31352 17060
rect 29920 16940 29972 16949
rect 31208 16940 31260 16992
rect 36636 17212 36688 17264
rect 33876 17144 33928 17196
rect 37924 17144 37976 17196
rect 38476 17187 38528 17196
rect 38476 17153 38485 17187
rect 38485 17153 38519 17187
rect 38519 17153 38528 17187
rect 38476 17144 38528 17153
rect 39212 17255 39264 17264
rect 33140 17076 33192 17128
rect 33508 17119 33560 17128
rect 33508 17085 33517 17119
rect 33517 17085 33551 17119
rect 33551 17085 33560 17119
rect 33508 17076 33560 17085
rect 33692 17076 33744 17128
rect 33784 17076 33836 17128
rect 39212 17221 39218 17255
rect 39218 17221 39252 17255
rect 39252 17221 39264 17255
rect 39212 17212 39264 17221
rect 32956 17008 33008 17060
rect 38752 17008 38804 17060
rect 40500 17119 40552 17128
rect 40500 17085 40509 17119
rect 40509 17085 40543 17119
rect 40543 17085 40552 17119
rect 40500 17076 40552 17085
rect 39488 17008 39540 17060
rect 33416 16940 33468 16992
rect 34152 16940 34204 16992
rect 34244 16940 34296 16992
rect 36268 16940 36320 16992
rect 38936 16983 38988 16992
rect 38936 16949 38945 16983
rect 38945 16949 38979 16983
rect 38979 16949 38988 16983
rect 38936 16940 38988 16949
rect 39396 16940 39448 16992
rect 41052 16983 41104 16992
rect 41052 16949 41061 16983
rect 41061 16949 41095 16983
rect 41095 16949 41104 16983
rect 41052 16940 41104 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 8668 16736 8720 16788
rect 8760 16736 8812 16788
rect 9312 16736 9364 16788
rect 15200 16736 15252 16788
rect 16028 16736 16080 16788
rect 16120 16736 16172 16788
rect 17776 16779 17828 16788
rect 17776 16745 17785 16779
rect 17785 16745 17819 16779
rect 17819 16745 17828 16779
rect 17776 16736 17828 16745
rect 21456 16736 21508 16788
rect 5080 16668 5132 16720
rect 4712 16643 4764 16652
rect 3792 16532 3844 16584
rect 4068 16575 4120 16584
rect 4068 16541 4077 16575
rect 4077 16541 4111 16575
rect 4111 16541 4120 16575
rect 4068 16532 4120 16541
rect 4344 16532 4396 16584
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 4620 16532 4672 16584
rect 4988 16532 5040 16584
rect 11520 16668 11572 16720
rect 16304 16668 16356 16720
rect 9404 16600 9456 16652
rect 5264 16507 5316 16516
rect 5264 16473 5273 16507
rect 5273 16473 5307 16507
rect 5307 16473 5316 16507
rect 5264 16464 5316 16473
rect 4528 16396 4580 16448
rect 7288 16532 7340 16584
rect 7932 16532 7984 16584
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 8300 16575 8352 16584
rect 8300 16541 8309 16575
rect 8309 16541 8343 16575
rect 8343 16541 8352 16575
rect 8300 16532 8352 16541
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 8484 16532 8536 16584
rect 9588 16600 9640 16652
rect 10784 16600 10836 16652
rect 5540 16464 5592 16516
rect 9772 16532 9824 16584
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 11704 16532 11756 16584
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 12256 16532 12308 16584
rect 12348 16575 12400 16584
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 12348 16532 12400 16541
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 13820 16600 13872 16652
rect 12992 16532 13044 16584
rect 5632 16396 5684 16448
rect 5724 16396 5776 16448
rect 7380 16396 7432 16448
rect 7656 16439 7708 16448
rect 7656 16405 7665 16439
rect 7665 16405 7699 16439
rect 7699 16405 7708 16439
rect 7656 16396 7708 16405
rect 10876 16396 10928 16448
rect 13452 16464 13504 16516
rect 15384 16532 15436 16584
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 19248 16668 19300 16720
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 17592 16600 17644 16652
rect 13268 16396 13320 16448
rect 15200 16396 15252 16448
rect 16028 16396 16080 16448
rect 17040 16532 17092 16584
rect 16488 16507 16540 16516
rect 16488 16473 16523 16507
rect 16523 16473 16540 16507
rect 16488 16464 16540 16473
rect 16764 16464 16816 16516
rect 17316 16464 17368 16516
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 18052 16532 18104 16584
rect 20444 16668 20496 16720
rect 20904 16668 20956 16720
rect 21364 16600 21416 16652
rect 20168 16532 20220 16584
rect 20260 16575 20312 16584
rect 20260 16541 20269 16575
rect 20269 16541 20303 16575
rect 20303 16541 20312 16575
rect 20260 16532 20312 16541
rect 20352 16532 20404 16584
rect 20812 16575 20864 16584
rect 20812 16541 20821 16575
rect 20821 16541 20855 16575
rect 20855 16541 20864 16575
rect 20812 16532 20864 16541
rect 21180 16575 21232 16584
rect 21180 16541 21189 16575
rect 21189 16541 21223 16575
rect 21223 16541 21232 16575
rect 21180 16532 21232 16541
rect 21824 16668 21876 16720
rect 21640 16600 21692 16652
rect 20536 16464 20588 16516
rect 20904 16507 20956 16516
rect 20904 16473 20913 16507
rect 20913 16473 20947 16507
rect 20947 16473 20956 16507
rect 22008 16532 22060 16584
rect 22928 16532 22980 16584
rect 23112 16736 23164 16788
rect 25504 16736 25556 16788
rect 25596 16736 25648 16788
rect 23848 16600 23900 16652
rect 24032 16600 24084 16652
rect 24400 16600 24452 16652
rect 26240 16668 26292 16720
rect 26516 16736 26568 16788
rect 23388 16575 23440 16584
rect 23388 16541 23398 16575
rect 23398 16541 23432 16575
rect 23432 16541 23440 16575
rect 23388 16532 23440 16541
rect 20904 16464 20956 16473
rect 21364 16464 21416 16516
rect 24308 16532 24360 16584
rect 26976 16600 27028 16652
rect 26332 16532 26384 16584
rect 26516 16575 26568 16584
rect 26516 16541 26525 16575
rect 26525 16541 26559 16575
rect 26559 16541 26568 16575
rect 26516 16532 26568 16541
rect 26700 16532 26752 16584
rect 24216 16464 24268 16516
rect 27712 16575 27764 16584
rect 27712 16541 27721 16575
rect 27721 16541 27755 16575
rect 27755 16541 27764 16575
rect 27712 16532 27764 16541
rect 28816 16600 28868 16652
rect 29460 16736 29512 16788
rect 29368 16668 29420 16720
rect 29552 16668 29604 16720
rect 22836 16396 22888 16448
rect 23480 16396 23532 16448
rect 25136 16439 25188 16448
rect 25136 16405 25145 16439
rect 25145 16405 25179 16439
rect 25179 16405 25188 16439
rect 25136 16396 25188 16405
rect 25596 16396 25648 16448
rect 26056 16439 26108 16448
rect 26056 16405 26065 16439
rect 26065 16405 26099 16439
rect 26099 16405 26108 16439
rect 26056 16396 26108 16405
rect 28172 16507 28224 16516
rect 28172 16473 28181 16507
rect 28181 16473 28215 16507
rect 28215 16473 28224 16507
rect 28172 16464 28224 16473
rect 28540 16575 28592 16584
rect 28540 16541 28552 16575
rect 28552 16541 28586 16575
rect 28586 16541 28592 16575
rect 28540 16532 28592 16541
rect 29644 16600 29696 16652
rect 30104 16600 30156 16652
rect 30196 16643 30248 16652
rect 30196 16609 30205 16643
rect 30205 16609 30239 16643
rect 30239 16609 30248 16643
rect 30196 16600 30248 16609
rect 31300 16600 31352 16652
rect 26792 16396 26844 16448
rect 28724 16396 28776 16448
rect 29000 16396 29052 16448
rect 30104 16464 30156 16516
rect 30932 16532 30984 16584
rect 31208 16575 31260 16584
rect 31208 16541 31217 16575
rect 31217 16541 31251 16575
rect 31251 16541 31260 16575
rect 31208 16532 31260 16541
rect 33140 16736 33192 16788
rect 34520 16736 34572 16788
rect 31024 16464 31076 16516
rect 32956 16575 33008 16584
rect 32956 16541 32965 16575
rect 32965 16541 32999 16575
rect 32999 16541 33008 16575
rect 32956 16532 33008 16541
rect 33600 16600 33652 16652
rect 33416 16575 33468 16584
rect 33416 16541 33447 16575
rect 33447 16541 33468 16575
rect 33416 16532 33468 16541
rect 33968 16532 34020 16584
rect 34612 16668 34664 16720
rect 35992 16532 36044 16584
rect 38476 16736 38528 16788
rect 38844 16736 38896 16788
rect 38936 16736 38988 16788
rect 39212 16779 39264 16788
rect 39212 16745 39221 16779
rect 39221 16745 39255 16779
rect 39255 16745 39264 16779
rect 39212 16736 39264 16745
rect 39304 16736 39356 16788
rect 37924 16668 37976 16720
rect 38660 16668 38712 16720
rect 38660 16532 38712 16584
rect 38936 16575 38988 16584
rect 38936 16541 38945 16575
rect 38945 16541 38979 16575
rect 38979 16541 38988 16575
rect 38936 16532 38988 16541
rect 39580 16600 39632 16652
rect 40592 16643 40644 16652
rect 40592 16609 40601 16643
rect 40601 16609 40635 16643
rect 40635 16609 40644 16643
rect 40592 16600 40644 16609
rect 39396 16575 39448 16584
rect 39396 16541 39405 16575
rect 39405 16541 39439 16575
rect 39439 16541 39448 16575
rect 39396 16532 39448 16541
rect 29460 16396 29512 16448
rect 29644 16396 29696 16448
rect 31300 16396 31352 16448
rect 31668 16439 31720 16448
rect 31668 16405 31677 16439
rect 31677 16405 31711 16439
rect 31711 16405 31720 16439
rect 31668 16396 31720 16405
rect 32312 16396 32364 16448
rect 33508 16396 33560 16448
rect 33784 16439 33836 16448
rect 33784 16405 33793 16439
rect 33793 16405 33827 16439
rect 33827 16405 33836 16439
rect 33784 16396 33836 16405
rect 33876 16396 33928 16448
rect 34428 16439 34480 16448
rect 34428 16405 34437 16439
rect 34437 16405 34471 16439
rect 34471 16405 34480 16439
rect 34428 16396 34480 16405
rect 34520 16396 34572 16448
rect 35900 16396 35952 16448
rect 36544 16396 36596 16448
rect 37740 16396 37792 16448
rect 38476 16396 38528 16448
rect 38660 16439 38712 16448
rect 38660 16405 38675 16439
rect 38675 16405 38709 16439
rect 38709 16405 38712 16439
rect 38660 16396 38712 16405
rect 39304 16464 39356 16516
rect 38844 16396 38896 16448
rect 39488 16439 39540 16448
rect 39488 16405 39497 16439
rect 39497 16405 39531 16439
rect 39531 16405 39540 16439
rect 39488 16396 39540 16405
rect 41052 16532 41104 16584
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 3792 16099 3844 16108
rect 3792 16065 3801 16099
rect 3801 16065 3835 16099
rect 3835 16065 3844 16099
rect 3792 16056 3844 16065
rect 4344 16192 4396 16244
rect 5264 16235 5316 16244
rect 5264 16201 5273 16235
rect 5273 16201 5307 16235
rect 5307 16201 5316 16235
rect 5264 16192 5316 16201
rect 5908 16192 5960 16244
rect 7380 16235 7432 16244
rect 7380 16201 7389 16235
rect 7389 16201 7423 16235
rect 7423 16201 7432 16235
rect 7380 16192 7432 16201
rect 7564 16192 7616 16244
rect 7656 16192 7708 16244
rect 9588 16192 9640 16244
rect 12348 16192 12400 16244
rect 15200 16192 15252 16244
rect 4160 16099 4212 16108
rect 4160 16065 4169 16099
rect 4169 16065 4203 16099
rect 4203 16065 4212 16099
rect 4160 16056 4212 16065
rect 4620 16056 4672 16108
rect 5724 16099 5776 16108
rect 4528 16031 4580 16040
rect 4528 15997 4537 16031
rect 4537 15997 4571 16031
rect 4571 15997 4580 16031
rect 4528 15988 4580 15997
rect 4896 15920 4948 15972
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 5632 15988 5684 16040
rect 6552 16056 6604 16108
rect 9036 16124 9088 16176
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 9220 16099 9272 16108
rect 9220 16065 9229 16099
rect 9229 16065 9263 16099
rect 9263 16065 9272 16099
rect 9220 16056 9272 16065
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 11060 16056 11112 16108
rect 11336 16056 11388 16108
rect 11428 16056 11480 16108
rect 14556 16124 14608 16176
rect 15476 16192 15528 16244
rect 15844 16192 15896 16244
rect 15936 16192 15988 16244
rect 16488 16192 16540 16244
rect 17224 16192 17276 16244
rect 17408 16192 17460 16244
rect 18144 16192 18196 16244
rect 20352 16192 20404 16244
rect 20904 16192 20956 16244
rect 21364 16124 21416 16176
rect 6460 15920 6512 15972
rect 6644 15920 6696 15972
rect 940 15852 992 15904
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 7472 15920 7524 15972
rect 11888 15988 11940 16040
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 12348 16099 12400 16108
rect 12348 16065 12357 16099
rect 12357 16065 12391 16099
rect 12391 16065 12400 16099
rect 12348 16056 12400 16065
rect 14004 16056 14056 16108
rect 15292 16056 15344 16108
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 15752 16056 15804 16108
rect 17776 16056 17828 16108
rect 18144 16097 18196 16108
rect 18144 16063 18153 16097
rect 18153 16063 18187 16097
rect 18187 16063 18196 16097
rect 18144 16056 18196 16063
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20812 16056 20864 16108
rect 20904 16099 20956 16108
rect 20904 16065 20913 16099
rect 20913 16065 20947 16099
rect 20947 16065 20956 16099
rect 20904 16056 20956 16065
rect 21088 16056 21140 16108
rect 22376 16056 22428 16108
rect 22744 16056 22796 16108
rect 17316 15988 17368 16040
rect 18420 15988 18472 16040
rect 20720 15988 20772 16040
rect 23664 16124 23716 16176
rect 25136 16192 25188 16244
rect 26240 16192 26292 16244
rect 26332 16192 26384 16244
rect 26792 16192 26844 16244
rect 23112 16099 23164 16108
rect 23112 16065 23121 16099
rect 23121 16065 23155 16099
rect 23155 16065 23164 16099
rect 23112 16056 23164 16065
rect 23388 16056 23440 16108
rect 21180 15988 21232 16040
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 8116 15852 8168 15904
rect 11796 15852 11848 15904
rect 17040 15895 17092 15904
rect 17040 15861 17049 15895
rect 17049 15861 17083 15895
rect 17083 15861 17092 15895
rect 17040 15852 17092 15861
rect 17224 15895 17276 15904
rect 17224 15861 17233 15895
rect 17233 15861 17267 15895
rect 17267 15861 17276 15895
rect 17224 15852 17276 15861
rect 18236 15852 18288 15904
rect 20168 15852 20220 15904
rect 20260 15895 20312 15904
rect 20260 15861 20269 15895
rect 20269 15861 20303 15895
rect 20303 15861 20312 15895
rect 20260 15852 20312 15861
rect 20904 15920 20956 15972
rect 21916 15920 21968 15972
rect 22928 16031 22980 16040
rect 22928 15997 22937 16031
rect 22937 15997 22971 16031
rect 22971 15997 22980 16031
rect 22928 15988 22980 15997
rect 24032 15988 24084 16040
rect 24308 15988 24360 16040
rect 24768 16056 24820 16108
rect 25688 16099 25740 16108
rect 25688 16065 25697 16099
rect 25697 16065 25731 16099
rect 25731 16065 25740 16099
rect 25688 16056 25740 16065
rect 29092 16124 29144 16176
rect 29184 16124 29236 16176
rect 26700 16056 26752 16108
rect 26792 16099 26844 16108
rect 26792 16065 26801 16099
rect 26801 16065 26835 16099
rect 26835 16065 26844 16099
rect 26792 16056 26844 16065
rect 22376 15852 22428 15904
rect 22560 15852 22612 15904
rect 22744 15852 22796 15904
rect 23664 15895 23716 15904
rect 23664 15861 23673 15895
rect 23673 15861 23707 15895
rect 23707 15861 23716 15895
rect 23664 15852 23716 15861
rect 24308 15852 24360 15904
rect 24768 15852 24820 15904
rect 26608 15920 26660 15972
rect 26700 15920 26752 15972
rect 27252 16099 27304 16108
rect 27252 16065 27261 16099
rect 27261 16065 27295 16099
rect 27295 16065 27304 16099
rect 27252 16056 27304 16065
rect 28540 16056 28592 16108
rect 29000 16099 29052 16108
rect 29000 16065 29009 16099
rect 29009 16065 29043 16099
rect 29043 16065 29052 16099
rect 29000 16056 29052 16065
rect 29828 16124 29880 16176
rect 30656 16124 30708 16176
rect 34520 16124 34572 16176
rect 29736 16056 29788 16108
rect 29920 16099 29972 16108
rect 29920 16065 29929 16099
rect 29929 16065 29963 16099
rect 29963 16065 29972 16099
rect 29920 16056 29972 16065
rect 32772 16056 32824 16108
rect 30932 15988 30984 16040
rect 32312 15988 32364 16040
rect 29644 15920 29696 15972
rect 33600 16099 33652 16108
rect 33600 16065 33609 16099
rect 33609 16065 33643 16099
rect 33643 16065 33652 16099
rect 33600 16056 33652 16065
rect 33876 16099 33928 16108
rect 33876 16065 33885 16099
rect 33885 16065 33919 16099
rect 33919 16065 33928 16099
rect 33876 16056 33928 16065
rect 33968 16099 34020 16108
rect 33968 16065 33977 16099
rect 33977 16065 34011 16099
rect 34011 16065 34020 16099
rect 33968 16056 34020 16065
rect 34244 16056 34296 16108
rect 34428 16056 34480 16108
rect 33416 15988 33468 16040
rect 28816 15852 28868 15904
rect 34244 15920 34296 15972
rect 34704 16056 34756 16108
rect 36820 16099 36872 16108
rect 36820 16065 36829 16099
rect 36829 16065 36863 16099
rect 36863 16065 36872 16099
rect 36820 16056 36872 16065
rect 37096 16056 37148 16108
rect 37832 16099 37884 16108
rect 37832 16065 37841 16099
rect 37841 16065 37875 16099
rect 37875 16065 37884 16099
rect 37832 16056 37884 16065
rect 38476 16056 38528 16108
rect 39212 16192 39264 16244
rect 39488 16192 39540 16244
rect 40500 16192 40552 16244
rect 40040 16124 40092 16176
rect 39028 15988 39080 16040
rect 36636 15963 36688 15972
rect 36636 15929 36645 15963
rect 36645 15929 36679 15963
rect 36679 15929 36688 15963
rect 36636 15920 36688 15929
rect 37372 15920 37424 15972
rect 33600 15852 33652 15904
rect 35348 15852 35400 15904
rect 39304 15852 39356 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1400 15648 1452 15700
rect 7104 15648 7156 15700
rect 7564 15648 7616 15700
rect 14004 15648 14056 15700
rect 14096 15648 14148 15700
rect 15660 15648 15712 15700
rect 17592 15691 17644 15700
rect 17592 15657 17601 15691
rect 17601 15657 17635 15691
rect 17635 15657 17644 15691
rect 17592 15648 17644 15657
rect 18144 15648 18196 15700
rect 18420 15648 18472 15700
rect 2688 15512 2740 15564
rect 3056 15444 3108 15496
rect 4804 15512 4856 15564
rect 10784 15623 10836 15632
rect 10784 15589 10793 15623
rect 10793 15589 10827 15623
rect 10827 15589 10836 15623
rect 10784 15580 10836 15589
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 10876 15512 10928 15564
rect 5080 15487 5132 15496
rect 5080 15453 5089 15487
rect 5089 15453 5123 15487
rect 5123 15453 5132 15487
rect 5080 15444 5132 15453
rect 5448 15444 5500 15496
rect 11980 15580 12032 15632
rect 11888 15512 11940 15564
rect 20904 15648 20956 15700
rect 21732 15648 21784 15700
rect 22008 15648 22060 15700
rect 22836 15648 22888 15700
rect 29644 15648 29696 15700
rect 32220 15648 32272 15700
rect 33416 15691 33468 15700
rect 33416 15657 33425 15691
rect 33425 15657 33459 15691
rect 33459 15657 33468 15691
rect 33416 15648 33468 15657
rect 17408 15512 17460 15564
rect 10232 15308 10284 15360
rect 11244 15444 11296 15496
rect 13360 15444 13412 15496
rect 13912 15444 13964 15496
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 11152 15308 11204 15360
rect 14648 15376 14700 15428
rect 17224 15376 17276 15428
rect 20168 15512 20220 15564
rect 22652 15580 22704 15632
rect 24216 15580 24268 15632
rect 34704 15648 34756 15700
rect 35348 15648 35400 15700
rect 18144 15487 18196 15496
rect 18144 15453 18153 15487
rect 18153 15453 18187 15487
rect 18187 15453 18196 15487
rect 18144 15444 18196 15453
rect 18420 15487 18472 15496
rect 18420 15453 18429 15487
rect 18429 15453 18463 15487
rect 18463 15453 18472 15487
rect 18420 15444 18472 15453
rect 16304 15308 16356 15360
rect 16856 15308 16908 15360
rect 18052 15376 18104 15428
rect 18144 15308 18196 15360
rect 18880 15444 18932 15496
rect 19432 15444 19484 15496
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 21732 15487 21784 15496
rect 21732 15453 21741 15487
rect 21741 15453 21775 15487
rect 21775 15453 21784 15487
rect 21732 15444 21784 15453
rect 21824 15419 21876 15428
rect 21824 15385 21833 15419
rect 21833 15385 21867 15419
rect 21867 15385 21876 15419
rect 21824 15376 21876 15385
rect 22284 15444 22336 15496
rect 22652 15444 22704 15496
rect 22928 15444 22980 15496
rect 23756 15512 23808 15564
rect 23940 15512 23992 15564
rect 27252 15512 27304 15564
rect 29184 15512 29236 15564
rect 30104 15555 30156 15564
rect 30104 15521 30113 15555
rect 30113 15521 30147 15555
rect 30147 15521 30156 15555
rect 30104 15512 30156 15521
rect 21364 15308 21416 15360
rect 23204 15376 23256 15428
rect 22100 15351 22152 15360
rect 22100 15317 22109 15351
rect 22109 15317 22143 15351
rect 22143 15317 22152 15351
rect 22100 15308 22152 15317
rect 22284 15308 22336 15360
rect 22836 15308 22888 15360
rect 23388 15419 23440 15428
rect 23388 15385 23397 15419
rect 23397 15385 23431 15419
rect 23431 15385 23440 15419
rect 23388 15376 23440 15385
rect 24124 15444 24176 15496
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 24584 15487 24636 15496
rect 24584 15453 24591 15487
rect 24591 15453 24636 15487
rect 24584 15444 24636 15453
rect 24860 15487 24912 15496
rect 24860 15453 24874 15487
rect 24874 15453 24908 15487
rect 24908 15453 24912 15487
rect 24860 15444 24912 15453
rect 29460 15444 29512 15496
rect 33692 15580 33744 15632
rect 34612 15580 34664 15632
rect 33968 15444 34020 15496
rect 34060 15444 34112 15496
rect 24768 15419 24820 15428
rect 24768 15385 24777 15419
rect 24777 15385 24811 15419
rect 24811 15385 24820 15419
rect 24768 15376 24820 15385
rect 25136 15376 25188 15428
rect 24216 15308 24268 15360
rect 24584 15308 24636 15360
rect 24952 15308 25004 15360
rect 31944 15376 31996 15428
rect 33784 15351 33836 15360
rect 33784 15317 33793 15351
rect 33793 15317 33827 15351
rect 33827 15317 33836 15351
rect 33784 15308 33836 15317
rect 35532 15308 35584 15360
rect 38660 15308 38712 15360
rect 39488 15308 39540 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 7472 15104 7524 15156
rect 6552 15036 6604 15088
rect 9220 15104 9272 15156
rect 10416 15104 10468 15156
rect 10784 15104 10836 15156
rect 10876 15104 10928 15156
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 5816 14968 5868 15020
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14968 7340 14977
rect 5908 14900 5960 14952
rect 8208 14900 8260 14952
rect 8852 15011 8904 15020
rect 8852 14977 8861 15011
rect 8861 14977 8895 15011
rect 8895 14977 8904 15011
rect 8852 14968 8904 14977
rect 9128 15011 9180 15020
rect 9128 14977 9163 15011
rect 9163 14977 9180 15011
rect 9128 14968 9180 14977
rect 9404 14968 9456 15020
rect 9956 15011 10008 15020
rect 9956 14977 9965 15011
rect 9965 14977 9999 15011
rect 9999 14977 10008 15011
rect 9956 14968 10008 14977
rect 10232 15011 10284 15020
rect 10232 14977 10241 15011
rect 10241 14977 10275 15011
rect 10275 14977 10284 15011
rect 10232 14968 10284 14977
rect 10876 15011 10928 15020
rect 10876 14977 10885 15011
rect 10885 14977 10919 15011
rect 10919 14977 10928 15011
rect 10876 14968 10928 14977
rect 11152 14968 11204 15020
rect 11336 15036 11388 15088
rect 11888 14968 11940 15020
rect 13912 15104 13964 15156
rect 16488 15104 16540 15156
rect 15660 15036 15712 15088
rect 9312 14943 9364 14952
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 6368 14832 6420 14884
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 14464 14900 14516 14952
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 16304 14968 16356 15020
rect 16764 14968 16816 15020
rect 17960 15104 18012 15156
rect 18052 15104 18104 15156
rect 18788 15104 18840 15156
rect 19800 15104 19852 15156
rect 23388 15104 23440 15156
rect 23480 15104 23532 15156
rect 15752 14900 15804 14952
rect 17408 14968 17460 15020
rect 23664 15036 23716 15088
rect 24400 15147 24452 15156
rect 24400 15113 24409 15147
rect 24409 15113 24443 15147
rect 24443 15113 24452 15147
rect 24400 15104 24452 15113
rect 26240 15104 26292 15156
rect 27712 15104 27764 15156
rect 28356 15104 28408 15156
rect 30012 15104 30064 15156
rect 30104 15104 30156 15156
rect 19340 14968 19392 15020
rect 17960 14943 18012 14952
rect 17960 14909 17969 14943
rect 17969 14909 18003 14943
rect 18003 14909 18012 14943
rect 17960 14900 18012 14909
rect 18236 14900 18288 14952
rect 19524 14968 19576 15020
rect 20168 15011 20220 15020
rect 20168 14977 20177 15011
rect 20177 14977 20211 15011
rect 20211 14977 20220 15011
rect 20168 14968 20220 14977
rect 20260 14968 20312 15020
rect 20720 14968 20772 15020
rect 20076 14900 20128 14952
rect 21180 14900 21232 14952
rect 21548 14900 21600 14952
rect 22928 14968 22980 15020
rect 23112 14968 23164 15020
rect 23756 14968 23808 15020
rect 15292 14832 15344 14884
rect 16488 14832 16540 14884
rect 18420 14832 18472 14884
rect 19432 14832 19484 14884
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 24860 15036 24912 15088
rect 26516 15036 26568 15088
rect 27252 15079 27304 15088
rect 27252 15045 27261 15079
rect 27261 15045 27295 15079
rect 27295 15045 27304 15079
rect 27252 15036 27304 15045
rect 25964 14968 26016 15020
rect 26056 14900 26108 14952
rect 26240 14900 26292 14952
rect 26700 14900 26752 14952
rect 27528 14968 27580 15020
rect 27712 14968 27764 15020
rect 27804 15011 27856 15020
rect 27804 14977 27813 15011
rect 27813 14977 27847 15011
rect 27847 14977 27856 15011
rect 27804 14968 27856 14977
rect 27896 15011 27948 15020
rect 27896 14977 27905 15011
rect 27905 14977 27939 15011
rect 27939 14977 27948 15011
rect 27896 14968 27948 14977
rect 28080 14968 28132 15020
rect 28264 14968 28316 15020
rect 7012 14764 7064 14816
rect 8024 14764 8076 14816
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 9864 14764 9916 14816
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 10692 14807 10744 14816
rect 10692 14773 10701 14807
rect 10701 14773 10735 14807
rect 10735 14773 10744 14807
rect 10692 14764 10744 14773
rect 10968 14764 11020 14816
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 16764 14764 16816 14816
rect 17040 14764 17092 14816
rect 27620 14832 27672 14884
rect 39764 15104 39816 15156
rect 31944 15036 31996 15088
rect 31392 15011 31444 15020
rect 31392 14977 31401 15011
rect 31401 14977 31435 15011
rect 31435 14977 31444 15011
rect 31392 14968 31444 14977
rect 31300 14900 31352 14952
rect 31576 15011 31628 15020
rect 31576 14977 31585 15011
rect 31585 14977 31619 15011
rect 31619 14977 31628 15011
rect 31576 14968 31628 14977
rect 33968 14968 34020 15020
rect 34704 14968 34756 15020
rect 35624 14968 35676 15020
rect 39304 14968 39356 15020
rect 31852 14943 31904 14952
rect 31852 14909 31861 14943
rect 31861 14909 31895 14943
rect 31895 14909 31904 14943
rect 31852 14900 31904 14909
rect 25044 14764 25096 14816
rect 27528 14807 27580 14816
rect 27528 14773 27537 14807
rect 27537 14773 27571 14807
rect 27571 14773 27580 14807
rect 27528 14764 27580 14773
rect 28172 14807 28224 14816
rect 28172 14773 28181 14807
rect 28181 14773 28215 14807
rect 28215 14773 28224 14807
rect 28172 14764 28224 14773
rect 29552 14807 29604 14816
rect 29552 14773 29561 14807
rect 29561 14773 29595 14807
rect 29595 14773 29604 14807
rect 29552 14764 29604 14773
rect 31116 14807 31168 14816
rect 31116 14773 31125 14807
rect 31125 14773 31159 14807
rect 31159 14773 31168 14807
rect 31116 14764 31168 14773
rect 32220 14832 32272 14884
rect 31300 14764 31352 14816
rect 31576 14764 31628 14816
rect 32036 14764 32088 14816
rect 35808 14832 35860 14884
rect 35440 14807 35492 14816
rect 35440 14773 35449 14807
rect 35449 14773 35483 14807
rect 35483 14773 35492 14807
rect 35440 14764 35492 14773
rect 38660 14764 38712 14816
rect 38844 14807 38896 14816
rect 38844 14773 38853 14807
rect 38853 14773 38887 14807
rect 38887 14773 38896 14807
rect 38844 14764 38896 14773
rect 39396 14832 39448 14884
rect 39580 14764 39632 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3424 14603 3476 14612
rect 3424 14569 3433 14603
rect 3433 14569 3467 14603
rect 3467 14569 3476 14603
rect 3424 14560 3476 14569
rect 5724 14560 5776 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 5908 14560 5960 14612
rect 4068 14356 4120 14408
rect 5080 14424 5132 14476
rect 5816 14424 5868 14476
rect 6184 14467 6236 14476
rect 6184 14433 6193 14467
rect 6193 14433 6227 14467
rect 6227 14433 6236 14467
rect 8668 14560 8720 14612
rect 9128 14560 9180 14612
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 10692 14560 10744 14612
rect 6184 14424 6236 14433
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 3608 14263 3660 14272
rect 3608 14229 3617 14263
rect 3617 14229 3651 14263
rect 3651 14229 3660 14263
rect 3608 14220 3660 14229
rect 4620 14220 4672 14272
rect 4896 14220 4948 14272
rect 5724 14356 5776 14408
rect 6276 14399 6328 14408
rect 6276 14365 6285 14399
rect 6285 14365 6319 14399
rect 6319 14365 6328 14399
rect 6276 14356 6328 14365
rect 7288 14492 7340 14544
rect 8024 14492 8076 14544
rect 8944 14492 8996 14544
rect 10876 14560 10928 14612
rect 12440 14560 12492 14612
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 8024 14399 8076 14408
rect 8024 14365 8033 14399
rect 8033 14365 8067 14399
rect 8067 14365 8076 14399
rect 8024 14356 8076 14365
rect 10416 14424 10468 14476
rect 6644 14288 6696 14340
rect 7012 14331 7064 14340
rect 7012 14297 7047 14331
rect 7047 14297 7064 14331
rect 7012 14288 7064 14297
rect 6736 14220 6788 14272
rect 8484 14288 8536 14340
rect 9220 14356 9272 14408
rect 8208 14220 8260 14272
rect 9036 14288 9088 14340
rect 10784 14424 10836 14476
rect 13912 14424 13964 14476
rect 11336 14399 11388 14408
rect 11336 14365 11346 14399
rect 11346 14365 11380 14399
rect 11380 14365 11388 14399
rect 11336 14356 11388 14365
rect 11888 14356 11940 14408
rect 11428 14288 11480 14340
rect 14924 14399 14976 14408
rect 14924 14365 14934 14399
rect 14934 14365 14968 14399
rect 14968 14365 14976 14399
rect 15200 14560 15252 14612
rect 17500 14560 17552 14612
rect 17776 14492 17828 14544
rect 14924 14356 14976 14365
rect 16028 14424 16080 14476
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 16212 14356 16264 14408
rect 9680 14220 9732 14272
rect 10600 14220 10652 14272
rect 15568 14331 15620 14340
rect 15568 14297 15577 14331
rect 15577 14297 15611 14331
rect 15611 14297 15620 14331
rect 15568 14288 15620 14297
rect 17040 14399 17092 14408
rect 17040 14365 17055 14399
rect 17055 14365 17089 14399
rect 17089 14365 17092 14399
rect 17040 14356 17092 14365
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 18144 14424 18196 14476
rect 18696 14492 18748 14544
rect 21916 14560 21968 14612
rect 24492 14560 24544 14612
rect 24584 14560 24636 14612
rect 26884 14560 26936 14612
rect 27528 14560 27580 14612
rect 20444 14492 20496 14544
rect 22744 14492 22796 14544
rect 18788 14356 18840 14408
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 14924 14220 14976 14272
rect 15108 14220 15160 14272
rect 15936 14220 15988 14272
rect 16120 14220 16172 14272
rect 16764 14220 16816 14272
rect 20996 14424 21048 14476
rect 19800 14356 19852 14408
rect 20444 14356 20496 14408
rect 20812 14356 20864 14408
rect 21548 14424 21600 14476
rect 22928 14467 22980 14476
rect 22928 14433 22937 14467
rect 22937 14433 22971 14467
rect 22971 14433 22980 14467
rect 22928 14424 22980 14433
rect 23020 14424 23072 14476
rect 24860 14424 24912 14476
rect 26148 14424 26200 14476
rect 26608 14424 26660 14476
rect 22284 14356 22336 14408
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 26332 14399 26384 14408
rect 26332 14365 26341 14399
rect 26341 14365 26375 14399
rect 26375 14365 26384 14399
rect 26332 14356 26384 14365
rect 26516 14399 26568 14408
rect 26516 14365 26525 14399
rect 26525 14365 26559 14399
rect 26559 14365 26568 14399
rect 26516 14356 26568 14365
rect 26700 14399 26752 14408
rect 26700 14365 26709 14399
rect 26709 14365 26743 14399
rect 26743 14365 26752 14399
rect 26700 14356 26752 14365
rect 27068 14356 27120 14408
rect 28172 14560 28224 14612
rect 29552 14560 29604 14612
rect 31300 14560 31352 14612
rect 31392 14560 31444 14612
rect 32220 14603 32272 14612
rect 32220 14569 32229 14603
rect 32229 14569 32263 14603
rect 32263 14569 32272 14603
rect 32220 14560 32272 14569
rect 35256 14560 35308 14612
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 17408 14220 17460 14229
rect 18788 14220 18840 14272
rect 21180 14220 21232 14272
rect 22100 14220 22152 14272
rect 22744 14220 22796 14272
rect 23664 14220 23716 14272
rect 25320 14288 25372 14340
rect 26608 14331 26660 14340
rect 26608 14297 26617 14331
rect 26617 14297 26651 14331
rect 26651 14297 26660 14331
rect 26608 14288 26660 14297
rect 27804 14399 27856 14408
rect 27804 14365 27813 14399
rect 27813 14365 27847 14399
rect 27847 14365 27856 14399
rect 27804 14356 27856 14365
rect 29276 14424 29328 14476
rect 31852 14492 31904 14544
rect 32128 14492 32180 14544
rect 33968 14492 34020 14544
rect 37188 14560 37240 14612
rect 28356 14356 28408 14408
rect 30840 14356 30892 14408
rect 33784 14424 33836 14476
rect 35348 14424 35400 14476
rect 35440 14424 35492 14476
rect 35808 14424 35860 14476
rect 31300 14356 31352 14408
rect 31484 14356 31536 14408
rect 26884 14263 26936 14272
rect 26884 14229 26893 14263
rect 26893 14229 26927 14263
rect 26927 14229 26936 14263
rect 26884 14220 26936 14229
rect 26976 14263 27028 14272
rect 26976 14229 26985 14263
rect 26985 14229 27019 14263
rect 27019 14229 27028 14263
rect 26976 14220 27028 14229
rect 27620 14263 27672 14272
rect 27620 14229 27629 14263
rect 27629 14229 27663 14263
rect 27663 14229 27672 14263
rect 27620 14220 27672 14229
rect 27712 14220 27764 14272
rect 31116 14288 31168 14340
rect 28172 14220 28224 14272
rect 31484 14220 31536 14272
rect 35532 14399 35584 14408
rect 35532 14365 35541 14399
rect 35541 14365 35575 14399
rect 35575 14365 35584 14399
rect 35532 14356 35584 14365
rect 36084 14356 36136 14408
rect 36176 14356 36228 14408
rect 33324 14220 33376 14272
rect 34520 14220 34572 14272
rect 35256 14288 35308 14340
rect 35900 14331 35952 14340
rect 35900 14297 35909 14331
rect 35909 14297 35943 14331
rect 35943 14297 35952 14331
rect 35900 14288 35952 14297
rect 38752 14492 38804 14544
rect 39488 14535 39540 14544
rect 39488 14501 39497 14535
rect 39497 14501 39531 14535
rect 39531 14501 39540 14535
rect 39488 14492 39540 14501
rect 39764 14424 39816 14476
rect 38660 14399 38712 14408
rect 38660 14365 38669 14399
rect 38669 14365 38703 14399
rect 38703 14365 38712 14399
rect 38660 14356 38712 14365
rect 38752 14399 38804 14408
rect 38752 14365 38761 14399
rect 38761 14365 38795 14399
rect 38795 14365 38804 14399
rect 38752 14356 38804 14365
rect 38292 14331 38344 14340
rect 38292 14297 38301 14331
rect 38301 14297 38335 14331
rect 38335 14297 38344 14331
rect 38292 14288 38344 14297
rect 39304 14399 39356 14408
rect 39304 14365 39313 14399
rect 39313 14365 39347 14399
rect 39347 14365 39356 14399
rect 39304 14356 39356 14365
rect 39396 14399 39448 14408
rect 39396 14365 39405 14399
rect 39405 14365 39439 14399
rect 39439 14365 39448 14399
rect 39396 14356 39448 14365
rect 39580 14399 39632 14408
rect 39580 14365 39589 14399
rect 39589 14365 39623 14399
rect 39623 14365 39632 14399
rect 39580 14356 39632 14365
rect 40500 14331 40552 14340
rect 40500 14297 40509 14331
rect 40509 14297 40543 14331
rect 40543 14297 40552 14331
rect 40500 14288 40552 14297
rect 39304 14220 39356 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 3608 14016 3660 14068
rect 3056 13948 3108 14000
rect 4528 14016 4580 14068
rect 8484 14016 8536 14068
rect 9220 14016 9272 14068
rect 9680 14016 9732 14068
rect 12072 14016 12124 14068
rect 12440 14016 12492 14068
rect 15016 14016 15068 14068
rect 15200 14016 15252 14068
rect 16856 14016 16908 14068
rect 6920 13880 6972 13932
rect 8116 13880 8168 13932
rect 11336 13880 11388 13932
rect 11888 13923 11940 13932
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 14372 13948 14424 14000
rect 15200 13880 15252 13932
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 15844 13948 15896 14000
rect 16948 13991 17000 14000
rect 16948 13957 16957 13991
rect 16957 13957 16991 13991
rect 16991 13957 17000 13991
rect 16948 13948 17000 13957
rect 18788 14059 18840 14068
rect 18788 14025 18797 14059
rect 18797 14025 18831 14059
rect 18831 14025 18840 14059
rect 18788 14016 18840 14025
rect 19984 14016 20036 14068
rect 2688 13855 2740 13864
rect 2688 13821 2697 13855
rect 2697 13821 2731 13855
rect 2731 13821 2740 13855
rect 2688 13812 2740 13821
rect 3700 13812 3752 13864
rect 7932 13812 7984 13864
rect 8668 13812 8720 13864
rect 11244 13812 11296 13864
rect 12348 13812 12400 13864
rect 15108 13812 15160 13864
rect 15384 13812 15436 13864
rect 15752 13812 15804 13864
rect 15936 13812 15988 13864
rect 16120 13812 16172 13864
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 17132 13880 17184 13932
rect 17408 13880 17460 13932
rect 17776 13923 17828 13932
rect 17776 13889 17785 13923
rect 17785 13889 17819 13923
rect 17819 13889 17828 13923
rect 17776 13880 17828 13889
rect 18052 13880 18104 13932
rect 18144 13923 18196 13930
rect 18144 13889 18153 13923
rect 18153 13889 18187 13923
rect 18187 13889 18196 13923
rect 18144 13878 18196 13889
rect 19708 13948 19760 14000
rect 17776 13744 17828 13796
rect 18236 13744 18288 13796
rect 18604 13923 18656 13932
rect 18604 13889 18618 13923
rect 18618 13889 18652 13923
rect 18652 13889 18656 13923
rect 18604 13880 18656 13889
rect 20076 13880 20128 13932
rect 20444 13880 20496 13932
rect 20904 13923 20956 13932
rect 20904 13889 20913 13923
rect 20913 13889 20947 13923
rect 20947 13889 20956 13923
rect 20904 13880 20956 13889
rect 21456 14016 21508 14068
rect 22284 14016 22336 14068
rect 23480 14016 23532 14068
rect 23848 14016 23900 14068
rect 21180 13948 21232 14000
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 21456 13923 21508 13932
rect 21456 13889 21465 13923
rect 21465 13889 21499 13923
rect 21499 13889 21508 13923
rect 21456 13880 21508 13889
rect 22376 13880 22428 13932
rect 22744 13923 22796 13932
rect 22744 13889 22753 13923
rect 22753 13889 22787 13923
rect 22787 13889 22796 13923
rect 22744 13880 22796 13889
rect 22836 13923 22888 13932
rect 22836 13889 22846 13923
rect 22846 13889 22880 13923
rect 22880 13889 22888 13923
rect 22836 13880 22888 13889
rect 23020 13923 23072 13932
rect 23020 13889 23029 13923
rect 23029 13889 23063 13923
rect 23063 13889 23072 13923
rect 23020 13880 23072 13889
rect 23480 13923 23532 13932
rect 23480 13889 23489 13923
rect 23489 13889 23523 13923
rect 23523 13889 23532 13923
rect 23480 13880 23532 13889
rect 23664 13923 23716 13932
rect 23664 13889 23673 13923
rect 23673 13889 23707 13923
rect 23707 13889 23716 13923
rect 23664 13880 23716 13889
rect 19524 13812 19576 13864
rect 18420 13744 18472 13796
rect 20260 13787 20312 13796
rect 20260 13753 20269 13787
rect 20269 13753 20303 13787
rect 20303 13753 20312 13787
rect 20260 13744 20312 13753
rect 21640 13855 21692 13864
rect 21640 13821 21649 13855
rect 21649 13821 21683 13855
rect 21683 13821 21692 13855
rect 21640 13812 21692 13821
rect 23756 13812 23808 13864
rect 24032 13812 24084 13864
rect 14556 13676 14608 13728
rect 15936 13676 15988 13728
rect 16028 13676 16080 13728
rect 17960 13676 18012 13728
rect 18144 13676 18196 13728
rect 21732 13676 21784 13728
rect 22560 13787 22612 13796
rect 22560 13753 22569 13787
rect 22569 13753 22603 13787
rect 22603 13753 22612 13787
rect 22560 13744 22612 13753
rect 24400 13880 24452 13932
rect 24584 13880 24636 13932
rect 25964 14016 26016 14068
rect 27252 14016 27304 14068
rect 27344 14016 27396 14068
rect 24676 13855 24728 13898
rect 24676 13846 24685 13855
rect 24685 13846 24719 13855
rect 24719 13846 24728 13855
rect 23388 13719 23440 13728
rect 23388 13685 23397 13719
rect 23397 13685 23431 13719
rect 23431 13685 23440 13719
rect 23388 13676 23440 13685
rect 23756 13676 23808 13728
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 25136 13923 25188 13932
rect 25136 13889 25145 13923
rect 25145 13889 25179 13923
rect 25179 13889 25188 13923
rect 25136 13880 25188 13889
rect 25320 13923 25372 13932
rect 25320 13889 25329 13923
rect 25329 13889 25363 13923
rect 25363 13889 25372 13923
rect 25320 13880 25372 13889
rect 25044 13744 25096 13796
rect 26884 13880 26936 13932
rect 27712 13880 27764 13932
rect 25780 13744 25832 13796
rect 26792 13744 26844 13796
rect 27344 13787 27396 13796
rect 27344 13753 27353 13787
rect 27353 13753 27387 13787
rect 27387 13753 27396 13787
rect 27344 13744 27396 13753
rect 28080 13812 28132 13864
rect 28264 13923 28316 13932
rect 28264 13889 28273 13923
rect 28273 13889 28307 13923
rect 28307 13889 28316 13923
rect 28264 13880 28316 13889
rect 31024 14016 31076 14068
rect 32956 14016 33008 14068
rect 33232 14016 33284 14068
rect 33968 14016 34020 14068
rect 31392 13948 31444 14000
rect 30196 13880 30248 13932
rect 31024 13923 31076 13932
rect 31024 13889 31033 13923
rect 31033 13889 31067 13923
rect 31067 13889 31076 13923
rect 31024 13880 31076 13889
rect 31576 13923 31628 13932
rect 31576 13889 31585 13923
rect 31585 13889 31619 13923
rect 31619 13889 31628 13923
rect 31576 13880 31628 13889
rect 28448 13812 28500 13864
rect 28356 13744 28408 13796
rect 32036 13880 32088 13932
rect 32128 13923 32180 13932
rect 32128 13889 32137 13923
rect 32137 13889 32171 13923
rect 32171 13889 32180 13923
rect 32128 13880 32180 13889
rect 32220 13880 32272 13932
rect 33140 13880 33192 13932
rect 33324 13923 33376 13932
rect 33324 13889 33330 13923
rect 33330 13889 33364 13923
rect 33364 13889 33376 13923
rect 33324 13880 33376 13889
rect 33600 13880 33652 13932
rect 34244 13948 34296 14000
rect 34704 14059 34756 14068
rect 34704 14025 34713 14059
rect 34713 14025 34747 14059
rect 34747 14025 34756 14059
rect 34704 14016 34756 14025
rect 34152 13923 34204 13932
rect 34152 13889 34161 13923
rect 34161 13889 34195 13923
rect 34195 13889 34204 13923
rect 34152 13880 34204 13889
rect 34336 13923 34388 13932
rect 34336 13889 34345 13923
rect 34345 13889 34379 13923
rect 34379 13889 34388 13923
rect 34336 13880 34388 13889
rect 34612 13923 34664 13932
rect 34612 13889 34621 13923
rect 34621 13889 34655 13923
rect 34655 13889 34664 13923
rect 34612 13880 34664 13889
rect 34704 13880 34756 13932
rect 34888 13880 34940 13932
rect 35348 13948 35400 14000
rect 35900 14016 35952 14068
rect 35532 13923 35584 13932
rect 35532 13889 35541 13923
rect 35541 13889 35575 13923
rect 35575 13889 35584 13923
rect 35532 13880 35584 13889
rect 25136 13676 25188 13728
rect 25320 13676 25372 13728
rect 26240 13676 26292 13728
rect 27252 13676 27304 13728
rect 31852 13676 31904 13728
rect 34796 13744 34848 13796
rect 33692 13719 33744 13728
rect 33692 13685 33701 13719
rect 33701 13685 33735 13719
rect 33735 13685 33744 13719
rect 33692 13676 33744 13685
rect 33968 13676 34020 13728
rect 35900 13812 35952 13864
rect 38660 13880 38712 13932
rect 36268 13744 36320 13796
rect 35992 13676 36044 13728
rect 38292 13812 38344 13864
rect 38476 13855 38528 13864
rect 38476 13821 38485 13855
rect 38485 13821 38519 13855
rect 38519 13821 38528 13855
rect 38476 13812 38528 13821
rect 38752 13812 38804 13864
rect 39396 14016 39448 14068
rect 39304 13991 39356 14000
rect 39304 13957 39313 13991
rect 39313 13957 39347 13991
rect 39347 13957 39356 13991
rect 39304 13948 39356 13957
rect 40040 13948 40092 14000
rect 39028 13855 39080 13864
rect 39028 13821 39037 13855
rect 39037 13821 39071 13855
rect 39071 13821 39080 13855
rect 39028 13812 39080 13821
rect 38384 13676 38436 13728
rect 38660 13676 38712 13728
rect 39764 13676 39816 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 6276 13472 6328 13524
rect 6736 13472 6788 13524
rect 8484 13472 8536 13524
rect 10968 13472 11020 13524
rect 11888 13472 11940 13524
rect 12808 13472 12860 13524
rect 16488 13472 16540 13524
rect 19340 13472 19392 13524
rect 5724 13336 5776 13388
rect 7380 13404 7432 13456
rect 6828 13336 6880 13388
rect 6736 13200 6788 13252
rect 8024 13268 8076 13320
rect 8392 13200 8444 13252
rect 16028 13404 16080 13456
rect 12716 13379 12768 13388
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 12992 13268 13044 13320
rect 13452 13336 13504 13388
rect 13544 13379 13596 13388
rect 13544 13345 13553 13379
rect 13553 13345 13587 13379
rect 13587 13345 13596 13379
rect 13544 13336 13596 13345
rect 13360 13200 13412 13252
rect 6920 13132 6972 13184
rect 8024 13175 8076 13184
rect 8024 13141 8033 13175
rect 8033 13141 8067 13175
rect 8067 13141 8076 13175
rect 8024 13132 8076 13141
rect 11704 13132 11756 13184
rect 12900 13175 12952 13184
rect 12900 13141 12909 13175
rect 12909 13141 12943 13175
rect 12943 13141 12952 13175
rect 12900 13132 12952 13141
rect 15844 13200 15896 13252
rect 20996 13404 21048 13456
rect 21824 13404 21876 13456
rect 17132 13336 17184 13388
rect 17224 13379 17276 13388
rect 17224 13345 17233 13379
rect 17233 13345 17267 13379
rect 17267 13345 17276 13379
rect 17224 13336 17276 13345
rect 17408 13379 17460 13388
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 18052 13336 18104 13388
rect 20168 13336 20220 13388
rect 23572 13472 23624 13524
rect 24584 13472 24636 13524
rect 22284 13404 22336 13456
rect 16304 13311 16356 13320
rect 16304 13277 16314 13311
rect 16314 13277 16348 13311
rect 16348 13277 16356 13311
rect 16304 13268 16356 13277
rect 18236 13268 18288 13320
rect 22192 13336 22244 13388
rect 16580 13243 16632 13252
rect 16580 13209 16589 13243
rect 16589 13209 16623 13243
rect 16623 13209 16632 13243
rect 16580 13200 16632 13209
rect 16948 13243 17000 13252
rect 16948 13209 16957 13243
rect 16957 13209 16991 13243
rect 16991 13209 17000 13243
rect 16948 13200 17000 13209
rect 21824 13268 21876 13320
rect 22284 13311 22336 13320
rect 22284 13277 22293 13311
rect 22293 13277 22327 13311
rect 22327 13277 22336 13311
rect 22284 13268 22336 13277
rect 16120 13132 16172 13184
rect 16764 13132 16816 13184
rect 21456 13200 21508 13252
rect 23388 13268 23440 13320
rect 22744 13200 22796 13252
rect 19064 13132 19116 13184
rect 19248 13132 19300 13184
rect 22100 13175 22152 13184
rect 22100 13141 22109 13175
rect 22109 13141 22143 13175
rect 22143 13141 22152 13175
rect 22100 13132 22152 13141
rect 22652 13132 22704 13184
rect 23480 13200 23532 13252
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 30104 13472 30156 13524
rect 24768 13336 24820 13388
rect 25136 13336 25188 13388
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 25780 13404 25832 13456
rect 25964 13404 26016 13456
rect 27712 13404 27764 13456
rect 25964 13311 26016 13320
rect 25964 13277 25973 13311
rect 25973 13277 26007 13311
rect 26007 13277 26016 13311
rect 25964 13268 26016 13277
rect 26424 13311 26476 13320
rect 26424 13277 26438 13311
rect 26438 13277 26472 13311
rect 26472 13277 26476 13311
rect 26424 13268 26476 13277
rect 26700 13268 26752 13320
rect 27068 13268 27120 13320
rect 31024 13404 31076 13456
rect 22928 13175 22980 13184
rect 22928 13141 22937 13175
rect 22937 13141 22971 13175
rect 22971 13141 22980 13175
rect 22928 13132 22980 13141
rect 24400 13175 24452 13184
rect 24400 13141 24409 13175
rect 24409 13141 24443 13175
rect 24443 13141 24452 13175
rect 24400 13132 24452 13141
rect 25044 13132 25096 13184
rect 25504 13132 25556 13184
rect 26332 13243 26384 13252
rect 26332 13209 26341 13243
rect 26341 13209 26375 13243
rect 26375 13209 26384 13243
rect 26332 13200 26384 13209
rect 26516 13200 26568 13252
rect 27344 13200 27396 13252
rect 26700 13175 26752 13184
rect 26700 13141 26709 13175
rect 26709 13141 26743 13175
rect 26743 13141 26752 13175
rect 26700 13132 26752 13141
rect 26792 13132 26844 13184
rect 32036 13404 32088 13456
rect 33140 13472 33192 13524
rect 35440 13472 35492 13524
rect 35624 13472 35676 13524
rect 35900 13472 35952 13524
rect 34704 13404 34756 13456
rect 36268 13404 36320 13456
rect 28356 13268 28408 13320
rect 31484 13311 31536 13320
rect 31484 13277 31493 13311
rect 31493 13277 31527 13311
rect 31527 13277 31536 13311
rect 31484 13268 31536 13277
rect 31576 13311 31628 13320
rect 31576 13277 31585 13311
rect 31585 13277 31619 13311
rect 31619 13277 31628 13311
rect 31576 13268 31628 13277
rect 31944 13311 31996 13320
rect 31944 13277 31953 13311
rect 31953 13277 31987 13311
rect 31987 13277 31996 13311
rect 31944 13268 31996 13277
rect 32956 13268 33008 13320
rect 34152 13268 34204 13320
rect 34428 13311 34480 13320
rect 34428 13277 34437 13311
rect 34437 13277 34471 13311
rect 34471 13277 34480 13311
rect 34428 13268 34480 13277
rect 34520 13311 34572 13320
rect 34520 13277 34529 13311
rect 34529 13277 34563 13311
rect 34563 13277 34572 13311
rect 35992 13336 36044 13388
rect 34520 13268 34572 13277
rect 35532 13268 35584 13320
rect 29000 13200 29052 13252
rect 35072 13200 35124 13252
rect 31300 13132 31352 13184
rect 32220 13175 32272 13184
rect 32220 13141 32229 13175
rect 32229 13141 32263 13175
rect 32263 13141 32272 13175
rect 32220 13132 32272 13141
rect 34704 13132 34756 13184
rect 35716 13200 35768 13252
rect 35900 13268 35952 13320
rect 38936 13472 38988 13524
rect 38568 13336 38620 13388
rect 36268 13200 36320 13252
rect 38384 13268 38436 13320
rect 38660 13311 38712 13320
rect 38660 13277 38669 13311
rect 38669 13277 38703 13311
rect 38703 13277 38712 13311
rect 38660 13268 38712 13277
rect 39120 13268 39172 13320
rect 39396 13268 39448 13320
rect 39764 13268 39816 13320
rect 36636 13200 36688 13252
rect 38752 13200 38804 13252
rect 39764 13132 39816 13184
rect 39856 13132 39908 13184
rect 41052 13175 41104 13184
rect 41052 13141 41061 13175
rect 41061 13141 41095 13175
rect 41095 13141 41104 13175
rect 41052 13132 41104 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 6092 12903 6144 12912
rect 6092 12869 6101 12903
rect 6101 12869 6135 12903
rect 6135 12869 6144 12903
rect 6092 12860 6144 12869
rect 6276 12860 6328 12912
rect 8024 12928 8076 12980
rect 8576 12928 8628 12980
rect 8760 12928 8812 12980
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7012 12792 7064 12844
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 7932 12792 7984 12844
rect 10784 12928 10836 12980
rect 11428 12928 11480 12980
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 5448 12656 5500 12708
rect 6828 12656 6880 12708
rect 8576 12835 8628 12844
rect 8576 12801 8585 12835
rect 8585 12801 8619 12835
rect 8619 12801 8628 12835
rect 8576 12792 8628 12801
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 9128 12792 9180 12844
rect 9588 12792 9640 12844
rect 12900 12928 12952 12980
rect 15292 12860 15344 12912
rect 16580 12928 16632 12980
rect 17132 12928 17184 12980
rect 17684 12928 17736 12980
rect 19524 12928 19576 12980
rect 20720 12928 20772 12980
rect 24952 12928 25004 12980
rect 25596 12928 25648 12980
rect 31392 12928 31444 12980
rect 31852 12928 31904 12980
rect 18604 12860 18656 12912
rect 9772 12724 9824 12776
rect 10784 12792 10836 12844
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12716 12792 12768 12844
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 14096 12792 14148 12844
rect 16948 12792 17000 12844
rect 17868 12792 17920 12844
rect 18236 12792 18288 12844
rect 18788 12792 18840 12844
rect 11060 12724 11112 12776
rect 12348 12724 12400 12776
rect 12624 12724 12676 12776
rect 17960 12724 18012 12776
rect 19340 12860 19392 12912
rect 19248 12792 19300 12844
rect 19984 12835 20036 12844
rect 19984 12801 19993 12835
rect 19993 12801 20027 12835
rect 20027 12801 20036 12835
rect 19984 12792 20036 12801
rect 20168 12835 20220 12844
rect 20168 12801 20177 12835
rect 20177 12801 20211 12835
rect 20211 12801 20220 12835
rect 20168 12792 20220 12801
rect 20260 12792 20312 12844
rect 23940 12860 23992 12912
rect 24216 12903 24268 12912
rect 24216 12869 24225 12903
rect 24225 12869 24259 12903
rect 24259 12869 24268 12903
rect 24216 12860 24268 12869
rect 25320 12860 25372 12912
rect 25688 12860 25740 12912
rect 28816 12903 28868 12912
rect 28816 12869 28825 12903
rect 28825 12869 28859 12903
rect 28859 12869 28868 12903
rect 28816 12860 28868 12869
rect 29000 12860 29052 12912
rect 29276 12860 29328 12912
rect 30748 12860 30800 12912
rect 21088 12792 21140 12844
rect 23480 12792 23532 12844
rect 23664 12792 23716 12844
rect 24584 12792 24636 12844
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 6368 12631 6420 12640
rect 6368 12597 6377 12631
rect 6377 12597 6411 12631
rect 6411 12597 6420 12631
rect 6368 12588 6420 12597
rect 8392 12631 8444 12640
rect 8392 12597 8401 12631
rect 8401 12597 8435 12631
rect 8435 12597 8444 12631
rect 8392 12588 8444 12597
rect 9036 12656 9088 12708
rect 10048 12656 10100 12708
rect 13544 12656 13596 12708
rect 16120 12656 16172 12708
rect 15016 12631 15068 12640
rect 15016 12597 15046 12631
rect 15046 12597 15068 12631
rect 15016 12588 15068 12597
rect 15384 12588 15436 12640
rect 15660 12588 15712 12640
rect 18880 12588 18932 12640
rect 19064 12656 19116 12708
rect 19156 12656 19208 12708
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 25044 12724 25096 12776
rect 28632 12724 28684 12776
rect 31300 12835 31352 12844
rect 31300 12801 31309 12835
rect 31309 12801 31343 12835
rect 31343 12801 31352 12835
rect 31300 12792 31352 12801
rect 32220 12860 32272 12912
rect 31760 12835 31812 12844
rect 31760 12801 31769 12835
rect 31769 12801 31803 12835
rect 31803 12801 31812 12835
rect 31760 12792 31812 12801
rect 36176 12928 36228 12980
rect 33232 12860 33284 12912
rect 33784 12860 33836 12912
rect 35072 12860 35124 12912
rect 36636 12860 36688 12912
rect 37464 12835 37516 12844
rect 37464 12801 37473 12835
rect 37473 12801 37507 12835
rect 37507 12801 37516 12835
rect 37464 12792 37516 12801
rect 31392 12724 31444 12776
rect 31668 12767 31720 12776
rect 31668 12733 31677 12767
rect 31677 12733 31711 12767
rect 31711 12733 31720 12767
rect 31668 12724 31720 12733
rect 34520 12724 34572 12776
rect 37372 12767 37424 12776
rect 37372 12733 37381 12767
rect 37381 12733 37415 12767
rect 37415 12733 37424 12767
rect 37372 12724 37424 12733
rect 38660 12928 38712 12980
rect 40040 12860 40092 12912
rect 38384 12792 38436 12844
rect 39580 12767 39632 12776
rect 39580 12733 39589 12767
rect 39589 12733 39623 12767
rect 39623 12733 39632 12767
rect 39580 12724 39632 12733
rect 23480 12656 23532 12708
rect 27068 12656 27120 12708
rect 32220 12656 32272 12708
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 23940 12588 23992 12640
rect 26608 12588 26660 12640
rect 32588 12588 32640 12640
rect 33048 12588 33100 12640
rect 39672 12588 39724 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6644 12384 6696 12436
rect 8208 12384 8260 12436
rect 8668 12384 8720 12436
rect 9312 12384 9364 12436
rect 9496 12384 9548 12436
rect 10784 12427 10836 12436
rect 10784 12393 10793 12427
rect 10793 12393 10827 12427
rect 10827 12393 10836 12427
rect 10784 12384 10836 12393
rect 11704 12384 11756 12436
rect 12992 12384 13044 12436
rect 3700 12248 3752 12300
rect 6092 12248 6144 12300
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 2964 12112 3016 12164
rect 4068 12155 4120 12164
rect 4068 12121 4077 12155
rect 4077 12121 4111 12155
rect 4111 12121 4120 12155
rect 4068 12112 4120 12121
rect 4712 12112 4764 12164
rect 6552 12180 6604 12232
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 2228 12044 2280 12096
rect 6460 12112 6512 12164
rect 7472 12180 7524 12232
rect 8300 12180 8352 12232
rect 7840 12112 7892 12164
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 9680 12248 9732 12300
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 5632 12087 5684 12096
rect 5632 12053 5641 12087
rect 5641 12053 5675 12087
rect 5675 12053 5684 12087
rect 5632 12044 5684 12053
rect 5724 12044 5776 12096
rect 6184 12044 6236 12096
rect 6828 12044 6880 12096
rect 8668 12044 8720 12096
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9036 12044 9088 12053
rect 9128 12044 9180 12096
rect 9220 12044 9272 12096
rect 12072 12248 12124 12300
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 12624 12291 12676 12300
rect 12624 12257 12633 12291
rect 12633 12257 12667 12291
rect 12667 12257 12676 12291
rect 12624 12248 12676 12257
rect 13360 12384 13412 12436
rect 15016 12384 15068 12436
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 12900 12180 12952 12232
rect 16396 12316 16448 12368
rect 18144 12316 18196 12368
rect 19340 12384 19392 12436
rect 22284 12384 22336 12436
rect 23204 12384 23256 12436
rect 20812 12316 20864 12368
rect 21456 12316 21508 12368
rect 15936 12291 15988 12300
rect 15936 12257 15945 12291
rect 15945 12257 15979 12291
rect 15979 12257 15988 12291
rect 15936 12248 15988 12257
rect 16120 12291 16172 12300
rect 16120 12257 16129 12291
rect 16129 12257 16163 12291
rect 16163 12257 16172 12291
rect 16120 12248 16172 12257
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 19616 12248 19668 12300
rect 19984 12248 20036 12300
rect 9588 12044 9640 12096
rect 10324 12044 10376 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 16580 12112 16632 12164
rect 18880 12180 18932 12232
rect 20168 12180 20220 12232
rect 21180 12223 21232 12232
rect 21180 12189 21189 12223
rect 21189 12189 21223 12223
rect 21223 12189 21232 12223
rect 21180 12180 21232 12189
rect 21640 12248 21692 12300
rect 21548 12223 21600 12232
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 14188 12044 14240 12096
rect 15476 12044 15528 12096
rect 15752 12044 15804 12096
rect 16304 12044 16356 12096
rect 18512 12044 18564 12096
rect 19156 12112 19208 12164
rect 20996 12112 21048 12164
rect 21272 12112 21324 12164
rect 21364 12155 21416 12164
rect 21364 12121 21373 12155
rect 21373 12121 21407 12155
rect 21407 12121 21416 12155
rect 21364 12112 21416 12121
rect 22744 12248 22796 12300
rect 23940 12291 23992 12300
rect 23940 12257 23949 12291
rect 23949 12257 23983 12291
rect 23983 12257 23992 12291
rect 23940 12248 23992 12257
rect 22376 12180 22428 12232
rect 28724 12384 28776 12436
rect 28908 12384 28960 12436
rect 30012 12384 30064 12436
rect 30288 12384 30340 12436
rect 24768 12316 24820 12368
rect 21824 12044 21876 12096
rect 22744 12044 22796 12096
rect 23112 12044 23164 12096
rect 23664 12112 23716 12164
rect 25320 12180 25372 12232
rect 25504 12180 25556 12232
rect 26148 12180 26200 12232
rect 26976 12180 27028 12232
rect 27068 12223 27120 12232
rect 27068 12189 27077 12223
rect 27077 12189 27111 12223
rect 27111 12189 27120 12223
rect 27068 12180 27120 12189
rect 27252 12223 27304 12232
rect 27252 12189 27261 12223
rect 27261 12189 27295 12223
rect 27295 12189 27304 12223
rect 27252 12180 27304 12189
rect 27344 12223 27396 12232
rect 27344 12189 27353 12223
rect 27353 12189 27387 12223
rect 27387 12189 27396 12223
rect 27344 12180 27396 12189
rect 30196 12291 30248 12300
rect 30196 12257 30205 12291
rect 30205 12257 30239 12291
rect 30239 12257 30248 12291
rect 30196 12248 30248 12257
rect 30288 12291 30340 12300
rect 30288 12257 30297 12291
rect 30297 12257 30331 12291
rect 30331 12257 30340 12291
rect 30288 12248 30340 12257
rect 29552 12180 29604 12232
rect 30656 12180 30708 12232
rect 31300 12316 31352 12368
rect 31760 12384 31812 12436
rect 39580 12384 39632 12436
rect 33048 12316 33100 12368
rect 31116 12180 31168 12232
rect 31392 12223 31444 12232
rect 31392 12189 31401 12223
rect 31401 12189 31435 12223
rect 31435 12189 31444 12223
rect 31392 12180 31444 12189
rect 31576 12291 31628 12300
rect 31576 12257 31585 12291
rect 31585 12257 31619 12291
rect 31619 12257 31628 12291
rect 31576 12248 31628 12257
rect 33692 12248 33744 12300
rect 35716 12248 35768 12300
rect 40592 12291 40644 12300
rect 40592 12257 40601 12291
rect 40601 12257 40635 12291
rect 40635 12257 40644 12291
rect 40592 12248 40644 12257
rect 31668 12223 31720 12232
rect 31668 12189 31677 12223
rect 31677 12189 31711 12223
rect 31711 12189 31720 12223
rect 31668 12180 31720 12189
rect 24584 12044 24636 12096
rect 24768 12044 24820 12096
rect 26516 12087 26568 12096
rect 26516 12053 26525 12087
rect 26525 12053 26559 12087
rect 26559 12053 26568 12087
rect 26516 12044 26568 12053
rect 26884 12087 26936 12096
rect 26884 12053 26893 12087
rect 26893 12053 26927 12087
rect 26927 12053 26936 12087
rect 26884 12044 26936 12053
rect 28540 12087 28592 12096
rect 28540 12053 28549 12087
rect 28549 12053 28583 12087
rect 28583 12053 28592 12087
rect 28540 12044 28592 12053
rect 30748 12155 30800 12164
rect 30748 12121 30757 12155
rect 30757 12121 30791 12155
rect 30791 12121 30800 12155
rect 30748 12112 30800 12121
rect 30840 12155 30892 12164
rect 30840 12121 30849 12155
rect 30849 12121 30883 12155
rect 30883 12121 30892 12155
rect 30840 12112 30892 12121
rect 31300 12112 31352 12164
rect 32036 12223 32088 12232
rect 32036 12189 32045 12223
rect 32045 12189 32079 12223
rect 32079 12189 32088 12223
rect 32036 12180 32088 12189
rect 32956 12180 33008 12232
rect 34612 12180 34664 12232
rect 38660 12223 38712 12232
rect 38660 12189 38669 12223
rect 38669 12189 38703 12223
rect 38703 12189 38712 12223
rect 38660 12180 38712 12189
rect 38476 12087 38528 12096
rect 38476 12053 38485 12087
rect 38485 12053 38519 12087
rect 38519 12053 38528 12087
rect 38476 12044 38528 12053
rect 41052 12180 41104 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4068 11840 4120 11892
rect 2228 11772 2280 11824
rect 3056 11704 3108 11756
rect 3700 11704 3752 11756
rect 4896 11704 4948 11756
rect 5632 11840 5684 11892
rect 6276 11840 6328 11892
rect 5172 11772 5224 11824
rect 5448 11772 5500 11824
rect 8576 11840 8628 11892
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 4620 11568 4672 11620
rect 1492 11500 1544 11552
rect 2964 11500 3016 11552
rect 5080 11500 5132 11552
rect 6644 11568 6696 11620
rect 6828 11568 6880 11620
rect 8300 11704 8352 11756
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 8760 11840 8812 11892
rect 9036 11840 9088 11892
rect 9128 11840 9180 11892
rect 10324 11840 10376 11892
rect 12808 11840 12860 11892
rect 12900 11840 12952 11892
rect 9128 11679 9180 11688
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 9128 11636 9180 11645
rect 9220 11568 9272 11620
rect 10508 11636 10560 11688
rect 11060 11636 11112 11688
rect 12072 11815 12124 11824
rect 12072 11781 12081 11815
rect 12081 11781 12115 11815
rect 12115 11781 12124 11815
rect 12072 11772 12124 11781
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 15384 11840 15436 11892
rect 16212 11840 16264 11892
rect 17040 11840 17092 11892
rect 18420 11840 18472 11892
rect 18512 11840 18564 11892
rect 20352 11840 20404 11892
rect 20904 11840 20956 11892
rect 21180 11840 21232 11892
rect 21916 11883 21968 11892
rect 21916 11849 21949 11883
rect 21949 11849 21968 11883
rect 21916 11840 21968 11849
rect 22100 11840 22152 11892
rect 24216 11840 24268 11892
rect 14188 11772 14240 11824
rect 15292 11772 15344 11824
rect 12992 11704 13044 11756
rect 14740 11704 14792 11756
rect 15200 11747 15252 11756
rect 15200 11713 15209 11747
rect 15209 11713 15243 11747
rect 15243 11713 15252 11747
rect 15200 11704 15252 11713
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 16028 11704 16080 11756
rect 20260 11772 20312 11824
rect 18144 11704 18196 11756
rect 12624 11636 12676 11688
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 17224 11636 17276 11688
rect 18512 11636 18564 11688
rect 15384 11568 15436 11620
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 6736 11500 6788 11552
rect 8208 11500 8260 11552
rect 8944 11500 8996 11552
rect 11612 11543 11664 11552
rect 11612 11509 11621 11543
rect 11621 11509 11655 11543
rect 11655 11509 11664 11543
rect 11612 11500 11664 11509
rect 12532 11500 12584 11552
rect 15568 11568 15620 11620
rect 16488 11568 16540 11620
rect 17960 11611 18012 11620
rect 17960 11577 17969 11611
rect 17969 11577 18003 11611
rect 18003 11577 18012 11611
rect 17960 11568 18012 11577
rect 18052 11568 18104 11620
rect 18880 11679 18932 11688
rect 18880 11645 18889 11679
rect 18889 11645 18923 11679
rect 18923 11645 18932 11679
rect 18880 11636 18932 11645
rect 20444 11747 20496 11756
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 20444 11704 20496 11713
rect 21272 11772 21324 11824
rect 21456 11772 21508 11824
rect 22008 11772 22060 11824
rect 23480 11772 23532 11824
rect 20904 11704 20956 11756
rect 21180 11747 21232 11756
rect 21180 11713 21189 11747
rect 21189 11713 21223 11747
rect 21223 11713 21232 11747
rect 21180 11704 21232 11713
rect 21272 11636 21324 11688
rect 22100 11704 22152 11756
rect 23204 11704 23256 11756
rect 17132 11500 17184 11552
rect 19892 11568 19944 11620
rect 20720 11568 20772 11620
rect 23664 11704 23716 11756
rect 24308 11772 24360 11824
rect 25044 11840 25096 11892
rect 24860 11815 24912 11824
rect 24860 11781 24869 11815
rect 24869 11781 24903 11815
rect 24903 11781 24912 11815
rect 24860 11772 24912 11781
rect 23848 11704 23900 11756
rect 25596 11840 25648 11892
rect 26516 11840 26568 11892
rect 26884 11840 26936 11892
rect 24768 11636 24820 11688
rect 24492 11568 24544 11620
rect 25688 11704 25740 11756
rect 26240 11704 26292 11756
rect 26332 11747 26384 11756
rect 26332 11713 26341 11747
rect 26341 11713 26375 11747
rect 26375 11713 26384 11747
rect 26332 11704 26384 11713
rect 26516 11747 26568 11756
rect 26516 11713 26530 11747
rect 26530 11713 26564 11747
rect 26564 11713 26568 11747
rect 26516 11704 26568 11713
rect 26976 11747 27028 11756
rect 26976 11713 26985 11747
rect 26985 11713 27019 11747
rect 27019 11713 27028 11747
rect 26976 11704 27028 11713
rect 27068 11704 27120 11756
rect 26792 11636 26844 11688
rect 26056 11568 26108 11620
rect 27344 11636 27396 11688
rect 28632 11840 28684 11892
rect 29276 11840 29328 11892
rect 30012 11840 30064 11892
rect 28540 11815 28592 11824
rect 28540 11781 28549 11815
rect 28549 11781 28583 11815
rect 28583 11781 28592 11815
rect 28540 11772 28592 11781
rect 30196 11772 30248 11824
rect 30472 11840 30524 11892
rect 35716 11772 35768 11824
rect 29644 11704 29696 11756
rect 35532 11636 35584 11688
rect 19616 11500 19668 11552
rect 21364 11500 21416 11552
rect 21824 11500 21876 11552
rect 23204 11500 23256 11552
rect 23756 11543 23808 11552
rect 23756 11509 23765 11543
rect 23765 11509 23799 11543
rect 23799 11509 23808 11543
rect 23756 11500 23808 11509
rect 33600 11568 33652 11620
rect 36084 11747 36136 11756
rect 36084 11713 36093 11747
rect 36093 11713 36127 11747
rect 36127 11713 36136 11747
rect 36084 11704 36136 11713
rect 38384 11772 38436 11824
rect 38844 11772 38896 11824
rect 37556 11636 37608 11688
rect 38476 11636 38528 11688
rect 26884 11500 26936 11552
rect 30472 11500 30524 11552
rect 35716 11543 35768 11552
rect 35716 11509 35725 11543
rect 35725 11509 35759 11543
rect 35759 11509 35768 11543
rect 35716 11500 35768 11509
rect 37464 11568 37516 11620
rect 35992 11500 36044 11552
rect 36544 11500 36596 11552
rect 36728 11500 36780 11552
rect 39856 11543 39908 11552
rect 39856 11509 39865 11543
rect 39865 11509 39899 11543
rect 39899 11509 39908 11543
rect 39856 11500 39908 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 940 11296 992 11348
rect 3056 11296 3108 11348
rect 4620 11296 4672 11348
rect 9036 11296 9088 11348
rect 9404 11296 9456 11348
rect 10876 11296 10928 11348
rect 11704 11228 11756 11280
rect 12072 11271 12124 11280
rect 12072 11237 12081 11271
rect 12081 11237 12115 11271
rect 12115 11237 12124 11271
rect 12072 11228 12124 11237
rect 5172 11160 5224 11212
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 5632 11092 5684 11144
rect 8392 11160 8444 11212
rect 9220 11160 9272 11212
rect 12532 11228 12584 11280
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 2872 11024 2924 11076
rect 6368 11092 6420 11144
rect 9956 11024 10008 11076
rect 12532 11067 12584 11076
rect 12532 11033 12541 11067
rect 12541 11033 12575 11067
rect 12575 11033 12584 11067
rect 12532 11024 12584 11033
rect 13268 11024 13320 11076
rect 13544 11296 13596 11348
rect 17040 11296 17092 11348
rect 18236 11296 18288 11348
rect 18880 11296 18932 11348
rect 19432 11339 19484 11348
rect 19432 11305 19441 11339
rect 19441 11305 19475 11339
rect 19475 11305 19484 11339
rect 19432 11296 19484 11305
rect 18052 11271 18104 11280
rect 18052 11237 18061 11271
rect 18061 11237 18095 11271
rect 18095 11237 18104 11271
rect 20812 11339 20864 11348
rect 20812 11305 20821 11339
rect 20821 11305 20855 11339
rect 20855 11305 20864 11339
rect 20812 11296 20864 11305
rect 21640 11296 21692 11348
rect 22376 11296 22428 11348
rect 23296 11296 23348 11348
rect 18052 11228 18104 11237
rect 14464 11160 14516 11212
rect 15016 11160 15068 11212
rect 14096 11092 14148 11144
rect 6092 10999 6144 11008
rect 6092 10965 6101 10999
rect 6101 10965 6135 10999
rect 6135 10965 6144 10999
rect 6092 10956 6144 10965
rect 6184 10956 6236 11008
rect 9404 10956 9456 11008
rect 9588 10956 9640 11008
rect 11888 10956 11940 11008
rect 13728 10999 13780 11008
rect 13728 10965 13737 10999
rect 13737 10965 13771 10999
rect 13771 10965 13780 10999
rect 13728 10956 13780 10965
rect 14464 10999 14516 11008
rect 14464 10965 14473 10999
rect 14473 10965 14507 10999
rect 14507 10965 14516 10999
rect 14464 10956 14516 10965
rect 14740 11024 14792 11076
rect 15936 11024 15988 11076
rect 16304 11024 16356 11076
rect 18788 11160 18840 11212
rect 17960 11092 18012 11144
rect 18144 11092 18196 11144
rect 16856 10999 16908 11008
rect 16856 10965 16865 10999
rect 16865 10965 16899 10999
rect 16899 10965 16908 10999
rect 16856 10956 16908 10965
rect 17040 11067 17092 11076
rect 17040 11033 17049 11067
rect 17049 11033 17083 11067
rect 17083 11033 17092 11067
rect 17040 11024 17092 11033
rect 18328 11024 18380 11076
rect 18512 11092 18564 11144
rect 19064 11160 19116 11212
rect 19616 11203 19668 11212
rect 19616 11169 19625 11203
rect 19625 11169 19659 11203
rect 19659 11169 19668 11203
rect 19616 11160 19668 11169
rect 18788 11024 18840 11076
rect 17224 10956 17276 11008
rect 18604 10999 18656 11008
rect 18604 10965 18613 10999
rect 18613 10965 18647 10999
rect 18647 10965 18656 10999
rect 18604 10956 18656 10965
rect 19432 11092 19484 11144
rect 22836 11271 22888 11280
rect 22836 11237 22845 11271
rect 22845 11237 22879 11271
rect 22879 11237 22888 11271
rect 22836 11228 22888 11237
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 21364 11203 21416 11212
rect 21364 11169 21373 11203
rect 21373 11169 21407 11203
rect 21407 11169 21416 11203
rect 21364 11160 21416 11169
rect 21456 11160 21508 11212
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 21548 11092 21600 11144
rect 21640 11135 21692 11144
rect 21640 11101 21649 11135
rect 21649 11101 21683 11135
rect 21683 11101 21692 11135
rect 21640 11092 21692 11101
rect 20168 11024 20220 11076
rect 20812 11024 20864 11076
rect 20904 11024 20956 11076
rect 21272 11067 21324 11076
rect 21272 11033 21281 11067
rect 21281 11033 21315 11067
rect 21315 11033 21324 11067
rect 21272 11024 21324 11033
rect 24676 11228 24728 11280
rect 32496 11296 32548 11348
rect 23756 11160 23808 11212
rect 22192 11092 22244 11144
rect 23204 11135 23256 11144
rect 23204 11101 23213 11135
rect 23213 11101 23247 11135
rect 23247 11101 23256 11135
rect 23204 11092 23256 11101
rect 23480 11092 23532 11144
rect 23664 11135 23716 11144
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 24492 11135 24544 11144
rect 24492 11101 24502 11135
rect 24502 11101 24536 11135
rect 24536 11101 24544 11135
rect 25596 11160 25648 11212
rect 25964 11228 26016 11280
rect 26148 11271 26200 11280
rect 26148 11237 26157 11271
rect 26157 11237 26191 11271
rect 26191 11237 26200 11271
rect 26148 11228 26200 11237
rect 26516 11228 26568 11280
rect 24492 11092 24544 11101
rect 24860 11135 24912 11144
rect 24860 11101 24874 11135
rect 24874 11101 24908 11135
rect 24908 11101 24912 11135
rect 24860 11092 24912 11101
rect 25688 11092 25740 11144
rect 22652 11024 22704 11076
rect 24584 11024 24636 11076
rect 22376 10956 22428 11008
rect 23204 10956 23256 11008
rect 25044 10956 25096 11008
rect 25964 11135 26016 11144
rect 25964 11101 25973 11135
rect 25973 11101 26007 11135
rect 26007 11101 26016 11135
rect 25964 11092 26016 11101
rect 26516 11092 26568 11144
rect 26240 11024 26292 11076
rect 26700 11024 26752 11076
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 26976 11135 27028 11144
rect 26976 11101 26986 11135
rect 26986 11101 27020 11135
rect 27020 11101 27028 11135
rect 26976 11092 27028 11101
rect 32588 11228 32640 11280
rect 32128 11160 32180 11212
rect 35716 11296 35768 11348
rect 38660 11296 38712 11348
rect 32772 11160 32824 11212
rect 33508 11160 33560 11212
rect 34796 11203 34848 11212
rect 34796 11169 34805 11203
rect 34805 11169 34839 11203
rect 34839 11169 34848 11203
rect 34796 11160 34848 11169
rect 35992 11160 36044 11212
rect 32680 11092 32732 11144
rect 25872 10956 25924 11008
rect 30656 10956 30708 11008
rect 33416 10956 33468 11008
rect 36084 11092 36136 11144
rect 35532 11024 35584 11076
rect 36728 11160 36780 11212
rect 38752 11160 38804 11212
rect 35256 10999 35308 11008
rect 35256 10965 35265 10999
rect 35265 10965 35299 10999
rect 35299 10965 35308 10999
rect 35256 10956 35308 10965
rect 38016 11092 38068 11144
rect 39856 11228 39908 11280
rect 39672 11160 39724 11212
rect 39028 11024 39080 11076
rect 36820 10999 36872 11008
rect 36820 10965 36829 10999
rect 36829 10965 36863 10999
rect 36863 10965 36872 10999
rect 36820 10956 36872 10965
rect 38660 10999 38712 11008
rect 38660 10965 38669 10999
rect 38669 10965 38703 10999
rect 38703 10965 38712 10999
rect 38660 10956 38712 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3976 10752 4028 10804
rect 7932 10752 7984 10804
rect 8852 10752 8904 10804
rect 8576 10616 8628 10668
rect 8760 10616 8812 10668
rect 9588 10752 9640 10804
rect 9864 10752 9916 10804
rect 13728 10752 13780 10804
rect 14464 10752 14516 10804
rect 15476 10752 15528 10804
rect 18236 10752 18288 10804
rect 18512 10795 18564 10804
rect 18512 10761 18530 10795
rect 18530 10761 18564 10795
rect 18512 10752 18564 10761
rect 18788 10752 18840 10804
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 8484 10591 8536 10600
rect 8484 10557 8493 10591
rect 8493 10557 8527 10591
rect 8527 10557 8536 10591
rect 8484 10548 8536 10557
rect 9312 10548 9364 10600
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11060 10616 11112 10668
rect 13176 10616 13228 10668
rect 15016 10616 15068 10668
rect 15568 10727 15620 10736
rect 15568 10693 15577 10727
rect 15577 10693 15611 10727
rect 15611 10693 15620 10727
rect 15568 10684 15620 10693
rect 17132 10727 17184 10736
rect 17132 10693 17141 10727
rect 17141 10693 17175 10727
rect 17175 10693 17184 10727
rect 17132 10684 17184 10693
rect 18052 10684 18104 10736
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 8116 10412 8168 10464
rect 9588 10412 9640 10464
rect 13636 10548 13688 10600
rect 14096 10548 14148 10600
rect 16856 10616 16908 10668
rect 19984 10752 20036 10804
rect 19432 10684 19484 10736
rect 20812 10684 20864 10736
rect 21824 10684 21876 10736
rect 23480 10727 23532 10736
rect 23480 10693 23489 10727
rect 23489 10693 23523 10727
rect 23523 10693 23532 10727
rect 23480 10684 23532 10693
rect 24676 10684 24728 10736
rect 25228 10684 25280 10736
rect 26516 10752 26568 10804
rect 26884 10752 26936 10804
rect 27436 10752 27488 10804
rect 32128 10752 32180 10804
rect 15844 10548 15896 10600
rect 16488 10548 16540 10600
rect 18604 10548 18656 10600
rect 22836 10616 22888 10668
rect 23204 10616 23256 10668
rect 20168 10548 20220 10600
rect 20260 10548 20312 10600
rect 24032 10616 24084 10668
rect 25688 10659 25740 10668
rect 25688 10625 25697 10659
rect 25697 10625 25731 10659
rect 25731 10625 25740 10659
rect 25688 10616 25740 10625
rect 10968 10480 11020 10532
rect 16948 10480 17000 10532
rect 11336 10412 11388 10464
rect 15844 10455 15896 10464
rect 15844 10421 15853 10455
rect 15853 10421 15887 10455
rect 15887 10421 15896 10455
rect 15844 10412 15896 10421
rect 18420 10412 18472 10464
rect 21088 10480 21140 10532
rect 20352 10412 20404 10464
rect 25412 10591 25464 10600
rect 25412 10557 25421 10591
rect 25421 10557 25455 10591
rect 25455 10557 25464 10591
rect 25412 10548 25464 10557
rect 25964 10659 26016 10668
rect 25964 10625 25973 10659
rect 25973 10625 26007 10659
rect 26007 10625 26016 10659
rect 25964 10616 26016 10625
rect 26056 10659 26108 10668
rect 26056 10625 26065 10659
rect 26065 10625 26099 10659
rect 26099 10625 26108 10659
rect 26056 10616 26108 10625
rect 26240 10616 26292 10668
rect 27344 10684 27396 10736
rect 30380 10684 30432 10736
rect 26700 10616 26752 10668
rect 26792 10616 26844 10668
rect 33232 10752 33284 10804
rect 33600 10752 33652 10804
rect 34796 10752 34848 10804
rect 35256 10752 35308 10804
rect 38660 10795 38712 10804
rect 38660 10761 38669 10795
rect 38669 10761 38703 10795
rect 38703 10761 38712 10795
rect 38660 10752 38712 10761
rect 38752 10752 38804 10804
rect 32588 10684 32640 10736
rect 30288 10591 30340 10600
rect 30288 10557 30297 10591
rect 30297 10557 30331 10591
rect 30331 10557 30340 10591
rect 30288 10548 30340 10557
rect 31392 10591 31444 10600
rect 31392 10557 31401 10591
rect 31401 10557 31435 10591
rect 31435 10557 31444 10591
rect 31392 10548 31444 10557
rect 33048 10659 33100 10668
rect 33048 10625 33057 10659
rect 33057 10625 33091 10659
rect 33091 10625 33100 10659
rect 33048 10616 33100 10625
rect 32864 10548 32916 10600
rect 31668 10480 31720 10532
rect 33600 10591 33652 10600
rect 33600 10557 33609 10591
rect 33609 10557 33643 10591
rect 33643 10557 33652 10591
rect 33600 10548 33652 10557
rect 33784 10659 33836 10668
rect 33784 10625 33793 10659
rect 33793 10625 33827 10659
rect 33827 10625 33836 10659
rect 33784 10616 33836 10625
rect 34612 10616 34664 10668
rect 36820 10684 36872 10736
rect 35992 10591 36044 10600
rect 35992 10557 36001 10591
rect 36001 10557 36035 10591
rect 36035 10557 36044 10591
rect 35992 10548 36044 10557
rect 39120 10591 39172 10600
rect 39120 10557 39129 10591
rect 39129 10557 39163 10591
rect 39163 10557 39172 10591
rect 39120 10548 39172 10557
rect 39304 10591 39356 10600
rect 39304 10557 39313 10591
rect 39313 10557 39347 10591
rect 39347 10557 39356 10591
rect 39304 10548 39356 10557
rect 25964 10412 26016 10464
rect 29736 10455 29788 10464
rect 29736 10421 29745 10455
rect 29745 10421 29779 10455
rect 29779 10421 29788 10455
rect 29736 10412 29788 10421
rect 33140 10412 33192 10464
rect 33508 10455 33560 10464
rect 33508 10421 33517 10455
rect 33517 10421 33551 10455
rect 33551 10421 33560 10455
rect 33508 10412 33560 10421
rect 34796 10412 34848 10464
rect 36084 10455 36136 10464
rect 36084 10421 36093 10455
rect 36093 10421 36127 10455
rect 36127 10421 36136 10455
rect 36084 10412 36136 10421
rect 38660 10412 38712 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 5172 10208 5224 10260
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 4620 9979 4672 9988
rect 4620 9945 4629 9979
rect 4629 9945 4663 9979
rect 4663 9945 4672 9979
rect 4620 9936 4672 9945
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 6736 10140 6788 10192
rect 6828 10140 6880 10192
rect 8392 10208 8444 10260
rect 9588 10208 9640 10260
rect 11612 10208 11664 10260
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 15844 10208 15896 10260
rect 18880 10251 18932 10260
rect 18880 10217 18889 10251
rect 18889 10217 18923 10251
rect 18923 10217 18932 10251
rect 18880 10208 18932 10217
rect 20720 10208 20772 10260
rect 23848 10208 23900 10260
rect 24032 10208 24084 10260
rect 24952 10208 25004 10260
rect 25504 10208 25556 10260
rect 25964 10208 26016 10260
rect 26424 10208 26476 10260
rect 29736 10208 29788 10260
rect 31392 10208 31444 10260
rect 33048 10208 33100 10260
rect 6276 10047 6328 10056
rect 5632 9936 5684 9988
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 7104 10072 7156 10124
rect 8116 10140 8168 10192
rect 8208 10140 8260 10192
rect 9128 10072 9180 10124
rect 5080 9911 5132 9920
rect 5080 9877 5089 9911
rect 5089 9877 5123 9911
rect 5123 9877 5132 9911
rect 5080 9868 5132 9877
rect 6552 9979 6604 9988
rect 6552 9945 6561 9979
rect 6561 9945 6595 9979
rect 6595 9945 6604 9979
rect 6552 9936 6604 9945
rect 6920 9936 6972 9988
rect 9496 10004 9548 10056
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 11336 10140 11388 10192
rect 11980 10072 12032 10124
rect 11152 10047 11204 10056
rect 11152 10013 11159 10047
rect 11159 10013 11204 10047
rect 11152 10004 11204 10013
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11428 10047 11480 10056
rect 11428 10013 11442 10047
rect 11442 10013 11476 10047
rect 11476 10013 11480 10047
rect 11428 10004 11480 10013
rect 11888 10047 11940 10056
rect 11888 10013 11897 10047
rect 11897 10013 11931 10047
rect 11931 10013 11940 10047
rect 11888 10004 11940 10013
rect 23480 10140 23532 10192
rect 21456 10072 21508 10124
rect 22376 10072 22428 10124
rect 8300 9936 8352 9988
rect 8392 9979 8444 9988
rect 8392 9945 8401 9979
rect 8401 9945 8435 9979
rect 8435 9945 8444 9979
rect 8392 9936 8444 9945
rect 7748 9868 7800 9920
rect 9220 9868 9272 9920
rect 10968 9868 11020 9920
rect 11612 9911 11664 9920
rect 11612 9877 11621 9911
rect 11621 9877 11655 9911
rect 11655 9877 11664 9911
rect 11612 9868 11664 9877
rect 15476 9868 15528 9920
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 18880 10004 18932 10056
rect 21732 10047 21784 10056
rect 21732 10013 21741 10047
rect 21741 10013 21775 10047
rect 21775 10013 21784 10047
rect 21732 10004 21784 10013
rect 22468 10004 22520 10056
rect 23204 10047 23256 10056
rect 19248 9936 19300 9988
rect 22008 9979 22060 9988
rect 22008 9945 22017 9979
rect 22017 9945 22051 9979
rect 22051 9945 22060 9979
rect 22008 9936 22060 9945
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 22744 9868 22796 9920
rect 25688 10072 25740 10124
rect 25228 10004 25280 10056
rect 25320 10004 25372 10056
rect 26976 10004 27028 10056
rect 27988 10047 28040 10056
rect 27988 10013 27997 10047
rect 27997 10013 28031 10047
rect 28031 10013 28040 10047
rect 27988 10004 28040 10013
rect 32588 10183 32640 10192
rect 32588 10149 32597 10183
rect 32597 10149 32631 10183
rect 32631 10149 32640 10183
rect 32588 10140 32640 10149
rect 31116 10072 31168 10124
rect 31300 10072 31352 10124
rect 35992 10208 36044 10260
rect 39120 10208 39172 10260
rect 34704 10140 34756 10192
rect 30656 10047 30708 10056
rect 30656 10013 30665 10047
rect 30665 10013 30699 10047
rect 30699 10013 30708 10047
rect 30656 10004 30708 10013
rect 32496 10047 32548 10056
rect 32496 10013 32505 10047
rect 32505 10013 32539 10047
rect 32539 10013 32548 10047
rect 32496 10004 32548 10013
rect 25872 9936 25924 9988
rect 30472 9936 30524 9988
rect 33048 10047 33100 10056
rect 33048 10013 33057 10047
rect 33057 10013 33091 10047
rect 33091 10013 33100 10047
rect 33048 10004 33100 10013
rect 33140 10047 33192 10056
rect 33140 10013 33149 10047
rect 33149 10013 33183 10047
rect 33183 10013 33192 10047
rect 33140 10004 33192 10013
rect 33784 9936 33836 9988
rect 34612 10004 34664 10056
rect 34796 10004 34848 10056
rect 39028 10115 39080 10124
rect 39028 10081 39037 10115
rect 39037 10081 39071 10115
rect 39071 10081 39080 10115
rect 39028 10072 39080 10081
rect 35256 9936 35308 9988
rect 39212 10047 39264 10056
rect 39212 10013 39221 10047
rect 39221 10013 39255 10047
rect 39255 10013 39264 10047
rect 39212 10004 39264 10013
rect 39396 10004 39448 10056
rect 39764 10072 39816 10124
rect 39856 10004 39908 10056
rect 27804 9911 27856 9920
rect 27804 9877 27813 9911
rect 27813 9877 27847 9911
rect 27847 9877 27856 9911
rect 27804 9868 27856 9877
rect 29184 9911 29236 9920
rect 29184 9877 29193 9911
rect 29193 9877 29227 9911
rect 29227 9877 29236 9911
rect 29184 9868 29236 9877
rect 32680 9868 32732 9920
rect 32772 9911 32824 9920
rect 32772 9877 32781 9911
rect 32781 9877 32815 9911
rect 32815 9877 32824 9911
rect 32772 9868 32824 9877
rect 34612 9868 34664 9920
rect 34796 9868 34848 9920
rect 39396 9911 39448 9920
rect 39396 9877 39405 9911
rect 39405 9877 39439 9911
rect 39439 9877 39448 9911
rect 39396 9868 39448 9877
rect 39580 9911 39632 9920
rect 39580 9877 39589 9911
rect 39589 9877 39623 9911
rect 39623 9877 39632 9911
rect 39580 9868 39632 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4896 9639 4948 9648
rect 4896 9605 4905 9639
rect 4905 9605 4939 9639
rect 4939 9605 4948 9639
rect 4896 9596 4948 9605
rect 5356 9596 5408 9648
rect 8024 9596 8076 9648
rect 8760 9596 8812 9648
rect 4620 9528 4672 9580
rect 4344 9392 4396 9444
rect 5080 9460 5132 9512
rect 4620 9392 4672 9444
rect 5172 9392 5224 9444
rect 5448 9324 5500 9376
rect 7748 9528 7800 9580
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 6460 9460 6512 9512
rect 6368 9367 6420 9376
rect 6368 9333 6377 9367
rect 6377 9333 6411 9367
rect 6411 9333 6420 9367
rect 6368 9324 6420 9333
rect 7104 9392 7156 9444
rect 9864 9571 9916 9580
rect 9864 9537 9873 9571
rect 9873 9537 9907 9571
rect 9907 9537 9916 9571
rect 9864 9528 9916 9537
rect 10784 9664 10836 9716
rect 11152 9664 11204 9716
rect 10508 9596 10560 9648
rect 15476 9664 15528 9716
rect 16304 9664 16356 9716
rect 21732 9664 21784 9716
rect 21916 9664 21968 9716
rect 25412 9664 25464 9716
rect 15200 9596 15252 9648
rect 15568 9596 15620 9648
rect 15936 9639 15988 9648
rect 15936 9605 15945 9639
rect 15945 9605 15979 9639
rect 15979 9605 15988 9639
rect 15936 9596 15988 9605
rect 19524 9596 19576 9648
rect 20076 9596 20128 9648
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 12072 9528 12124 9580
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 7932 9324 7984 9376
rect 16580 9528 16632 9580
rect 16764 9528 16816 9580
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 17132 9528 17184 9580
rect 16120 9503 16172 9512
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 19340 9460 19392 9512
rect 20720 9528 20772 9580
rect 20444 9460 20496 9512
rect 22928 9596 22980 9648
rect 23020 9596 23072 9648
rect 17592 9392 17644 9444
rect 15476 9367 15528 9376
rect 15476 9333 15485 9367
rect 15485 9333 15519 9367
rect 15519 9333 15528 9367
rect 15476 9324 15528 9333
rect 15568 9324 15620 9376
rect 22008 9528 22060 9580
rect 25228 9571 25280 9580
rect 25228 9537 25237 9571
rect 25237 9537 25271 9571
rect 25271 9537 25280 9571
rect 25228 9528 25280 9537
rect 25320 9528 25372 9580
rect 21456 9460 21508 9512
rect 25688 9571 25740 9580
rect 25688 9537 25697 9571
rect 25697 9537 25731 9571
rect 25731 9537 25740 9571
rect 25688 9528 25740 9537
rect 25964 9528 26016 9580
rect 26424 9528 26476 9580
rect 26608 9528 26660 9580
rect 27160 9528 27212 9580
rect 27528 9528 27580 9580
rect 25872 9392 25924 9444
rect 26884 9460 26936 9512
rect 30380 9707 30432 9716
rect 30380 9673 30389 9707
rect 30389 9673 30423 9707
rect 30423 9673 30432 9707
rect 30380 9664 30432 9673
rect 31116 9707 31168 9716
rect 31116 9673 31125 9707
rect 31125 9673 31159 9707
rect 31159 9673 31168 9707
rect 31116 9664 31168 9673
rect 32680 9664 32732 9716
rect 32864 9664 32916 9716
rect 35256 9664 35308 9716
rect 38568 9664 38620 9716
rect 29184 9596 29236 9648
rect 29644 9596 29696 9648
rect 28540 9528 28592 9580
rect 28632 9571 28684 9580
rect 28632 9537 28641 9571
rect 28641 9537 28675 9571
rect 28675 9537 28684 9571
rect 28632 9528 28684 9537
rect 32772 9596 32824 9648
rect 36176 9596 36228 9648
rect 37096 9596 37148 9648
rect 37188 9596 37240 9648
rect 39212 9664 39264 9716
rect 39856 9707 39908 9716
rect 39856 9673 39865 9707
rect 39865 9673 39899 9707
rect 39899 9673 39908 9707
rect 39856 9664 39908 9673
rect 32588 9528 32640 9580
rect 27896 9503 27948 9512
rect 27896 9469 27905 9503
rect 27905 9469 27939 9503
rect 27939 9469 27948 9503
rect 27896 9460 27948 9469
rect 27988 9460 28040 9512
rect 30656 9503 30708 9512
rect 30656 9469 30665 9503
rect 30665 9469 30699 9503
rect 30699 9469 30708 9503
rect 30656 9460 30708 9469
rect 37372 9528 37424 9580
rect 37924 9571 37976 9580
rect 37924 9537 37933 9571
rect 37933 9537 37967 9571
rect 37967 9537 37976 9571
rect 37924 9528 37976 9537
rect 39396 9528 39448 9580
rect 38568 9460 38620 9512
rect 38660 9392 38712 9444
rect 39580 9571 39632 9580
rect 39580 9537 39589 9571
rect 39589 9537 39623 9571
rect 39623 9537 39632 9571
rect 39580 9528 39632 9537
rect 39764 9392 39816 9444
rect 18972 9367 19024 9376
rect 18972 9333 18981 9367
rect 18981 9333 19015 9367
rect 19015 9333 19024 9367
rect 18972 9324 19024 9333
rect 19340 9324 19392 9376
rect 21456 9367 21508 9376
rect 21456 9333 21465 9367
rect 21465 9333 21499 9367
rect 21499 9333 21508 9367
rect 21456 9324 21508 9333
rect 22008 9367 22060 9376
rect 22008 9333 22017 9367
rect 22017 9333 22051 9367
rect 22051 9333 22060 9367
rect 22008 9324 22060 9333
rect 26148 9324 26200 9376
rect 26332 9367 26384 9376
rect 26332 9333 26341 9367
rect 26341 9333 26375 9367
rect 26375 9333 26384 9367
rect 26332 9324 26384 9333
rect 26792 9324 26844 9376
rect 32220 9367 32272 9376
rect 32220 9333 32229 9367
rect 32229 9333 32263 9367
rect 32263 9333 32272 9367
rect 32220 9324 32272 9333
rect 33140 9324 33192 9376
rect 36452 9324 36504 9376
rect 36912 9324 36964 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4804 9120 4856 9172
rect 5448 9120 5500 9172
rect 8576 9163 8628 9172
rect 8576 9129 8585 9163
rect 8585 9129 8619 9163
rect 8619 9129 8628 9163
rect 8576 9120 8628 9129
rect 10968 9120 11020 9172
rect 13912 9120 13964 9172
rect 15476 9120 15528 9172
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 19524 9163 19576 9172
rect 19524 9129 19533 9163
rect 19533 9129 19567 9163
rect 19567 9129 19576 9163
rect 19524 9120 19576 9129
rect 4896 8984 4948 9036
rect 8300 9052 8352 9104
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 6092 8916 6144 8968
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 7748 8984 7800 9036
rect 9128 8984 9180 9036
rect 9312 8984 9364 9036
rect 9496 8984 9548 9036
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 9588 8916 9640 8968
rect 8484 8848 8536 8900
rect 11612 8916 11664 8968
rect 19984 9052 20036 9104
rect 16212 8916 16264 8968
rect 16764 8984 16816 9036
rect 17960 8984 18012 9036
rect 21456 8984 21508 9036
rect 16488 8959 16540 8968
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 16856 8916 16908 8968
rect 17040 8916 17092 8968
rect 18972 8916 19024 8968
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 22008 9120 22060 9172
rect 22468 9120 22520 9172
rect 23112 9120 23164 9172
rect 26700 9120 26752 9172
rect 25596 9052 25648 9104
rect 27620 9120 27672 9172
rect 28632 9120 28684 9172
rect 28540 9052 28592 9104
rect 22008 8984 22060 9036
rect 23756 8916 23808 8968
rect 25320 8916 25372 8968
rect 26332 8916 26384 8968
rect 17132 8891 17184 8900
rect 17132 8857 17141 8891
rect 17141 8857 17175 8891
rect 17175 8857 17184 8891
rect 17132 8848 17184 8857
rect 26884 9027 26936 9036
rect 26884 8993 26893 9027
rect 26893 8993 26927 9027
rect 26927 8993 26936 9027
rect 26884 8984 26936 8993
rect 26976 9027 27028 9036
rect 26976 8993 26985 9027
rect 26985 8993 27019 9027
rect 27019 8993 27028 9027
rect 26976 8984 27028 8993
rect 27160 8984 27212 9036
rect 32312 9052 32364 9104
rect 33876 9052 33928 9104
rect 33140 8984 33192 9036
rect 26792 8959 26844 8968
rect 26792 8925 26801 8959
rect 26801 8925 26835 8959
rect 26835 8925 26844 8959
rect 26792 8916 26844 8925
rect 28632 8916 28684 8968
rect 29644 8916 29696 8968
rect 30288 8916 30340 8968
rect 31668 8916 31720 8968
rect 7656 8780 7708 8832
rect 10232 8780 10284 8832
rect 14096 8780 14148 8832
rect 15016 8780 15068 8832
rect 16580 8780 16632 8832
rect 16764 8780 16816 8832
rect 18420 8780 18472 8832
rect 23480 8780 23532 8832
rect 25136 8780 25188 8832
rect 26424 8823 26476 8832
rect 26424 8789 26433 8823
rect 26433 8789 26467 8823
rect 26467 8789 26476 8823
rect 26424 8780 26476 8789
rect 27436 8848 27488 8900
rect 27804 8848 27856 8900
rect 31760 8848 31812 8900
rect 33232 8916 33284 8968
rect 34520 9120 34572 9172
rect 33600 8848 33652 8900
rect 31116 8780 31168 8832
rect 33048 8823 33100 8832
rect 33048 8789 33057 8823
rect 33057 8789 33091 8823
rect 33091 8789 33100 8823
rect 34612 8916 34664 8968
rect 34060 8848 34112 8900
rect 35808 8916 35860 8968
rect 36084 8916 36136 8968
rect 36452 9027 36504 9036
rect 36452 8993 36461 9027
rect 36461 8993 36495 9027
rect 36495 8993 36504 9027
rect 36452 8984 36504 8993
rect 36912 8984 36964 9036
rect 33048 8780 33100 8789
rect 34520 8780 34572 8832
rect 37096 8959 37148 8968
rect 37096 8925 37110 8959
rect 37110 8925 37144 8959
rect 37144 8925 37148 8959
rect 37096 8916 37148 8925
rect 37372 8959 37424 8968
rect 37372 8925 37381 8959
rect 37381 8925 37415 8959
rect 37415 8925 37424 8959
rect 37372 8916 37424 8925
rect 37924 8916 37976 8968
rect 38568 9027 38620 9036
rect 38568 8993 38577 9027
rect 38577 8993 38611 9027
rect 38611 8993 38620 9027
rect 38568 8984 38620 8993
rect 38660 8984 38712 9036
rect 37280 8823 37332 8832
rect 37280 8789 37289 8823
rect 37289 8789 37323 8823
rect 37323 8789 37332 8823
rect 37280 8780 37332 8789
rect 37464 8780 37516 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 3884 8576 3936 8628
rect 4896 8576 4948 8628
rect 10048 8576 10100 8628
rect 10416 8576 10468 8628
rect 4620 8508 4672 8560
rect 4620 8236 4672 8288
rect 6552 8372 6604 8424
rect 8208 8372 8260 8424
rect 9404 8440 9456 8492
rect 13728 8508 13780 8560
rect 14096 8508 14148 8560
rect 14280 8576 14332 8628
rect 15292 8576 15344 8628
rect 16580 8508 16632 8560
rect 17132 8576 17184 8628
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 14832 8483 14884 8492
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 15016 8440 15068 8492
rect 16212 8440 16264 8492
rect 9496 8372 9548 8424
rect 9680 8372 9732 8424
rect 10600 8372 10652 8424
rect 12440 8372 12492 8424
rect 13820 8415 13872 8424
rect 13820 8381 13829 8415
rect 13829 8381 13863 8415
rect 13863 8381 13872 8415
rect 13820 8372 13872 8381
rect 5540 8304 5592 8356
rect 10048 8304 10100 8356
rect 5724 8236 5776 8288
rect 7932 8236 7984 8288
rect 17316 8508 17368 8560
rect 18420 8576 18472 8628
rect 20168 8576 20220 8628
rect 23296 8576 23348 8628
rect 24124 8619 24176 8628
rect 24124 8585 24133 8619
rect 24133 8585 24167 8619
rect 24167 8585 24176 8619
rect 24124 8576 24176 8585
rect 26424 8576 26476 8628
rect 27620 8576 27672 8628
rect 27896 8576 27948 8628
rect 30656 8576 30708 8628
rect 31392 8576 31444 8628
rect 32220 8576 32272 8628
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 19340 8440 19392 8492
rect 25504 8508 25556 8560
rect 17040 8372 17092 8424
rect 16948 8304 17000 8356
rect 18696 8372 18748 8424
rect 19432 8372 19484 8424
rect 19892 8304 19944 8356
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 20168 8483 20220 8492
rect 20168 8449 20177 8483
rect 20177 8449 20211 8483
rect 20211 8449 20220 8483
rect 20168 8440 20220 8449
rect 20352 8440 20404 8492
rect 21548 8440 21600 8492
rect 22192 8440 22244 8492
rect 23756 8440 23808 8492
rect 24952 8483 25004 8492
rect 24952 8449 24961 8483
rect 24961 8449 24995 8483
rect 24995 8449 25004 8483
rect 24952 8440 25004 8449
rect 28632 8508 28684 8560
rect 30104 8508 30156 8560
rect 21180 8372 21232 8424
rect 17408 8236 17460 8288
rect 19708 8236 19760 8288
rect 22284 8304 22336 8356
rect 25228 8372 25280 8424
rect 24492 8304 24544 8356
rect 23296 8236 23348 8288
rect 30288 8483 30340 8492
rect 30288 8449 30297 8483
rect 30297 8449 30331 8483
rect 30331 8449 30340 8483
rect 30288 8440 30340 8449
rect 31116 8551 31168 8560
rect 31116 8517 31125 8551
rect 31125 8517 31159 8551
rect 31159 8517 31168 8551
rect 31116 8508 31168 8517
rect 30564 8372 30616 8424
rect 31668 8440 31720 8492
rect 33600 8508 33652 8560
rect 34060 8619 34112 8628
rect 34060 8585 34069 8619
rect 34069 8585 34103 8619
rect 34103 8585 34112 8619
rect 34060 8576 34112 8585
rect 31116 8236 31168 8288
rect 32036 8372 32088 8424
rect 33876 8483 33928 8492
rect 33876 8449 33885 8483
rect 33885 8449 33919 8483
rect 33919 8449 33928 8483
rect 33876 8440 33928 8449
rect 34520 8508 34572 8560
rect 34428 8440 34480 8492
rect 34704 8440 34756 8492
rect 35808 8576 35860 8628
rect 37188 8576 37240 8628
rect 37280 8576 37332 8628
rect 37464 8508 37516 8560
rect 37648 8508 37700 8560
rect 38844 8508 38896 8560
rect 33692 8304 33744 8356
rect 31392 8236 31444 8288
rect 31484 8279 31536 8288
rect 31484 8245 31493 8279
rect 31493 8245 31527 8279
rect 31527 8245 31536 8279
rect 31484 8236 31536 8245
rect 32220 8236 32272 8288
rect 37188 8440 37240 8492
rect 40684 8483 40736 8492
rect 40684 8449 40693 8483
rect 40693 8449 40727 8483
rect 40727 8449 40736 8483
rect 40684 8440 40736 8449
rect 35532 8415 35584 8424
rect 35532 8381 35541 8415
rect 35541 8381 35575 8415
rect 35575 8381 35584 8415
rect 35532 8372 35584 8381
rect 36176 8372 36228 8424
rect 37280 8415 37332 8424
rect 37280 8381 37289 8415
rect 37289 8381 37323 8415
rect 37323 8381 37332 8415
rect 37280 8372 37332 8381
rect 41052 8304 41104 8356
rect 35440 8279 35492 8288
rect 35440 8245 35449 8279
rect 35449 8245 35483 8279
rect 35483 8245 35492 8279
rect 35440 8236 35492 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 12440 8032 12492 8084
rect 15660 8032 15712 8084
rect 16396 8032 16448 8084
rect 16856 8032 16908 8084
rect 20904 8075 20956 8084
rect 20904 8041 20913 8075
rect 20913 8041 20947 8075
rect 20947 8041 20956 8075
rect 20904 8032 20956 8041
rect 21088 8032 21140 8084
rect 21824 8032 21876 8084
rect 22192 8032 22244 8084
rect 24768 8032 24820 8084
rect 26056 8032 26108 8084
rect 4620 7896 4672 7948
rect 5724 7896 5776 7948
rect 940 7828 992 7880
rect 6368 7828 6420 7880
rect 4068 7760 4120 7812
rect 4712 7760 4764 7812
rect 7564 7760 7616 7812
rect 7656 7760 7708 7812
rect 8668 7828 8720 7880
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 14556 7964 14608 8016
rect 13544 7939 13596 7948
rect 13544 7905 13553 7939
rect 13553 7905 13587 7939
rect 13587 7905 13596 7939
rect 13544 7896 13596 7905
rect 16672 7964 16724 8016
rect 11336 7828 11388 7880
rect 11704 7803 11756 7812
rect 11704 7769 11713 7803
rect 11713 7769 11747 7803
rect 11747 7769 11756 7803
rect 11704 7760 11756 7769
rect 5724 7735 5776 7744
rect 5724 7701 5733 7735
rect 5733 7701 5767 7735
rect 5767 7701 5776 7735
rect 5724 7692 5776 7701
rect 7104 7692 7156 7744
rect 7932 7692 7984 7744
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 9496 7692 9548 7744
rect 10140 7692 10192 7744
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 13820 7828 13872 7880
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 16396 7828 16448 7880
rect 16488 7828 16540 7880
rect 16580 7828 16632 7880
rect 16764 7828 16816 7880
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 17408 7828 17460 7880
rect 22744 7896 22796 7948
rect 22928 7939 22980 7948
rect 22928 7905 22937 7939
rect 22937 7905 22971 7939
rect 22971 7905 22980 7939
rect 22928 7896 22980 7905
rect 25596 7896 25648 7948
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 14740 7760 14792 7812
rect 14924 7803 14976 7812
rect 14924 7769 14933 7803
rect 14933 7769 14967 7803
rect 14967 7769 14976 7803
rect 14924 7760 14976 7769
rect 15200 7760 15252 7812
rect 15752 7803 15804 7812
rect 15752 7769 15761 7803
rect 15761 7769 15795 7803
rect 15795 7769 15804 7803
rect 15752 7760 15804 7769
rect 18604 7760 18656 7812
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 19984 7828 20036 7880
rect 21088 7871 21140 7880
rect 21088 7837 21097 7871
rect 21097 7837 21131 7871
rect 21131 7837 21140 7871
rect 21088 7828 21140 7837
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 21364 7871 21416 7880
rect 21364 7837 21373 7871
rect 21373 7837 21407 7871
rect 21407 7837 21416 7871
rect 21364 7828 21416 7837
rect 21640 7828 21692 7880
rect 22008 7828 22060 7880
rect 23296 7828 23348 7880
rect 25136 7828 25188 7880
rect 25228 7871 25280 7880
rect 25228 7837 25237 7871
rect 25237 7837 25271 7871
rect 25271 7837 25280 7871
rect 25228 7828 25280 7837
rect 25320 7871 25372 7880
rect 25320 7837 25329 7871
rect 25329 7837 25363 7871
rect 25363 7837 25372 7871
rect 25320 7828 25372 7837
rect 25688 7871 25740 7880
rect 25688 7837 25697 7871
rect 25697 7837 25731 7871
rect 25731 7837 25740 7871
rect 25688 7828 25740 7837
rect 28080 7964 28132 8016
rect 34612 8032 34664 8084
rect 30564 7939 30616 7948
rect 30564 7905 30573 7939
rect 30573 7905 30607 7939
rect 30607 7905 30616 7939
rect 30564 7896 30616 7905
rect 31116 7939 31168 7948
rect 31116 7905 31125 7939
rect 31125 7905 31159 7939
rect 31159 7905 31168 7939
rect 31116 7896 31168 7905
rect 34612 7896 34664 7948
rect 35532 7964 35584 8016
rect 25964 7871 26016 7880
rect 25964 7837 25973 7871
rect 25973 7837 26007 7871
rect 26007 7837 26016 7871
rect 25964 7828 26016 7837
rect 26148 7871 26200 7880
rect 26148 7837 26162 7871
rect 26162 7837 26196 7871
rect 26196 7837 26200 7871
rect 26148 7828 26200 7837
rect 13452 7692 13504 7744
rect 14280 7692 14332 7744
rect 16120 7735 16172 7744
rect 16120 7701 16129 7735
rect 16129 7701 16163 7735
rect 16163 7701 16172 7735
rect 16120 7692 16172 7701
rect 17224 7735 17276 7744
rect 17224 7701 17233 7735
rect 17233 7701 17267 7735
rect 17267 7701 17276 7735
rect 17224 7692 17276 7701
rect 19064 7692 19116 7744
rect 21180 7692 21232 7744
rect 22652 7692 22704 7744
rect 22744 7735 22796 7744
rect 22744 7701 22753 7735
rect 22753 7701 22787 7735
rect 22787 7701 22796 7735
rect 22744 7692 22796 7701
rect 24216 7692 24268 7744
rect 26056 7803 26108 7812
rect 26056 7769 26065 7803
rect 26065 7769 26099 7803
rect 26099 7769 26108 7803
rect 26056 7760 26108 7769
rect 31484 7828 31536 7880
rect 33048 7828 33100 7880
rect 33692 7871 33744 7880
rect 33692 7837 33701 7871
rect 33701 7837 33735 7871
rect 33735 7837 33744 7871
rect 33692 7828 33744 7837
rect 34060 7828 34112 7880
rect 34520 7871 34572 7880
rect 34520 7837 34529 7871
rect 34529 7837 34563 7871
rect 34563 7837 34572 7871
rect 34520 7828 34572 7837
rect 32220 7760 32272 7812
rect 37832 7896 37884 7948
rect 26332 7735 26384 7744
rect 26332 7701 26341 7735
rect 26341 7701 26375 7735
rect 26375 7701 26384 7735
rect 26332 7692 26384 7701
rect 26976 7692 27028 7744
rect 27528 7692 27580 7744
rect 32036 7692 32088 7744
rect 33600 7692 33652 7744
rect 38016 7828 38068 7880
rect 40684 7828 40736 7880
rect 39120 7692 39172 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 5724 7488 5776 7540
rect 9680 7488 9732 7540
rect 8024 7463 8076 7472
rect 8024 7429 8033 7463
rect 8033 7429 8067 7463
rect 8067 7429 8076 7463
rect 8024 7420 8076 7429
rect 8116 7420 8168 7472
rect 10140 7488 10192 7540
rect 15292 7488 15344 7540
rect 15844 7488 15896 7540
rect 16120 7488 16172 7540
rect 21272 7488 21324 7540
rect 21364 7488 21416 7540
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 8116 7284 8168 7336
rect 11796 7420 11848 7472
rect 14556 7420 14608 7472
rect 14832 7352 14884 7404
rect 15016 7352 15068 7404
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 15752 7395 15804 7404
rect 15752 7361 15761 7395
rect 15761 7361 15795 7395
rect 15795 7361 15804 7395
rect 15752 7352 15804 7361
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 14280 7216 14332 7268
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 17224 7352 17276 7404
rect 18328 7420 18380 7472
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 19248 7352 19300 7404
rect 20260 7352 20312 7404
rect 21088 7395 21140 7404
rect 21088 7361 21098 7395
rect 21098 7361 21132 7395
rect 21132 7361 21140 7395
rect 21088 7352 21140 7361
rect 21272 7395 21324 7404
rect 21272 7361 21281 7395
rect 21281 7361 21315 7395
rect 21315 7361 21324 7395
rect 21272 7352 21324 7361
rect 21364 7395 21416 7404
rect 21364 7361 21373 7395
rect 21373 7361 21407 7395
rect 21407 7361 21416 7395
rect 21364 7352 21416 7361
rect 21548 7352 21600 7404
rect 21824 7395 21876 7404
rect 21824 7361 21833 7395
rect 21833 7361 21867 7395
rect 21867 7361 21876 7395
rect 21824 7352 21876 7361
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 22652 7420 22704 7472
rect 24768 7420 24820 7472
rect 24952 7531 25004 7540
rect 24952 7497 24961 7531
rect 24961 7497 24995 7531
rect 24995 7497 25004 7531
rect 24952 7488 25004 7497
rect 25228 7488 25280 7540
rect 25596 7488 25648 7540
rect 26700 7488 26752 7540
rect 31760 7488 31812 7540
rect 33048 7488 33100 7540
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 9496 7148 9548 7157
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 15292 7148 15344 7200
rect 19064 7148 19116 7200
rect 19156 7191 19208 7200
rect 19156 7157 19165 7191
rect 19165 7157 19199 7191
rect 19199 7157 19208 7191
rect 19156 7148 19208 7157
rect 22468 7216 22520 7268
rect 24400 7352 24452 7404
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 25228 7395 25280 7404
rect 25228 7361 25237 7395
rect 25237 7361 25271 7395
rect 25271 7361 25280 7395
rect 25228 7352 25280 7361
rect 26332 7420 26384 7472
rect 40684 7488 40736 7540
rect 24952 7216 25004 7268
rect 25136 7216 25188 7268
rect 25688 7352 25740 7404
rect 25964 7352 26016 7404
rect 26240 7395 26292 7404
rect 26240 7361 26254 7395
rect 26254 7361 26288 7395
rect 26288 7361 26292 7395
rect 26240 7352 26292 7361
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 26608 7216 26660 7268
rect 38844 7420 38896 7472
rect 34612 7352 34664 7404
rect 29092 7284 29144 7336
rect 35440 7284 35492 7336
rect 35532 7284 35584 7336
rect 37280 7284 37332 7336
rect 39120 7327 39172 7336
rect 39120 7293 39129 7327
rect 39129 7293 39163 7327
rect 39163 7293 39172 7327
rect 39120 7284 39172 7293
rect 28540 7191 28592 7200
rect 28540 7157 28549 7191
rect 28549 7157 28583 7191
rect 28583 7157 28592 7191
rect 28540 7148 28592 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 5540 6987 5592 6996
rect 5540 6953 5570 6987
rect 5570 6953 5592 6987
rect 5540 6944 5592 6953
rect 7104 6944 7156 6996
rect 9036 6944 9088 6996
rect 13452 6944 13504 6996
rect 13544 6876 13596 6928
rect 4068 6808 4120 6860
rect 5080 6808 5132 6860
rect 7748 6740 7800 6792
rect 8852 6740 8904 6792
rect 12532 6808 12584 6860
rect 4712 6672 4764 6724
rect 6000 6672 6052 6724
rect 9956 6715 10008 6724
rect 9956 6681 9965 6715
rect 9965 6681 9999 6715
rect 9999 6681 10008 6715
rect 12164 6783 12216 6792
rect 12164 6749 12173 6783
rect 12173 6749 12207 6783
rect 12207 6749 12216 6783
rect 12164 6740 12216 6749
rect 15384 6808 15436 6860
rect 16028 6808 16080 6860
rect 16580 6808 16632 6860
rect 17040 6808 17092 6860
rect 9956 6672 10008 6681
rect 12440 6715 12492 6724
rect 12440 6681 12449 6715
rect 12449 6681 12483 6715
rect 12483 6681 12492 6715
rect 12440 6672 12492 6681
rect 13820 6672 13872 6724
rect 9588 6604 9640 6656
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 10968 6647 11020 6656
rect 10968 6613 10977 6647
rect 10977 6613 11011 6647
rect 11011 6613 11020 6647
rect 10968 6604 11020 6613
rect 11336 6647 11388 6656
rect 11336 6613 11345 6647
rect 11345 6613 11379 6647
rect 11379 6613 11388 6647
rect 11336 6604 11388 6613
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 15936 6740 15988 6792
rect 17684 6740 17736 6792
rect 19248 6944 19300 6996
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 20444 6876 20496 6928
rect 21272 6944 21324 6996
rect 21640 6944 21692 6996
rect 22560 6944 22612 6996
rect 22928 6944 22980 6996
rect 26608 6944 26660 6996
rect 27436 6944 27488 6996
rect 20168 6808 20220 6860
rect 19156 6672 19208 6724
rect 14924 6604 14976 6656
rect 15844 6604 15896 6656
rect 17868 6604 17920 6656
rect 18880 6647 18932 6656
rect 18880 6613 18889 6647
rect 18889 6613 18923 6647
rect 18923 6613 18932 6647
rect 18880 6604 18932 6613
rect 20444 6740 20496 6792
rect 21548 6808 21600 6860
rect 24400 6876 24452 6928
rect 26148 6876 26200 6928
rect 26332 6876 26384 6928
rect 21364 6647 21416 6656
rect 21364 6613 21373 6647
rect 21373 6613 21407 6647
rect 21407 6613 21416 6647
rect 21364 6604 21416 6613
rect 21640 6715 21692 6724
rect 21640 6681 21649 6715
rect 21649 6681 21683 6715
rect 21683 6681 21692 6715
rect 21640 6672 21692 6681
rect 21732 6715 21784 6724
rect 21732 6681 21741 6715
rect 21741 6681 21775 6715
rect 21775 6681 21784 6715
rect 21732 6672 21784 6681
rect 21824 6604 21876 6656
rect 22192 6808 22244 6860
rect 23388 6808 23440 6860
rect 25320 6851 25372 6860
rect 25320 6817 25329 6851
rect 25329 6817 25363 6851
rect 25363 6817 25372 6851
rect 25320 6808 25372 6817
rect 26700 6851 26752 6860
rect 26700 6817 26709 6851
rect 26709 6817 26743 6851
rect 26743 6817 26752 6851
rect 26700 6808 26752 6817
rect 27344 6808 27396 6860
rect 27436 6808 27488 6860
rect 24492 6783 24544 6792
rect 24492 6749 24501 6783
rect 24501 6749 24535 6783
rect 24535 6749 24544 6783
rect 24492 6740 24544 6749
rect 24860 6740 24912 6792
rect 25136 6783 25188 6792
rect 25136 6749 25145 6783
rect 25145 6749 25179 6783
rect 25179 6749 25188 6783
rect 25136 6740 25188 6749
rect 26608 6783 26660 6792
rect 26608 6749 26617 6783
rect 26617 6749 26651 6783
rect 26651 6749 26660 6783
rect 26608 6740 26660 6749
rect 27068 6783 27120 6792
rect 27068 6749 27077 6783
rect 27077 6749 27111 6783
rect 27111 6749 27120 6783
rect 27068 6740 27120 6749
rect 28632 6740 28684 6792
rect 29552 6808 29604 6860
rect 26148 6672 26200 6724
rect 24400 6604 24452 6656
rect 24676 6604 24728 6656
rect 26240 6647 26292 6656
rect 26240 6613 26249 6647
rect 26249 6613 26283 6647
rect 26283 6613 26292 6647
rect 26240 6604 26292 6613
rect 26976 6672 27028 6724
rect 28356 6672 28408 6724
rect 31116 6740 31168 6792
rect 36636 6783 36688 6792
rect 36636 6749 36645 6783
rect 36645 6749 36679 6783
rect 36679 6749 36688 6783
rect 36636 6740 36688 6749
rect 37280 6672 37332 6724
rect 29184 6647 29236 6656
rect 29184 6613 29193 6647
rect 29193 6613 29227 6647
rect 29227 6613 29236 6647
rect 29184 6604 29236 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4896 6443 4948 6452
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 4988 6332 5040 6384
rect 6460 6332 6512 6384
rect 8116 6400 8168 6452
rect 9772 6400 9824 6452
rect 11244 6400 11296 6452
rect 11336 6400 11388 6452
rect 12440 6400 12492 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 14096 6400 14148 6452
rect 6000 6264 6052 6316
rect 4988 6239 5040 6248
rect 4988 6205 4997 6239
rect 4997 6205 5031 6239
rect 5031 6205 5040 6239
rect 4988 6196 5040 6205
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 4988 6060 5040 6112
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 9588 6264 9640 6316
rect 11704 6239 11756 6248
rect 11704 6205 11713 6239
rect 11713 6205 11747 6239
rect 11747 6205 11756 6239
rect 11704 6196 11756 6205
rect 13728 6307 13780 6316
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 15844 6443 15896 6452
rect 15844 6409 15853 6443
rect 15853 6409 15887 6443
rect 15887 6409 15896 6443
rect 15844 6400 15896 6409
rect 15936 6443 15988 6452
rect 15936 6409 15945 6443
rect 15945 6409 15979 6443
rect 15979 6409 15988 6443
rect 15936 6400 15988 6409
rect 17960 6400 18012 6452
rect 18052 6264 18104 6316
rect 20168 6400 20220 6452
rect 21364 6400 21416 6452
rect 22376 6400 22428 6452
rect 26148 6400 26200 6452
rect 26240 6400 26292 6452
rect 26976 6443 27028 6452
rect 26976 6409 26985 6443
rect 26985 6409 27019 6443
rect 27019 6409 27028 6443
rect 26976 6400 27028 6409
rect 19984 6264 20036 6316
rect 21180 6264 21232 6316
rect 8392 6128 8444 6180
rect 13084 6128 13136 6180
rect 7748 6060 7800 6112
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 8944 6103 8996 6112
rect 8944 6069 8953 6103
rect 8953 6069 8987 6103
rect 8987 6069 8996 6103
rect 8944 6060 8996 6069
rect 12164 6060 12216 6112
rect 14188 6060 14240 6112
rect 15016 6060 15068 6112
rect 16028 6239 16080 6248
rect 16028 6205 16037 6239
rect 16037 6205 16071 6239
rect 16071 6205 16080 6239
rect 16028 6196 16080 6205
rect 17040 6239 17092 6248
rect 17040 6205 17049 6239
rect 17049 6205 17083 6239
rect 17083 6205 17092 6239
rect 17040 6196 17092 6205
rect 18880 6239 18932 6248
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 18604 6128 18656 6180
rect 21824 6128 21876 6180
rect 22100 6128 22152 6180
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 22560 6239 22612 6248
rect 22560 6205 22569 6239
rect 22569 6205 22603 6239
rect 22603 6205 22612 6239
rect 22560 6196 22612 6205
rect 24584 6264 24636 6316
rect 24676 6264 24728 6316
rect 28540 6400 28592 6452
rect 29092 6443 29144 6452
rect 29092 6409 29101 6443
rect 29101 6409 29135 6443
rect 29135 6409 29144 6443
rect 29092 6400 29144 6409
rect 29184 6400 29236 6452
rect 38844 6332 38896 6384
rect 28724 6264 28776 6316
rect 29276 6307 29328 6316
rect 29276 6273 29285 6307
rect 29285 6273 29319 6307
rect 29319 6273 29328 6307
rect 29276 6264 29328 6273
rect 24860 6239 24912 6248
rect 24860 6205 24869 6239
rect 24869 6205 24903 6239
rect 24903 6205 24912 6239
rect 24860 6196 24912 6205
rect 22928 6060 22980 6112
rect 23756 6060 23808 6112
rect 25504 6103 25556 6112
rect 25504 6069 25513 6103
rect 25513 6069 25547 6103
rect 25547 6069 25556 6103
rect 25504 6060 25556 6069
rect 26516 6060 26568 6112
rect 27068 6060 27120 6112
rect 28356 6196 28408 6248
rect 34612 6264 34664 6316
rect 37096 6307 37148 6316
rect 37096 6273 37105 6307
rect 37105 6273 37139 6307
rect 37139 6273 37148 6307
rect 37096 6264 37148 6273
rect 37280 6239 37332 6248
rect 37280 6205 37289 6239
rect 37289 6205 37323 6239
rect 37323 6205 37332 6239
rect 37280 6196 37332 6205
rect 40684 6196 40736 6248
rect 29276 6128 29328 6180
rect 31116 6060 31168 6112
rect 39764 6103 39816 6112
rect 39764 6069 39773 6103
rect 39773 6069 39807 6103
rect 39807 6069 39816 6103
rect 39764 6060 39816 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 7380 5856 7432 5908
rect 8944 5856 8996 5908
rect 10968 5856 11020 5908
rect 13176 5856 13228 5908
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 10600 5720 10652 5772
rect 16580 5856 16632 5908
rect 17040 5856 17092 5908
rect 11612 5652 11664 5704
rect 11796 5652 11848 5704
rect 5632 5584 5684 5636
rect 6000 5584 6052 5636
rect 13544 5720 13596 5772
rect 14188 5720 14240 5772
rect 15016 5720 15068 5772
rect 17868 5720 17920 5772
rect 20076 5720 20128 5772
rect 21180 5652 21232 5704
rect 21456 5856 21508 5908
rect 22560 5856 22612 5908
rect 37096 5856 37148 5908
rect 39764 5856 39816 5908
rect 13820 5584 13872 5636
rect 14556 5584 14608 5636
rect 6736 5516 6788 5568
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 13912 5516 13964 5568
rect 20168 5584 20220 5636
rect 29276 5788 29328 5840
rect 23112 5720 23164 5772
rect 17960 5516 18012 5568
rect 22284 5559 22336 5568
rect 22284 5525 22293 5559
rect 22293 5525 22327 5559
rect 22327 5525 22336 5559
rect 22284 5516 22336 5525
rect 23756 5516 23808 5568
rect 23848 5559 23900 5568
rect 23848 5525 23857 5559
rect 23857 5525 23891 5559
rect 23891 5525 23900 5559
rect 23848 5516 23900 5525
rect 24584 5720 24636 5772
rect 25780 5720 25832 5772
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 30472 5720 30524 5772
rect 31300 5763 31352 5772
rect 31300 5729 31309 5763
rect 31309 5729 31343 5763
rect 31343 5729 31352 5763
rect 31300 5720 31352 5729
rect 32864 5788 32916 5840
rect 25504 5652 25556 5704
rect 28816 5652 28868 5704
rect 33048 5720 33100 5772
rect 25044 5584 25096 5636
rect 31760 5584 31812 5636
rect 31852 5627 31904 5636
rect 31852 5593 31861 5627
rect 31861 5593 31895 5627
rect 31895 5593 31904 5627
rect 31852 5584 31904 5593
rect 34796 5720 34848 5772
rect 34704 5652 34756 5704
rect 35624 5720 35676 5772
rect 37832 5720 37884 5772
rect 34520 5516 34572 5568
rect 36268 5652 36320 5704
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3884 5312 3936 5364
rect 5632 5355 5684 5364
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 6000 5244 6052 5296
rect 5080 5176 5132 5228
rect 8392 5312 8444 5364
rect 12716 5312 12768 5364
rect 13912 5355 13964 5364
rect 13912 5321 13921 5355
rect 13921 5321 13955 5355
rect 13955 5321 13964 5355
rect 13912 5312 13964 5321
rect 17316 5312 17368 5364
rect 20168 5312 20220 5364
rect 20536 5312 20588 5364
rect 22284 5312 22336 5364
rect 6460 5244 6512 5296
rect 13820 5244 13872 5296
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 5540 4972 5592 5024
rect 6736 4972 6788 5024
rect 12164 5219 12216 5228
rect 12164 5185 12173 5219
rect 12173 5185 12207 5219
rect 12207 5185 12216 5219
rect 12164 5176 12216 5185
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 20904 5176 20956 5228
rect 23112 5244 23164 5296
rect 23848 5312 23900 5364
rect 24676 5244 24728 5296
rect 24952 5312 25004 5364
rect 25136 5312 25188 5364
rect 27712 5312 27764 5364
rect 31852 5312 31904 5364
rect 22928 5219 22980 5228
rect 22928 5185 22937 5219
rect 22937 5185 22971 5219
rect 22971 5185 22980 5219
rect 22928 5176 22980 5185
rect 24952 5219 25004 5228
rect 24952 5185 24961 5219
rect 24961 5185 24995 5219
rect 24995 5185 25004 5219
rect 24952 5176 25004 5185
rect 26608 5176 26660 5228
rect 28356 5176 28408 5228
rect 31760 5176 31812 5228
rect 34520 5312 34572 5364
rect 34612 5312 34664 5364
rect 38844 5244 38896 5296
rect 23296 5108 23348 5160
rect 24860 5108 24912 5160
rect 25320 5108 25372 5160
rect 26516 5108 26568 5160
rect 21364 5040 21416 5092
rect 21916 5040 21968 5092
rect 11336 4972 11388 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 36268 5015 36320 5024
rect 36268 4981 36277 5015
rect 36277 4981 36311 5015
rect 36311 4981 36320 5015
rect 36268 4972 36320 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 11520 4768 11572 4820
rect 12440 4768 12492 4820
rect 18328 4811 18380 4820
rect 18328 4777 18337 4811
rect 18337 4777 18371 4811
rect 18371 4777 18380 4811
rect 18328 4768 18380 4777
rect 24952 4768 25004 4820
rect 26516 4768 26568 4820
rect 28080 4768 28132 4820
rect 36268 4768 36320 4820
rect 11336 4700 11388 4752
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 12164 4632 12216 4684
rect 26240 4700 26292 4752
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 21732 4632 21784 4684
rect 22008 4632 22060 4684
rect 25044 4632 25096 4684
rect 11612 4564 11664 4616
rect 13084 4564 13136 4616
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 17960 4564 18012 4616
rect 19064 4564 19116 4616
rect 20996 4564 21048 4616
rect 25136 4607 25188 4616
rect 25136 4573 25145 4607
rect 25145 4573 25179 4607
rect 25179 4573 25188 4607
rect 25136 4564 25188 4573
rect 25964 4632 26016 4684
rect 26332 4632 26384 4684
rect 37464 4700 37516 4752
rect 37740 4632 37792 4684
rect 37832 4632 37884 4684
rect 28356 4564 28408 4616
rect 16856 4539 16908 4548
rect 16856 4505 16865 4539
rect 16865 4505 16899 4539
rect 16899 4505 16908 4539
rect 16856 4496 16908 4505
rect 18420 4428 18472 4480
rect 20352 4471 20404 4480
rect 20352 4437 20361 4471
rect 20361 4437 20395 4471
rect 20395 4437 20404 4471
rect 20352 4428 20404 4437
rect 26700 4539 26752 4548
rect 26700 4505 26709 4539
rect 26709 4505 26743 4539
rect 26743 4505 26752 4539
rect 26700 4496 26752 4505
rect 28080 4496 28132 4548
rect 39028 4564 39080 4616
rect 41052 4428 41104 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 14188 4224 14240 4276
rect 15016 4224 15068 4276
rect 15568 4267 15620 4276
rect 15568 4233 15577 4267
rect 15577 4233 15611 4267
rect 15611 4233 15620 4267
rect 15568 4224 15620 4233
rect 16488 4224 16540 4276
rect 16764 4224 16816 4276
rect 16856 4224 16908 4276
rect 17316 4267 17368 4276
rect 17316 4233 17325 4267
rect 17325 4233 17359 4267
rect 17359 4233 17368 4267
rect 17316 4224 17368 4233
rect 18420 4224 18472 4276
rect 13728 4088 13780 4140
rect 14556 4156 14608 4208
rect 16580 4156 16632 4208
rect 18696 4224 18748 4276
rect 21088 4224 21140 4276
rect 21364 4267 21416 4276
rect 21364 4233 21373 4267
rect 21373 4233 21407 4267
rect 21407 4233 21416 4267
rect 21364 4224 21416 4233
rect 22100 4224 22152 4276
rect 24032 4224 24084 4276
rect 26240 4224 26292 4276
rect 26700 4224 26752 4276
rect 19064 4156 19116 4208
rect 14096 4063 14148 4072
rect 14096 4029 14105 4063
rect 14105 4029 14139 4063
rect 14139 4029 14148 4063
rect 14096 4020 14148 4029
rect 16948 4131 17000 4140
rect 16948 4097 16957 4131
rect 16957 4097 16991 4131
rect 16991 4097 17000 4131
rect 16948 4088 17000 4097
rect 17316 4088 17368 4140
rect 17684 4088 17736 4140
rect 18328 4131 18380 4140
rect 18328 4097 18337 4131
rect 18337 4097 18371 4131
rect 18371 4097 18380 4131
rect 18328 4088 18380 4097
rect 20076 4020 20128 4072
rect 15108 3884 15160 3936
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16764 3927 16816 3936
rect 16764 3893 16773 3927
rect 16773 3893 16807 3927
rect 16807 3893 16816 3927
rect 16764 3884 16816 3893
rect 18420 3884 18472 3936
rect 20444 4088 20496 4140
rect 22836 4088 22888 4140
rect 24124 4131 24176 4140
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 24124 4088 24176 4097
rect 25228 4088 25280 4140
rect 25688 4088 25740 4140
rect 37464 4156 37516 4208
rect 38844 4156 38896 4208
rect 37280 4131 37332 4140
rect 37280 4097 37289 4131
rect 37289 4097 37323 4131
rect 37323 4097 37332 4131
rect 37280 4088 37332 4097
rect 24676 4020 24728 4072
rect 22008 3952 22060 4004
rect 25596 3952 25648 4004
rect 26608 3952 26660 4004
rect 20812 3927 20864 3936
rect 20812 3893 20821 3927
rect 20821 3893 20855 3927
rect 20855 3893 20864 3927
rect 20812 3884 20864 3893
rect 20904 3927 20956 3936
rect 20904 3893 20913 3927
rect 20913 3893 20947 3927
rect 20947 3893 20956 3927
rect 20904 3884 20956 3893
rect 21824 3927 21876 3936
rect 21824 3893 21833 3927
rect 21833 3893 21867 3927
rect 21867 3893 21876 3927
rect 21824 3884 21876 3893
rect 23848 3884 23900 3936
rect 24768 3884 24820 3936
rect 39028 3927 39080 3936
rect 39028 3893 39037 3927
rect 39037 3893 39071 3927
rect 39071 3893 39080 3927
rect 39028 3884 39080 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 13544 3680 13596 3732
rect 14096 3680 14148 3732
rect 14556 3680 14608 3732
rect 15476 3680 15528 3732
rect 15660 3680 15712 3732
rect 16948 3680 17000 3732
rect 17684 3680 17736 3732
rect 15108 3612 15160 3664
rect 5540 3476 5592 3528
rect 940 3340 992 3392
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 14372 3340 14424 3392
rect 14832 3476 14884 3528
rect 15016 3408 15068 3460
rect 17684 3544 17736 3596
rect 17776 3587 17828 3596
rect 17776 3553 17785 3587
rect 17785 3553 17819 3587
rect 17819 3553 17828 3587
rect 17776 3544 17828 3553
rect 17868 3587 17920 3596
rect 17868 3553 17877 3587
rect 17877 3553 17911 3587
rect 17911 3553 17920 3587
rect 17868 3544 17920 3553
rect 18696 3680 18748 3732
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 15292 3383 15344 3392
rect 15292 3349 15301 3383
rect 15301 3349 15335 3383
rect 15335 3349 15344 3383
rect 15292 3340 15344 3349
rect 16580 3451 16632 3460
rect 16580 3417 16589 3451
rect 16589 3417 16623 3451
rect 16623 3417 16632 3451
rect 16580 3408 16632 3417
rect 20812 3680 20864 3732
rect 21088 3680 21140 3732
rect 20076 3544 20128 3596
rect 24032 3723 24084 3732
rect 24032 3689 24041 3723
rect 24041 3689 24075 3723
rect 24075 3689 24084 3723
rect 24032 3680 24084 3689
rect 24124 3680 24176 3732
rect 24768 3680 24820 3732
rect 25320 3680 25372 3732
rect 26056 3680 26108 3732
rect 23296 3544 23348 3596
rect 24584 3544 24636 3596
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 20168 3383 20220 3392
rect 20168 3349 20177 3383
rect 20177 3349 20211 3383
rect 20211 3349 20220 3383
rect 20168 3340 20220 3349
rect 20720 3451 20772 3460
rect 20720 3417 20729 3451
rect 20729 3417 20763 3451
rect 20763 3417 20772 3451
rect 20720 3408 20772 3417
rect 20996 3408 21048 3460
rect 22560 3451 22612 3460
rect 22560 3417 22569 3451
rect 22569 3417 22603 3451
rect 22603 3417 22612 3451
rect 22560 3408 22612 3417
rect 24676 3476 24728 3528
rect 24584 3408 24636 3460
rect 25596 3544 25648 3596
rect 26608 3476 26660 3528
rect 24860 3383 24912 3392
rect 24860 3349 24869 3383
rect 24869 3349 24903 3383
rect 24903 3349 24912 3383
rect 24860 3340 24912 3349
rect 25872 3340 25924 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 13728 3136 13780 3188
rect 12900 3068 12952 3120
rect 14372 3068 14424 3120
rect 13728 2932 13780 2984
rect 16580 3136 16632 3188
rect 15292 3068 15344 3120
rect 15476 3068 15528 3120
rect 16764 3136 16816 3188
rect 20076 3136 20128 3188
rect 21272 3179 21324 3188
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 21824 3136 21876 3188
rect 17960 3068 18012 3120
rect 21180 3068 21232 3120
rect 22560 3136 22612 3188
rect 25228 3179 25280 3188
rect 25228 3145 25237 3179
rect 25237 3145 25271 3179
rect 25271 3145 25280 3179
rect 25228 3136 25280 3145
rect 25688 3179 25740 3188
rect 25688 3145 25697 3179
rect 25697 3145 25731 3179
rect 25731 3145 25740 3179
rect 25688 3136 25740 3145
rect 25964 3136 26016 3188
rect 26056 3179 26108 3188
rect 26056 3145 26065 3179
rect 26065 3145 26099 3179
rect 26099 3145 26108 3179
rect 26056 3136 26108 3145
rect 23848 3068 23900 3120
rect 24768 3068 24820 3120
rect 23296 3000 23348 3052
rect 14556 2864 14608 2916
rect 16488 2907 16540 2916
rect 16488 2873 16497 2907
rect 16497 2873 16531 2907
rect 16531 2873 16540 2907
rect 16488 2864 16540 2873
rect 14832 2796 14884 2848
rect 17684 2796 17736 2848
rect 20168 2932 20220 2984
rect 25320 3000 25372 3052
rect 27528 2932 27580 2984
rect 24860 2796 24912 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 14280 2592 14332 2644
rect 20720 2592 20772 2644
rect 11980 2456 12032 2508
rect 8852 2388 8904 2440
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 17684 2388 17736 2440
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 20812 2388 20864 2440
rect 31116 2431 31168 2440
rect 31116 2397 31125 2431
rect 31125 2397 31159 2431
rect 31159 2397 31168 2431
rect 31116 2388 31168 2397
rect 34612 2388 34664 2440
rect 39028 2388 39080 2440
rect 40684 2431 40736 2440
rect 40684 2397 40693 2431
rect 40693 2397 40727 2431
rect 40727 2397 40736 2431
rect 40684 2388 40736 2397
rect 20 2320 72 2372
rect 4988 2320 5040 2372
rect 20628 2320 20680 2372
rect 3976 2252 4028 2304
rect 7748 2252 7800 2304
rect 11612 2252 11664 2304
rect 15476 2252 15528 2304
rect 19340 2252 19392 2304
rect 23296 2252 23348 2304
rect 27068 2252 27120 2304
rect 30932 2252 30984 2304
rect 34796 2252 34848 2304
rect 38660 2252 38712 2304
rect 39948 2252 40000 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 2778 44296 2834 44305
rect 2778 44231 2834 44240
rect 2792 42294 2820 44231
rect 3238 43864 3294 44664
rect 7102 43864 7158 44664
rect 10966 43864 11022 44664
rect 14830 43864 14886 44664
rect 18694 43864 18750 44664
rect 22558 43864 22614 44664
rect 26422 43864 26478 44664
rect 30286 43864 30342 44664
rect 34150 44010 34206 44664
rect 38014 44010 38070 44664
rect 34150 43982 34468 44010
rect 34150 43864 34206 43982
rect 2780 42288 2832 42294
rect 2780 42230 2832 42236
rect 3252 42226 3280 43864
rect 7116 42294 7144 43864
rect 10876 42560 10928 42566
rect 10876 42502 10928 42508
rect 7104 42288 7156 42294
rect 7104 42230 7156 42236
rect 1492 42220 1544 42226
rect 1492 42162 1544 42168
rect 3240 42220 3292 42226
rect 3240 42162 3292 42168
rect 940 40520 992 40526
rect 940 40462 992 40468
rect 952 40225 980 40462
rect 938 40216 994 40225
rect 938 40151 994 40160
rect 938 36136 994 36145
rect 938 36071 994 36080
rect 952 36038 980 36071
rect 940 36032 992 36038
rect 940 35974 992 35980
rect 940 32224 992 32230
rect 940 32166 992 32172
rect 952 32065 980 32166
rect 938 32056 994 32065
rect 938 31991 994 32000
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 938 27976 994 27985
rect 938 27911 940 27920
rect 992 27911 994 27920
rect 940 27882 992 27888
rect 940 24064 992 24070
rect 940 24006 992 24012
rect 952 23905 980 24006
rect 938 23896 994 23905
rect 938 23831 994 23840
rect 1412 23322 1440 28018
rect 1400 23316 1452 23322
rect 1400 23258 1452 23264
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 938 19816 994 19825
rect 938 19751 940 19760
rect 992 19751 994 19760
rect 940 19722 992 19728
rect 1412 18290 1440 21422
rect 1504 18426 1532 42162
rect 10888 42090 10916 42502
rect 10980 42378 11008 43864
rect 14556 42560 14608 42566
rect 14556 42502 14608 42508
rect 10980 42362 11100 42378
rect 10980 42356 11112 42362
rect 10980 42350 11060 42356
rect 11060 42298 11112 42304
rect 10876 42084 10928 42090
rect 10876 42026 10928 42032
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 7196 41540 7248 41546
rect 7196 41482 7248 41488
rect 7208 41414 7236 41482
rect 10600 41472 10652 41478
rect 10888 41449 10916 42026
rect 14004 42016 14056 42022
rect 14004 41958 14056 41964
rect 14016 41750 14044 41958
rect 14568 41818 14596 42502
rect 14844 42226 14872 43864
rect 18708 42362 18736 43864
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 18696 42356 18748 42362
rect 18696 42298 18748 42304
rect 22572 42226 22600 43864
rect 14648 42220 14700 42226
rect 14648 42162 14700 42168
rect 14832 42220 14884 42226
rect 14832 42162 14884 42168
rect 16028 42220 16080 42226
rect 16028 42162 16080 42168
rect 22560 42220 22612 42226
rect 22560 42162 22612 42168
rect 14660 41857 14688 42162
rect 16040 42090 16068 42162
rect 16028 42084 16080 42090
rect 16028 42026 16080 42032
rect 23480 42084 23532 42090
rect 23480 42026 23532 42032
rect 24400 42084 24452 42090
rect 24400 42026 24452 42032
rect 20720 42016 20772 42022
rect 20720 41958 20772 41964
rect 14646 41848 14702 41857
rect 14556 41812 14608 41818
rect 19430 41848 19486 41857
rect 14646 41783 14702 41792
rect 17776 41812 17828 41818
rect 14556 41754 14608 41760
rect 19430 41783 19486 41792
rect 17776 41754 17828 41760
rect 14004 41744 14056 41750
rect 14004 41686 14056 41692
rect 11060 41676 11112 41682
rect 11060 41618 11112 41624
rect 12716 41676 12768 41682
rect 12716 41618 12768 41624
rect 10600 41414 10652 41420
rect 10874 41440 10930 41449
rect 7208 41386 7328 41414
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 1676 40520 1728 40526
rect 1676 40462 1728 40468
rect 1688 26382 1716 40462
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 6920 38888 6972 38894
rect 6920 38830 6972 38836
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 6932 37806 6960 38830
rect 6920 37800 6972 37806
rect 6920 37742 6972 37748
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 6828 36236 6880 36242
rect 6932 36224 6960 37742
rect 6880 36196 6960 36224
rect 6828 36178 6880 36184
rect 6000 36168 6052 36174
rect 6000 36110 6052 36116
rect 4804 36100 4856 36106
rect 4804 36042 4856 36048
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4620 32224 4672 32230
rect 4620 32166 4672 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 31278 4660 32166
rect 4816 31754 4844 36042
rect 6012 35630 6040 36110
rect 7104 36032 7156 36038
rect 7104 35974 7156 35980
rect 7116 35766 7144 35974
rect 7104 35760 7156 35766
rect 7104 35702 7156 35708
rect 6000 35624 6052 35630
rect 6000 35566 6052 35572
rect 6736 35624 6788 35630
rect 6736 35566 6788 35572
rect 5540 34672 5592 34678
rect 4724 31726 4844 31754
rect 5368 34620 5540 34626
rect 5368 34614 5592 34620
rect 5368 34598 5580 34614
rect 4620 31272 4672 31278
rect 4620 31214 4672 31220
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4528 30796 4580 30802
rect 4632 30784 4660 31214
rect 4580 30756 4660 30784
rect 4528 30738 4580 30744
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3792 29096 3844 29102
rect 3792 29038 3844 29044
rect 3804 28014 3832 29038
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3792 28008 3844 28014
rect 3792 27950 3844 27956
rect 3804 27470 3832 27950
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 3804 25838 3832 27406
rect 4068 27396 4120 27402
rect 4068 27338 4120 27344
rect 4080 27130 4108 27338
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3792 25832 3844 25838
rect 3792 25774 3844 25780
rect 3804 25362 3832 25774
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4724 25498 4752 31726
rect 5264 29572 5316 29578
rect 5264 29514 5316 29520
rect 5276 28762 5304 29514
rect 5264 28756 5316 28762
rect 5264 28698 5316 28704
rect 5368 28082 5396 34598
rect 6012 34542 6040 35566
rect 6748 35290 6776 35566
rect 6736 35284 6788 35290
rect 6736 35226 6788 35232
rect 6826 34776 6882 34785
rect 6826 34711 6882 34720
rect 6840 34678 6868 34711
rect 6828 34672 6880 34678
rect 6828 34614 6880 34620
rect 6000 34536 6052 34542
rect 6000 34478 6052 34484
rect 6012 33454 6040 34478
rect 7116 33590 7144 35702
rect 7104 33584 7156 33590
rect 7104 33526 7156 33532
rect 6000 33448 6052 33454
rect 6000 33390 6052 33396
rect 6736 33448 6788 33454
rect 6736 33390 6788 33396
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 5632 32564 5684 32570
rect 5632 32506 5684 32512
rect 5448 30728 5500 30734
rect 5448 30670 5500 30676
rect 5460 29170 5488 30670
rect 5448 29164 5500 29170
rect 5448 29106 5500 29112
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 4712 25492 4764 25498
rect 4712 25434 4764 25440
rect 3792 25356 3844 25362
rect 3792 25298 3844 25304
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 4080 24954 4108 25162
rect 4724 24954 4752 25434
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4724 24138 4752 24686
rect 4712 24132 4764 24138
rect 4712 24074 4764 24080
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1872 22234 1900 23054
rect 1860 22228 1912 22234
rect 1860 22170 1912 22176
rect 4080 22098 4108 23598
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 23734
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22092 4120 22098
rect 4816 22094 4844 28018
rect 5172 27872 5224 27878
rect 5172 27814 5224 27820
rect 5184 26926 5212 27814
rect 5460 27470 5488 29106
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5552 28014 5580 28494
rect 5540 28008 5592 28014
rect 5540 27950 5592 27956
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 4988 26920 5040 26926
rect 4988 26862 5040 26868
rect 5172 26920 5224 26926
rect 5172 26862 5224 26868
rect 5000 26353 5028 26862
rect 4986 26344 5042 26353
rect 4986 26279 5042 26288
rect 5080 26240 5132 26246
rect 5080 26182 5132 26188
rect 5092 26042 5120 26182
rect 5080 26036 5132 26042
rect 5080 25978 5132 25984
rect 5460 25974 5488 27406
rect 5552 26994 5580 27950
rect 5644 27674 5672 32506
rect 5920 32026 5948 32846
rect 6012 32230 6040 33390
rect 6748 33114 6776 33390
rect 6736 33108 6788 33114
rect 6736 33050 6788 33056
rect 6092 32904 6144 32910
rect 6090 32872 6092 32881
rect 6276 32904 6328 32910
rect 6144 32872 6146 32881
rect 6276 32846 6328 32852
rect 6090 32807 6146 32816
rect 6000 32224 6052 32230
rect 6000 32166 6052 32172
rect 5908 32020 5960 32026
rect 5908 31962 5960 31968
rect 5722 31920 5778 31929
rect 5722 31855 5778 31864
rect 5736 31822 5764 31855
rect 5724 31816 5776 31822
rect 5724 31758 5776 31764
rect 6000 31816 6052 31822
rect 6000 31758 6052 31764
rect 5736 29646 5764 31758
rect 5816 31748 5868 31754
rect 5816 31690 5868 31696
rect 5828 31346 5856 31690
rect 6012 31346 6040 31758
rect 6104 31346 6132 32807
rect 6288 32570 6316 32846
rect 6460 32836 6512 32842
rect 6460 32778 6512 32784
rect 6472 32570 6500 32778
rect 6276 32564 6328 32570
rect 6276 32506 6328 32512
rect 6460 32564 6512 32570
rect 6460 32506 6512 32512
rect 7116 32502 7144 33526
rect 7104 32496 7156 32502
rect 7104 32438 7156 32444
rect 6368 32428 6420 32434
rect 6368 32370 6420 32376
rect 6184 32360 6236 32366
rect 6184 32302 6236 32308
rect 6196 32026 6224 32302
rect 6184 32020 6236 32026
rect 6184 31962 6236 31968
rect 6380 31754 6408 32370
rect 7300 31754 7328 41386
rect 10612 41138 10640 41414
rect 10874 41375 10930 41384
rect 11072 41274 11100 41618
rect 11428 41608 11480 41614
rect 11428 41550 11480 41556
rect 11440 41274 11468 41550
rect 12440 41540 12492 41546
rect 12440 41482 12492 41488
rect 11060 41268 11112 41274
rect 11060 41210 11112 41216
rect 11428 41268 11480 41274
rect 11428 41210 11480 41216
rect 10600 41132 10652 41138
rect 10600 41074 10652 41080
rect 10876 41132 10928 41138
rect 10876 41074 10928 41080
rect 9496 41064 9548 41070
rect 9496 41006 9548 41012
rect 9508 40730 9536 41006
rect 10232 40928 10284 40934
rect 10232 40870 10284 40876
rect 9496 40724 9548 40730
rect 9496 40666 9548 40672
rect 10244 40526 10272 40870
rect 10232 40520 10284 40526
rect 10232 40462 10284 40468
rect 10416 40520 10468 40526
rect 10416 40462 10468 40468
rect 8484 40044 8536 40050
rect 8484 39986 8536 39992
rect 9588 40044 9640 40050
rect 9588 39986 9640 39992
rect 8300 39840 8352 39846
rect 8300 39782 8352 39788
rect 8312 39098 8340 39782
rect 8496 39642 8524 39986
rect 9220 39840 9272 39846
rect 9220 39782 9272 39788
rect 9312 39840 9364 39846
rect 9312 39782 9364 39788
rect 8484 39636 8536 39642
rect 8484 39578 8536 39584
rect 9232 39574 9260 39782
rect 9220 39568 9272 39574
rect 9220 39510 9272 39516
rect 8300 39092 8352 39098
rect 8300 39034 8352 39040
rect 9036 38820 9088 38826
rect 9036 38762 9088 38768
rect 9048 37942 9076 38762
rect 9036 37936 9088 37942
rect 8772 37896 9036 37924
rect 7564 37800 7616 37806
rect 7564 37742 7616 37748
rect 8576 37800 8628 37806
rect 8576 37742 8628 37748
rect 7576 37466 7604 37742
rect 7564 37460 7616 37466
rect 7564 37402 7616 37408
rect 8588 36854 8616 37742
rect 8668 37256 8720 37262
rect 8668 37198 8720 37204
rect 8680 36922 8708 37198
rect 8668 36916 8720 36922
rect 8668 36858 8720 36864
rect 8576 36848 8628 36854
rect 8576 36790 8628 36796
rect 8024 35556 8076 35562
rect 8024 35498 8076 35504
rect 8036 35290 8064 35498
rect 8024 35284 8076 35290
rect 8024 35226 8076 35232
rect 8680 35222 8708 36858
rect 8772 36854 8800 37896
rect 9036 37878 9088 37884
rect 9036 37664 9088 37670
rect 9036 37606 9088 37612
rect 9048 37262 9076 37606
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 8760 36848 8812 36854
rect 8760 36790 8812 36796
rect 8772 36174 8800 36790
rect 8760 36168 8812 36174
rect 8760 36110 8812 36116
rect 8852 36100 8904 36106
rect 8852 36042 8904 36048
rect 8668 35216 8720 35222
rect 8668 35158 8720 35164
rect 8668 35080 8720 35086
rect 8668 35022 8720 35028
rect 7378 34640 7434 34649
rect 7378 34575 7434 34584
rect 6380 31726 6500 31754
rect 6380 31686 6408 31726
rect 6368 31680 6420 31686
rect 6368 31622 6420 31628
rect 5816 31340 5868 31346
rect 5816 31282 5868 31288
rect 5908 31340 5960 31346
rect 5908 31282 5960 31288
rect 6000 31340 6052 31346
rect 6000 31282 6052 31288
rect 6092 31340 6144 31346
rect 6092 31282 6144 31288
rect 5724 29640 5776 29646
rect 5724 29582 5776 29588
rect 5736 29238 5764 29582
rect 5724 29232 5776 29238
rect 5724 29174 5776 29180
rect 5920 28422 5948 31282
rect 6012 30784 6040 31282
rect 6472 31142 6500 31726
rect 7208 31726 7328 31754
rect 6460 31136 6512 31142
rect 6460 31078 6512 31084
rect 6184 30796 6236 30802
rect 6012 30756 6184 30784
rect 6104 29646 6132 30756
rect 6184 30738 6236 30744
rect 6472 30734 6500 31078
rect 7208 30734 7236 31726
rect 7288 31408 7340 31414
rect 7288 31350 7340 31356
rect 7300 30938 7328 31350
rect 7288 30932 7340 30938
rect 7288 30874 7340 30880
rect 6276 30728 6328 30734
rect 6276 30670 6328 30676
rect 6460 30728 6512 30734
rect 6460 30670 6512 30676
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 6184 30660 6236 30666
rect 6184 30602 6236 30608
rect 6196 29646 6224 30602
rect 6092 29640 6144 29646
rect 6092 29582 6144 29588
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 6000 29504 6052 29510
rect 6000 29446 6052 29452
rect 6012 29034 6040 29446
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 6000 28620 6052 28626
rect 6104 28608 6132 29582
rect 6052 28580 6132 28608
rect 6000 28562 6052 28568
rect 5908 28416 5960 28422
rect 5908 28358 5960 28364
rect 5632 27668 5684 27674
rect 5632 27610 5684 27616
rect 6104 27606 6132 28580
rect 6184 28484 6236 28490
rect 6184 28426 6236 28432
rect 6092 27600 6144 27606
rect 6092 27542 6144 27548
rect 6196 27538 6224 28426
rect 6184 27532 6236 27538
rect 6184 27474 6236 27480
rect 6288 27470 6316 30670
rect 6472 29646 6500 30670
rect 6460 29640 6512 29646
rect 6460 29582 6512 29588
rect 6472 27470 6500 29582
rect 7300 28558 7328 30874
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 6736 27600 6788 27606
rect 6736 27542 6788 27548
rect 6748 27470 6776 27542
rect 6276 27464 6328 27470
rect 6276 27406 6328 27412
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 6288 27130 6316 27270
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 6748 26450 6776 27406
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6840 26586 6868 27338
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6932 27130 6960 27270
rect 6920 27124 6972 27130
rect 6920 27066 6972 27072
rect 7300 27062 7328 28494
rect 7288 27056 7340 27062
rect 7288 26998 7340 27004
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6920 26308 6972 26314
rect 6920 26250 6972 26256
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 5448 25968 5500 25974
rect 5448 25910 5500 25916
rect 5460 25294 5488 25910
rect 6564 25838 6592 26182
rect 6932 26042 6960 26250
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 6552 25832 6604 25838
rect 6552 25774 6604 25780
rect 6564 25498 6592 25774
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7300 25498 7328 25638
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 6826 25392 6882 25401
rect 6826 25327 6882 25336
rect 6840 25294 6868 25327
rect 5448 25288 5500 25294
rect 6828 25288 6880 25294
rect 5500 25236 5580 25242
rect 5448 25230 5580 25236
rect 6828 25230 6880 25236
rect 5460 25214 5580 25230
rect 4896 24744 4948 24750
rect 4896 24686 4948 24692
rect 4908 24410 4936 24686
rect 4896 24404 4948 24410
rect 4948 24364 5120 24392
rect 4896 24346 4948 24352
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4068 22034 4120 22040
rect 4724 22066 4844 22094
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 4724 21978 4752 22066
rect 2240 21486 2268 21966
rect 4528 21956 4580 21962
rect 4724 21950 4844 21978
rect 4528 21898 4580 21904
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 2976 21486 3004 21830
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 2228 21480 2280 21486
rect 2228 21422 2280 21428
rect 2964 21480 3016 21486
rect 2964 21422 3016 21428
rect 1674 19816 1730 19825
rect 1674 19751 1676 19760
rect 1728 19751 1730 19760
rect 1676 19722 1728 19728
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 3896 18834 3924 19110
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 1492 18420 1544 18426
rect 1492 18362 1544 18368
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1504 17746 1532 18362
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 17882 1716 18158
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1492 17740 1544 17746
rect 1492 17682 1544 17688
rect 2884 17734 3004 17762
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 952 15745 980 15846
rect 938 15736 994 15745
rect 1412 15706 1440 16050
rect 938 15671 994 15680
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2700 13870 2728 15506
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2884 12238 2912 17734
rect 2976 17678 3004 17734
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 3068 15502 3096 18294
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3068 14006 3096 15438
rect 3436 14618 3464 16934
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3804 16114 3832 16526
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 14074 3648 14214
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3712 12306 3740 13806
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2240 11830 2268 12038
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 952 11354 980 11591
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 940 11348 992 11354
rect 940 11290 992 11296
rect 1504 11150 1532 11494
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 2884 11082 2912 12174
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2976 11558 3004 12106
rect 3712 11762 3740 12242
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 3068 11354 3096 11698
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 3896 8634 3924 18566
rect 4080 18426 4108 21490
rect 4448 21332 4476 21830
rect 4540 21593 4568 21898
rect 4526 21584 4582 21593
rect 4816 21554 4844 21950
rect 4526 21519 4528 21528
rect 4580 21519 4582 21528
rect 4804 21548 4856 21554
rect 4528 21490 4580 21496
rect 4804 21490 4856 21496
rect 4908 21486 4936 22510
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4448 21304 4660 21332
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21146 4660 21304
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4724 19378 4752 19654
rect 4816 19446 4844 19790
rect 4908 19514 4936 20266
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 5000 19514 5028 19654
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4344 19304 4396 19310
rect 4528 19304 4580 19310
rect 4396 19252 4528 19258
rect 4632 19281 4660 19314
rect 4344 19246 4580 19252
rect 4618 19272 4674 19281
rect 4356 19230 4568 19246
rect 4618 19207 4674 19216
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4540 18834 4568 18906
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4344 18760 4396 18766
rect 4342 18728 4344 18737
rect 4396 18728 4398 18737
rect 4342 18663 4398 18672
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4540 18086 4568 18770
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 4080 16590 4108 17750
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16590 4660 19110
rect 4816 18714 4844 19110
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4724 18686 4844 18714
rect 4724 17678 4752 18686
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4724 16658 4752 17614
rect 4816 17218 4844 18022
rect 4908 17338 4936 18770
rect 5000 18630 5028 19450
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18426 5028 18566
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4816 17190 4936 17218
rect 4908 17134 4936 17190
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4080 16096 4108 16526
rect 4356 16250 4384 16526
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4160 16108 4212 16114
rect 4080 16068 4160 16096
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3988 10810 4016 15438
rect 4080 14414 4108 16068
rect 4160 16050 4212 16056
rect 4540 16046 4568 16390
rect 4632 16114 4660 16526
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4908 15978 4936 17070
rect 5000 16590 5028 18226
rect 5092 17354 5120 24364
rect 5552 23866 5580 25214
rect 6368 25152 6420 25158
rect 6368 25094 6420 25100
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6104 23866 6132 24142
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5552 22234 5580 22578
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 5368 21622 5396 22034
rect 5552 21894 5580 22170
rect 5736 22094 5764 22374
rect 5644 22066 5764 22094
rect 6380 22094 6408 25094
rect 7392 24342 7420 34575
rect 7932 34128 7984 34134
rect 7932 34070 7984 34076
rect 7656 32972 7708 32978
rect 7656 32914 7708 32920
rect 7668 31482 7696 32914
rect 7944 32858 7972 34070
rect 8208 33924 8260 33930
rect 8208 33866 8260 33872
rect 8024 33856 8076 33862
rect 8024 33798 8076 33804
rect 8036 33658 8064 33798
rect 8220 33697 8248 33866
rect 8206 33688 8262 33697
rect 8024 33652 8076 33658
rect 8206 33623 8262 33632
rect 8024 33594 8076 33600
rect 8220 33522 8248 33623
rect 8208 33516 8260 33522
rect 8208 33458 8260 33464
rect 7840 32836 7892 32842
rect 7944 32830 8064 32858
rect 8220 32842 8248 33458
rect 8300 33108 8352 33114
rect 8300 33050 8352 33056
rect 7840 32778 7892 32784
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7564 30796 7616 30802
rect 7564 30738 7616 30744
rect 7576 29306 7604 30738
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 7668 29850 7696 30194
rect 7656 29844 7708 29850
rect 7656 29786 7708 29792
rect 7852 29306 7880 32778
rect 8036 32774 8064 32830
rect 8208 32836 8260 32842
rect 8208 32778 8260 32784
rect 8024 32768 8076 32774
rect 8024 32710 8076 32716
rect 7930 32056 7986 32065
rect 7930 31991 7932 32000
rect 7984 31991 7986 32000
rect 7932 31962 7984 31968
rect 8036 31414 8064 32710
rect 8312 32450 8340 33050
rect 8390 33008 8446 33017
rect 8390 32943 8446 32952
rect 8484 32972 8536 32978
rect 8404 32910 8432 32943
rect 8484 32914 8536 32920
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 8496 32570 8524 32914
rect 8576 32836 8628 32842
rect 8576 32778 8628 32784
rect 8484 32564 8536 32570
rect 8484 32506 8536 32512
rect 8496 32450 8524 32506
rect 8220 32434 8340 32450
rect 8208 32428 8340 32434
rect 8260 32422 8340 32428
rect 8208 32370 8260 32376
rect 8116 32224 8168 32230
rect 8116 32166 8168 32172
rect 8128 31822 8156 32166
rect 8116 31816 8168 31822
rect 8116 31758 8168 31764
rect 8024 31408 8076 31414
rect 8312 31385 8340 32422
rect 8404 32422 8524 32450
rect 8588 32434 8616 32778
rect 8680 32570 8708 35022
rect 8760 34128 8812 34134
rect 8760 34070 8812 34076
rect 8772 32978 8800 34070
rect 8864 32994 8892 36042
rect 8942 35728 8998 35737
rect 8942 35663 8944 35672
rect 8996 35663 8998 35672
rect 8944 35634 8996 35640
rect 9048 35630 9076 37198
rect 9324 36922 9352 39782
rect 9600 39098 9628 39986
rect 9864 39908 9916 39914
rect 9864 39850 9916 39856
rect 9876 39658 9904 39850
rect 9784 39642 9904 39658
rect 9772 39636 9904 39642
rect 9824 39630 9904 39636
rect 9772 39578 9824 39584
rect 9680 39432 9732 39438
rect 9680 39374 9732 39380
rect 9588 39092 9640 39098
rect 9588 39034 9640 39040
rect 9600 38706 9628 39034
rect 9508 38678 9628 38706
rect 9312 36916 9364 36922
rect 9312 36858 9364 36864
rect 9312 36168 9364 36174
rect 9312 36110 9364 36116
rect 9128 36032 9180 36038
rect 9128 35974 9180 35980
rect 9036 35624 9088 35630
rect 9036 35566 9088 35572
rect 9048 34406 9076 35566
rect 9036 34400 9088 34406
rect 9036 34342 9088 34348
rect 9036 33312 9088 33318
rect 9036 33254 9088 33260
rect 8760 32972 8812 32978
rect 8864 32966 8984 32994
rect 8760 32914 8812 32920
rect 8852 32836 8904 32842
rect 8852 32778 8904 32784
rect 8668 32564 8720 32570
rect 8668 32506 8720 32512
rect 8576 32428 8628 32434
rect 8024 31350 8076 31356
rect 8298 31376 8354 31385
rect 8036 30784 8064 31350
rect 8298 31311 8354 31320
rect 7944 30756 8064 30784
rect 7944 30190 7972 30756
rect 8312 30682 8340 31311
rect 8036 30654 8340 30682
rect 7932 30184 7984 30190
rect 7932 30126 7984 30132
rect 8036 29714 8064 30654
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 8404 29646 8432 32422
rect 8576 32370 8628 32376
rect 8576 32292 8628 32298
rect 8576 32234 8628 32240
rect 8484 32224 8536 32230
rect 8484 32166 8536 32172
rect 8496 32026 8524 32166
rect 8484 32020 8536 32026
rect 8484 31962 8536 31968
rect 8588 31872 8616 32234
rect 8496 31844 8616 31872
rect 8496 31754 8524 31844
rect 8484 31748 8536 31754
rect 8484 31690 8536 31696
rect 8496 30394 8524 31690
rect 8576 31680 8628 31686
rect 8680 31668 8708 32506
rect 8760 32020 8812 32026
rect 8760 31962 8812 31968
rect 8772 31793 8800 31962
rect 8758 31784 8814 31793
rect 8758 31719 8814 31728
rect 8864 31686 8892 32778
rect 8956 32774 8984 32966
rect 8944 32768 8996 32774
rect 8944 32710 8996 32716
rect 8956 31890 8984 32710
rect 9048 32366 9076 33254
rect 9036 32360 9088 32366
rect 9036 32302 9088 32308
rect 9140 32298 9168 35974
rect 9324 35494 9352 36110
rect 9508 35834 9536 38678
rect 9692 38570 9720 39374
rect 9876 39098 9904 39630
rect 9956 39364 10008 39370
rect 9956 39306 10008 39312
rect 9968 39098 9996 39306
rect 9864 39092 9916 39098
rect 9864 39034 9916 39040
rect 9956 39092 10008 39098
rect 9956 39034 10008 39040
rect 10428 38962 10456 40462
rect 10612 39370 10640 41074
rect 10888 40118 10916 41074
rect 11072 40594 11100 41210
rect 11704 41064 11756 41070
rect 11704 41006 11756 41012
rect 11716 40934 11744 41006
rect 11704 40928 11756 40934
rect 11704 40870 11756 40876
rect 11060 40588 11112 40594
rect 11060 40530 11112 40536
rect 10968 40452 11020 40458
rect 10968 40394 11020 40400
rect 10980 40202 11008 40394
rect 10980 40174 11100 40202
rect 11072 40118 11100 40174
rect 10876 40112 10928 40118
rect 10968 40112 11020 40118
rect 10876 40054 10928 40060
rect 10966 40080 10968 40089
rect 11060 40112 11112 40118
rect 11020 40080 11022 40089
rect 11060 40054 11112 40060
rect 10966 40015 11022 40024
rect 10968 39976 11020 39982
rect 10968 39918 11020 39924
rect 10980 39574 11008 39918
rect 10968 39568 11020 39574
rect 10968 39510 11020 39516
rect 10600 39364 10652 39370
rect 10600 39306 10652 39312
rect 10416 38956 10468 38962
rect 10416 38898 10468 38904
rect 10612 38826 10640 39306
rect 10980 38962 11008 39510
rect 11612 39500 11664 39506
rect 11612 39442 11664 39448
rect 10968 38956 11020 38962
rect 10968 38898 11020 38904
rect 11428 38956 11480 38962
rect 11428 38898 11480 38904
rect 10600 38820 10652 38826
rect 10600 38762 10652 38768
rect 9600 38542 9720 38570
rect 9600 38418 9628 38542
rect 9588 38412 9640 38418
rect 9588 38354 9640 38360
rect 9600 37806 9628 38354
rect 10612 37942 10640 38762
rect 11440 38418 11468 38898
rect 11428 38412 11480 38418
rect 11428 38354 11480 38360
rect 10600 37936 10652 37942
rect 10600 37878 10652 37884
rect 9588 37800 9640 37806
rect 9588 37742 9640 37748
rect 10324 37664 10376 37670
rect 10324 37606 10376 37612
rect 10336 37330 10364 37606
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 11336 37256 11388 37262
rect 11336 37198 11388 37204
rect 11152 37188 11204 37194
rect 11152 37130 11204 37136
rect 10782 37088 10838 37097
rect 10782 37023 10838 37032
rect 9586 36816 9642 36825
rect 10796 36786 10824 37023
rect 11164 36854 11192 37130
rect 11152 36848 11204 36854
rect 11152 36790 11204 36796
rect 11348 36786 11376 37198
rect 11440 36786 11468 38354
rect 11520 37800 11572 37806
rect 11520 37742 11572 37748
rect 11532 37466 11560 37742
rect 11520 37460 11572 37466
rect 11520 37402 11572 37408
rect 11520 37324 11572 37330
rect 11520 37266 11572 37272
rect 11532 36922 11560 37266
rect 11520 36916 11572 36922
rect 11520 36858 11572 36864
rect 9586 36751 9642 36760
rect 9772 36780 9824 36786
rect 9496 35828 9548 35834
rect 9496 35770 9548 35776
rect 9312 35488 9364 35494
rect 9312 35430 9364 35436
rect 9220 35284 9272 35290
rect 9220 35226 9272 35232
rect 9232 34678 9260 35226
rect 9220 34672 9272 34678
rect 9220 34614 9272 34620
rect 9324 34542 9352 35430
rect 9508 35154 9536 35770
rect 9600 35222 9628 36751
rect 9772 36722 9824 36728
rect 10784 36780 10836 36786
rect 10784 36722 10836 36728
rect 11336 36780 11388 36786
rect 11336 36722 11388 36728
rect 11428 36780 11480 36786
rect 11428 36722 11480 36728
rect 11520 36780 11572 36786
rect 11520 36722 11572 36728
rect 9784 36582 9812 36722
rect 10048 36644 10100 36650
rect 10048 36586 10100 36592
rect 9772 36576 9824 36582
rect 9772 36518 9824 36524
rect 9588 35216 9640 35222
rect 9588 35158 9640 35164
rect 9496 35148 9548 35154
rect 9496 35090 9548 35096
rect 9600 35057 9628 35158
rect 9586 35048 9642 35057
rect 9404 35012 9456 35018
rect 9586 34983 9642 34992
rect 9404 34954 9456 34960
rect 9416 34746 9444 34954
rect 9588 34944 9640 34950
rect 9588 34886 9640 34892
rect 9404 34740 9456 34746
rect 9404 34682 9456 34688
rect 9312 34536 9364 34542
rect 9312 34478 9364 34484
rect 9220 33448 9272 33454
rect 9220 33390 9272 33396
rect 9128 32292 9180 32298
rect 9128 32234 9180 32240
rect 9232 32178 9260 33390
rect 9324 32570 9352 34478
rect 9404 34400 9456 34406
rect 9404 34342 9456 34348
rect 9416 34134 9444 34342
rect 9404 34128 9456 34134
rect 9404 34070 9456 34076
rect 9496 33856 9548 33862
rect 9496 33798 9548 33804
rect 9508 33522 9536 33798
rect 9600 33658 9628 34886
rect 9680 34400 9732 34406
rect 9680 34342 9732 34348
rect 9692 34202 9720 34342
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 9588 33652 9640 33658
rect 9588 33594 9640 33600
rect 9496 33516 9548 33522
rect 9496 33458 9548 33464
rect 9312 32564 9364 32570
rect 9312 32506 9364 32512
rect 9324 32298 9352 32506
rect 9312 32292 9364 32298
rect 9312 32234 9364 32240
rect 9496 32292 9548 32298
rect 9496 32234 9548 32240
rect 9048 32150 9260 32178
rect 9310 32192 9366 32201
rect 8944 31884 8996 31890
rect 8944 31826 8996 31832
rect 8852 31680 8904 31686
rect 8680 31640 8800 31668
rect 8576 31622 8628 31628
rect 8484 30388 8536 30394
rect 8484 30330 8536 30336
rect 7932 29640 7984 29646
rect 7932 29582 7984 29588
rect 8208 29640 8260 29646
rect 8208 29582 8260 29588
rect 8392 29640 8444 29646
rect 8392 29582 8444 29588
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 7564 29300 7616 29306
rect 7564 29242 7616 29248
rect 7840 29300 7892 29306
rect 7840 29242 7892 29248
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 7576 28762 7604 29106
rect 7944 29102 7972 29582
rect 7932 29096 7984 29102
rect 7932 29038 7984 29044
rect 8116 29096 8168 29102
rect 8116 29038 8168 29044
rect 8128 28994 8156 29038
rect 8220 29034 8248 29582
rect 8300 29504 8352 29510
rect 8300 29446 8352 29452
rect 8036 28966 8156 28994
rect 8208 29028 8260 29034
rect 8208 28970 8260 28976
rect 7564 28756 7616 28762
rect 7564 28698 7616 28704
rect 8036 28082 8064 28966
rect 8024 28076 8076 28082
rect 8024 28018 8076 28024
rect 8220 27062 8248 28970
rect 8312 28150 8340 29446
rect 8496 29306 8524 29582
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 8588 29186 8616 31622
rect 8772 31346 8800 31640
rect 8852 31622 8904 31628
rect 8852 31476 8904 31482
rect 8852 31418 8904 31424
rect 8760 31340 8812 31346
rect 8760 31282 8812 31288
rect 8668 31204 8720 31210
rect 8668 31146 8720 31152
rect 8680 29578 8708 31146
rect 8760 30184 8812 30190
rect 8760 30126 8812 30132
rect 8668 29572 8720 29578
rect 8668 29514 8720 29520
rect 8772 29306 8800 30126
rect 8864 30122 8892 31418
rect 8956 31346 8984 31826
rect 9048 31754 9076 32150
rect 9310 32127 9366 32136
rect 9324 32008 9352 32127
rect 9232 31980 9352 32008
rect 9128 31952 9180 31958
rect 9128 31894 9180 31900
rect 9036 31748 9088 31754
rect 9036 31690 9088 31696
rect 8944 31340 8996 31346
rect 8944 31282 8996 31288
rect 9048 30666 9076 31690
rect 9036 30660 9088 30666
rect 9036 30602 9088 30608
rect 8944 30592 8996 30598
rect 8944 30534 8996 30540
rect 8852 30116 8904 30122
rect 8852 30058 8904 30064
rect 8956 29714 8984 30534
rect 8944 29708 8996 29714
rect 8944 29650 8996 29656
rect 8852 29572 8904 29578
rect 8852 29514 8904 29520
rect 8760 29300 8812 29306
rect 8760 29242 8812 29248
rect 8496 29158 8616 29186
rect 8300 28144 8352 28150
rect 8300 28086 8352 28092
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 8208 27056 8260 27062
rect 8208 26998 8260 27004
rect 8220 26382 8248 26998
rect 8312 26790 8340 27950
rect 8496 27538 8524 29158
rect 8772 28558 8800 29242
rect 8760 28552 8812 28558
rect 8760 28494 8812 28500
rect 8576 28144 8628 28150
rect 8576 28086 8628 28092
rect 8484 27532 8536 27538
rect 8484 27474 8536 27480
rect 8300 26784 8352 26790
rect 8300 26726 8352 26732
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8114 26208 8170 26217
rect 8114 26143 8170 26152
rect 8024 25968 8076 25974
rect 8024 25910 8076 25916
rect 8036 25294 8064 25910
rect 8128 25294 8156 26143
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 8024 25288 8076 25294
rect 8024 25230 8076 25236
rect 8116 25288 8168 25294
rect 8116 25230 8168 25236
rect 8220 24750 8248 25298
rect 8312 24954 8340 26726
rect 8392 26444 8444 26450
rect 8392 26386 8444 26392
rect 8404 25226 8432 26386
rect 8496 26246 8524 27474
rect 8484 26240 8536 26246
rect 8484 26182 8536 26188
rect 8496 26042 8524 26182
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 8588 25906 8616 28086
rect 8864 27614 8892 29514
rect 8956 28218 8984 29650
rect 9036 29504 9088 29510
rect 9140 29492 9168 31894
rect 9232 31686 9260 31980
rect 9508 31872 9536 32234
rect 9600 32201 9628 33594
rect 9678 32328 9734 32337
rect 9678 32263 9734 32272
rect 9586 32192 9642 32201
rect 9586 32127 9642 32136
rect 9692 32026 9720 32263
rect 9784 32026 9812 36518
rect 10060 36174 10088 36586
rect 11440 36242 11468 36722
rect 11532 36582 11560 36722
rect 11520 36576 11572 36582
rect 11520 36518 11572 36524
rect 11428 36236 11480 36242
rect 11428 36178 11480 36184
rect 10048 36168 10100 36174
rect 10048 36110 10100 36116
rect 10508 36100 10560 36106
rect 10508 36042 10560 36048
rect 10692 36100 10744 36106
rect 10692 36042 10744 36048
rect 11336 36100 11388 36106
rect 11336 36042 11388 36048
rect 10232 35828 10284 35834
rect 10232 35770 10284 35776
rect 10046 35728 10102 35737
rect 10046 35663 10102 35672
rect 10060 35494 10088 35663
rect 10140 35624 10192 35630
rect 10140 35566 10192 35572
rect 9864 35488 9916 35494
rect 9864 35430 9916 35436
rect 10048 35488 10100 35494
rect 10048 35430 10100 35436
rect 9876 35290 9904 35430
rect 9864 35284 9916 35290
rect 9916 35244 9996 35272
rect 9864 35226 9916 35232
rect 9968 34066 9996 35244
rect 10046 34640 10102 34649
rect 10152 34610 10180 35566
rect 10244 35494 10272 35770
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 10244 35290 10272 35430
rect 10232 35284 10284 35290
rect 10232 35226 10284 35232
rect 10324 35216 10376 35222
rect 10376 35176 10456 35204
rect 10324 35158 10376 35164
rect 10232 35080 10284 35086
rect 10232 35022 10284 35028
rect 10046 34575 10102 34584
rect 10140 34604 10192 34610
rect 10060 34474 10088 34575
rect 10140 34546 10192 34552
rect 10048 34468 10100 34474
rect 10048 34410 10100 34416
rect 10244 34134 10272 35022
rect 10232 34128 10284 34134
rect 10232 34070 10284 34076
rect 9956 34060 10008 34066
rect 9956 34002 10008 34008
rect 9864 33992 9916 33998
rect 9864 33934 9916 33940
rect 9876 33522 9904 33934
rect 10324 33924 10376 33930
rect 10324 33866 10376 33872
rect 9956 33856 10008 33862
rect 9956 33798 10008 33804
rect 9864 33516 9916 33522
rect 9864 33458 9916 33464
rect 9864 33380 9916 33386
rect 9864 33322 9916 33328
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9772 32020 9824 32026
rect 9772 31962 9824 31968
rect 9876 31906 9904 33322
rect 9416 31844 9536 31872
rect 9784 31878 9904 31906
rect 9220 31680 9272 31686
rect 9220 31622 9272 31628
rect 9416 31634 9444 31844
rect 9784 31804 9812 31878
rect 9586 31784 9642 31793
rect 9586 31719 9642 31728
rect 9692 31776 9812 31804
rect 9600 31686 9628 31719
rect 9588 31680 9640 31686
rect 9232 31482 9260 31622
rect 9416 31606 9536 31634
rect 9588 31622 9640 31628
rect 9402 31512 9458 31521
rect 9220 31476 9272 31482
rect 9402 31447 9458 31456
rect 9220 31418 9272 31424
rect 9416 31414 9444 31447
rect 9404 31408 9456 31414
rect 9404 31350 9456 31356
rect 9404 31204 9456 31210
rect 9404 31146 9456 31152
rect 9220 30048 9272 30054
rect 9220 29990 9272 29996
rect 9088 29464 9168 29492
rect 9036 29446 9088 29452
rect 9128 29028 9180 29034
rect 9128 28970 9180 28976
rect 9140 28694 9168 28970
rect 9128 28688 9180 28694
rect 9128 28630 9180 28636
rect 8944 28212 8996 28218
rect 8944 28154 8996 28160
rect 9126 28112 9182 28121
rect 9126 28047 9128 28056
rect 9180 28047 9182 28056
rect 9128 28018 9180 28024
rect 8944 27940 8996 27946
rect 8944 27882 8996 27888
rect 8772 27586 8892 27614
rect 8956 27606 8984 27882
rect 9036 27668 9088 27674
rect 9036 27610 9088 27616
rect 8944 27600 8996 27606
rect 8668 26308 8720 26314
rect 8668 26250 8720 26256
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8392 25220 8444 25226
rect 8392 25162 8444 25168
rect 8496 24954 8524 25230
rect 8588 24954 8616 25842
rect 8300 24948 8352 24954
rect 8300 24890 8352 24896
rect 8484 24948 8536 24954
rect 8484 24890 8536 24896
rect 8576 24948 8628 24954
rect 8576 24890 8628 24896
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8208 24744 8260 24750
rect 8404 24721 8432 24754
rect 8208 24686 8260 24692
rect 8390 24712 8446 24721
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7380 24336 7432 24342
rect 7380 24278 7432 24284
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 6840 23118 6868 24006
rect 7024 23662 7052 24006
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 7116 23322 7144 24142
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 7852 23186 7880 24550
rect 8220 24274 8248 24686
rect 8390 24647 8446 24656
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8496 23497 8524 24890
rect 8680 24818 8708 26250
rect 8772 26042 8800 27586
rect 8944 27542 8996 27548
rect 8852 27464 8904 27470
rect 8850 27432 8852 27441
rect 8904 27432 8906 27441
rect 8850 27367 8906 27376
rect 8864 27062 8892 27367
rect 8852 27056 8904 27062
rect 8852 26998 8904 27004
rect 9048 26994 9076 27610
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 8760 26036 8812 26042
rect 8760 25978 8812 25984
rect 8864 25906 8892 26726
rect 9034 26344 9090 26353
rect 9034 26279 9090 26288
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 8852 25900 8904 25906
rect 8852 25842 8904 25848
rect 8772 25498 8800 25842
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 9048 25430 9076 26279
rect 9036 25424 9088 25430
rect 9036 25366 9088 25372
rect 9140 25362 9168 28018
rect 9232 27606 9260 29990
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9220 27600 9272 27606
rect 9220 27542 9272 27548
rect 9232 26382 9260 27542
rect 9220 26376 9272 26382
rect 9220 26318 9272 26324
rect 9324 25702 9352 29582
rect 9416 29510 9444 31146
rect 9508 29866 9536 31606
rect 9588 31408 9640 31414
rect 9586 31376 9588 31385
rect 9692 31396 9720 31776
rect 9772 31680 9824 31686
rect 9772 31622 9824 31628
rect 9640 31376 9720 31396
rect 9642 31368 9720 31376
rect 9586 31311 9642 31320
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 9600 30938 9628 31214
rect 9588 30932 9640 30938
rect 9588 30874 9640 30880
rect 9588 30660 9640 30666
rect 9784 30648 9812 31622
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9640 30620 9812 30648
rect 9588 30602 9640 30608
rect 9600 30122 9628 30602
rect 9680 30388 9732 30394
rect 9680 30330 9732 30336
rect 9588 30116 9640 30122
rect 9588 30058 9640 30064
rect 9508 29838 9628 29866
rect 9496 29776 9548 29782
rect 9496 29718 9548 29724
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9416 29306 9444 29446
rect 9404 29300 9456 29306
rect 9404 29242 9456 29248
rect 9404 29164 9456 29170
rect 9404 29106 9456 29112
rect 9416 28558 9444 29106
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9508 28014 9536 29718
rect 9600 29714 9628 29838
rect 9692 29782 9720 30330
rect 9772 30048 9824 30054
rect 9772 29990 9824 29996
rect 9680 29776 9732 29782
rect 9680 29718 9732 29724
rect 9588 29708 9640 29714
rect 9588 29650 9640 29656
rect 9784 29646 9812 29990
rect 9680 29640 9732 29646
rect 9680 29582 9732 29588
rect 9772 29640 9824 29646
rect 9772 29582 9824 29588
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 9600 29238 9628 29514
rect 9588 29232 9640 29238
rect 9588 29174 9640 29180
rect 9692 29170 9720 29582
rect 9784 29170 9812 29582
rect 9680 29164 9732 29170
rect 9680 29106 9732 29112
rect 9772 29164 9824 29170
rect 9772 29106 9824 29112
rect 9678 29064 9734 29073
rect 9678 28999 9680 29008
rect 9732 28999 9734 29008
rect 9772 29028 9824 29034
rect 9680 28970 9732 28976
rect 9772 28970 9824 28976
rect 9496 28008 9548 28014
rect 9496 27950 9548 27956
rect 9508 27538 9536 27950
rect 9404 27532 9456 27538
rect 9404 27474 9456 27480
rect 9496 27532 9548 27538
rect 9496 27474 9548 27480
rect 9416 27062 9444 27474
rect 9588 27464 9640 27470
rect 9586 27432 9588 27441
rect 9640 27432 9642 27441
rect 9586 27367 9642 27376
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9508 27062 9536 27270
rect 9404 27056 9456 27062
rect 9404 26998 9456 27004
rect 9496 27056 9548 27062
rect 9496 26998 9548 27004
rect 9416 26625 9444 26998
rect 9692 26874 9720 28970
rect 9784 27470 9812 28970
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9784 26994 9812 27406
rect 9876 26994 9904 31078
rect 9968 30802 9996 33798
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 10060 31890 10088 32710
rect 10140 32360 10192 32366
rect 10140 32302 10192 32308
rect 10048 31884 10100 31890
rect 10048 31826 10100 31832
rect 10048 31748 10100 31754
rect 10048 31690 10100 31696
rect 10060 31482 10088 31690
rect 10048 31476 10100 31482
rect 10048 31418 10100 31424
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 9956 30592 10008 30598
rect 9956 30534 10008 30540
rect 9968 29782 9996 30534
rect 9956 29776 10008 29782
rect 9956 29718 10008 29724
rect 10060 29646 10088 31078
rect 10152 30054 10180 32302
rect 10232 31952 10284 31958
rect 10232 31894 10284 31900
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 10048 29640 10100 29646
rect 10048 29582 10100 29588
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9968 28994 9996 29446
rect 10060 29170 10088 29582
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 9968 28966 10088 28994
rect 10060 27470 10088 28966
rect 10152 28937 10180 29582
rect 10138 28928 10194 28937
rect 10138 28863 10194 28872
rect 10048 27464 10100 27470
rect 10048 27406 10100 27412
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9864 26988 9916 26994
rect 9864 26930 9916 26936
rect 9508 26846 9720 26874
rect 9402 26616 9458 26625
rect 9402 26551 9458 26560
rect 9508 26518 9536 26846
rect 9784 26790 9812 26930
rect 9956 26852 10008 26858
rect 9956 26794 10008 26800
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9496 26512 9548 26518
rect 9496 26454 9548 26460
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 9416 26217 9444 26318
rect 9402 26208 9458 26217
rect 9402 26143 9458 26152
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9232 25362 9260 25638
rect 9128 25356 9180 25362
rect 9128 25298 9180 25304
rect 9220 25356 9272 25362
rect 9220 25298 9272 25304
rect 9416 25294 9444 25842
rect 9508 25294 9536 26454
rect 9692 25974 9720 26726
rect 9784 26450 9812 26726
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 9968 26382 9996 26794
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 9862 25936 9918 25945
rect 9588 25832 9640 25838
rect 9586 25800 9588 25809
rect 9640 25800 9642 25809
rect 9586 25735 9642 25744
rect 9588 25696 9640 25702
rect 9588 25638 9640 25644
rect 9600 25430 9628 25638
rect 9588 25424 9640 25430
rect 9588 25366 9640 25372
rect 9692 25294 9720 25910
rect 9968 25906 9996 26318
rect 10060 25974 10088 27406
rect 10152 27062 10180 28863
rect 10244 28762 10272 31894
rect 10336 29646 10364 33866
rect 10428 32230 10456 35176
rect 10520 35154 10548 36042
rect 10508 35148 10560 35154
rect 10508 35090 10560 35096
rect 10704 34785 10732 36042
rect 10874 35728 10930 35737
rect 10784 35692 10836 35698
rect 10874 35663 10930 35672
rect 10784 35634 10836 35640
rect 10796 35018 10824 35634
rect 10888 35562 10916 35663
rect 10876 35556 10928 35562
rect 10876 35498 10928 35504
rect 10876 35080 10928 35086
rect 10876 35022 10928 35028
rect 10784 35012 10836 35018
rect 10784 34954 10836 34960
rect 10690 34776 10746 34785
rect 10690 34711 10746 34720
rect 10784 34128 10836 34134
rect 10784 34070 10836 34076
rect 10508 33992 10560 33998
rect 10508 33934 10560 33940
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10428 31890 10456 32166
rect 10416 31884 10468 31890
rect 10416 31826 10468 31832
rect 10428 31142 10456 31826
rect 10520 31754 10548 33934
rect 10600 32564 10652 32570
rect 10600 32506 10652 32512
rect 10612 32366 10640 32506
rect 10600 32360 10652 32366
rect 10600 32302 10652 32308
rect 10508 31748 10560 31754
rect 10508 31690 10560 31696
rect 10520 31482 10548 31690
rect 10508 31476 10560 31482
rect 10508 31418 10560 31424
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10428 30258 10456 30534
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10520 30190 10548 31078
rect 10612 30240 10640 32302
rect 10796 32230 10824 34070
rect 10888 33998 10916 35022
rect 11060 34944 11112 34950
rect 11060 34886 11112 34892
rect 11072 34649 11100 34886
rect 11058 34640 11114 34649
rect 11058 34575 11114 34584
rect 11152 34128 11204 34134
rect 11152 34070 11204 34076
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 11060 33856 11112 33862
rect 11060 33798 11112 33804
rect 11072 33318 11100 33798
rect 11060 33312 11112 33318
rect 11060 33254 11112 33260
rect 11072 32434 11100 33254
rect 11164 32473 11192 34070
rect 11348 33810 11376 36042
rect 11624 35494 11652 39442
rect 11716 38654 11744 40870
rect 12452 40526 12480 41482
rect 12624 40588 12676 40594
rect 12624 40530 12676 40536
rect 12440 40520 12492 40526
rect 12440 40462 12492 40468
rect 12636 40186 12664 40530
rect 12624 40180 12676 40186
rect 12624 40122 12676 40128
rect 12440 40112 12492 40118
rect 12440 40054 12492 40060
rect 12164 39296 12216 39302
rect 12164 39238 12216 39244
rect 12176 39098 12204 39238
rect 12164 39092 12216 39098
rect 12164 39034 12216 39040
rect 11716 38626 11928 38654
rect 11796 38276 11848 38282
rect 11796 38218 11848 38224
rect 11808 38010 11836 38218
rect 11796 38004 11848 38010
rect 11796 37946 11848 37952
rect 11796 36780 11848 36786
rect 11796 36722 11848 36728
rect 11808 36038 11836 36722
rect 11900 36666 11928 38626
rect 12256 38412 12308 38418
rect 12256 38354 12308 38360
rect 11980 37936 12032 37942
rect 11980 37878 12032 37884
rect 11992 37194 12020 37878
rect 12164 37664 12216 37670
rect 12164 37606 12216 37612
rect 11980 37188 12032 37194
rect 11980 37130 12032 37136
rect 11992 36786 12020 37130
rect 12072 36916 12124 36922
rect 12072 36858 12124 36864
rect 11980 36780 12032 36786
rect 11980 36722 12032 36728
rect 11900 36638 12020 36666
rect 11796 36032 11848 36038
rect 11796 35974 11848 35980
rect 11704 35556 11756 35562
rect 11704 35498 11756 35504
rect 11888 35556 11940 35562
rect 11888 35498 11940 35504
rect 11612 35488 11664 35494
rect 11612 35430 11664 35436
rect 11520 35080 11572 35086
rect 11624 35068 11652 35430
rect 11716 35154 11744 35498
rect 11704 35148 11756 35154
rect 11704 35090 11756 35096
rect 11796 35148 11848 35154
rect 11796 35090 11848 35096
rect 11572 35040 11652 35068
rect 11520 35022 11572 35028
rect 11520 34944 11572 34950
rect 11520 34886 11572 34892
rect 11428 34536 11480 34542
rect 11428 34478 11480 34484
rect 11256 33782 11376 33810
rect 11150 32464 11206 32473
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 11060 32428 11112 32434
rect 11150 32399 11206 32408
rect 11060 32370 11112 32376
rect 10784 32224 10836 32230
rect 10784 32166 10836 32172
rect 10690 32056 10746 32065
rect 10888 32042 10916 32370
rect 11152 32360 11204 32366
rect 11152 32302 11204 32308
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 10746 32014 10916 32042
rect 10690 31991 10746 32000
rect 10784 31952 10836 31958
rect 10784 31894 10836 31900
rect 10796 31793 10824 31894
rect 10782 31784 10838 31793
rect 10782 31719 10838 31728
rect 10690 31648 10746 31657
rect 10690 31583 10746 31592
rect 10704 30870 10732 31583
rect 10692 30864 10744 30870
rect 10692 30806 10744 30812
rect 10796 30802 10824 31719
rect 10968 31680 11020 31686
rect 10968 31622 11020 31628
rect 10980 31278 11008 31622
rect 10968 31272 11020 31278
rect 10968 31214 11020 31220
rect 10980 30938 11008 31214
rect 10968 30932 11020 30938
rect 10968 30874 11020 30880
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 10980 30433 11008 30670
rect 10966 30424 11022 30433
rect 11072 30394 11100 32166
rect 11164 31385 11192 32302
rect 11150 31376 11206 31385
rect 11150 31311 11206 31320
rect 10966 30359 11022 30368
rect 11060 30388 11112 30394
rect 11060 30330 11112 30336
rect 10692 30252 10744 30258
rect 10612 30212 10692 30240
rect 10692 30194 10744 30200
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 10520 29889 10548 30126
rect 10600 30116 10652 30122
rect 10600 30058 10652 30064
rect 10506 29880 10562 29889
rect 10506 29815 10562 29824
rect 10520 29646 10548 29815
rect 10324 29640 10376 29646
rect 10324 29582 10376 29588
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10520 29238 10548 29582
rect 10508 29232 10560 29238
rect 10506 29200 10508 29209
rect 10560 29200 10562 29209
rect 10506 29135 10562 29144
rect 10414 29064 10470 29073
rect 10414 28999 10470 29008
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10244 27674 10272 28698
rect 10428 28626 10456 28999
rect 10416 28620 10468 28626
rect 10416 28562 10468 28568
rect 10612 28014 10640 30058
rect 10600 28008 10652 28014
rect 10600 27950 10652 27956
rect 10232 27668 10284 27674
rect 10232 27610 10284 27616
rect 10612 27334 10640 27950
rect 10600 27328 10652 27334
rect 10322 27296 10378 27305
rect 10600 27270 10652 27276
rect 10322 27231 10378 27240
rect 10140 27056 10192 27062
rect 10140 26998 10192 27004
rect 10140 26920 10192 26926
rect 10138 26888 10140 26897
rect 10232 26920 10284 26926
rect 10192 26888 10194 26897
rect 10232 26862 10284 26868
rect 10138 26823 10194 26832
rect 10048 25968 10100 25974
rect 10048 25910 10100 25916
rect 9862 25871 9918 25880
rect 9956 25900 10008 25906
rect 9770 25800 9826 25809
rect 9770 25735 9826 25744
rect 9784 25498 9812 25735
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9404 25288 9456 25294
rect 9034 25256 9090 25265
rect 9496 25288 9548 25294
rect 9404 25230 9456 25236
rect 9494 25256 9496 25265
rect 9680 25288 9732 25294
rect 9548 25256 9550 25265
rect 9090 25200 9168 25208
rect 9034 25191 9036 25200
rect 9088 25180 9168 25200
rect 9680 25230 9732 25236
rect 9494 25191 9550 25200
rect 9036 25162 9088 25168
rect 9140 24818 9168 25180
rect 9404 25152 9456 25158
rect 9876 25106 9904 25871
rect 9956 25842 10008 25848
rect 9956 25764 10008 25770
rect 9956 25706 10008 25712
rect 9456 25100 9904 25106
rect 9404 25094 9904 25100
rect 9416 25078 9904 25094
rect 9218 24848 9274 24857
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 9128 24812 9180 24818
rect 9218 24783 9274 24792
rect 9128 24754 9180 24760
rect 8772 23866 8800 24754
rect 8864 24206 8892 24754
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 8760 23860 8812 23866
rect 8760 23802 8812 23808
rect 9140 23526 9168 24550
rect 8852 23520 8904 23526
rect 8482 23488 8538 23497
rect 8852 23462 8904 23468
rect 9128 23520 9180 23526
rect 9128 23462 9180 23468
rect 8482 23423 8538 23432
rect 8864 23186 8892 23462
rect 9232 23254 9260 24783
rect 9312 24744 9364 24750
rect 9310 24712 9312 24721
rect 9364 24712 9366 24721
rect 9968 24682 9996 25706
rect 10060 24886 10088 25910
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 9310 24647 9366 24656
rect 9956 24676 10008 24682
rect 9956 24618 10008 24624
rect 10152 24206 10180 26823
rect 10244 26314 10272 26862
rect 10232 26308 10284 26314
rect 10232 26250 10284 26256
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9220 23248 9272 23254
rect 9218 23216 9220 23225
rect 9272 23216 9274 23225
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 8852 23180 8904 23186
rect 9218 23151 9274 23160
rect 8852 23122 8904 23128
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 9324 23050 9352 24142
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 8024 23044 8076 23050
rect 8024 22986 8076 22992
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6380 22066 6500 22094
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5184 20777 5212 21490
rect 5644 20942 5672 22066
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5828 21554 5856 21830
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5828 20874 5856 21286
rect 5920 21146 5948 21286
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 6472 21010 6500 22066
rect 6564 21622 6592 22510
rect 7116 21622 7144 22578
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 6552 21616 6604 21622
rect 7104 21616 7156 21622
rect 6552 21558 6604 21564
rect 7102 21584 7104 21593
rect 7156 21584 7158 21593
rect 7102 21519 7158 21528
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 6656 21146 6684 21422
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 5816 20868 5868 20874
rect 5816 20810 5868 20816
rect 5170 20768 5226 20777
rect 5170 20703 5226 20712
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5184 19174 5212 19790
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5184 18426 5212 19110
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5092 17326 5212 17354
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 5092 16726 5120 17138
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 4988 16584 5040 16590
rect 5184 16538 5212 17326
rect 5276 17218 5304 20198
rect 6656 20058 6684 20878
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5460 18850 5488 19314
rect 6000 19304 6052 19310
rect 5814 19272 5870 19281
rect 6000 19246 6052 19252
rect 5814 19207 5816 19216
rect 5868 19207 5870 19216
rect 5816 19178 5868 19184
rect 5828 18902 5856 19178
rect 5816 18896 5868 18902
rect 5356 18828 5408 18834
rect 5460 18822 5580 18850
rect 5816 18838 5868 18844
rect 5356 18770 5408 18776
rect 5368 18086 5396 18770
rect 5552 18766 5580 18822
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5460 18358 5488 18702
rect 5552 18426 5580 18702
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17678 5396 18022
rect 5460 17746 5488 18294
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5552 17678 5580 18158
rect 5828 17678 5856 18838
rect 6012 18426 6040 19246
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 18834 6408 19110
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6380 18698 6408 18770
rect 6564 18698 6592 19790
rect 6644 19372 6696 19378
rect 6748 19360 6776 21082
rect 6920 21072 6972 21078
rect 6920 21014 6972 21020
rect 6932 20942 6960 21014
rect 6920 20936 6972 20942
rect 6840 20884 6920 20890
rect 6840 20878 6972 20884
rect 6840 20862 6960 20878
rect 6840 19854 6868 20862
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 19922 6960 20742
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6828 19848 6880 19854
rect 6880 19796 6960 19802
rect 6828 19790 6960 19796
rect 6840 19774 6960 19790
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6840 19514 6868 19654
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6696 19332 6776 19360
rect 6644 19314 6696 19320
rect 6368 18692 6420 18698
rect 6368 18634 6420 18640
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5276 17202 5396 17218
rect 5276 17196 5408 17202
rect 5276 17190 5356 17196
rect 5356 17138 5408 17144
rect 4988 16526 5040 16532
rect 5092 16510 5212 16538
rect 5264 16516 5316 16522
rect 5092 16402 5120 16510
rect 5264 16458 5316 16464
rect 5000 16374 5120 16402
rect 4896 15972 4948 15978
rect 4896 15914 4948 15920
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4540 14074 4568 14350
rect 4632 14278 4660 15846
rect 4816 15570 4844 15846
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4080 11898 4108 12106
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4632 11626 4660 14214
rect 4908 12646 4936 14214
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11354 4660 11562
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4632 9586 4660 9930
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4356 9450 4660 9466
rect 4344 9444 4672 9450
rect 4396 9438 4620 9444
rect 4344 9386 4396 9392
rect 4620 9386 4672 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 8974 4660 9386
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 4632 8566 4660 8910
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7954 4660 8230
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 940 7880 992 7886
rect 940 7822 992 7828
rect 952 7585 980 7822
rect 4724 7818 4752 12106
rect 4908 11762 4936 12582
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4816 9178 4844 9998
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4908 9042 4936 9590
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 938 7576 994 7585
rect 938 7511 994 7520
rect 4080 6866 4108 7754
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4724 6730 4752 7754
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4908 6458 4936 8570
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 5000 6390 5028 16374
rect 5276 16250 5304 16458
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5092 14482 5120 15438
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5262 13696 5318 13705
rect 5262 13631 5318 13640
rect 5276 12850 5304 13631
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5092 11558 5120 12786
rect 5184 11830 5212 12786
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5184 11218 5212 11766
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 10266 5212 11154
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5092 9518 5120 9862
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5184 9450 5212 9998
rect 5368 9654 5396 17138
rect 5552 17134 5580 17478
rect 5828 17270 5856 17614
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 6012 17202 6040 18362
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5552 16522 5580 17070
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 15201 5488 15438
rect 5446 15192 5502 15201
rect 5552 15162 5580 16458
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5644 16046 5672 16390
rect 5736 16114 5764 16390
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5446 15127 5502 15136
rect 5540 15156 5592 15162
rect 5460 14498 5488 15127
rect 5540 15098 5592 15104
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5828 14618 5856 14962
rect 5920 14958 5948 16186
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5920 14618 5948 14894
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5460 14470 5580 14498
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5460 11830 5488 12650
rect 5552 12186 5580 14470
rect 5736 14414 5764 14554
rect 5816 14476 5868 14482
rect 6184 14476 6236 14482
rect 5868 14436 6184 14464
rect 5816 14418 5868 14424
rect 6184 14418 6236 14424
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 5736 13394 5764 14350
rect 6288 13530 6316 14350
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 6092 12912 6144 12918
rect 6092 12854 6144 12860
rect 6276 12912 6328 12918
rect 6380 12900 6408 14826
rect 6328 12872 6408 12900
rect 6276 12854 6328 12860
rect 6104 12306 6132 12854
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6276 12300 6328 12306
rect 6380 12288 6408 12582
rect 6328 12260 6408 12288
rect 6276 12242 6328 12248
rect 5552 12158 5764 12186
rect 6472 12170 6500 15914
rect 6564 15094 6592 16050
rect 6656 15978 6684 19314
rect 6932 18970 6960 19774
rect 7024 19174 7052 21422
rect 7196 19984 7248 19990
rect 7196 19926 7248 19932
rect 7208 19854 7236 19926
rect 7392 19854 7420 22170
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7944 21146 7972 21830
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 7562 21040 7618 21049
rect 7562 20975 7564 20984
rect 7616 20975 7618 20984
rect 7564 20946 7616 20952
rect 7196 19848 7248 19854
rect 7380 19848 7432 19854
rect 7248 19808 7328 19836
rect 7196 19790 7248 19796
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6840 18698 6868 18838
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 7208 18630 7236 19654
rect 7300 19378 7328 19808
rect 7380 19790 7432 19796
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7392 19258 7420 19790
rect 7300 19230 7420 19258
rect 7300 18766 7328 19230
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18766 7788 19110
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7380 18760 7432 18766
rect 7748 18760 7800 18766
rect 7380 18702 7432 18708
rect 7470 18728 7526 18737
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 6748 17202 6776 18566
rect 7208 18290 7236 18566
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7208 17338 7236 18226
rect 7300 18086 7328 18702
rect 7392 18358 7420 18702
rect 7748 18702 7800 18708
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7470 18663 7472 18672
rect 7524 18663 7526 18672
rect 7472 18634 7524 18640
rect 7944 18426 7972 18702
rect 8036 18426 8064 22986
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8128 22098 8156 22918
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 8574 22400 8630 22409
rect 8574 22335 8630 22344
rect 8588 22098 8616 22335
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8128 21486 8156 22034
rect 8206 21992 8262 22001
rect 8206 21927 8208 21936
rect 8260 21927 8262 21936
rect 8208 21898 8260 21904
rect 8390 21584 8446 21593
rect 8390 21519 8392 21528
rect 8444 21519 8446 21528
rect 8392 21490 8444 21496
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8588 20466 8616 22034
rect 9140 21894 9168 22510
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 9232 21622 9260 22714
rect 9220 21616 9272 21622
rect 9220 21558 9272 21564
rect 9232 21078 9260 21558
rect 9220 21072 9272 21078
rect 9220 21014 9272 21020
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8208 19780 8260 19786
rect 8208 19722 8260 19728
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8220 18902 8248 19722
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8588 18630 8616 19246
rect 8680 18902 8708 19246
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 7932 18148 7984 18154
rect 7932 18090 7984 18096
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7944 17202 7972 18090
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15706 7144 15846
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 7300 15026 7328 16526
rect 7392 16454 7420 17002
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 16250 7420 16390
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7484 16114 7512 16934
rect 7944 16590 7972 17138
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 8128 16590 8156 16934
rect 8312 16590 8340 18022
rect 8404 16590 8432 18226
rect 8956 17626 8984 19722
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9416 19378 9444 19654
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 18290 9168 19246
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18902 9260 19110
rect 9220 18896 9272 18902
rect 9220 18838 9272 18844
rect 9324 18698 9352 19314
rect 9312 18692 9364 18698
rect 9312 18634 9364 18640
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9416 17762 9444 19314
rect 9508 19258 9536 24074
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 10060 23118 10088 24006
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10152 22030 10180 22374
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 9784 21690 9812 21966
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 10244 21010 10272 21966
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10336 19990 10364 27231
rect 10612 27010 10640 27270
rect 10520 26982 10640 27010
rect 10520 26466 10548 26982
rect 10520 26450 10640 26466
rect 10520 26444 10652 26450
rect 10520 26438 10600 26444
rect 10600 26386 10652 26392
rect 10704 26382 10732 30194
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11072 29850 11100 29990
rect 11060 29844 11112 29850
rect 11060 29786 11112 29792
rect 11060 29572 11112 29578
rect 11060 29514 11112 29520
rect 11072 29481 11100 29514
rect 11058 29472 11114 29481
rect 11058 29407 11114 29416
rect 11060 29096 11112 29102
rect 11060 29038 11112 29044
rect 10784 28960 10836 28966
rect 10784 28902 10836 28908
rect 10796 28558 10824 28902
rect 10968 28620 11020 28626
rect 10968 28562 11020 28568
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 10876 28416 10928 28422
rect 10876 28358 10928 28364
rect 10888 28121 10916 28358
rect 10980 28218 11008 28562
rect 11072 28218 11100 29038
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10874 28112 10930 28121
rect 11164 28098 11192 31311
rect 11256 31142 11284 33782
rect 11336 33652 11388 33658
rect 11336 33594 11388 33600
rect 11348 33454 11376 33594
rect 11336 33448 11388 33454
rect 11336 33390 11388 33396
rect 11440 32910 11468 34478
rect 11532 33522 11560 34886
rect 11612 33992 11664 33998
rect 11612 33934 11664 33940
rect 11624 33522 11652 33934
rect 11520 33516 11572 33522
rect 11520 33458 11572 33464
rect 11612 33516 11664 33522
rect 11612 33458 11664 33464
rect 11716 33402 11744 35090
rect 11808 34678 11836 35090
rect 11900 35086 11928 35498
rect 11888 35080 11940 35086
rect 11992 35068 12020 36638
rect 12084 36378 12112 36858
rect 12072 36372 12124 36378
rect 12072 36314 12124 36320
rect 12176 35222 12204 37606
rect 12268 36106 12296 38354
rect 12452 37942 12480 40054
rect 12728 38962 12756 41618
rect 14016 41614 14044 41686
rect 15016 41676 15068 41682
rect 15016 41618 15068 41624
rect 13452 41608 13504 41614
rect 13452 41550 13504 41556
rect 13544 41608 13596 41614
rect 14004 41608 14056 41614
rect 13596 41568 13860 41596
rect 13544 41550 13596 41556
rect 13464 41478 13492 41550
rect 13268 41472 13320 41478
rect 13268 41414 13320 41420
rect 13452 41472 13504 41478
rect 13452 41414 13504 41420
rect 13280 41154 13308 41414
rect 13464 41256 13492 41414
rect 13832 41274 13860 41568
rect 14004 41550 14056 41556
rect 15028 41274 15056 41618
rect 17500 41540 17552 41546
rect 17500 41482 17552 41488
rect 15108 41472 15160 41478
rect 15108 41414 15160 41420
rect 13820 41268 13872 41274
rect 13464 41228 13584 41256
rect 13280 41138 13492 41154
rect 13280 41132 13504 41138
rect 13280 41126 13452 41132
rect 13452 41074 13504 41080
rect 12808 41064 12860 41070
rect 12806 41032 12808 41041
rect 12992 41064 13044 41070
rect 12860 41032 12862 41041
rect 12992 41006 13044 41012
rect 12806 40967 12862 40976
rect 13004 39846 13032 41006
rect 13464 40594 13492 41074
rect 13452 40588 13504 40594
rect 13452 40530 13504 40536
rect 12992 39840 13044 39846
rect 12992 39782 13044 39788
rect 13358 39128 13414 39137
rect 13358 39063 13414 39072
rect 12716 38956 12768 38962
rect 12716 38898 12768 38904
rect 12992 38480 13044 38486
rect 12992 38422 13044 38428
rect 12440 37936 12492 37942
rect 12440 37878 12492 37884
rect 13004 37874 13032 38422
rect 13084 38004 13136 38010
rect 13084 37946 13136 37952
rect 13096 37874 13124 37946
rect 12992 37868 13044 37874
rect 12992 37810 13044 37816
rect 13084 37868 13136 37874
rect 13084 37810 13136 37816
rect 12440 37800 12492 37806
rect 12440 37742 12492 37748
rect 12256 36100 12308 36106
rect 12256 36042 12308 36048
rect 12348 36100 12400 36106
rect 12348 36042 12400 36048
rect 12360 35834 12388 36042
rect 12348 35828 12400 35834
rect 12348 35770 12400 35776
rect 12164 35216 12216 35222
rect 12164 35158 12216 35164
rect 12072 35080 12124 35086
rect 11992 35040 12072 35068
rect 11888 35022 11940 35028
rect 12124 35028 12204 35034
rect 12072 35022 12204 35028
rect 12084 35006 12204 35022
rect 12072 34944 12124 34950
rect 12072 34886 12124 34892
rect 11796 34672 11848 34678
rect 11796 34614 11848 34620
rect 11888 34604 11940 34610
rect 11888 34546 11940 34552
rect 11900 34066 11928 34546
rect 12084 34134 12112 34886
rect 12072 34128 12124 34134
rect 12072 34070 12124 34076
rect 11888 34060 11940 34066
rect 11888 34002 11940 34008
rect 11888 33924 11940 33930
rect 11888 33866 11940 33872
rect 11900 33658 11928 33866
rect 12072 33856 12124 33862
rect 11992 33816 12072 33844
rect 11888 33652 11940 33658
rect 11888 33594 11940 33600
rect 11624 33374 11744 33402
rect 11428 32904 11480 32910
rect 11428 32846 11480 32852
rect 11440 31142 11468 32846
rect 11624 32434 11652 33374
rect 11704 33312 11756 33318
rect 11704 33254 11756 33260
rect 11612 32428 11664 32434
rect 11612 32370 11664 32376
rect 11520 32224 11572 32230
rect 11520 32166 11572 32172
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11428 31136 11480 31142
rect 11428 31078 11480 31084
rect 11532 30920 11560 32166
rect 11612 31748 11664 31754
rect 11612 31690 11664 31696
rect 10874 28047 10930 28056
rect 11072 28070 11192 28098
rect 11256 30892 11560 30920
rect 10888 27946 10916 28047
rect 10876 27940 10928 27946
rect 10876 27882 10928 27888
rect 11072 27588 11100 28070
rect 11152 28008 11204 28014
rect 11152 27950 11204 27956
rect 10980 27560 11100 27588
rect 10784 27396 10836 27402
rect 10784 27338 10836 27344
rect 10796 26926 10824 27338
rect 10876 27056 10928 27062
rect 10876 26998 10928 27004
rect 10784 26920 10836 26926
rect 10784 26862 10836 26868
rect 10692 26376 10744 26382
rect 10692 26318 10744 26324
rect 10508 26308 10560 26314
rect 10508 26250 10560 26256
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 10428 23866 10456 25638
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 9588 19984 9640 19990
rect 9588 19926 9640 19932
rect 10048 19984 10100 19990
rect 10048 19926 10100 19932
rect 10324 19984 10376 19990
rect 10324 19926 10376 19932
rect 9600 19378 9628 19926
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9508 19230 9904 19258
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9508 17882 9536 18634
rect 9600 18290 9628 19110
rect 9876 18902 9904 19230
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9586 17776 9642 17785
rect 9416 17734 9536 17762
rect 9312 17672 9364 17678
rect 8956 17598 9168 17626
rect 9312 17614 9364 17620
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 8496 17066 8524 17206
rect 9048 17202 9076 17478
rect 9140 17202 9168 17598
rect 9324 17270 9352 17614
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8496 16590 8524 17002
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 16794 8708 16934
rect 8772 16794 8800 17138
rect 8864 17066 8892 17138
rect 8852 17060 8904 17066
rect 8852 17002 8904 17008
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7668 16250 7696 16390
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7576 16114 7604 16186
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7484 15978 7512 16050
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7484 15162 7512 15914
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 6736 15020 6788 15026
rect 6656 14980 6736 15008
rect 6656 14346 6684 14980
rect 6736 14962 6788 14968
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6828 14408 6880 14414
rect 6880 14356 6960 14362
rect 6828 14350 6960 14356
rect 6644 14340 6696 14346
rect 6840 14334 6960 14350
rect 7024 14346 7052 14758
rect 7300 14550 7328 14962
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 6644 14282 6696 14288
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 13530 6776 14214
rect 6932 13938 6960 14334
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6748 12850 6776 13194
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6656 12442 6684 12786
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 5736 12102 5764 12158
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 5644 11898 5672 12038
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 9994 5672 11086
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 9178 5488 9318
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5552 8090 5580 8298
rect 5736 8294 5764 12038
rect 6196 11014 6224 12038
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6104 8974 6132 10950
rect 6288 10062 6316 11834
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11150 6408 11494
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6472 9518 6500 12106
rect 6564 9994 6592 12174
rect 6656 11626 6684 12174
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6748 11558 6776 12786
rect 6840 12714 6868 13330
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6932 12850 6960 13126
rect 7392 12850 7420 13398
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6840 12102 6868 12650
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6840 10198 6868 11562
rect 7024 11121 7052 12786
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7484 11762 7512 12174
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7010 11112 7066 11121
rect 7010 11047 7066 11056
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5736 7954 5764 8230
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 6380 7886 6408 9318
rect 6748 8974 6776 10134
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6932 8974 6960 9930
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6564 8430 6592 8910
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7546 5764 7686
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 7002 5580 7142
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 5000 6254 5028 6326
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 3896 5370 3924 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 5000 5030 5028 6054
rect 5092 5710 5120 6802
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 6012 6322 6040 6666
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5092 5234 5120 5646
rect 6012 5642 6040 6258
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 5644 5370 5672 5578
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 6012 5302 6040 5578
rect 6472 5302 6500 6326
rect 7024 5710 7052 11047
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7116 9450 7144 10066
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7576 7818 7604 15642
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8036 14550 8064 14758
rect 8024 14544 8076 14550
rect 8024 14486 8076 14492
rect 8036 14414 8064 14486
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 7944 13870 7972 14350
rect 8128 13938 8156 15846
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8220 14278 8248 14894
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 8024 13320 8076 13326
rect 7944 13280 8024 13308
rect 7944 12850 7972 13280
rect 8024 13262 8076 13268
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12986 8064 13126
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7852 12753 7880 12786
rect 7838 12744 7894 12753
rect 7838 12679 7894 12688
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7852 11762 7880 12106
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 8128 11540 8156 13874
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8220 12050 8248 12378
rect 8312 12238 8340 16526
rect 8404 13258 8432 16526
rect 8864 15026 8892 17002
rect 9048 16182 9076 17138
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9140 15026 9168 17138
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9324 16794 9352 17070
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9416 16658 9444 17206
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9232 15162 9260 16050
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9416 15026 9444 16050
rect 8852 15020 8904 15026
rect 9128 15020 9180 15026
rect 8904 14980 9076 15008
rect 8852 14962 8904 14968
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8680 14618 8708 14758
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8944 14544 8996 14550
rect 8864 14492 8944 14498
rect 8864 14486 8996 14492
rect 9048 14498 9076 14980
rect 9128 14962 9180 14968
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9140 14618 9168 14962
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9324 14618 9352 14894
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 8864 14470 8984 14486
rect 9048 14470 9168 14498
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8496 14074 8524 14282
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8496 13954 8524 14010
rect 8496 13926 8616 13954
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8392 12640 8444 12646
rect 8496 12594 8524 13466
rect 8588 12986 8616 13926
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8588 12850 8616 12922
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8444 12588 8524 12594
rect 8392 12582 8524 12588
rect 8404 12566 8524 12582
rect 8496 12238 8524 12566
rect 8680 12442 8708 13806
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8300 12232 8352 12238
rect 8484 12232 8536 12238
rect 8352 12192 8432 12220
rect 8300 12174 8352 12180
rect 8404 12050 8432 12192
rect 8484 12174 8536 12180
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8220 12022 8340 12050
rect 8404 12022 8524 12050
rect 8312 11914 8340 12022
rect 8312 11886 8432 11914
rect 8404 11762 8432 11886
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8208 11552 8260 11558
rect 8128 11512 8208 11540
rect 8208 11494 8260 11500
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7760 9586 7788 9862
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 9042 7788 9522
rect 7944 9382 7972 10746
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8036 9654 8064 10406
rect 8128 10198 8156 10406
rect 8220 10198 8248 11494
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8312 10146 8340 11698
rect 8404 11218 8432 11698
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8496 10606 8524 12022
rect 8588 11898 8616 12174
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8404 10266 8432 10542
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 8128 9586 8156 10134
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7668 7818 7696 8774
rect 8220 8430 8248 10134
rect 8312 10118 8432 10146
rect 8404 9994 8432 10118
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8392 9988 8444 9994
rect 8444 9948 8524 9976
rect 8392 9930 8444 9936
rect 8312 9110 8340 9930
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8496 8906 8524 9948
rect 8588 9178 8616 10610
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7944 7750 7972 8230
rect 8680 7886 8708 12038
rect 8772 11898 8800 12922
rect 8864 12850 8892 14470
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8944 12844 8996 12850
rect 9048 12832 9076 14282
rect 9140 12850 9168 14470
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9232 14074 9260 14350
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 8996 12804 9076 12832
rect 9128 12844 9180 12850
rect 8944 12786 8996 12792
rect 9128 12786 9180 12792
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8864 10810 8892 12786
rect 8956 11558 8984 12786
rect 9034 12744 9090 12753
rect 9034 12679 9036 12688
rect 9088 12679 9090 12688
rect 9036 12650 9088 12656
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9324 12238 9352 12378
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9048 11898 9076 12038
rect 9140 11898 9168 12038
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8772 9654 8800 10610
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7116 7002 7144 7686
rect 8036 7478 8064 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7760 6798 7788 7346
rect 8128 7342 8156 7414
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5914 7420 6190
rect 7760 6118 7788 6734
rect 8128 6458 8156 7278
rect 9048 7002 9076 11290
rect 9140 10130 9168 11630
rect 9232 11626 9260 12038
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9416 11354 9444 14962
rect 9508 12442 9536 17734
rect 9586 17711 9588 17720
rect 9640 17711 9642 17720
rect 9588 17682 9640 17688
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 16658 9628 17138
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9600 16250 9628 16594
rect 9784 16590 9812 16934
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9968 15026 9996 19382
rect 10060 17678 10088 19926
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10152 17882 10180 19450
rect 10336 19378 10364 19790
rect 10428 19514 10456 23462
rect 10520 22642 10548 26250
rect 10888 25702 10916 26998
rect 10980 26314 11008 27560
rect 11060 26512 11112 26518
rect 11060 26454 11112 26460
rect 10968 26308 11020 26314
rect 10968 26250 11020 26256
rect 11072 26042 11100 26454
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 11164 25906 11192 27950
rect 11256 26790 11284 30892
rect 11428 30796 11480 30802
rect 11428 30738 11480 30744
rect 11336 30728 11388 30734
rect 11336 30670 11388 30676
rect 11348 30598 11376 30670
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 11348 29850 11376 30534
rect 11336 29844 11388 29850
rect 11336 29786 11388 29792
rect 11336 28416 11388 28422
rect 11336 28358 11388 28364
rect 11348 28218 11376 28358
rect 11336 28212 11388 28218
rect 11336 28154 11388 28160
rect 11440 27577 11468 30738
rect 11520 30184 11572 30190
rect 11520 30126 11572 30132
rect 11532 29714 11560 30126
rect 11624 30025 11652 31690
rect 11610 30016 11666 30025
rect 11610 29951 11666 29960
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 11520 28484 11572 28490
rect 11520 28426 11572 28432
rect 11532 28257 11560 28426
rect 11518 28248 11574 28257
rect 11518 28183 11574 28192
rect 11532 27878 11560 28183
rect 11610 27976 11666 27985
rect 11610 27911 11666 27920
rect 11520 27872 11572 27878
rect 11520 27814 11572 27820
rect 11426 27568 11482 27577
rect 11426 27503 11482 27512
rect 11624 27130 11652 27911
rect 11716 27130 11744 33254
rect 11794 32872 11850 32881
rect 11794 32807 11850 32816
rect 11808 32774 11836 32807
rect 11796 32768 11848 32774
rect 11796 32710 11848 32716
rect 11808 32065 11836 32710
rect 11886 32464 11942 32473
rect 11886 32399 11888 32408
rect 11940 32399 11942 32408
rect 11888 32370 11940 32376
rect 11888 32292 11940 32298
rect 11888 32234 11940 32240
rect 11794 32056 11850 32065
rect 11794 31991 11850 32000
rect 11900 31890 11928 32234
rect 11888 31884 11940 31890
rect 11888 31826 11940 31832
rect 11796 31136 11848 31142
rect 11796 31078 11848 31084
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11704 27124 11756 27130
rect 11704 27066 11756 27072
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11716 26450 11744 27066
rect 11704 26444 11756 26450
rect 11704 26386 11756 26392
rect 11428 26036 11480 26042
rect 11428 25978 11480 25984
rect 11152 25900 11204 25906
rect 11152 25842 11204 25848
rect 10876 25696 10928 25702
rect 10782 25664 10838 25673
rect 10876 25638 10928 25644
rect 10782 25599 10838 25608
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 10598 23760 10654 23769
rect 10598 23695 10654 23704
rect 10612 23662 10640 23695
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10612 23254 10640 23598
rect 10600 23248 10652 23254
rect 10600 23190 10652 23196
rect 10704 23118 10732 24006
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 10796 22574 10824 25599
rect 11164 25294 11192 25842
rect 11244 25832 11296 25838
rect 11244 25774 11296 25780
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 10968 24200 11020 24206
rect 11072 24177 11100 24686
rect 11256 24410 11284 25774
rect 11334 25256 11390 25265
rect 11334 25191 11390 25200
rect 11244 24404 11296 24410
rect 11244 24346 11296 24352
rect 11244 24200 11296 24206
rect 10968 24142 11020 24148
rect 11058 24168 11114 24177
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10520 20942 10548 21830
rect 10612 21690 10640 21966
rect 10796 21729 10824 22510
rect 10980 22166 11008 24142
rect 11244 24142 11296 24148
rect 11058 24103 11114 24112
rect 11256 23594 11284 24142
rect 11244 23588 11296 23594
rect 11244 23530 11296 23536
rect 11348 23526 11376 25191
rect 11440 24818 11468 25978
rect 11520 25288 11572 25294
rect 11520 25230 11572 25236
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11532 24954 11560 25230
rect 11520 24948 11572 24954
rect 11520 24890 11572 24896
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 11612 24676 11664 24682
rect 11612 24618 11664 24624
rect 11518 24440 11574 24449
rect 11440 24398 11518 24426
rect 11440 24206 11468 24398
rect 11518 24375 11574 24384
rect 11520 24336 11572 24342
rect 11520 24278 11572 24284
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11428 23316 11480 23322
rect 11428 23258 11480 23264
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10876 21956 10928 21962
rect 10876 21898 10928 21904
rect 10782 21720 10838 21729
rect 10600 21684 10652 21690
rect 10782 21655 10838 21664
rect 10600 21626 10652 21632
rect 10888 21554 10916 21898
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10612 21457 10640 21490
rect 10598 21448 10654 21457
rect 10598 21383 10654 21392
rect 10704 21146 10732 21490
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10520 19394 10548 20878
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10612 19514 10640 19858
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10324 19372 10376 19378
rect 10520 19366 10640 19394
rect 10324 19314 10376 19320
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10428 18698 10456 19110
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10506 18320 10562 18329
rect 10506 18255 10508 18264
rect 10560 18255 10562 18264
rect 10508 18226 10560 18232
rect 10612 18222 10640 19366
rect 10980 19310 11008 22102
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10600 18216 10652 18222
rect 10598 18184 10600 18193
rect 10652 18184 10654 18193
rect 10598 18119 10654 18128
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10060 17066 10088 17614
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10152 17338 10180 17546
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10796 15638 10824 16594
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 15026 10272 15302
rect 10796 15162 10824 15574
rect 10888 15570 10916 16390
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10888 15162 10916 15506
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 14074 9720 14214
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9600 12322 9628 12786
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9508 12294 9628 12322
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9232 9926 9260 11154
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9058 9260 9862
rect 9140 9042 9260 9058
rect 9324 9042 9352 10542
rect 9128 9036 9260 9042
rect 9180 9030 9260 9036
rect 9312 9036 9364 9042
rect 9128 8978 9180 8984
rect 9312 8978 9364 8984
rect 9416 8498 9444 10950
rect 9508 10062 9536 12294
rect 9600 12288 9628 12294
rect 9680 12300 9732 12306
rect 9600 12260 9680 12288
rect 9680 12242 9732 12248
rect 9588 12096 9640 12102
rect 9784 12084 9812 12718
rect 9640 12056 9812 12084
rect 9588 12038 9640 12044
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10810 9628 10950
rect 9876 10810 9904 14758
rect 10428 14482 10456 15098
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10612 14278 10640 14758
rect 10704 14618 10732 14758
rect 10888 14618 10916 14962
rect 10980 14822 11008 18566
rect 11072 18358 11100 22918
rect 11440 22817 11468 23258
rect 11426 22808 11482 22817
rect 11426 22743 11482 22752
rect 11440 22094 11468 22743
rect 11348 22066 11468 22094
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 21690 11284 21830
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10796 12986 10824 14418
rect 10980 13530 11008 14758
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10266 9628 10406
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9600 10062 9628 10202
rect 9496 10056 9548 10062
rect 9494 10024 9496 10033
rect 9588 10056 9640 10062
rect 9548 10024 9550 10033
rect 9588 9998 9640 10004
rect 9494 9959 9550 9968
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9508 8430 9536 8978
rect 9600 8974 9628 9998
rect 9876 9586 9904 10746
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7206 9536 7686
rect 9692 7546 9720 8366
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9586 6760 9642 6769
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7760 5778 7788 6054
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 6748 5030 6776 5510
rect 8404 5370 8432 6122
rect 8864 6118 8892 6734
rect 9968 6730 9996 11018
rect 10060 8634 10088 12650
rect 10796 12442 10824 12786
rect 11072 12782 11100 16050
rect 11164 15994 11192 20878
rect 11348 19802 11376 22066
rect 11532 22030 11560 24278
rect 11624 24206 11652 24618
rect 11716 24410 11744 25230
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 11808 24290 11836 31078
rect 11992 30376 12020 33816
rect 12072 33798 12124 33804
rect 12176 33674 12204 35006
rect 12348 34128 12400 34134
rect 12084 33646 12204 33674
rect 12268 34088 12348 34116
rect 12084 33590 12112 33646
rect 12072 33584 12124 33590
rect 12072 33526 12124 33532
rect 11900 30348 12020 30376
rect 11900 30258 11928 30348
rect 12084 30308 12112 33526
rect 12164 32768 12216 32774
rect 12164 32710 12216 32716
rect 12176 32434 12204 32710
rect 12164 32428 12216 32434
rect 12164 32370 12216 32376
rect 12268 32314 12296 34088
rect 12348 34070 12400 34076
rect 12348 33312 12400 33318
rect 12348 33254 12400 33260
rect 11992 30280 12112 30308
rect 12176 32286 12296 32314
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11900 29306 11928 29990
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11888 28552 11940 28558
rect 11992 28540 12020 30280
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 12084 28994 12112 30126
rect 12176 29322 12204 32286
rect 12256 32224 12308 32230
rect 12256 32166 12308 32172
rect 12268 32026 12296 32166
rect 12360 32026 12388 33254
rect 12452 32774 12480 37742
rect 12532 37392 12584 37398
rect 12532 37334 12584 37340
rect 12900 37392 12952 37398
rect 12900 37334 12952 37340
rect 12544 36854 12572 37334
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 12532 36848 12584 36854
rect 12532 36790 12584 36796
rect 12728 36310 12756 37062
rect 12716 36304 12768 36310
rect 12716 36246 12768 36252
rect 12808 36032 12860 36038
rect 12808 35974 12860 35980
rect 12820 35766 12848 35974
rect 12808 35760 12860 35766
rect 12808 35702 12860 35708
rect 12624 35488 12676 35494
rect 12624 35430 12676 35436
rect 12716 35488 12768 35494
rect 12716 35430 12768 35436
rect 12636 35086 12664 35430
rect 12624 35080 12676 35086
rect 12624 35022 12676 35028
rect 12728 34610 12756 35430
rect 12808 35012 12860 35018
rect 12808 34954 12860 34960
rect 12716 34604 12768 34610
rect 12716 34546 12768 34552
rect 12624 34400 12676 34406
rect 12624 34342 12676 34348
rect 12636 33658 12664 34342
rect 12728 33862 12756 34546
rect 12716 33856 12768 33862
rect 12716 33798 12768 33804
rect 12624 33652 12676 33658
rect 12624 33594 12676 33600
rect 12532 33448 12584 33454
rect 12530 33416 12532 33425
rect 12584 33416 12586 33425
rect 12530 33351 12586 33360
rect 12440 32768 12492 32774
rect 12440 32710 12492 32716
rect 12530 32736 12586 32745
rect 12256 32020 12308 32026
rect 12256 31962 12308 31968
rect 12348 32020 12400 32026
rect 12348 31962 12400 31968
rect 12360 31906 12388 31962
rect 12268 31878 12388 31906
rect 12268 31210 12296 31878
rect 12256 31204 12308 31210
rect 12256 31146 12308 31152
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 12360 30938 12388 31078
rect 12348 30932 12400 30938
rect 12348 30874 12400 30880
rect 12256 30320 12308 30326
rect 12256 30262 12308 30268
rect 12268 29850 12296 30262
rect 12256 29844 12308 29850
rect 12256 29786 12308 29792
rect 12452 29646 12480 32710
rect 12530 32671 12586 32680
rect 12544 32570 12572 32671
rect 12532 32564 12584 32570
rect 12532 32506 12584 32512
rect 12532 32428 12584 32434
rect 12532 32370 12584 32376
rect 12544 32201 12572 32370
rect 12530 32192 12586 32201
rect 12530 32127 12586 32136
rect 12636 31906 12664 33594
rect 12544 31878 12664 31906
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 12440 29504 12492 29510
rect 12438 29472 12440 29481
rect 12492 29472 12494 29481
rect 12438 29407 12494 29416
rect 12176 29294 12480 29322
rect 12084 28966 12204 28994
rect 12176 28801 12204 28966
rect 12162 28792 12218 28801
rect 12162 28727 12218 28736
rect 12256 28756 12308 28762
rect 12256 28698 12308 28704
rect 11940 28512 12020 28540
rect 12164 28552 12216 28558
rect 11888 28494 11940 28500
rect 12268 28540 12296 28698
rect 12216 28512 12296 28540
rect 12164 28494 12216 28500
rect 12072 28484 12124 28490
rect 12072 28426 12124 28432
rect 11888 27668 11940 27674
rect 11888 27610 11940 27616
rect 11900 27130 11928 27610
rect 11888 27124 11940 27130
rect 11888 27066 11940 27072
rect 12084 26994 12112 28426
rect 12176 27402 12204 28494
rect 12452 28422 12480 29294
rect 12544 28558 12572 31878
rect 12624 31680 12676 31686
rect 12624 31622 12676 31628
rect 12636 31346 12664 31622
rect 12728 31346 12756 33798
rect 12624 31340 12676 31346
rect 12624 31282 12676 31288
rect 12716 31340 12768 31346
rect 12716 31282 12768 31288
rect 12624 31204 12676 31210
rect 12624 31146 12676 31152
rect 12636 29073 12664 31146
rect 12728 30938 12756 31282
rect 12716 30932 12768 30938
rect 12716 30874 12768 30880
rect 12820 30734 12848 34954
rect 12912 34649 12940 37334
rect 13004 37126 13032 37810
rect 13096 37262 13124 37810
rect 13084 37256 13136 37262
rect 13084 37198 13136 37204
rect 12992 37120 13044 37126
rect 12992 37062 13044 37068
rect 13176 37120 13228 37126
rect 13176 37062 13228 37068
rect 12992 35760 13044 35766
rect 12992 35702 13044 35708
rect 13004 35562 13032 35702
rect 12992 35556 13044 35562
rect 12992 35498 13044 35504
rect 13188 35290 13216 37062
rect 13372 36922 13400 39063
rect 13556 39030 13584 41228
rect 13820 41210 13872 41216
rect 15016 41268 15068 41274
rect 15016 41210 15068 41216
rect 14740 41064 14792 41070
rect 14740 41006 14792 41012
rect 14752 40730 14780 41006
rect 14740 40724 14792 40730
rect 14740 40666 14792 40672
rect 15120 40526 15148 41414
rect 15660 41268 15712 41274
rect 15660 41210 15712 41216
rect 15672 41138 15700 41210
rect 17316 41200 17368 41206
rect 17368 41160 17448 41188
rect 17316 41142 17368 41148
rect 15384 41132 15436 41138
rect 15384 41074 15436 41080
rect 15660 41132 15712 41138
rect 15660 41074 15712 41080
rect 15752 41132 15804 41138
rect 15752 41074 15804 41080
rect 16764 41132 16816 41138
rect 16764 41074 16816 41080
rect 17132 41132 17184 41138
rect 17132 41074 17184 41080
rect 15200 40928 15252 40934
rect 15200 40870 15252 40876
rect 15212 40662 15240 40870
rect 15200 40656 15252 40662
rect 15200 40598 15252 40604
rect 14556 40520 14608 40526
rect 14556 40462 14608 40468
rect 15108 40520 15160 40526
rect 15108 40462 15160 40468
rect 13728 40384 13780 40390
rect 13728 40326 13780 40332
rect 14188 40384 14240 40390
rect 14188 40326 14240 40332
rect 14464 40384 14516 40390
rect 14464 40326 14516 40332
rect 13740 40186 13768 40326
rect 13728 40180 13780 40186
rect 13728 40122 13780 40128
rect 13636 39840 13688 39846
rect 13636 39782 13688 39788
rect 13648 39098 13676 39782
rect 13636 39092 13688 39098
rect 13636 39034 13688 39040
rect 13544 39024 13596 39030
rect 13464 38984 13544 39012
rect 13464 38350 13492 38984
rect 13544 38966 13596 38972
rect 13452 38344 13504 38350
rect 13452 38286 13504 38292
rect 13464 36922 13492 38286
rect 13544 38276 13596 38282
rect 13544 38218 13596 38224
rect 13556 37806 13584 38218
rect 13636 37868 13688 37874
rect 13636 37810 13688 37816
rect 13544 37800 13596 37806
rect 13544 37742 13596 37748
rect 13648 37194 13676 37810
rect 13636 37188 13688 37194
rect 13636 37130 13688 37136
rect 13360 36916 13412 36922
rect 13360 36858 13412 36864
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 14200 36106 14228 40326
rect 14476 40186 14504 40326
rect 14464 40180 14516 40186
rect 14464 40122 14516 40128
rect 14372 40044 14424 40050
rect 14372 39986 14424 39992
rect 14384 39642 14412 39986
rect 14372 39636 14424 39642
rect 14372 39578 14424 39584
rect 14568 39506 14596 40462
rect 15106 40216 15162 40225
rect 15106 40151 15108 40160
rect 15160 40151 15162 40160
rect 15108 40122 15160 40128
rect 15106 40080 15162 40089
rect 15162 40038 15332 40066
rect 15106 40015 15108 40024
rect 15160 40015 15162 40024
rect 15108 39986 15160 39992
rect 15200 39908 15252 39914
rect 15200 39850 15252 39856
rect 14556 39500 14608 39506
rect 14556 39442 14608 39448
rect 14568 39098 14596 39442
rect 14556 39092 14608 39098
rect 14556 39034 14608 39040
rect 14278 38040 14334 38049
rect 14278 37975 14334 37984
rect 14292 37942 14320 37975
rect 14280 37936 14332 37942
rect 14280 37878 14332 37884
rect 15016 37868 15068 37874
rect 15016 37810 15068 37816
rect 15028 37262 15056 37810
rect 15016 37256 15068 37262
rect 15016 37198 15068 37204
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 14292 36854 14320 37062
rect 14280 36848 14332 36854
rect 14280 36790 14332 36796
rect 15028 36582 15056 37062
rect 15212 36922 15240 39850
rect 15304 39642 15332 40038
rect 15396 39846 15424 41074
rect 15672 40662 15700 41074
rect 15764 40934 15792 41074
rect 16210 41032 16266 41041
rect 16210 40967 16212 40976
rect 16264 40967 16266 40976
rect 16212 40938 16264 40944
rect 15752 40928 15804 40934
rect 15752 40870 15804 40876
rect 16672 40928 16724 40934
rect 16672 40870 16724 40876
rect 15660 40656 15712 40662
rect 15660 40598 15712 40604
rect 15476 40588 15528 40594
rect 15476 40530 15528 40536
rect 15488 40390 15516 40530
rect 15568 40452 15620 40458
rect 15568 40394 15620 40400
rect 15476 40384 15528 40390
rect 15476 40326 15528 40332
rect 15580 39982 15608 40394
rect 15568 39976 15620 39982
rect 15568 39918 15620 39924
rect 15384 39840 15436 39846
rect 15384 39782 15436 39788
rect 15292 39636 15344 39642
rect 15292 39578 15344 39584
rect 15292 39296 15344 39302
rect 15292 39238 15344 39244
rect 15304 38894 15332 39238
rect 15292 38888 15344 38894
rect 15292 38830 15344 38836
rect 15304 37369 15332 38830
rect 15396 37806 15424 39782
rect 15580 39302 15608 39918
rect 15660 39636 15712 39642
rect 15660 39578 15712 39584
rect 15568 39296 15620 39302
rect 15568 39238 15620 39244
rect 15672 38298 15700 39578
rect 15764 38654 15792 40870
rect 16578 40760 16634 40769
rect 16578 40695 16634 40704
rect 16592 40662 16620 40695
rect 16580 40656 16632 40662
rect 16580 40598 16632 40604
rect 15936 40520 15988 40526
rect 16028 40520 16080 40526
rect 15936 40462 15988 40468
rect 16026 40488 16028 40497
rect 16580 40520 16632 40526
rect 16080 40488 16082 40497
rect 15844 40384 15896 40390
rect 15844 40326 15896 40332
rect 15856 39982 15884 40326
rect 15948 40186 15976 40462
rect 16684 40474 16712 40870
rect 16776 40662 16804 41074
rect 17144 41041 17172 41074
rect 17316 41064 17368 41070
rect 17130 41032 17186 41041
rect 16960 40990 17130 41018
rect 16764 40656 16816 40662
rect 16764 40598 16816 40604
rect 16960 40594 16988 40990
rect 17316 41006 17368 41012
rect 17130 40967 17186 40976
rect 17222 40896 17278 40905
rect 17144 40854 17222 40882
rect 17144 40610 17172 40854
rect 17222 40831 17278 40840
rect 17328 40730 17356 41006
rect 17316 40724 17368 40730
rect 17316 40666 17368 40672
rect 17052 40594 17172 40610
rect 16948 40588 17000 40594
rect 16948 40530 17000 40536
rect 17052 40588 17184 40594
rect 17052 40582 17132 40588
rect 16632 40468 16712 40474
rect 16580 40462 16712 40468
rect 16026 40423 16082 40432
rect 16488 40452 16540 40458
rect 15936 40180 15988 40186
rect 15936 40122 15988 40128
rect 15948 40050 15976 40122
rect 15936 40044 15988 40050
rect 15936 39986 15988 39992
rect 15844 39976 15896 39982
rect 15844 39918 15896 39924
rect 15856 39506 15884 39918
rect 15948 39658 15976 39986
rect 16040 39914 16068 40423
rect 16592 40446 16712 40462
rect 16488 40394 16540 40400
rect 16500 40361 16528 40394
rect 16486 40352 16542 40361
rect 16486 40287 16542 40296
rect 16120 40180 16172 40186
rect 16120 40122 16172 40128
rect 16028 39908 16080 39914
rect 16028 39850 16080 39856
rect 15948 39630 16068 39658
rect 15936 39568 15988 39574
rect 15936 39510 15988 39516
rect 15844 39500 15896 39506
rect 15844 39442 15896 39448
rect 15764 38626 15884 38654
rect 15672 38270 15792 38298
rect 15764 38214 15792 38270
rect 15568 38208 15620 38214
rect 15568 38150 15620 38156
rect 15660 38208 15712 38214
rect 15660 38150 15712 38156
rect 15752 38208 15804 38214
rect 15752 38150 15804 38156
rect 15580 37874 15608 38150
rect 15672 37942 15700 38150
rect 15660 37936 15712 37942
rect 15660 37878 15712 37884
rect 15568 37868 15620 37874
rect 15568 37810 15620 37816
rect 15384 37800 15436 37806
rect 15764 37754 15792 38150
rect 15856 37806 15884 38626
rect 15948 38418 15976 39510
rect 15936 38412 15988 38418
rect 15936 38354 15988 38360
rect 16040 37874 16068 39630
rect 16132 38049 16160 40122
rect 16212 39908 16264 39914
rect 16212 39850 16264 39856
rect 16224 39438 16252 39850
rect 16500 39642 16528 40287
rect 16762 40216 16818 40225
rect 16762 40151 16818 40160
rect 16580 40112 16632 40118
rect 16580 40054 16632 40060
rect 16592 39642 16620 40054
rect 16488 39636 16540 39642
rect 16488 39578 16540 39584
rect 16580 39636 16632 39642
rect 16580 39578 16632 39584
rect 16304 39500 16356 39506
rect 16304 39442 16356 39448
rect 16580 39500 16632 39506
rect 16580 39442 16632 39448
rect 16212 39432 16264 39438
rect 16212 39374 16264 39380
rect 16118 38040 16174 38049
rect 16118 37975 16174 37984
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 16120 37868 16172 37874
rect 16120 37810 16172 37816
rect 15384 37742 15436 37748
rect 15290 37360 15346 37369
rect 15290 37295 15346 37304
rect 15304 37262 15332 37295
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 15396 37126 15424 37742
rect 15672 37726 15792 37754
rect 15844 37800 15896 37806
rect 15844 37742 15896 37748
rect 15476 37664 15528 37670
rect 15476 37606 15528 37612
rect 15488 37330 15516 37606
rect 15476 37324 15528 37330
rect 15476 37266 15528 37272
rect 15672 37194 15700 37726
rect 15752 37664 15804 37670
rect 15752 37606 15804 37612
rect 15764 37466 15792 37606
rect 15752 37460 15804 37466
rect 15752 37402 15804 37408
rect 16040 37262 16068 37810
rect 16132 37369 16160 37810
rect 16316 37806 16344 39442
rect 16396 39432 16448 39438
rect 16396 39374 16448 39380
rect 16408 37874 16436 39374
rect 16488 39296 16540 39302
rect 16488 39238 16540 39244
rect 16500 39098 16528 39238
rect 16488 39092 16540 39098
rect 16488 39034 16540 39040
rect 16500 38214 16528 39034
rect 16592 38214 16620 39442
rect 16776 38214 16804 40151
rect 16948 40112 17000 40118
rect 16946 40080 16948 40089
rect 17000 40080 17002 40089
rect 16946 40015 17002 40024
rect 17052 38654 17080 40582
rect 17132 40530 17184 40536
rect 17132 40452 17184 40458
rect 17132 40394 17184 40400
rect 17144 40186 17172 40394
rect 17420 40390 17448 41160
rect 17512 41070 17540 41482
rect 17592 41132 17644 41138
rect 17592 41074 17644 41080
rect 17500 41064 17552 41070
rect 17500 41006 17552 41012
rect 17316 40384 17368 40390
rect 17316 40326 17368 40332
rect 17408 40384 17460 40390
rect 17408 40326 17460 40332
rect 17328 40186 17356 40326
rect 17132 40180 17184 40186
rect 17132 40122 17184 40128
rect 17316 40180 17368 40186
rect 17604 40168 17632 41074
rect 17788 40526 17816 41754
rect 19444 41750 19472 41783
rect 19432 41744 19484 41750
rect 18970 41712 19026 41721
rect 18696 41676 18748 41682
rect 20260 41744 20312 41750
rect 19432 41686 19484 41692
rect 19904 41682 20208 41698
rect 20732 41721 20760 41958
rect 20260 41686 20312 41692
rect 20718 41712 20774 41721
rect 18970 41647 19026 41656
rect 19064 41676 19116 41682
rect 18696 41618 18748 41624
rect 17960 41472 18012 41478
rect 17960 41414 18012 41420
rect 17972 41138 18000 41414
rect 18052 41200 18104 41206
rect 18328 41200 18380 41206
rect 18104 41148 18184 41154
rect 18052 41142 18184 41148
rect 18328 41142 18380 41148
rect 18418 41168 18474 41177
rect 17868 41132 17920 41138
rect 17868 41074 17920 41080
rect 17960 41132 18012 41138
rect 18064 41126 18184 41142
rect 17960 41074 18012 41080
rect 17880 40594 17908 41074
rect 17868 40588 17920 40594
rect 17868 40530 17920 40536
rect 17776 40520 17828 40526
rect 17316 40122 17368 40128
rect 17512 40140 17632 40168
rect 17696 40480 17776 40508
rect 17512 39914 17540 40140
rect 17696 40089 17724 40480
rect 17776 40462 17828 40468
rect 17776 40384 17828 40390
rect 17776 40326 17828 40332
rect 17682 40080 17738 40089
rect 17592 40044 17644 40050
rect 17682 40015 17738 40024
rect 17592 39986 17644 39992
rect 17500 39908 17552 39914
rect 17500 39850 17552 39856
rect 16960 38626 17080 38654
rect 17512 38654 17540 39850
rect 17604 39846 17632 39986
rect 17592 39840 17644 39846
rect 17592 39782 17644 39788
rect 17604 39506 17632 39782
rect 17684 39568 17736 39574
rect 17684 39510 17736 39516
rect 17592 39500 17644 39506
rect 17592 39442 17644 39448
rect 17592 38752 17644 38758
rect 17592 38694 17644 38700
rect 17604 38654 17632 38694
rect 17512 38626 17632 38654
rect 16488 38208 16540 38214
rect 16488 38150 16540 38156
rect 16580 38208 16632 38214
rect 16580 38150 16632 38156
rect 16672 38208 16724 38214
rect 16672 38150 16724 38156
rect 16764 38208 16816 38214
rect 16764 38150 16816 38156
rect 16396 37868 16448 37874
rect 16396 37810 16448 37816
rect 16304 37800 16356 37806
rect 16304 37742 16356 37748
rect 16316 37466 16344 37742
rect 16304 37460 16356 37466
rect 16304 37402 16356 37408
rect 16118 37360 16174 37369
rect 16118 37295 16174 37304
rect 15752 37256 15804 37262
rect 15752 37198 15804 37204
rect 15936 37256 15988 37262
rect 15936 37198 15988 37204
rect 16028 37256 16080 37262
rect 16028 37198 16080 37204
rect 15660 37188 15712 37194
rect 15660 37130 15712 37136
rect 15384 37120 15436 37126
rect 15384 37062 15436 37068
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15764 36854 15792 37198
rect 15948 37097 15976 37198
rect 15934 37088 15990 37097
rect 15934 37023 15990 37032
rect 16212 36916 16264 36922
rect 16212 36858 16264 36864
rect 15752 36848 15804 36854
rect 15752 36790 15804 36796
rect 15384 36780 15436 36786
rect 15384 36722 15436 36728
rect 15396 36689 15424 36722
rect 15382 36680 15438 36689
rect 15382 36615 15438 36624
rect 15016 36576 15068 36582
rect 15016 36518 15068 36524
rect 15028 36106 15056 36518
rect 16224 36281 16252 36858
rect 16316 36718 16344 37402
rect 16408 36854 16436 37810
rect 16592 37482 16620 38150
rect 16684 37806 16712 38150
rect 16960 37874 16988 38626
rect 17224 38344 17276 38350
rect 17224 38286 17276 38292
rect 17236 38010 17264 38286
rect 17224 38004 17276 38010
rect 17224 37946 17276 37952
rect 16948 37868 17000 37874
rect 16948 37810 17000 37816
rect 16672 37800 16724 37806
rect 16672 37742 16724 37748
rect 16500 37454 16620 37482
rect 16500 37330 16528 37454
rect 16488 37324 16540 37330
rect 16488 37266 16540 37272
rect 16580 37256 16632 37262
rect 16580 37198 16632 37204
rect 16396 36848 16448 36854
rect 16396 36790 16448 36796
rect 16592 36786 16620 37198
rect 16488 36780 16540 36786
rect 16488 36722 16540 36728
rect 16580 36780 16632 36786
rect 16580 36722 16632 36728
rect 16304 36712 16356 36718
rect 16304 36654 16356 36660
rect 16500 36378 16528 36722
rect 16592 36417 16620 36722
rect 16684 36582 16712 37742
rect 16762 36816 16818 36825
rect 16762 36751 16764 36760
rect 16816 36751 16818 36760
rect 16764 36722 16816 36728
rect 16776 36650 16804 36722
rect 16764 36644 16816 36650
rect 16764 36586 16816 36592
rect 16672 36576 16724 36582
rect 16672 36518 16724 36524
rect 16578 36408 16634 36417
rect 16488 36372 16540 36378
rect 16578 36343 16634 36352
rect 16488 36314 16540 36320
rect 16210 36272 16266 36281
rect 16210 36207 16266 36216
rect 15844 36168 15896 36174
rect 15844 36110 15896 36116
rect 14188 36100 14240 36106
rect 14188 36042 14240 36048
rect 15016 36100 15068 36106
rect 15016 36042 15068 36048
rect 13542 36000 13598 36009
rect 13542 35935 13598 35944
rect 13360 35488 13412 35494
rect 13360 35430 13412 35436
rect 13176 35284 13228 35290
rect 13176 35226 13228 35232
rect 13268 35284 13320 35290
rect 13268 35226 13320 35232
rect 13280 35086 13308 35226
rect 13268 35080 13320 35086
rect 13174 35048 13230 35057
rect 13268 35022 13320 35028
rect 13174 34983 13176 34992
rect 13228 34983 13230 34992
rect 13176 34954 13228 34960
rect 13176 34672 13228 34678
rect 12898 34640 12954 34649
rect 13176 34614 13228 34620
rect 12898 34575 12954 34584
rect 12992 33992 13044 33998
rect 12992 33934 13044 33940
rect 13004 33289 13032 33934
rect 12990 33280 13046 33289
rect 12990 33215 13046 33224
rect 12900 32836 12952 32842
rect 12900 32778 12952 32784
rect 12912 32570 12940 32778
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 12900 32428 12952 32434
rect 12952 32388 13032 32416
rect 12900 32370 12952 32376
rect 12898 31920 12954 31929
rect 12898 31855 12954 31864
rect 12912 31822 12940 31855
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 12820 30258 12848 30670
rect 12808 30252 12860 30258
rect 12808 30194 12860 30200
rect 12622 29064 12678 29073
rect 12622 28999 12678 29008
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12348 28416 12400 28422
rect 12254 28384 12310 28393
rect 12348 28358 12400 28364
rect 12440 28416 12492 28422
rect 12440 28358 12492 28364
rect 12254 28319 12310 28328
rect 12268 27674 12296 28319
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 12164 27396 12216 27402
rect 12164 27338 12216 27344
rect 12072 26988 12124 26994
rect 11900 26948 12072 26976
rect 11900 25226 11928 26948
rect 12072 26930 12124 26936
rect 12164 26852 12216 26858
rect 12164 26794 12216 26800
rect 11980 26784 12032 26790
rect 12176 26761 12204 26794
rect 11980 26726 12032 26732
rect 12162 26752 12218 26761
rect 11888 25220 11940 25226
rect 11888 25162 11940 25168
rect 11716 24262 11836 24290
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11716 23322 11744 24262
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11808 23730 11836 24142
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11808 22778 11836 23666
rect 11900 22982 11928 25162
rect 11992 24698 12020 26726
rect 12162 26687 12218 26696
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 12176 25770 12204 26250
rect 12164 25764 12216 25770
rect 12164 25706 12216 25712
rect 12176 24954 12204 25706
rect 12256 25152 12308 25158
rect 12256 25094 12308 25100
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 11992 24670 12204 24698
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 11992 24206 12020 24550
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11992 23730 12020 24006
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11900 22778 11928 22918
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11520 22024 11572 22030
rect 11572 21984 11652 22012
rect 11520 21966 11572 21972
rect 11428 21888 11480 21894
rect 11426 21856 11428 21865
rect 11520 21888 11572 21894
rect 11480 21856 11482 21865
rect 11520 21830 11572 21836
rect 11426 21791 11482 21800
rect 11532 21146 11560 21830
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11426 19952 11482 19961
rect 11426 19887 11482 19896
rect 11256 19786 11376 19802
rect 11440 19786 11468 19887
rect 11244 19780 11376 19786
rect 11296 19774 11376 19780
rect 11244 19722 11296 19728
rect 11348 19446 11376 19774
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11336 19440 11388 19446
rect 11336 19382 11388 19388
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11256 16561 11284 18362
rect 11348 18290 11376 19110
rect 11532 18970 11560 21082
rect 11624 19990 11652 21984
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 12084 21622 12112 21830
rect 12072 21616 12124 21622
rect 12072 21558 12124 21564
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 12084 20942 12112 21286
rect 12176 21010 12204 24670
rect 12268 21010 12296 25094
rect 12360 21962 12388 28358
rect 12452 28082 12480 28358
rect 12532 28144 12584 28150
rect 12530 28112 12532 28121
rect 12584 28112 12586 28121
rect 12440 28076 12492 28082
rect 12530 28047 12586 28056
rect 12440 28018 12492 28024
rect 12532 28008 12584 28014
rect 12532 27950 12584 27956
rect 12544 27674 12572 27950
rect 12532 27668 12584 27674
rect 12532 27610 12584 27616
rect 12440 27600 12492 27606
rect 12440 27542 12492 27548
rect 12452 27130 12480 27542
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12544 26858 12572 27338
rect 12532 26852 12584 26858
rect 12532 26794 12584 26800
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12452 24818 12480 25638
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12544 24886 12572 25094
rect 12532 24880 12584 24886
rect 12532 24822 12584 24828
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12532 24744 12584 24750
rect 12530 24712 12532 24721
rect 12584 24712 12586 24721
rect 12530 24647 12586 24656
rect 12532 24336 12584 24342
rect 12532 24278 12584 24284
rect 12544 23905 12572 24278
rect 12530 23896 12586 23905
rect 12452 23854 12530 23882
rect 12452 23186 12480 23854
rect 12530 23831 12586 23840
rect 12636 23730 12664 28999
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12728 26489 12756 26998
rect 12714 26480 12770 26489
rect 12714 26415 12770 26424
rect 12716 25832 12768 25838
rect 12716 25774 12768 25780
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22778 12480 23122
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12544 22094 12572 23462
rect 12728 22545 12756 25774
rect 12714 22536 12770 22545
rect 12624 22500 12676 22506
rect 12714 22471 12770 22480
rect 12624 22442 12676 22448
rect 12636 22098 12664 22442
rect 12452 22066 12572 22094
rect 12624 22092 12676 22098
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 11612 19984 11664 19990
rect 11612 19926 11664 19932
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11808 19242 11836 19722
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11520 18964 11572 18970
rect 11520 18906 11572 18912
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11242 16552 11298 16561
rect 11242 16487 11298 16496
rect 11348 16114 11376 18022
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11532 17270 11560 17750
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11624 17338 11652 17614
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11520 17264 11572 17270
rect 11520 17206 11572 17212
rect 11716 17082 11744 17614
rect 11532 17054 11744 17082
rect 11532 16726 11560 17054
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11440 16153 11468 16526
rect 11426 16144 11482 16153
rect 11336 16108 11388 16114
rect 11426 16079 11428 16088
rect 11336 16050 11388 16056
rect 11480 16079 11482 16088
rect 11428 16050 11480 16056
rect 11164 15966 11376 15994
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11164 15026 11192 15302
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11256 13870 11284 15438
rect 11348 15094 11376 15966
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 13938 11376 14350
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11440 12986 11468 14282
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10508 12232 10560 12238
rect 10600 12232 10652 12238
rect 10508 12174 10560 12180
rect 10598 12200 10600 12209
rect 10652 12200 10654 12209
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10336 11898 10364 12038
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10520 11694 10548 12174
rect 10598 12135 10654 12144
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10888 11354 10916 11698
rect 11072 11694 11100 12718
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11072 10674 11100 11630
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10796 9722 10824 10610
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10980 9926 11008 10474
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10198 11376 10406
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11348 10062 11376 10134
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11336 10056 11388 10062
rect 11428 10056 11480 10062
rect 11336 9998 11388 10004
rect 11426 10024 11428 10033
rect 11480 10024 11482 10033
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 10060 7886 10088 8298
rect 10244 7886 10272 8774
rect 10520 8650 10548 9590
rect 10980 9178 11008 9862
rect 11164 9722 11192 9998
rect 11426 9959 11482 9968
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10428 8634 10548 8650
rect 10416 8628 10548 8634
rect 10468 8622 10548 8628
rect 10416 8570 10468 8576
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10152 7546 10180 7686
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 9586 6695 9642 6704
rect 9956 6724 10008 6730
rect 9600 6662 9628 6695
rect 9956 6666 10008 6672
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9600 6322 9628 6598
rect 9784 6458 9812 6598
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 952 3398 980 3431
rect 940 3392 992 3398
rect 940 3334 992 3340
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 3896 2366 4016 2394
rect 5000 2378 5028 4966
rect 5552 3534 5580 4966
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 8864 2446 8892 6054
rect 8956 5914 8984 6054
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 10612 5778 10640 8366
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11348 7206 11376 7822
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11532 6914 11560 16662
rect 11716 16590 11744 16934
rect 11808 16590 11836 17682
rect 11900 17354 11928 19110
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 18426 12020 18566
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 12084 17814 12112 20878
rect 12176 20466 12204 20946
rect 12268 20466 12296 20946
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12346 20088 12402 20097
rect 12346 20023 12402 20032
rect 12360 19446 12388 20023
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12452 18766 12480 22066
rect 12820 22094 12848 30194
rect 12912 29764 12940 31282
rect 13004 30258 13032 32388
rect 13082 32328 13138 32337
rect 13188 32298 13216 34614
rect 13372 34610 13400 35430
rect 13360 34604 13412 34610
rect 13360 34546 13412 34552
rect 13452 34400 13504 34406
rect 13452 34342 13504 34348
rect 13464 33436 13492 34342
rect 13556 33833 13584 35935
rect 14004 35828 14056 35834
rect 14004 35770 14056 35776
rect 15200 35828 15252 35834
rect 15200 35770 15252 35776
rect 13912 35556 13964 35562
rect 13912 35498 13964 35504
rect 13924 35086 13952 35498
rect 14016 35154 14044 35770
rect 14740 35624 14792 35630
rect 14740 35566 14792 35572
rect 14094 35184 14150 35193
rect 14004 35148 14056 35154
rect 14094 35119 14150 35128
rect 14004 35090 14056 35096
rect 14108 35086 14136 35119
rect 13912 35080 13964 35086
rect 13912 35022 13964 35028
rect 14096 35080 14148 35086
rect 14096 35022 14148 35028
rect 14280 35080 14332 35086
rect 14280 35022 14332 35028
rect 13636 35012 13688 35018
rect 13636 34954 13688 34960
rect 13728 35012 13780 35018
rect 13728 34954 13780 34960
rect 13648 33969 13676 34954
rect 13740 34610 13768 34954
rect 13728 34604 13780 34610
rect 13728 34546 13780 34552
rect 13634 33960 13690 33969
rect 13634 33895 13690 33904
rect 13820 33924 13872 33930
rect 13820 33866 13872 33872
rect 13636 33856 13688 33862
rect 13542 33824 13598 33833
rect 13636 33798 13688 33804
rect 13542 33759 13598 33768
rect 13544 33448 13596 33454
rect 13464 33408 13544 33436
rect 13544 33390 13596 33396
rect 13556 33114 13584 33390
rect 13648 33114 13676 33798
rect 13544 33108 13596 33114
rect 13544 33050 13596 33056
rect 13636 33108 13688 33114
rect 13636 33050 13688 33056
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 13082 32263 13138 32272
rect 13176 32292 13228 32298
rect 13096 31890 13124 32263
rect 13176 32234 13228 32240
rect 13188 32008 13216 32234
rect 13188 31980 13308 32008
rect 13084 31884 13136 31890
rect 13084 31826 13136 31832
rect 13176 31680 13228 31686
rect 13176 31622 13228 31628
rect 13188 31482 13216 31622
rect 13176 31476 13228 31482
rect 13176 31418 13228 31424
rect 13082 30288 13138 30297
rect 12992 30252 13044 30258
rect 13082 30223 13138 30232
rect 12992 30194 13044 30200
rect 12912 29736 13032 29764
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12912 29306 12940 29582
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 13004 29209 13032 29736
rect 12990 29200 13046 29209
rect 12990 29135 13046 29144
rect 12900 29096 12952 29102
rect 12900 29038 12952 29044
rect 12912 28558 12940 29038
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 12900 27872 12952 27878
rect 12900 27814 12952 27820
rect 12912 27130 12940 27814
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 12898 26616 12954 26625
rect 12898 26551 12954 26560
rect 12912 25838 12940 26551
rect 13004 25906 13032 29135
rect 13096 27062 13124 30223
rect 13174 30016 13230 30025
rect 13174 29951 13230 29960
rect 13188 29646 13216 29951
rect 13176 29640 13228 29646
rect 13176 29582 13228 29588
rect 13280 28994 13308 31980
rect 13372 31736 13400 32710
rect 13556 32609 13584 33050
rect 13636 32904 13688 32910
rect 13636 32846 13688 32852
rect 13832 32858 13860 33866
rect 13924 33522 13952 35022
rect 14096 34944 14148 34950
rect 14148 34904 14228 34932
rect 14096 34886 14148 34892
rect 14004 34740 14056 34746
rect 14004 34682 14056 34688
rect 14016 33862 14044 34682
rect 14096 34536 14148 34542
rect 14096 34478 14148 34484
rect 14108 34202 14136 34478
rect 14200 34474 14228 34904
rect 14188 34468 14240 34474
rect 14188 34410 14240 34416
rect 14096 34196 14148 34202
rect 14096 34138 14148 34144
rect 14004 33856 14056 33862
rect 14004 33798 14056 33804
rect 13912 33516 13964 33522
rect 13912 33458 13964 33464
rect 13924 33114 13952 33458
rect 14004 33312 14056 33318
rect 14004 33254 14056 33260
rect 13912 33108 13964 33114
rect 13912 33050 13964 33056
rect 14016 33017 14044 33254
rect 14108 33114 14136 34138
rect 14200 33930 14228 34410
rect 14188 33924 14240 33930
rect 14188 33866 14240 33872
rect 14200 33522 14228 33866
rect 14188 33516 14240 33522
rect 14188 33458 14240 33464
rect 14096 33108 14148 33114
rect 14096 33050 14148 33056
rect 14002 33008 14058 33017
rect 14002 32943 14058 32952
rect 13542 32600 13598 32609
rect 13542 32535 13598 32544
rect 13556 32502 13584 32535
rect 13544 32496 13596 32502
rect 13544 32438 13596 32444
rect 13544 32360 13596 32366
rect 13544 32302 13596 32308
rect 13556 31890 13584 32302
rect 13544 31884 13596 31890
rect 13544 31826 13596 31832
rect 13452 31748 13504 31754
rect 13372 31708 13452 31736
rect 13372 31482 13400 31708
rect 13452 31690 13504 31696
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13372 29617 13400 31418
rect 13648 31346 13676 32846
rect 13832 32830 13952 32858
rect 13820 32768 13872 32774
rect 13820 32710 13872 32716
rect 13832 32434 13860 32710
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 13820 32292 13872 32298
rect 13820 32234 13872 32240
rect 13832 31414 13860 32234
rect 13924 31929 13952 32830
rect 13910 31920 13966 31929
rect 13910 31855 13912 31864
rect 13964 31855 13966 31864
rect 13912 31826 13964 31832
rect 13820 31408 13872 31414
rect 13820 31350 13872 31356
rect 13636 31340 13688 31346
rect 13636 31282 13688 31288
rect 14016 31226 14044 32943
rect 14200 32434 14228 33458
rect 14188 32428 14240 32434
rect 14188 32370 14240 32376
rect 14096 32292 14148 32298
rect 14096 32234 14148 32240
rect 14108 32026 14136 32234
rect 14292 32026 14320 35022
rect 14556 34944 14608 34950
rect 14556 34886 14608 34892
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 14372 33924 14424 33930
rect 14372 33866 14424 33872
rect 14384 33658 14412 33866
rect 14372 33652 14424 33658
rect 14372 33594 14424 33600
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 14384 32910 14412 33254
rect 14372 32904 14424 32910
rect 14372 32846 14424 32852
rect 14372 32768 14424 32774
rect 14372 32710 14424 32716
rect 14096 32020 14148 32026
rect 14280 32020 14332 32026
rect 14096 31962 14148 31968
rect 14200 31980 14280 32008
rect 14096 31816 14148 31822
rect 14096 31758 14148 31764
rect 14108 31346 14136 31758
rect 14096 31340 14148 31346
rect 14096 31282 14148 31288
rect 14016 31198 14136 31226
rect 13728 30728 13780 30734
rect 13728 30670 13780 30676
rect 13634 30560 13690 30569
rect 13634 30495 13690 30504
rect 13452 30252 13504 30258
rect 13504 30212 13584 30240
rect 13452 30194 13504 30200
rect 13358 29608 13414 29617
rect 13358 29543 13414 29552
rect 13556 29306 13584 30212
rect 13544 29300 13596 29306
rect 13544 29242 13596 29248
rect 13556 28994 13584 29242
rect 13648 29102 13676 30495
rect 13740 30326 13768 30670
rect 14004 30388 14056 30394
rect 14004 30330 14056 30336
rect 13728 30320 13780 30326
rect 14016 30297 14044 30330
rect 13728 30262 13780 30268
rect 14002 30288 14058 30297
rect 14002 30223 14058 30232
rect 14004 30184 14056 30190
rect 14004 30126 14056 30132
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 13188 28966 13308 28994
rect 13464 28966 13584 28994
rect 13740 28966 13768 29582
rect 13912 29504 13964 29510
rect 13912 29446 13964 29452
rect 13820 29164 13872 29170
rect 13820 29106 13872 29112
rect 13188 27674 13216 28966
rect 13464 28744 13492 28966
rect 13728 28960 13780 28966
rect 13728 28902 13780 28908
rect 13280 28716 13492 28744
rect 13176 27668 13228 27674
rect 13176 27610 13228 27616
rect 13188 27402 13216 27610
rect 13280 27606 13308 28716
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 13268 27600 13320 27606
rect 13268 27542 13320 27548
rect 13280 27402 13308 27542
rect 13176 27396 13228 27402
rect 13176 27338 13228 27344
rect 13268 27396 13320 27402
rect 13268 27338 13320 27344
rect 13084 27056 13136 27062
rect 13280 27033 13308 27338
rect 13084 26998 13136 27004
rect 13266 27024 13322 27033
rect 13266 26959 13322 26968
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 13268 26784 13320 26790
rect 13268 26726 13320 26732
rect 13096 25974 13124 26726
rect 13280 26586 13308 26726
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 13174 26072 13230 26081
rect 13174 26007 13176 26016
rect 13228 26007 13230 26016
rect 13176 25978 13228 25984
rect 13084 25968 13136 25974
rect 13084 25910 13136 25916
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 12900 25832 12952 25838
rect 12900 25774 12952 25780
rect 13268 25832 13320 25838
rect 13268 25774 13320 25780
rect 12900 25696 12952 25702
rect 12900 25638 12952 25644
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 12912 23322 12940 25638
rect 13004 24449 13032 25638
rect 13174 24984 13230 24993
rect 13174 24919 13230 24928
rect 13188 24818 13216 24919
rect 13280 24834 13308 25774
rect 13372 25294 13400 28562
rect 13544 28484 13596 28490
rect 13544 28426 13596 28432
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 13452 27396 13504 27402
rect 13452 27338 13504 27344
rect 13464 26926 13492 27338
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 13556 25906 13584 28426
rect 13636 28008 13688 28014
rect 13740 27985 13768 28426
rect 13636 27950 13688 27956
rect 13726 27976 13782 27985
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13648 25537 13676 27950
rect 13726 27911 13782 27920
rect 13832 27878 13860 29106
rect 13924 27946 13952 29446
rect 14016 29345 14044 30126
rect 14002 29336 14058 29345
rect 14002 29271 14058 29280
rect 14016 28762 14044 29271
rect 14108 28762 14136 31198
rect 14200 28994 14228 31980
rect 14280 31962 14332 31968
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14292 30734 14320 31282
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14182 28966 14228 28994
rect 14004 28756 14056 28762
rect 14004 28698 14056 28704
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 13912 27940 13964 27946
rect 13912 27882 13964 27888
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13634 25528 13690 25537
rect 13634 25463 13690 25472
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13464 24954 13492 25094
rect 13452 24948 13504 24954
rect 13452 24890 13504 24896
rect 13648 24886 13676 25094
rect 13636 24880 13688 24886
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13176 24812 13228 24818
rect 13280 24806 13492 24834
rect 13636 24822 13688 24828
rect 13176 24754 13228 24760
rect 12990 24440 13046 24449
rect 12990 24375 13046 24384
rect 13004 24206 13032 24375
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 23316 12952 23322
rect 12900 23258 12952 23264
rect 13004 22710 13032 23666
rect 13096 23186 13124 24754
rect 13193 24698 13221 24754
rect 13188 24670 13221 24698
rect 13188 24410 13216 24670
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 13280 24206 13308 24550
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13372 23798 13400 24550
rect 13464 23905 13492 24806
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13450 23896 13506 23905
rect 13450 23831 13506 23840
rect 13360 23792 13412 23798
rect 13360 23734 13412 23740
rect 13268 23656 13320 23662
rect 13268 23598 13320 23604
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 13096 23050 13124 23122
rect 13280 23050 13308 23598
rect 13084 23044 13136 23050
rect 13084 22986 13136 22992
rect 13268 23044 13320 23050
rect 13268 22986 13320 22992
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 13096 22642 13124 22986
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13082 22264 13138 22273
rect 12992 22228 13044 22234
rect 13082 22199 13138 22208
rect 12992 22170 13044 22176
rect 13004 22137 13032 22170
rect 12990 22128 13046 22137
rect 12820 22066 12940 22094
rect 12624 22034 12676 22040
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12544 21350 12572 21966
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12544 20466 12572 20946
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12636 20466 12664 20878
rect 12728 20602 12756 21830
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 12530 20224 12586 20233
rect 12530 20159 12586 20168
rect 12544 19514 12572 20159
rect 12636 19854 12664 20402
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12728 19378 12756 20538
rect 12820 19854 12848 21830
rect 12912 20806 12940 22066
rect 12990 22063 13046 22072
rect 12990 21856 13046 21865
rect 12990 21791 13046 21800
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12898 20632 12954 20641
rect 12898 20567 12954 20576
rect 12912 20466 12940 20567
rect 13004 20534 13032 21791
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12912 19854 12940 20402
rect 13096 20058 13124 22199
rect 13188 22030 13216 22578
rect 13280 22030 13308 22986
rect 13556 22692 13584 24346
rect 13740 24342 13768 27338
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 13728 23860 13780 23866
rect 13832 23848 13860 27814
rect 13912 27328 13964 27334
rect 13912 27270 13964 27276
rect 13924 24721 13952 27270
rect 14016 27010 14044 28698
rect 14108 27538 14136 28698
rect 14182 28540 14210 28966
rect 14182 28512 14228 28540
rect 14096 27532 14148 27538
rect 14096 27474 14148 27480
rect 14016 26982 14136 27010
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14016 24818 14044 26862
rect 14108 26586 14136 26982
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 14096 25968 14148 25974
rect 14096 25910 14148 25916
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 13910 24712 13966 24721
rect 13910 24647 13966 24656
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14016 24274 14044 24550
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 13780 23820 13860 23848
rect 13728 23802 13780 23808
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13464 22664 13584 22692
rect 13464 22234 13492 22664
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13360 22160 13412 22166
rect 13358 22128 13360 22137
rect 13412 22128 13414 22137
rect 13358 22063 13414 22072
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 13464 21554 13492 21898
rect 13648 21672 13676 23598
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13728 22704 13780 22710
rect 13728 22646 13780 22652
rect 13556 21644 13676 21672
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13556 21146 13584 21644
rect 13636 21548 13688 21554
rect 13740 21536 13768 22646
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13832 21622 13860 21966
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13688 21508 13768 21536
rect 13636 21490 13688 21496
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13832 21146 13860 21354
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13924 21078 13952 23054
rect 14108 22658 14136 25910
rect 14200 24818 14228 28512
rect 14292 26790 14320 30670
rect 14384 29850 14412 32710
rect 14476 30258 14504 34478
rect 14568 34406 14596 34886
rect 14556 34400 14608 34406
rect 14556 34342 14608 34348
rect 14648 34400 14700 34406
rect 14648 34342 14700 34348
rect 14556 33380 14608 33386
rect 14556 33322 14608 33328
rect 14568 32910 14596 33322
rect 14556 32904 14608 32910
rect 14556 32846 14608 32852
rect 14556 32496 14608 32502
rect 14556 32438 14608 32444
rect 14568 31210 14596 32438
rect 14556 31204 14608 31210
rect 14556 31146 14608 31152
rect 14556 30796 14608 30802
rect 14556 30738 14608 30744
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14384 29238 14412 29582
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 14384 29050 14412 29174
rect 14384 29022 14504 29050
rect 14476 27614 14504 29022
rect 14568 28994 14596 30738
rect 14660 29238 14688 34342
rect 14752 34202 14780 35566
rect 14832 35556 14884 35562
rect 14832 35498 14884 35504
rect 14844 35086 14872 35498
rect 15016 35488 15068 35494
rect 15016 35430 15068 35436
rect 15028 35086 15056 35430
rect 14832 35080 14884 35086
rect 14832 35022 14884 35028
rect 15016 35080 15068 35086
rect 15016 35022 15068 35028
rect 14844 34542 14872 35022
rect 14832 34536 14884 34542
rect 14832 34478 14884 34484
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 15028 33522 15056 35022
rect 15212 34474 15240 35770
rect 15384 35080 15436 35086
rect 15382 35048 15384 35057
rect 15436 35048 15438 35057
rect 15382 34983 15438 34992
rect 15752 34944 15804 34950
rect 15752 34886 15804 34892
rect 15200 34468 15252 34474
rect 15200 34410 15252 34416
rect 15106 33960 15162 33969
rect 15106 33895 15162 33904
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 14924 32836 14976 32842
rect 14924 32778 14976 32784
rect 14832 32360 14884 32366
rect 14832 32302 14884 32308
rect 14844 32042 14872 32302
rect 14752 32014 14872 32042
rect 14752 30122 14780 32014
rect 14936 31346 14964 32778
rect 15014 32328 15070 32337
rect 15014 32263 15070 32272
rect 15028 32026 15056 32263
rect 15016 32020 15068 32026
rect 15016 31962 15068 31968
rect 15016 31680 15068 31686
rect 15016 31622 15068 31628
rect 14924 31340 14976 31346
rect 14924 31282 14976 31288
rect 14936 30802 14964 31282
rect 14924 30796 14976 30802
rect 14924 30738 14976 30744
rect 15028 30598 15056 31622
rect 15120 30870 15148 33895
rect 15212 32910 15240 34410
rect 15476 33992 15528 33998
rect 15476 33934 15528 33940
rect 15292 33312 15344 33318
rect 15292 33254 15344 33260
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15304 32230 15332 33254
rect 15488 33114 15516 33934
rect 15764 33930 15792 34886
rect 15752 33924 15804 33930
rect 15752 33866 15804 33872
rect 15476 33108 15528 33114
rect 15476 33050 15528 33056
rect 15384 33040 15436 33046
rect 15384 32982 15436 32988
rect 15396 32434 15424 32982
rect 15660 32768 15712 32774
rect 15660 32710 15712 32716
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 15568 32428 15620 32434
rect 15568 32370 15620 32376
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15292 32224 15344 32230
rect 15292 32166 15344 32172
rect 15108 30864 15160 30870
rect 15108 30806 15160 30812
rect 15016 30592 15068 30598
rect 15016 30534 15068 30540
rect 14740 30116 14792 30122
rect 14740 30058 14792 30064
rect 14752 29850 14780 30058
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 14740 29844 14792 29850
rect 14740 29786 14792 29792
rect 14844 29560 14872 29990
rect 14936 29714 14964 29990
rect 14924 29708 14976 29714
rect 14924 29650 14976 29656
rect 14924 29572 14976 29578
rect 14844 29532 14924 29560
rect 14924 29514 14976 29520
rect 14738 29336 14794 29345
rect 14936 29306 14964 29514
rect 14738 29271 14794 29280
rect 14924 29300 14976 29306
rect 14648 29232 14700 29238
rect 14648 29174 14700 29180
rect 14752 29170 14780 29271
rect 14924 29242 14976 29248
rect 14740 29164 14792 29170
rect 14740 29106 14792 29112
rect 14648 29096 14700 29102
rect 14832 29096 14884 29102
rect 14700 29044 14832 29050
rect 14648 29038 14884 29044
rect 14660 29022 14872 29038
rect 15028 28994 15056 30534
rect 15106 29608 15162 29617
rect 15106 29543 15162 29552
rect 14568 28966 14780 28994
rect 14646 27976 14702 27985
rect 14556 27940 14608 27946
rect 14646 27911 14648 27920
rect 14556 27882 14608 27888
rect 14700 27911 14702 27920
rect 14752 27928 14780 28966
rect 14844 28966 15056 28994
rect 14844 28082 14872 28966
rect 15120 28642 15148 29543
rect 15028 28614 15148 28642
rect 14832 28076 14884 28082
rect 14832 28018 14884 28024
rect 14924 28076 14976 28082
rect 14924 28018 14976 28024
rect 14832 27940 14884 27946
rect 14752 27900 14832 27928
rect 14648 27882 14700 27888
rect 14832 27882 14884 27888
rect 14384 27586 14504 27614
rect 14384 27130 14412 27586
rect 14568 27470 14596 27882
rect 14936 27674 14964 28018
rect 14924 27668 14976 27674
rect 14924 27610 14976 27616
rect 14648 27600 14700 27606
rect 14646 27568 14648 27577
rect 14700 27568 14702 27577
rect 14646 27503 14702 27512
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14372 27124 14424 27130
rect 14372 27066 14424 27072
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14292 26314 14320 26726
rect 14280 26308 14332 26314
rect 14280 26250 14332 26256
rect 14384 26024 14412 27066
rect 14476 26042 14504 27406
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14292 25996 14412 26024
rect 14464 26036 14516 26042
rect 14292 25158 14320 25996
rect 14464 25978 14516 25984
rect 14568 25838 14596 27270
rect 14646 27160 14702 27169
rect 14646 27095 14702 27104
rect 14660 26926 14688 27095
rect 14648 26920 14700 26926
rect 14648 26862 14700 26868
rect 14556 25832 14608 25838
rect 14556 25774 14608 25780
rect 14372 25696 14424 25702
rect 14372 25638 14424 25644
rect 14384 25226 14412 25638
rect 14554 25528 14610 25537
rect 14554 25463 14610 25472
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 14280 25152 14332 25158
rect 14280 25094 14332 25100
rect 14292 24818 14320 25094
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14188 24132 14240 24138
rect 14188 24074 14240 24080
rect 14200 23866 14228 24074
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14004 22636 14056 22642
rect 14108 22630 14228 22658
rect 14004 22578 14056 22584
rect 14016 22234 14044 22578
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 14200 22094 14228 22630
rect 14292 22438 14320 22918
rect 14280 22432 14332 22438
rect 14384 22420 14412 25162
rect 14568 24070 14596 25463
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14568 23633 14596 24006
rect 14554 23624 14610 23633
rect 14554 23559 14610 23568
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22522 14504 22918
rect 14660 22642 14688 26862
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14752 22556 14780 26726
rect 14844 25294 14872 27406
rect 15028 26926 15056 28614
rect 15108 28416 15160 28422
rect 15108 28358 15160 28364
rect 15120 27674 15148 28358
rect 15212 28082 15240 32166
rect 15396 30138 15424 32370
rect 15580 31414 15608 32370
rect 15672 31822 15700 32710
rect 15660 31816 15712 31822
rect 15660 31758 15712 31764
rect 15568 31408 15620 31414
rect 15568 31350 15620 31356
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15580 30326 15608 30670
rect 15660 30388 15712 30394
rect 15660 30330 15712 30336
rect 15568 30320 15620 30326
rect 15568 30262 15620 30268
rect 15396 30110 15516 30138
rect 15384 30048 15436 30054
rect 15384 29990 15436 29996
rect 15292 29776 15344 29782
rect 15396 29753 15424 29990
rect 15292 29718 15344 29724
rect 15382 29744 15438 29753
rect 15304 29102 15332 29718
rect 15382 29679 15438 29688
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15120 27062 15148 27610
rect 15396 27606 15424 29582
rect 15488 29170 15516 30110
rect 15568 29504 15620 29510
rect 15568 29446 15620 29452
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15488 28082 15516 29106
rect 15580 29102 15608 29446
rect 15672 29238 15700 30330
rect 15660 29232 15712 29238
rect 15660 29174 15712 29180
rect 15568 29096 15620 29102
rect 15568 29038 15620 29044
rect 15660 28960 15712 28966
rect 15660 28902 15712 28908
rect 15672 28762 15700 28902
rect 15660 28756 15712 28762
rect 15660 28698 15712 28704
rect 15660 28144 15712 28150
rect 15764 28132 15792 33866
rect 15856 31754 15884 36110
rect 16592 36009 16620 36343
rect 16684 36106 16712 36518
rect 16960 36378 16988 37810
rect 17224 37188 17276 37194
rect 17224 37130 17276 37136
rect 16948 36372 17000 36378
rect 16948 36314 17000 36320
rect 17236 36145 17264 37130
rect 17604 36242 17632 38626
rect 17696 38418 17724 39510
rect 17788 38962 17816 40326
rect 17972 40186 18000 41074
rect 18052 41064 18104 41070
rect 18050 41032 18052 41041
rect 18104 41032 18106 41041
rect 18156 41002 18184 41126
rect 18050 40967 18106 40976
rect 18144 40996 18196 41002
rect 18144 40938 18196 40944
rect 18052 40724 18104 40730
rect 18052 40666 18104 40672
rect 17960 40180 18012 40186
rect 17960 40122 18012 40128
rect 17960 39432 18012 39438
rect 17880 39380 17960 39386
rect 17880 39374 18012 39380
rect 17880 39358 18000 39374
rect 17776 38956 17828 38962
rect 17776 38898 17828 38904
rect 17788 38418 17816 38898
rect 17880 38554 17908 39358
rect 17960 39296 18012 39302
rect 17958 39264 17960 39273
rect 18012 39264 18014 39273
rect 17958 39199 18014 39208
rect 17960 39024 18012 39030
rect 17960 38966 18012 38972
rect 17972 38554 18000 38966
rect 18064 38962 18092 40666
rect 18340 40662 18368 41142
rect 18418 41103 18474 41112
rect 18512 41132 18564 41138
rect 18432 41070 18460 41103
rect 18512 41074 18564 41080
rect 18604 41132 18656 41138
rect 18604 41074 18656 41080
rect 18420 41064 18472 41070
rect 18420 41006 18472 41012
rect 18328 40656 18380 40662
rect 18328 40598 18380 40604
rect 18144 40520 18196 40526
rect 18142 40488 18144 40497
rect 18196 40488 18198 40497
rect 18142 40423 18198 40432
rect 18340 40390 18368 40598
rect 18328 40384 18380 40390
rect 18328 40326 18380 40332
rect 18144 40112 18196 40118
rect 18144 40054 18196 40060
rect 18156 39030 18184 40054
rect 18340 39964 18368 40326
rect 18432 40089 18460 41006
rect 18524 40662 18552 41074
rect 18512 40656 18564 40662
rect 18616 40633 18644 41074
rect 18708 40934 18736 41618
rect 18984 41546 19012 41647
rect 19064 41618 19116 41624
rect 19892 41676 20220 41682
rect 19944 41670 20168 41676
rect 19892 41618 19944 41624
rect 20168 41618 20220 41624
rect 18972 41540 19024 41546
rect 18972 41482 19024 41488
rect 19076 41120 19104 41618
rect 20076 41608 20128 41614
rect 19996 41568 20076 41596
rect 19996 41562 20024 41568
rect 19352 41534 20024 41562
rect 20076 41550 20128 41556
rect 20168 41540 20220 41546
rect 19156 41132 19208 41138
rect 19076 41092 19156 41120
rect 18878 41032 18934 41041
rect 18878 40967 18934 40976
rect 18696 40928 18748 40934
rect 18696 40870 18748 40876
rect 18512 40598 18564 40604
rect 18602 40624 18658 40633
rect 18418 40080 18474 40089
rect 18418 40015 18474 40024
rect 18340 39936 18460 39964
rect 18236 39432 18288 39438
rect 18236 39374 18288 39380
rect 18144 39024 18196 39030
rect 18144 38966 18196 38972
rect 18052 38956 18104 38962
rect 18052 38898 18104 38904
rect 17868 38548 17920 38554
rect 17868 38490 17920 38496
rect 17960 38548 18012 38554
rect 17960 38490 18012 38496
rect 17684 38412 17736 38418
rect 17684 38354 17736 38360
rect 17776 38412 17828 38418
rect 17776 38354 17828 38360
rect 17880 38010 17908 38490
rect 17868 38004 17920 38010
rect 17868 37946 17920 37952
rect 17776 37188 17828 37194
rect 17776 37130 17828 37136
rect 17684 36848 17736 36854
rect 17684 36790 17736 36796
rect 17592 36236 17644 36242
rect 17592 36178 17644 36184
rect 17222 36136 17278 36145
rect 16672 36100 16724 36106
rect 17222 36071 17278 36080
rect 16672 36042 16724 36048
rect 16578 36000 16634 36009
rect 16578 35935 16634 35944
rect 17696 35873 17724 36790
rect 17788 36174 17816 37130
rect 17960 37120 18012 37126
rect 17960 37062 18012 37068
rect 17972 36718 18000 37062
rect 18064 36854 18092 38898
rect 18156 37262 18184 38966
rect 18248 38554 18276 39374
rect 18328 39364 18380 39370
rect 18328 39306 18380 39312
rect 18340 39137 18368 39306
rect 18326 39128 18382 39137
rect 18326 39063 18382 39072
rect 18236 38548 18288 38554
rect 18236 38490 18288 38496
rect 18432 38418 18460 39936
rect 18524 39642 18552 40598
rect 18602 40559 18658 40568
rect 18616 40361 18644 40559
rect 18708 40526 18736 40870
rect 18696 40520 18748 40526
rect 18696 40462 18748 40468
rect 18602 40352 18658 40361
rect 18602 40287 18658 40296
rect 18604 40044 18656 40050
rect 18604 39986 18656 39992
rect 18512 39636 18564 39642
rect 18512 39578 18564 39584
rect 18420 38412 18472 38418
rect 18420 38354 18472 38360
rect 18236 38344 18288 38350
rect 18236 38286 18288 38292
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18052 36848 18104 36854
rect 18052 36790 18104 36796
rect 18144 36780 18196 36786
rect 18144 36722 18196 36728
rect 17960 36712 18012 36718
rect 17960 36654 18012 36660
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 18156 36530 18184 36722
rect 18248 36689 18276 38286
rect 18524 37738 18552 39578
rect 18616 39438 18644 39986
rect 18696 39636 18748 39642
rect 18696 39578 18748 39584
rect 18604 39432 18656 39438
rect 18602 39400 18604 39409
rect 18656 39400 18658 39409
rect 18602 39335 18658 39344
rect 18708 39302 18736 39578
rect 18788 39432 18840 39438
rect 18788 39374 18840 39380
rect 18800 39302 18828 39374
rect 18696 39296 18748 39302
rect 18696 39238 18748 39244
rect 18788 39296 18840 39302
rect 18788 39238 18840 39244
rect 18892 39098 18920 40967
rect 19076 40730 19104 41092
rect 19156 41074 19208 41080
rect 19352 41070 19380 41534
rect 20168 41482 20220 41488
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 20180 41313 20208 41482
rect 20166 41304 20222 41313
rect 20166 41239 20222 41248
rect 19800 41132 19852 41138
rect 19628 41092 19800 41120
rect 19248 41064 19300 41070
rect 19248 41006 19300 41012
rect 19340 41064 19392 41070
rect 19340 41006 19392 41012
rect 19260 40905 19288 41006
rect 19246 40896 19302 40905
rect 19246 40831 19302 40840
rect 19064 40724 19116 40730
rect 19064 40666 19116 40672
rect 18972 39432 19024 39438
rect 18972 39374 19024 39380
rect 18984 39273 19012 39374
rect 18970 39264 19026 39273
rect 18970 39199 19026 39208
rect 18880 39092 18932 39098
rect 18880 39034 18932 39040
rect 18892 38654 18920 39034
rect 18892 38626 19012 38654
rect 18880 37868 18932 37874
rect 18880 37810 18932 37816
rect 18420 37732 18472 37738
rect 18420 37674 18472 37680
rect 18512 37732 18564 37738
rect 18512 37674 18564 37680
rect 18328 37460 18380 37466
rect 18328 37402 18380 37408
rect 18234 36680 18290 36689
rect 18234 36615 18236 36624
rect 18288 36615 18290 36624
rect 18236 36586 18288 36592
rect 18340 36530 18368 37402
rect 17776 36168 17828 36174
rect 17776 36110 17828 36116
rect 17972 36106 18000 36518
rect 18156 36502 18368 36530
rect 18432 36242 18460 37674
rect 18892 37670 18920 37810
rect 18788 37664 18840 37670
rect 18788 37606 18840 37612
rect 18880 37664 18932 37670
rect 18880 37606 18932 37612
rect 18604 37120 18656 37126
rect 18604 37062 18656 37068
rect 18510 36952 18566 36961
rect 18616 36922 18644 37062
rect 18510 36887 18512 36896
rect 18564 36887 18566 36896
rect 18604 36916 18656 36922
rect 18512 36858 18564 36864
rect 18604 36858 18656 36864
rect 18512 36780 18564 36786
rect 18512 36722 18564 36728
rect 18144 36236 18196 36242
rect 18144 36178 18196 36184
rect 18420 36236 18472 36242
rect 18420 36178 18472 36184
rect 17960 36100 18012 36106
rect 17960 36042 18012 36048
rect 17682 35864 17738 35873
rect 17682 35799 17738 35808
rect 18156 35222 18184 36178
rect 18524 36009 18552 36722
rect 18616 36700 18644 36858
rect 18616 36672 18736 36700
rect 18708 36038 18736 36672
rect 18800 36582 18828 37606
rect 18892 37398 18920 37606
rect 18880 37392 18932 37398
rect 18880 37334 18932 37340
rect 18880 37120 18932 37126
rect 18880 37062 18932 37068
rect 18892 36961 18920 37062
rect 18878 36952 18934 36961
rect 18878 36887 18934 36896
rect 18984 36666 19012 38626
rect 19076 36825 19104 40666
rect 19628 40662 19656 41092
rect 19800 41074 19852 41080
rect 20076 41132 20128 41138
rect 20076 41074 20128 41080
rect 20168 41132 20220 41138
rect 20168 41074 20220 41080
rect 19708 40996 19760 41002
rect 19892 40996 19944 41002
rect 19760 40956 19892 40984
rect 19708 40938 19760 40944
rect 19892 40938 19944 40944
rect 19616 40656 19668 40662
rect 20088 40610 20116 41074
rect 20180 40730 20208 41074
rect 20168 40724 20220 40730
rect 20168 40666 20220 40672
rect 19616 40598 19668 40604
rect 19996 40582 20116 40610
rect 19248 40520 19300 40526
rect 19248 40462 19300 40468
rect 19708 40520 19760 40526
rect 19996 40508 20024 40582
rect 19760 40480 20024 40508
rect 20076 40520 20128 40526
rect 19708 40462 19760 40468
rect 20076 40462 20128 40468
rect 19260 40186 19288 40462
rect 19616 40384 19668 40390
rect 19338 40352 19394 40361
rect 19668 40361 20024 40372
rect 19668 40352 20038 40361
rect 19668 40344 19982 40352
rect 19616 40326 19668 40332
rect 19338 40287 19394 40296
rect 19248 40180 19300 40186
rect 19248 40122 19300 40128
rect 19156 39432 19208 39438
rect 19154 39400 19156 39409
rect 19208 39400 19210 39409
rect 19154 39335 19210 39344
rect 19156 37324 19208 37330
rect 19156 37266 19208 37272
rect 19062 36816 19118 36825
rect 19168 36786 19196 37266
rect 19260 36854 19288 40122
rect 19352 39302 19380 40287
rect 19574 40284 19882 40293
rect 19982 40287 20038 40296
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 20088 40186 20116 40462
rect 20272 40458 20300 41686
rect 20718 41647 20774 41656
rect 23296 41676 23348 41682
rect 23296 41618 23348 41624
rect 20536 41608 20588 41614
rect 22652 41608 22704 41614
rect 20536 41550 20588 41556
rect 20352 41200 20404 41206
rect 20352 41142 20404 41148
rect 20260 40452 20312 40458
rect 20260 40394 20312 40400
rect 20166 40216 20222 40225
rect 20076 40180 20128 40186
rect 20272 40186 20300 40394
rect 20166 40151 20222 40160
rect 20260 40180 20312 40186
rect 20076 40122 20128 40128
rect 20180 39914 20208 40151
rect 20260 40122 20312 40128
rect 20364 40118 20392 41142
rect 20444 41132 20496 41138
rect 20444 41074 20496 41080
rect 20456 40662 20484 41074
rect 20548 40730 20576 41550
rect 22204 41546 22508 41562
rect 22652 41550 22704 41556
rect 23202 41576 23258 41585
rect 21456 41540 21508 41546
rect 21456 41482 21508 41488
rect 22100 41540 22152 41546
rect 22100 41482 22152 41488
rect 22204 41540 22520 41546
rect 22204 41534 22468 41540
rect 20812 41472 20864 41478
rect 20812 41414 20864 41420
rect 20824 41138 20852 41414
rect 20812 41132 20864 41138
rect 20812 41074 20864 41080
rect 21088 41132 21140 41138
rect 21088 41074 21140 41080
rect 20536 40724 20588 40730
rect 20536 40666 20588 40672
rect 20444 40656 20496 40662
rect 20444 40598 20496 40604
rect 20824 40526 20852 41074
rect 21100 40934 21128 41074
rect 21468 41070 21496 41482
rect 21836 41386 22048 41414
rect 21638 41304 21694 41313
rect 21638 41239 21694 41248
rect 21732 41268 21784 41274
rect 21456 41064 21508 41070
rect 21456 41006 21508 41012
rect 21088 40928 21140 40934
rect 21088 40870 21140 40876
rect 20812 40520 20864 40526
rect 20812 40462 20864 40468
rect 20720 40384 20772 40390
rect 20720 40326 20772 40332
rect 20444 40180 20496 40186
rect 20444 40122 20496 40128
rect 20352 40112 20404 40118
rect 20352 40054 20404 40060
rect 19800 39908 19852 39914
rect 19800 39850 19852 39856
rect 20168 39908 20220 39914
rect 20168 39850 20220 39856
rect 19812 39817 19840 39850
rect 19892 39840 19944 39846
rect 19798 39808 19854 39817
rect 19892 39782 19944 39788
rect 19798 39743 19854 39752
rect 19904 39438 19932 39782
rect 19892 39432 19944 39438
rect 19892 39374 19944 39380
rect 20260 39432 20312 39438
rect 20260 39374 20312 39380
rect 19432 39364 19484 39370
rect 19432 39306 19484 39312
rect 20168 39364 20220 39370
rect 20168 39306 20220 39312
rect 19340 39296 19392 39302
rect 19340 39238 19392 39244
rect 19444 38962 19472 39306
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19800 39092 19852 39098
rect 19800 39034 19852 39040
rect 19432 38956 19484 38962
rect 19432 38898 19484 38904
rect 19432 38412 19484 38418
rect 19432 38354 19484 38360
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19352 37806 19380 38150
rect 19444 38010 19472 38354
rect 19812 38350 19840 39034
rect 20088 38962 20116 39238
rect 20180 38978 20208 39306
rect 20272 39098 20300 39374
rect 20260 39092 20312 39098
rect 20260 39034 20312 39040
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 20076 38956 20128 38962
rect 20180 38950 20300 38978
rect 20076 38898 20128 38904
rect 19800 38344 19852 38350
rect 19800 38286 19852 38292
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19996 38010 20024 38898
rect 20168 38888 20220 38894
rect 20088 38836 20168 38842
rect 20088 38830 20220 38836
rect 20088 38814 20208 38830
rect 19432 38004 19484 38010
rect 19432 37946 19484 37952
rect 19984 38004 20036 38010
rect 19984 37946 20036 37952
rect 19340 37800 19392 37806
rect 19340 37742 19392 37748
rect 19444 37262 19472 37946
rect 20088 37890 20116 38814
rect 19996 37874 20116 37890
rect 19984 37868 20116 37874
rect 20036 37862 20116 37868
rect 19984 37810 20036 37816
rect 20076 37800 20128 37806
rect 20272 37777 20300 38950
rect 20076 37742 20128 37748
rect 20258 37768 20314 37777
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19248 36848 19300 36854
rect 19248 36790 19300 36796
rect 19892 36848 19944 36854
rect 19892 36790 19944 36796
rect 19062 36751 19064 36760
rect 19116 36751 19118 36760
rect 19156 36780 19208 36786
rect 19064 36722 19116 36728
rect 19156 36722 19208 36728
rect 18984 36650 19104 36666
rect 18880 36644 18932 36650
rect 18984 36644 19116 36650
rect 18984 36638 19064 36644
rect 18880 36586 18932 36592
rect 19064 36586 19116 36592
rect 18788 36576 18840 36582
rect 18788 36518 18840 36524
rect 18892 36310 18920 36586
rect 19156 36576 19208 36582
rect 19260 36553 19288 36790
rect 19524 36712 19576 36718
rect 19524 36654 19576 36660
rect 19432 36576 19484 36582
rect 19156 36518 19208 36524
rect 19246 36544 19302 36553
rect 19168 36378 19196 36518
rect 19246 36479 19302 36488
rect 19352 36536 19432 36564
rect 19156 36372 19208 36378
rect 19156 36314 19208 36320
rect 18880 36304 18932 36310
rect 18880 36246 18932 36252
rect 19248 36236 19300 36242
rect 19248 36178 19300 36184
rect 19260 36106 19288 36178
rect 19352 36145 19380 36536
rect 19432 36518 19484 36524
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 19444 36174 19472 36314
rect 19432 36168 19484 36174
rect 19338 36136 19394 36145
rect 19064 36100 19116 36106
rect 19064 36042 19116 36048
rect 19248 36100 19300 36106
rect 19536 36145 19564 36654
rect 19904 36378 19932 36790
rect 19984 36712 20036 36718
rect 19984 36654 20036 36660
rect 19892 36372 19944 36378
rect 19892 36314 19944 36320
rect 19432 36110 19484 36116
rect 19522 36136 19578 36145
rect 19338 36071 19394 36080
rect 19522 36071 19578 36080
rect 19248 36042 19300 36048
rect 18696 36032 18748 36038
rect 18510 36000 18566 36009
rect 18696 35974 18748 35980
rect 18510 35935 18566 35944
rect 19076 35494 19104 36042
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35714 20024 36654
rect 19904 35698 20024 35714
rect 19892 35692 20024 35698
rect 19944 35686 20024 35692
rect 19892 35634 19944 35640
rect 19890 35592 19946 35601
rect 19890 35527 19946 35536
rect 19904 35494 19932 35527
rect 19064 35488 19116 35494
rect 19064 35430 19116 35436
rect 19892 35488 19944 35494
rect 19892 35430 19944 35436
rect 15936 35216 15988 35222
rect 15936 35158 15988 35164
rect 16488 35216 16540 35222
rect 16672 35216 16724 35222
rect 16488 35158 16540 35164
rect 16670 35184 16672 35193
rect 18144 35216 18196 35222
rect 16724 35184 16726 35193
rect 15948 34649 15976 35158
rect 16028 35012 16080 35018
rect 16028 34954 16080 34960
rect 16040 34678 16068 34954
rect 16028 34672 16080 34678
rect 15934 34640 15990 34649
rect 16028 34614 16080 34620
rect 15934 34575 15990 34584
rect 16120 33924 16172 33930
rect 16120 33866 16172 33872
rect 16212 33924 16264 33930
rect 16212 33866 16264 33872
rect 16026 33144 16082 33153
rect 16026 33079 16082 33088
rect 16040 32910 16068 33079
rect 16132 32910 16160 33866
rect 16224 33697 16252 33866
rect 16210 33688 16266 33697
rect 16210 33623 16266 33632
rect 16396 33584 16448 33590
rect 16396 33526 16448 33532
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16304 33312 16356 33318
rect 16304 33254 16356 33260
rect 16224 32910 16252 33254
rect 16028 32904 16080 32910
rect 16028 32846 16080 32852
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 16212 32904 16264 32910
rect 16212 32846 16264 32852
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15948 32570 15976 32778
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 15936 32564 15988 32570
rect 15936 32506 15988 32512
rect 16040 32434 16068 32710
rect 16028 32428 16080 32434
rect 16028 32370 16080 32376
rect 16132 32298 16160 32846
rect 16316 32552 16344 33254
rect 16408 32570 16436 33526
rect 16224 32524 16344 32552
rect 16396 32564 16448 32570
rect 16120 32292 16172 32298
rect 16120 32234 16172 32240
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15948 32026 15976 32166
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 15936 31816 15988 31822
rect 15936 31758 15988 31764
rect 16120 31816 16172 31822
rect 16120 31758 16172 31764
rect 15844 31748 15896 31754
rect 15844 31690 15896 31696
rect 15948 31686 15976 31758
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 16028 31680 16080 31686
rect 16028 31622 16080 31628
rect 15936 31408 15988 31414
rect 15856 31368 15936 31396
rect 15856 30938 15884 31368
rect 15936 31350 15988 31356
rect 15936 31204 15988 31210
rect 15936 31146 15988 31152
rect 15844 30932 15896 30938
rect 15844 30874 15896 30880
rect 15856 29866 15884 30874
rect 15948 30666 15976 31146
rect 15936 30660 15988 30666
rect 15936 30602 15988 30608
rect 15948 30054 15976 30602
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15856 29838 15976 29866
rect 16040 29850 16068 31622
rect 16132 31346 16160 31758
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 16120 31136 16172 31142
rect 16120 31078 16172 31084
rect 16132 30326 16160 31078
rect 16120 30320 16172 30326
rect 16120 30262 16172 30268
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 15712 28104 15792 28132
rect 15856 28121 15884 29446
rect 15842 28112 15898 28121
rect 15660 28086 15712 28092
rect 15476 28076 15528 28082
rect 15842 28047 15898 28056
rect 15476 28018 15528 28024
rect 15948 27962 15976 29838
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 16132 29782 16160 30262
rect 16224 30258 16252 32524
rect 16396 32506 16448 32512
rect 16304 32428 16356 32434
rect 16304 32370 16356 32376
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 16316 31346 16344 32370
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16408 30938 16436 32370
rect 16500 31278 16528 35158
rect 18144 35158 18196 35164
rect 16670 35119 16726 35128
rect 17592 35148 17644 35154
rect 17592 35090 17644 35096
rect 17040 35080 17092 35086
rect 17040 35022 17092 35028
rect 16764 34944 16816 34950
rect 16764 34886 16816 34892
rect 16776 34610 16804 34886
rect 16764 34604 16816 34610
rect 16764 34546 16816 34552
rect 17052 34406 17080 35022
rect 17604 34610 17632 35090
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 17788 34746 18184 34762
rect 17776 34740 18184 34746
rect 17828 34734 18184 34740
rect 17776 34682 17828 34688
rect 17132 34604 17184 34610
rect 17132 34546 17184 34552
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17592 34604 17644 34610
rect 17592 34546 17644 34552
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 18052 34604 18104 34610
rect 18052 34546 18104 34552
rect 16672 34400 16724 34406
rect 16672 34342 16724 34348
rect 17040 34400 17092 34406
rect 17040 34342 17092 34348
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 16592 31890 16620 33798
rect 16684 33658 16712 34342
rect 17052 34202 17080 34342
rect 17040 34196 17092 34202
rect 17040 34138 17092 34144
rect 17052 33998 17080 34138
rect 17040 33992 17092 33998
rect 17040 33934 17092 33940
rect 16764 33924 16816 33930
rect 16764 33866 16816 33872
rect 16672 33652 16724 33658
rect 16672 33594 16724 33600
rect 16776 32881 16804 33866
rect 17040 33856 17092 33862
rect 16868 33816 17040 33844
rect 16762 32872 16818 32881
rect 16762 32807 16818 32816
rect 16868 32756 16896 33816
rect 17040 33798 17092 33804
rect 17038 33008 17094 33017
rect 17038 32943 17094 32952
rect 17052 32910 17080 32943
rect 17040 32904 17092 32910
rect 17040 32846 17092 32852
rect 16776 32728 16896 32756
rect 16948 32768 17000 32774
rect 16672 32224 16724 32230
rect 16672 32166 16724 32172
rect 16684 32026 16712 32166
rect 16672 32020 16724 32026
rect 16672 31962 16724 31968
rect 16776 31906 16804 32728
rect 16948 32710 17000 32716
rect 16960 32450 16988 32710
rect 16868 32434 16988 32450
rect 16856 32428 16988 32434
rect 16908 32422 16988 32428
rect 16856 32370 16908 32376
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16684 31878 16804 31906
rect 16684 31793 16712 31878
rect 16670 31784 16726 31793
rect 16580 31748 16632 31754
rect 16670 31719 16726 31728
rect 16580 31690 16632 31696
rect 16488 31272 16540 31278
rect 16488 31214 16540 31220
rect 16396 30932 16448 30938
rect 16396 30874 16448 30880
rect 16488 30728 16540 30734
rect 16316 30676 16488 30682
rect 16316 30670 16540 30676
rect 16316 30654 16528 30670
rect 16316 30433 16344 30654
rect 16396 30592 16448 30598
rect 16592 30580 16620 31690
rect 16396 30534 16448 30540
rect 16500 30552 16620 30580
rect 16302 30424 16358 30433
rect 16408 30394 16436 30534
rect 16302 30359 16358 30368
rect 16396 30388 16448 30394
rect 16396 30330 16448 30336
rect 16302 30288 16358 30297
rect 16212 30252 16264 30258
rect 16500 30240 16528 30552
rect 16302 30223 16358 30232
rect 16212 30194 16264 30200
rect 16212 30048 16264 30054
rect 16212 29990 16264 29996
rect 16120 29776 16172 29782
rect 16120 29718 16172 29724
rect 16028 29504 16080 29510
rect 16026 29472 16028 29481
rect 16120 29504 16172 29510
rect 16080 29472 16082 29481
rect 16120 29446 16172 29452
rect 16026 29407 16082 29416
rect 16132 29170 16160 29446
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16120 29028 16172 29034
rect 16120 28970 16172 28976
rect 16026 28792 16082 28801
rect 16026 28727 16082 28736
rect 15856 27934 15976 27962
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15764 27606 15792 27814
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15752 27600 15804 27606
rect 15752 27542 15804 27548
rect 15200 27464 15252 27470
rect 15198 27432 15200 27441
rect 15252 27432 15254 27441
rect 15856 27418 15884 27934
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 15198 27367 15254 27376
rect 15764 27390 15884 27418
rect 15764 27334 15792 27390
rect 15752 27328 15804 27334
rect 15752 27270 15804 27276
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 15108 27056 15160 27062
rect 15108 26998 15160 27004
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15120 26772 15148 26998
rect 15028 26744 15148 26772
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 14936 25906 14964 26318
rect 14924 25900 14976 25906
rect 14924 25842 14976 25848
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14936 25498 14964 25638
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 14832 25288 14884 25294
rect 14832 25230 14884 25236
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14844 24857 14872 24890
rect 14830 24848 14886 24857
rect 14830 24783 14886 24792
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 14936 24698 14964 25094
rect 15028 24993 15056 26744
rect 15382 26480 15438 26489
rect 15200 26444 15252 26450
rect 15382 26415 15384 26424
rect 15200 26386 15252 26392
rect 15436 26415 15438 26424
rect 15384 26386 15436 26392
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 15014 24984 15070 24993
rect 15014 24919 15070 24928
rect 15028 24818 15056 24919
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 14844 24585 14872 24686
rect 14936 24670 15056 24698
rect 14924 24608 14976 24614
rect 14830 24576 14886 24585
rect 14924 24550 14976 24556
rect 14830 24511 14886 24520
rect 14844 24342 14872 24511
rect 14832 24336 14884 24342
rect 14832 24278 14884 24284
rect 14832 24064 14884 24070
rect 14832 24006 14884 24012
rect 14844 22710 14872 24006
rect 14832 22704 14884 22710
rect 14832 22646 14884 22652
rect 14936 22642 14964 24550
rect 15028 23474 15056 24670
rect 15120 23730 15148 25774
rect 15212 25498 15240 26386
rect 15292 26376 15344 26382
rect 15382 26344 15438 26353
rect 15344 26324 15382 26330
rect 15292 26318 15382 26324
rect 15304 26302 15382 26318
rect 15382 26279 15438 26288
rect 15292 26240 15344 26246
rect 15292 26182 15344 26188
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15304 25294 15332 26182
rect 15488 25537 15516 26182
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15660 25900 15712 25906
rect 15660 25842 15712 25848
rect 15474 25528 15530 25537
rect 15580 25498 15608 25842
rect 15474 25463 15530 25472
rect 15568 25492 15620 25498
rect 15384 25356 15436 25362
rect 15488 25344 15516 25463
rect 15568 25434 15620 25440
rect 15672 25362 15700 25842
rect 15764 25498 15792 27270
rect 15856 26994 15884 27270
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15856 26489 15884 26930
rect 15948 26858 15976 27814
rect 16040 27402 16068 28727
rect 16132 28393 16160 28970
rect 16118 28384 16174 28393
rect 16118 28319 16174 28328
rect 16120 28008 16172 28014
rect 16120 27950 16172 27956
rect 16028 27396 16080 27402
rect 16028 27338 16080 27344
rect 15936 26852 15988 26858
rect 15936 26794 15988 26800
rect 15842 26480 15898 26489
rect 15842 26415 15844 26424
rect 15896 26415 15898 26424
rect 15844 26386 15896 26392
rect 15844 26240 15896 26246
rect 15844 26182 15896 26188
rect 15856 25838 15884 26182
rect 15844 25832 15896 25838
rect 15844 25774 15896 25780
rect 15752 25492 15804 25498
rect 15752 25434 15804 25440
rect 15948 25378 15976 26794
rect 16040 26450 16068 27338
rect 16028 26444 16080 26450
rect 16028 26386 16080 26392
rect 16132 25974 16160 27950
rect 16120 25968 16172 25974
rect 16120 25910 16172 25916
rect 16026 25528 16082 25537
rect 16026 25463 16082 25472
rect 15436 25316 15516 25344
rect 15660 25356 15712 25362
rect 15384 25298 15436 25304
rect 15660 25298 15712 25304
rect 15764 25350 15976 25378
rect 16040 25362 16068 25463
rect 16028 25356 16080 25362
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15580 24886 15608 25094
rect 15568 24880 15620 24886
rect 15660 24880 15712 24886
rect 15568 24822 15620 24828
rect 15658 24848 15660 24857
rect 15712 24848 15714 24857
rect 15292 24812 15344 24818
rect 15658 24783 15714 24792
rect 15292 24754 15344 24760
rect 15200 24744 15252 24750
rect 15198 24712 15200 24721
rect 15252 24712 15254 24721
rect 15198 24647 15254 24656
rect 15198 24440 15254 24449
rect 15304 24410 15332 24754
rect 15198 24375 15200 24384
rect 15252 24375 15254 24384
rect 15292 24404 15344 24410
rect 15200 24346 15252 24352
rect 15292 24346 15344 24352
rect 15658 24032 15714 24041
rect 15658 23967 15714 23976
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 15384 23520 15436 23526
rect 15028 23446 15240 23474
rect 15384 23462 15436 23468
rect 15568 23520 15620 23526
rect 15568 23462 15620 23468
rect 15014 23352 15070 23361
rect 15014 23287 15070 23296
rect 15028 23118 15056 23287
rect 15212 23225 15240 23446
rect 15198 23216 15254 23225
rect 15198 23151 15254 23160
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15292 23112 15344 23118
rect 15396 23100 15424 23462
rect 15580 23254 15608 23462
rect 15568 23248 15620 23254
rect 15568 23190 15620 23196
rect 15344 23072 15424 23100
rect 15292 23054 15344 23060
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15106 22672 15162 22681
rect 14924 22636 14976 22642
rect 15106 22607 15162 22616
rect 14924 22578 14976 22584
rect 14752 22528 14872 22556
rect 14476 22494 14688 22522
rect 14556 22432 14608 22438
rect 14384 22392 14504 22420
rect 14280 22374 14332 22380
rect 14476 22098 14504 22392
rect 14556 22374 14608 22380
rect 14200 22066 14412 22094
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 14292 21486 14320 21898
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13280 20058 13308 20198
rect 13556 20058 13584 20402
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13832 19854 13860 20946
rect 14002 20360 14058 20369
rect 14002 20295 14058 20304
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13832 19446 13860 19790
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12636 18766 12664 19110
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12268 18290 12296 18634
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 11900 17326 12020 17354
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11808 15910 11836 16526
rect 11900 16046 11928 17206
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11992 15638 12020 17326
rect 12176 17066 12204 18090
rect 12268 17678 12296 18226
rect 12452 17882 12480 18226
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 13004 17746 13032 19314
rect 13924 18766 13952 19926
rect 14016 19854 14044 20295
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14016 19378 14044 19790
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12268 17202 12296 17614
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 12268 16590 12296 17138
rect 13004 16590 13032 17682
rect 13096 17218 13124 18566
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13188 17338 13216 17546
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17338 13308 17478
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13174 17232 13230 17241
rect 13096 17190 13174 17218
rect 13174 17167 13230 17176
rect 13188 17134 13216 17167
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12256 16584 12308 16590
rect 12070 16552 12126 16561
rect 12256 16526 12308 16532
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12070 16487 12126 16496
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11702 15192 11758 15201
rect 11702 15127 11704 15136
rect 11756 15127 11758 15136
rect 11704 15098 11756 15104
rect 11900 15026 11928 15506
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14414 11928 14962
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 12084 14074 12112 16487
rect 12268 16114 12296 16526
rect 12360 16250 12388 16526
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12346 16144 12402 16153
rect 12256 16108 12308 16114
rect 12346 16079 12348 16088
rect 12256 16050 12308 16056
rect 12400 16079 12402 16088
rect 12348 16050 12400 16056
rect 12162 14512 12218 14521
rect 12162 14447 12218 14456
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 13530 11928 13874
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11716 12850 11744 13126
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11704 12436 11756 12442
rect 11900 12434 11928 12922
rect 11900 12406 12020 12434
rect 11704 12378 11756 12384
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 10266 11652 11494
rect 11716 11286 11744 12378
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11624 8974 11652 9862
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11716 7818 11744 11222
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10062 11928 10950
rect 11992 10130 12020 12406
rect 12072 12300 12124 12306
rect 12176 12288 12204 14447
rect 12360 13870 12388 16050
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14618 12480 14894
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12360 12782 12388 13806
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12452 12306 12480 14010
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12728 12850 12756 13330
rect 12820 12850 12848 13466
rect 13004 13326 13032 16526
rect 12992 13320 13044 13326
rect 13096 13297 13124 16594
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 12992 13262 13044 13268
rect 13082 13288 13138 13297
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12912 12986 12940 13126
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12636 12306 12664 12718
rect 12124 12260 12204 12288
rect 12440 12300 12492 12306
rect 12072 12242 12124 12248
rect 12440 12242 12492 12248
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12084 11830 12112 12242
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12636 11694 12664 12242
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 11286 12572 11494
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12084 10266 12112 11222
rect 12636 11218 12664 11630
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11992 9586 12020 10066
rect 12084 9586 12112 10202
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12452 8090 12480 8366
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 7478 11836 7686
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 11256 6886 11560 6914
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10980 5914 11008 6598
rect 11256 6458 11284 6886
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 6458 11376 6598
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11348 4758 11376 4966
rect 11532 4826 11560 4966
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11624 4622 11652 5646
rect 11716 5556 11744 6190
rect 11808 5710 11836 7414
rect 12544 6866 12572 11018
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12176 6118 12204 6734
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12452 6458 12480 6666
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11980 5568 12032 5574
rect 11716 5528 11980 5556
rect 11980 5510 12032 5516
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11808 2446 11836 4694
rect 11992 2514 12020 5510
rect 12176 5234 12204 6054
rect 12728 5370 12756 12786
rect 13004 12594 13032 13262
rect 13082 13223 13138 13232
rect 12912 12566 13032 12594
rect 12912 12238 12940 12566
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11898 12848 12038
rect 12912 11898 12940 12174
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 13004 11762 13032 12378
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13096 6186 13124 13223
rect 13280 11082 13308 16390
rect 13372 15502 13400 17750
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 16658 13860 17614
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13464 13394 13492 16458
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 14016 15706 14044 16050
rect 14108 15706 14136 21354
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14200 20330 14228 20810
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14292 19922 14320 20198
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14200 19446 14228 19654
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14292 19242 14320 19858
rect 14384 19802 14412 22066
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14568 22030 14596 22374
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14384 19774 14504 19802
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14384 18290 14412 19654
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14186 17368 14242 17377
rect 14186 17303 14242 17312
rect 14200 17270 14228 17303
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13924 15162 13952 15438
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14482 13952 14758
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13372 12442 13400 13194
rect 13556 12714 13584 13330
rect 14108 12850 14136 15438
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13372 12050 13400 12378
rect 13372 12022 13492 12050
rect 13464 11898 13492 12022
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13634 11792 13690 11801
rect 13634 11727 13690 11736
rect 13648 11694 13676 11727
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 13188 5914 13216 10610
rect 13556 7954 13584 11290
rect 14108 11150 14136 12786
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11830 14228 12038
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10810 13768 10950
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 14108 10606 14136 11086
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 13648 9586 13676 10542
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13924 9178 13952 9454
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14108 8566 14136 8774
rect 14292 8634 14320 16934
rect 14476 14958 14504 19774
rect 14660 19334 14688 22494
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14752 21321 14780 21626
rect 14738 21312 14794 21321
rect 14738 21247 14794 21256
rect 14844 20466 14872 22528
rect 15120 22438 15148 22607
rect 15488 22438 15516 22918
rect 15580 22710 15608 22918
rect 15568 22704 15620 22710
rect 15568 22646 15620 22652
rect 15672 22642 15700 23967
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15304 21894 15332 22374
rect 15660 21956 15712 21962
rect 15660 21898 15712 21904
rect 15292 21888 15344 21894
rect 15672 21865 15700 21898
rect 15292 21830 15344 21836
rect 15658 21856 15714 21865
rect 15658 21791 15714 21800
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 15028 19446 15056 20538
rect 15764 20466 15792 25350
rect 16028 25298 16080 25304
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15856 24750 15884 25230
rect 15948 25158 15976 25230
rect 16028 25220 16080 25226
rect 16028 25162 16080 25168
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15948 24410 15976 24550
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 15934 24304 15990 24313
rect 15934 24239 15990 24248
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15856 23866 15884 24142
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15948 23730 15976 24239
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 16040 23610 16068 25162
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 15844 23588 15896 23594
rect 15844 23530 15896 23536
rect 15948 23582 16068 23610
rect 15856 22234 15884 23530
rect 15948 22964 15976 23582
rect 16026 23488 16082 23497
rect 16026 23423 16082 23432
rect 16040 23254 16068 23423
rect 16028 23248 16080 23254
rect 16028 23190 16080 23196
rect 16040 23118 16068 23190
rect 16028 23112 16080 23118
rect 16132 23089 16160 24142
rect 16028 23054 16080 23060
rect 16118 23080 16174 23089
rect 16118 23015 16174 23024
rect 15948 22936 16068 22964
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15844 22228 15896 22234
rect 15844 22170 15896 22176
rect 15948 21554 15976 22374
rect 16040 22166 16068 22936
rect 16132 22817 16160 23015
rect 16118 22808 16174 22817
rect 16118 22743 16174 22752
rect 16028 22160 16080 22166
rect 16028 22102 16080 22108
rect 16224 22094 16252 29990
rect 16316 29646 16344 30223
rect 16408 30212 16528 30240
rect 16408 29850 16436 30212
rect 16486 30152 16542 30161
rect 16486 30087 16542 30096
rect 16396 29844 16448 29850
rect 16396 29786 16448 29792
rect 16408 29646 16436 29786
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16396 29640 16448 29646
rect 16396 29582 16448 29588
rect 16500 29238 16528 30087
rect 16578 29880 16634 29889
rect 16578 29815 16634 29824
rect 16592 29646 16620 29815
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 16684 29306 16712 31719
rect 16868 30258 16896 32370
rect 17038 32328 17094 32337
rect 17038 32263 17094 32272
rect 17052 31958 17080 32263
rect 17040 31952 17092 31958
rect 17144 31929 17172 34546
rect 17040 31894 17092 31900
rect 17130 31920 17186 31929
rect 17130 31855 17186 31864
rect 17144 31822 17172 31855
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 16948 30932 17000 30938
rect 16948 30874 17000 30880
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16856 30048 16908 30054
rect 16856 29990 16908 29996
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16488 29232 16540 29238
rect 16488 29174 16540 29180
rect 16304 29164 16356 29170
rect 16672 29164 16724 29170
rect 16304 29106 16356 29112
rect 16592 29124 16672 29152
rect 16316 28966 16344 29106
rect 16304 28960 16356 28966
rect 16356 28920 16436 28948
rect 16304 28902 16356 28908
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 16316 26994 16344 27270
rect 16408 27130 16436 28920
rect 16486 27432 16542 27441
rect 16486 27367 16542 27376
rect 16500 27334 16528 27367
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16396 27124 16448 27130
rect 16396 27066 16448 27072
rect 16304 26988 16356 26994
rect 16304 26930 16356 26936
rect 16304 26580 16356 26586
rect 16304 26522 16356 26528
rect 16316 25362 16344 26522
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16408 22710 16436 27066
rect 16500 26382 16528 27270
rect 16592 26874 16620 29124
rect 16672 29106 16724 29112
rect 16764 28484 16816 28490
rect 16764 28426 16816 28432
rect 16670 27704 16726 27713
rect 16670 27639 16726 27648
rect 16684 27538 16712 27639
rect 16672 27532 16724 27538
rect 16672 27474 16724 27480
rect 16776 27402 16804 28426
rect 16764 27396 16816 27402
rect 16764 27338 16816 27344
rect 16592 26846 16712 26874
rect 16488 26376 16540 26382
rect 16486 26344 16488 26353
rect 16540 26344 16542 26353
rect 16486 26279 16542 26288
rect 16684 25673 16712 26846
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16776 26586 16804 26726
rect 16764 26580 16816 26586
rect 16764 26522 16816 26528
rect 16868 25906 16896 29990
rect 16960 29209 16988 30874
rect 17236 30870 17264 34546
rect 17684 34536 17736 34542
rect 17684 34478 17736 34484
rect 17696 33862 17724 34478
rect 17684 33856 17736 33862
rect 17684 33798 17736 33804
rect 17684 33652 17736 33658
rect 17684 33594 17736 33600
rect 17316 33516 17368 33522
rect 17316 33458 17368 33464
rect 17328 33289 17356 33458
rect 17314 33280 17370 33289
rect 17314 33215 17370 33224
rect 17328 32570 17356 33215
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 17420 32348 17448 33050
rect 17696 32910 17724 33594
rect 17880 33114 17908 34546
rect 17960 34400 18012 34406
rect 17960 34342 18012 34348
rect 17868 33108 17920 33114
rect 17868 33050 17920 33056
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 17500 32360 17552 32366
rect 17328 32320 17500 32348
rect 17224 30864 17276 30870
rect 17224 30806 17276 30812
rect 17040 30048 17092 30054
rect 17040 29990 17092 29996
rect 17052 29646 17080 29990
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 16946 29200 17002 29209
rect 16946 29135 17002 29144
rect 17040 29164 17092 29170
rect 16960 27470 16988 29135
rect 17040 29106 17092 29112
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 16960 27305 16988 27406
rect 16946 27296 17002 27305
rect 16946 27231 17002 27240
rect 17052 27062 17080 29106
rect 17144 28966 17172 29582
rect 17328 29510 17356 32320
rect 17500 32302 17552 32308
rect 17592 32360 17644 32366
rect 17592 32302 17644 32308
rect 17406 31920 17462 31929
rect 17406 31855 17408 31864
rect 17460 31855 17462 31864
rect 17408 31826 17460 31832
rect 17408 31476 17460 31482
rect 17408 31418 17460 31424
rect 17420 31278 17448 31418
rect 17408 31272 17460 31278
rect 17408 31214 17460 31220
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 17316 29300 17368 29306
rect 17316 29242 17368 29248
rect 17132 28960 17184 28966
rect 17328 28937 17356 29242
rect 17314 28928 17370 28937
rect 17132 28902 17184 28908
rect 17236 28886 17314 28914
rect 17236 28490 17264 28886
rect 17314 28863 17370 28872
rect 17224 28484 17276 28490
rect 17224 28426 17276 28432
rect 17132 28416 17184 28422
rect 17132 28358 17184 28364
rect 17144 27674 17172 28358
rect 17132 27668 17184 27674
rect 17132 27610 17184 27616
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17040 27056 17092 27062
rect 17040 26998 17092 27004
rect 17052 26761 17080 26998
rect 17144 26858 17172 27270
rect 17132 26852 17184 26858
rect 17132 26794 17184 26800
rect 17038 26752 17094 26761
rect 17038 26687 17094 26696
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16670 25664 16726 25673
rect 16670 25599 16726 25608
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16488 25220 16540 25226
rect 16488 25162 16540 25168
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16224 22066 16344 22094
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 16026 21176 16082 21185
rect 16026 21111 16082 21120
rect 16120 21140 16172 21146
rect 16040 21010 16068 21111
rect 16120 21082 16172 21088
rect 16028 21004 16080 21010
rect 16028 20946 16080 20952
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15856 20466 15884 20810
rect 15948 20602 15976 20878
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19553 15976 20198
rect 15934 19544 15990 19553
rect 15934 19479 15990 19488
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 14568 19306 14688 19334
rect 14568 17746 14596 19306
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14660 18426 14688 19110
rect 14844 18766 14872 19382
rect 15028 18766 15056 19382
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 15120 17678 15148 18090
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14844 17202 14872 17546
rect 15212 17542 15240 18906
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15304 18290 15332 18634
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15488 18426 15516 18566
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15396 17678 15424 18294
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15212 17202 15240 17478
rect 15304 17218 15332 17614
rect 15384 17332 15436 17338
rect 15488 17320 15516 18362
rect 15580 18290 15608 19110
rect 16040 18970 16068 20946
rect 16132 20058 16160 21082
rect 16316 21010 16344 22066
rect 16408 21690 16436 22646
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16224 20398 16252 20742
rect 16316 20398 16344 20946
rect 16500 20942 16528 25162
rect 16592 24818 16620 25434
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16684 24154 16712 25599
rect 16762 25528 16818 25537
rect 16868 25498 16896 25842
rect 16762 25463 16818 25472
rect 16856 25492 16908 25498
rect 16776 25430 16804 25463
rect 16856 25434 16908 25440
rect 16764 25424 16816 25430
rect 16816 25372 16896 25378
rect 16764 25366 16896 25372
rect 16776 25350 16896 25366
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 16776 24206 16804 25230
rect 16592 24126 16712 24154
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16592 22794 16620 24126
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16684 23905 16712 24006
rect 16670 23896 16726 23905
rect 16670 23831 16726 23840
rect 16684 22982 16712 23831
rect 16776 23798 16804 24142
rect 16764 23792 16816 23798
rect 16764 23734 16816 23740
rect 16868 23526 16896 25350
rect 16960 25294 16988 26386
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 17052 25906 17080 26182
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17040 25764 17092 25770
rect 17040 25706 17092 25712
rect 17052 25362 17080 25706
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16960 25158 16988 25230
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 17038 25120 17094 25129
rect 17038 25055 17094 25064
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 16960 23780 16988 24550
rect 17052 24449 17080 25055
rect 17144 24886 17172 26318
rect 17132 24880 17184 24886
rect 17132 24822 17184 24828
rect 17038 24440 17094 24449
rect 17038 24375 17094 24384
rect 17052 24342 17080 24375
rect 17236 24342 17264 28426
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 17328 27470 17356 28018
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17328 27169 17356 27406
rect 17314 27160 17370 27169
rect 17314 27095 17370 27104
rect 17420 26382 17448 31214
rect 17500 30728 17552 30734
rect 17500 30670 17552 30676
rect 17512 29170 17540 30670
rect 17604 30569 17632 32302
rect 17696 30802 17724 32846
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17880 32434 17908 32710
rect 17972 32570 18000 34342
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 18064 32484 18092 34546
rect 18156 34474 18184 34734
rect 18524 34610 18552 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19156 34740 19208 34746
rect 19156 34682 19208 34688
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 18604 34604 18656 34610
rect 18604 34546 18656 34552
rect 18144 34468 18196 34474
rect 18144 34410 18196 34416
rect 18616 34202 18644 34546
rect 18972 34400 19024 34406
rect 18972 34342 19024 34348
rect 18604 34196 18656 34202
rect 18604 34138 18656 34144
rect 18616 34048 18644 34138
rect 18984 34066 19012 34342
rect 18432 34020 18644 34048
rect 18972 34060 19024 34066
rect 18432 33658 18460 34020
rect 18972 34002 19024 34008
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18604 33856 18656 33862
rect 18604 33798 18656 33804
rect 18696 33856 18748 33862
rect 18696 33798 18748 33804
rect 18420 33652 18472 33658
rect 18420 33594 18472 33600
rect 18524 33454 18552 33798
rect 18512 33448 18564 33454
rect 18512 33390 18564 33396
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 18524 33114 18552 33254
rect 18236 33108 18288 33114
rect 18236 33050 18288 33056
rect 18512 33108 18564 33114
rect 18512 33050 18564 33056
rect 18144 32496 18196 32502
rect 18064 32456 18144 32484
rect 18144 32438 18196 32444
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 17774 32056 17830 32065
rect 17774 31991 17830 32000
rect 17684 30796 17736 30802
rect 17684 30738 17736 30744
rect 17788 30598 17816 31991
rect 17880 31958 17908 32370
rect 17868 31952 17920 31958
rect 17868 31894 17920 31900
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 17972 30705 18000 31758
rect 18156 31113 18184 32438
rect 18248 31958 18276 33050
rect 18616 32994 18644 33798
rect 18708 33522 18736 33798
rect 18696 33516 18748 33522
rect 18696 33458 18748 33464
rect 18984 33318 19012 34002
rect 19064 33584 19116 33590
rect 19064 33526 19116 33532
rect 18972 33312 19024 33318
rect 18972 33254 19024 33260
rect 18524 32966 18644 32994
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 18432 32745 18460 32846
rect 18418 32736 18474 32745
rect 18418 32671 18474 32680
rect 18418 32600 18474 32609
rect 18418 32535 18474 32544
rect 18432 32502 18460 32535
rect 18420 32496 18472 32502
rect 18420 32438 18472 32444
rect 18236 31952 18288 31958
rect 18236 31894 18288 31900
rect 18142 31104 18198 31113
rect 18142 31039 18198 31048
rect 18248 30784 18276 31894
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 18340 30938 18368 31758
rect 18524 31346 18552 32966
rect 18972 32904 19024 32910
rect 18972 32846 19024 32852
rect 18696 32836 18748 32842
rect 18696 32778 18748 32784
rect 18604 32428 18656 32434
rect 18604 32370 18656 32376
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18328 30932 18380 30938
rect 18328 30874 18380 30880
rect 18064 30756 18276 30784
rect 17958 30696 18014 30705
rect 17958 30631 18014 30640
rect 17776 30592 17828 30598
rect 17590 30560 17646 30569
rect 17776 30534 17828 30540
rect 17590 30495 17646 30504
rect 18064 30274 18092 30756
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 18248 30394 18276 30602
rect 18236 30388 18288 30394
rect 18236 30330 18288 30336
rect 17972 30246 18092 30274
rect 17868 29776 17920 29782
rect 17868 29718 17920 29724
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17604 28994 17632 29582
rect 17776 29028 17828 29034
rect 17604 28966 17724 28994
rect 17776 28970 17828 28976
rect 17684 28960 17736 28966
rect 17684 28902 17736 28908
rect 17590 28792 17646 28801
rect 17590 28727 17646 28736
rect 17604 27946 17632 28727
rect 17592 27940 17644 27946
rect 17592 27882 17644 27888
rect 17592 27668 17644 27674
rect 17592 27610 17644 27616
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17314 26208 17370 26217
rect 17314 26143 17370 26152
rect 17328 25974 17356 26143
rect 17316 25968 17368 25974
rect 17368 25916 17448 25922
rect 17316 25910 17448 25916
rect 17328 25894 17448 25910
rect 17316 25764 17368 25770
rect 17316 25706 17368 25712
rect 17040 24336 17092 24342
rect 17040 24278 17092 24284
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17130 24032 17186 24041
rect 17130 23967 17186 23976
rect 17040 23792 17092 23798
rect 16960 23752 17040 23780
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16776 23254 16804 23462
rect 16764 23248 16816 23254
rect 16764 23190 16816 23196
rect 16960 23118 16988 23752
rect 17040 23734 17092 23740
rect 17144 23662 17172 23967
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 17144 23322 17172 23462
rect 17132 23316 17184 23322
rect 17132 23258 17184 23264
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16946 22944 17002 22953
rect 16946 22879 17002 22888
rect 16592 22766 16804 22794
rect 16580 22704 16632 22710
rect 16580 22646 16632 22652
rect 16592 22506 16620 22646
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16132 19922 16160 19994
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 16224 18766 16252 19722
rect 16408 19242 16436 20878
rect 16500 20466 16528 20878
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16486 20360 16542 20369
rect 16486 20295 16542 20304
rect 16500 19514 16528 20295
rect 16684 20058 16712 22374
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16592 19689 16620 19790
rect 16578 19680 16634 19689
rect 16578 19615 16634 19624
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16776 19360 16804 22766
rect 16960 22642 16988 22879
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 16868 20874 16896 22578
rect 17236 22080 17264 24074
rect 17144 22052 17264 22080
rect 17144 20942 17172 22052
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17236 21690 17264 21898
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16868 20754 16896 20810
rect 17040 20800 17092 20806
rect 16868 20748 17040 20754
rect 16868 20742 17092 20748
rect 16868 20726 17080 20742
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16868 20058 16896 20198
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16960 19922 16988 20402
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16960 19378 16988 19858
rect 16948 19372 17000 19378
rect 16776 19332 16896 19360
rect 16762 19272 16818 19281
rect 16396 19236 16448 19242
rect 16868 19258 16896 19332
rect 16948 19314 17000 19320
rect 17052 19310 17080 20726
rect 17328 20618 17356 25706
rect 17420 25294 17448 25894
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17420 23497 17448 24210
rect 17406 23488 17462 23497
rect 17406 23423 17462 23432
rect 17408 23248 17460 23254
rect 17408 23190 17460 23196
rect 17420 22681 17448 23190
rect 17406 22672 17462 22681
rect 17406 22607 17462 22616
rect 17512 22094 17540 26726
rect 17604 25838 17632 27610
rect 17592 25832 17644 25838
rect 17592 25774 17644 25780
rect 17604 25158 17632 25774
rect 17592 25152 17644 25158
rect 17592 25094 17644 25100
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17604 22817 17632 24550
rect 17696 23866 17724 28902
rect 17788 28121 17816 28970
rect 17774 28112 17830 28121
rect 17774 28047 17830 28056
rect 17776 27872 17828 27878
rect 17880 27849 17908 29718
rect 17972 28014 18000 30246
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18052 29844 18104 29850
rect 18052 29786 18104 29792
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 17776 27814 17828 27820
rect 17866 27840 17922 27849
rect 17788 24138 17816 27814
rect 17866 27775 17922 27784
rect 17972 27470 18000 27950
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17958 26888 18014 26897
rect 17958 26823 18014 26832
rect 17972 26382 18000 26823
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 17880 26217 17908 26250
rect 17866 26208 17922 26217
rect 17866 26143 17922 26152
rect 17972 25906 18000 26318
rect 18064 26246 18092 29786
rect 18248 29782 18276 29990
rect 18236 29776 18288 29782
rect 18236 29718 18288 29724
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 18248 29510 18276 29582
rect 18144 29504 18196 29510
rect 18144 29446 18196 29452
rect 18236 29504 18288 29510
rect 18236 29446 18288 29452
rect 18156 29102 18184 29446
rect 18340 29102 18368 30126
rect 18432 30054 18460 30670
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18144 29096 18196 29102
rect 18144 29038 18196 29044
rect 18328 29096 18380 29102
rect 18328 29038 18380 29044
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 18248 28257 18276 28426
rect 18234 28248 18290 28257
rect 18234 28183 18290 28192
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18156 27334 18184 27950
rect 18236 27872 18288 27878
rect 18236 27814 18288 27820
rect 18248 27713 18276 27814
rect 18234 27704 18290 27713
rect 18234 27639 18290 27648
rect 18236 27396 18288 27402
rect 18236 27338 18288 27344
rect 18144 27328 18196 27334
rect 18144 27270 18196 27276
rect 18156 27062 18184 27270
rect 18248 27062 18276 27338
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 18236 27056 18288 27062
rect 18236 26998 18288 27004
rect 18236 26308 18288 26314
rect 18156 26268 18236 26296
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17880 25537 17908 25774
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 17866 25528 17922 25537
rect 17866 25463 17922 25472
rect 18064 25362 18092 25638
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17880 24410 17908 24550
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17684 23656 17736 23662
rect 17684 23598 17736 23604
rect 17696 23186 17724 23598
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17590 22808 17646 22817
rect 17590 22743 17646 22752
rect 17590 22672 17646 22681
rect 17590 22607 17646 22616
rect 17604 22273 17632 22607
rect 17590 22264 17646 22273
rect 17590 22199 17646 22208
rect 17512 22066 17632 22094
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17144 20590 17356 20618
rect 17040 19304 17092 19310
rect 16868 19230 16988 19258
rect 17040 19246 17092 19252
rect 16762 19207 16818 19216
rect 16396 19178 16448 19184
rect 16578 18864 16634 18873
rect 16396 18828 16448 18834
rect 16578 18799 16580 18808
rect 16396 18770 16448 18776
rect 16632 18799 16634 18808
rect 16672 18828 16724 18834
rect 16580 18770 16632 18776
rect 16776 18816 16804 19207
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16724 18788 16804 18816
rect 16672 18770 16724 18776
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15580 17746 15608 18226
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15672 17882 15700 18022
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15672 17338 15700 17818
rect 15436 17292 15516 17320
rect 15384 17274 15436 17280
rect 15304 17202 15424 17218
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15292 17196 15424 17202
rect 15344 17190 15424 17196
rect 15292 17138 15344 17144
rect 15290 16824 15346 16833
rect 15200 16788 15252 16794
rect 15290 16759 15346 16768
rect 15200 16730 15252 16736
rect 15212 16454 15240 16730
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14568 14958 14596 16118
rect 14648 15428 14700 15434
rect 14648 15370 14700 15376
rect 14660 15178 14688 15370
rect 14922 15192 14978 15201
rect 14660 15150 14780 15178
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7002 13492 7686
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13556 6934 13584 7890
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13556 5778 13584 6870
rect 13740 6322 13768 8502
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13832 7886 13860 8366
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 7274 14320 7686
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14384 7154 14412 13942
rect 14476 11218 14504 14894
rect 14568 13734 14596 14894
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14752 11762 14780 15150
rect 14922 15127 14978 15136
rect 14936 14414 14964 15127
rect 15106 14784 15162 14793
rect 15028 14742 15106 14770
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14924 14272 14976 14278
rect 14922 14240 14924 14249
rect 14976 14240 14978 14249
rect 14922 14175 14978 14184
rect 15028 14074 15056 14742
rect 15106 14719 15162 14728
rect 15212 14618 15240 16186
rect 15304 16114 15332 16759
rect 15396 16590 15424 17190
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15488 16250 15516 17292
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15580 17134 15608 17274
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15660 16584 15712 16590
rect 15566 16552 15622 16561
rect 15660 16526 15712 16532
rect 15566 16487 15622 16496
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15120 13870 15148 14214
rect 15212 14074 15240 14554
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15028 12442 15056 12582
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15212 11762 15240 13874
rect 15304 12918 15332 14826
rect 15488 14362 15516 16050
rect 15396 14334 15516 14362
rect 15580 14346 15608 16487
rect 15672 15706 15700 16526
rect 15764 16114 15792 18090
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 16026 18048 16082 18057
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15948 16250 15976 18022
rect 16026 17983 16082 17992
rect 16040 16794 16068 17983
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 16132 16794 16160 17002
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16316 16726 16344 17546
rect 16304 16720 16356 16726
rect 16304 16662 16356 16668
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15568 14340 15620 14346
rect 15396 13954 15424 14334
rect 15568 14282 15620 14288
rect 15396 13926 15516 13954
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15396 12764 15424 13806
rect 15304 12736 15424 12764
rect 15304 11830 15332 12736
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15396 11898 15424 12582
rect 15488 12102 15516 13926
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15580 12434 15608 13874
rect 15672 12646 15700 15030
rect 15764 14958 15792 16050
rect 15842 15600 15898 15609
rect 15842 15535 15898 15544
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15764 13870 15792 14894
rect 15856 14006 15884 15535
rect 16040 14482 16068 16390
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16316 15026 16344 15302
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16118 14920 16174 14929
rect 16118 14855 16174 14864
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16132 14414 16160 14855
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15856 13569 15884 13942
rect 15948 13870 15976 14214
rect 16132 13870 16160 14214
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15842 13560 15898 13569
rect 15842 13495 15898 13504
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15580 12406 15700 12434
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14752 11082 14780 11698
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14740 11076 14792 11082
rect 14740 11018 14792 11024
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14476 10810 14504 10950
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 15028 10674 15056 11154
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15028 9674 15056 10610
rect 15028 9654 15240 9674
rect 15028 9648 15252 9654
rect 15028 9646 15200 9648
rect 15028 8838 15056 9646
rect 15200 9590 15252 9596
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15304 8650 15332 11766
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 14752 8634 15332 8650
rect 14752 8628 15344 8634
rect 14752 8622 15292 8628
rect 14752 8498 14780 8622
rect 15292 8570 15344 8576
rect 15014 8528 15070 8537
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14832 8492 14884 8498
rect 15014 8463 15016 8472
rect 14832 8434 14884 8440
rect 15068 8463 15070 8472
rect 15016 8434 15068 8440
rect 14568 8022 14596 8434
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14568 7478 14596 7958
rect 14752 7818 14780 8434
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14844 7410 14872 8434
rect 15028 7886 15056 8434
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14936 7392 14964 7754
rect 15016 7404 15068 7410
rect 14936 7364 15016 7392
rect 14292 7126 14412 7154
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13832 6458 13860 6666
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6458 14136 6598
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12176 4690 12204 5170
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12452 4826 12480 5102
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 13096 4622 13124 5510
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13556 3738 13584 5714
rect 13832 5642 13860 6394
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5778 14228 6054
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5302 13860 5578
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13924 5370 13952 5510
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 14200 4282 14228 5714
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3126 12940 3334
rect 13740 3194 13768 4082
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14108 3738 14136 4014
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 13740 2990 13768 3130
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 14292 2650 14320 7126
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14568 4214 14596 5578
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14568 3738 14596 4150
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14384 3126 14412 3334
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 14568 2922 14596 3674
rect 14844 3534 14872 7346
rect 14936 6662 14964 7364
rect 15016 7346 15068 7352
rect 15108 7404 15160 7410
rect 15212 7392 15240 7754
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15160 7364 15240 7392
rect 15108 7346 15160 7352
rect 15304 7206 15332 7482
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15396 6866 15424 11562
rect 15488 10810 15516 11698
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15580 10742 15608 11562
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15488 9722 15516 9862
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15580 9382 15608 9590
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15488 9178 15516 9318
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15672 8090 15700 12406
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15764 10112 15792 12038
rect 15856 10606 15884 13194
rect 15948 12481 15976 13670
rect 16040 13462 16068 13670
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16132 12714 16160 13126
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 15934 12472 15990 12481
rect 15934 12407 15990 12416
rect 15948 12306 15976 12407
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 10266 15884 10406
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15764 10084 15884 10112
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15856 7886 15884 10084
rect 15948 9654 15976 11018
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 16040 8537 16068 11698
rect 16132 9518 16160 12242
rect 16224 11898 16252 14350
rect 16316 13326 16344 14962
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16408 12374 16436 18770
rect 16592 18290 16620 18770
rect 16776 18290 16804 18788
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16500 16250 16528 16458
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16500 15162 16528 16186
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16500 13530 16528 14826
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16592 13002 16620 13194
rect 16500 12986 16620 13002
rect 16500 12980 16632 12986
rect 16500 12974 16580 12980
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16304 12232 16356 12238
rect 16500 12220 16528 12974
rect 16580 12922 16632 12928
rect 16356 12192 16528 12220
rect 16304 12174 16356 12180
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16304 12096 16356 12102
rect 16592 12050 16620 12106
rect 16304 12038 16356 12044
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16316 11082 16344 12038
rect 16500 12022 16620 12050
rect 16500 11626 16528 12022
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9722 16344 9862
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16026 8528 16082 8537
rect 16026 8463 16082 8472
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15936 7880 15988 7886
rect 16132 7834 16160 9454
rect 16500 8974 16528 10542
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16592 8974 16620 9522
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16224 8498 16252 8910
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16408 7886 16436 8026
rect 16500 7886 16528 8910
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16592 8566 16620 8774
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16592 7886 16620 8502
rect 16684 8022 16712 16594
rect 16776 16522 16804 17070
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16868 15450 16896 19110
rect 16960 18068 16988 19230
rect 17144 18272 17172 20590
rect 17408 20528 17460 20534
rect 17408 20470 17460 20476
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17236 19922 17264 20402
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17222 19816 17278 19825
rect 17328 19802 17356 20402
rect 17420 19854 17448 20470
rect 17278 19774 17356 19802
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17222 19751 17278 19760
rect 17420 19514 17448 19790
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17512 19258 17540 21082
rect 17328 19230 17540 19258
rect 17144 18244 17264 18272
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 17040 18080 17092 18086
rect 16960 18040 17040 18068
rect 17040 18022 17092 18028
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17052 15910 17080 16526
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 16868 15422 16988 15450
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16776 14822 16804 14962
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 14278 16804 14758
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16868 14074 16896 15302
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16960 14006 16988 15422
rect 17038 15056 17094 15065
rect 17038 14991 17094 15000
rect 17052 14822 17080 14991
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 17038 14648 17094 14657
rect 17038 14583 17094 14592
rect 17052 14414 17080 14583
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17144 14056 17172 18090
rect 17236 17202 17264 18244
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17328 16998 17356 19230
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17512 18766 17540 19110
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17116 17448 18022
rect 17512 17218 17540 18566
rect 17604 17338 17632 22066
rect 17788 22030 17816 22918
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17788 21554 17816 21830
rect 17880 21554 17908 23802
rect 17972 22273 18000 25298
rect 18156 24392 18184 26268
rect 18236 26250 18288 26256
rect 18340 26058 18368 29038
rect 18432 28218 18460 29990
rect 18524 28422 18552 31282
rect 18616 29889 18644 32370
rect 18708 32366 18736 32778
rect 18696 32360 18748 32366
rect 18696 32302 18748 32308
rect 18696 32224 18748 32230
rect 18696 32166 18748 32172
rect 18708 31822 18736 32166
rect 18696 31816 18748 31822
rect 18696 31758 18748 31764
rect 18788 31680 18840 31686
rect 18788 31622 18840 31628
rect 18696 30728 18748 30734
rect 18696 30670 18748 30676
rect 18602 29880 18658 29889
rect 18602 29815 18658 29824
rect 18616 29170 18644 29815
rect 18708 29714 18736 30670
rect 18800 30326 18828 31622
rect 18880 30796 18932 30802
rect 18880 30738 18932 30744
rect 18788 30320 18840 30326
rect 18788 30262 18840 30268
rect 18788 30184 18840 30190
rect 18788 30126 18840 30132
rect 18696 29708 18748 29714
rect 18696 29650 18748 29656
rect 18696 29504 18748 29510
rect 18696 29446 18748 29452
rect 18708 29186 18736 29446
rect 18800 29306 18828 30126
rect 18788 29300 18840 29306
rect 18788 29242 18840 29248
rect 18604 29164 18656 29170
rect 18708 29158 18828 29186
rect 18604 29106 18656 29112
rect 18604 28756 18656 28762
rect 18604 28698 18656 28704
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 18420 27940 18472 27946
rect 18420 27882 18472 27888
rect 18248 26030 18368 26058
rect 18248 24857 18276 26030
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18340 24954 18368 25842
rect 18432 25106 18460 27882
rect 18512 27668 18564 27674
rect 18616 27656 18644 28698
rect 18564 27628 18644 27656
rect 18512 27610 18564 27616
rect 18524 27470 18552 27610
rect 18602 27568 18658 27577
rect 18602 27503 18658 27512
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18616 27130 18644 27503
rect 18604 27124 18656 27130
rect 18800 27112 18828 29158
rect 18892 29102 18920 30738
rect 18984 29646 19012 32846
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 18880 29096 18932 29102
rect 18880 29038 18932 29044
rect 18972 28484 19024 28490
rect 18972 28426 19024 28432
rect 18880 28416 18932 28422
rect 18880 28358 18932 28364
rect 18892 28218 18920 28358
rect 18880 28212 18932 28218
rect 18880 28154 18932 28160
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18892 27656 18920 28018
rect 18984 27826 19012 28426
rect 19076 28218 19104 33526
rect 19168 30122 19196 34682
rect 19352 34462 19656 34490
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19260 33590 19288 33934
rect 19248 33584 19300 33590
rect 19248 33526 19300 33532
rect 19248 32564 19300 32570
rect 19248 32506 19300 32512
rect 19260 32026 19288 32506
rect 19248 32020 19300 32026
rect 19248 31962 19300 31968
rect 19352 31249 19380 34462
rect 19524 34400 19576 34406
rect 19524 34342 19576 34348
rect 19432 34060 19484 34066
rect 19432 34002 19484 34008
rect 19444 33969 19472 34002
rect 19430 33960 19486 33969
rect 19430 33895 19486 33904
rect 19536 33844 19564 34342
rect 19628 33998 19656 34462
rect 20088 34406 20116 37742
rect 20258 37703 20314 37712
rect 20364 36650 20392 40054
rect 20456 37942 20484 40122
rect 20536 39840 20588 39846
rect 20536 39782 20588 39788
rect 20548 39098 20576 39782
rect 20536 39092 20588 39098
rect 20536 39034 20588 39040
rect 20626 38992 20682 39001
rect 20536 38956 20588 38962
rect 20732 38962 20760 40326
rect 20824 40050 20852 40462
rect 21100 40390 21128 40870
rect 21468 40662 21496 41006
rect 21456 40656 21508 40662
rect 21652 40633 21680 41239
rect 21732 41210 21784 41216
rect 21744 41177 21772 41210
rect 21730 41168 21786 41177
rect 21730 41103 21786 41112
rect 21836 41041 21864 41386
rect 22020 41274 22048 41386
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 22112 41154 22140 41482
rect 21928 41126 22140 41154
rect 21822 41032 21878 41041
rect 21822 40967 21878 40976
rect 21928 40730 21956 41126
rect 22100 40928 22152 40934
rect 22100 40870 22152 40876
rect 21916 40724 21968 40730
rect 21916 40666 21968 40672
rect 21456 40598 21508 40604
rect 21638 40624 21694 40633
rect 21928 40594 21956 40666
rect 22006 40624 22062 40633
rect 21638 40559 21694 40568
rect 21916 40588 21968 40594
rect 22006 40559 22008 40568
rect 21916 40530 21968 40536
rect 22060 40559 22062 40568
rect 22008 40530 22060 40536
rect 21456 40452 21508 40458
rect 21456 40394 21508 40400
rect 21088 40384 21140 40390
rect 21088 40326 21140 40332
rect 20904 40112 20956 40118
rect 20904 40054 20956 40060
rect 20812 40044 20864 40050
rect 20812 39986 20864 39992
rect 20824 39846 20852 39986
rect 20812 39840 20864 39846
rect 20812 39782 20864 39788
rect 20812 39568 20864 39574
rect 20812 39510 20864 39516
rect 20626 38927 20682 38936
rect 20720 38956 20772 38962
rect 20536 38898 20588 38904
rect 20548 38486 20576 38898
rect 20640 38826 20668 38927
rect 20720 38898 20772 38904
rect 20628 38820 20680 38826
rect 20628 38762 20680 38768
rect 20536 38480 20588 38486
rect 20536 38422 20588 38428
rect 20444 37936 20496 37942
rect 20444 37878 20496 37884
rect 20548 37262 20576 38422
rect 20732 37874 20760 38898
rect 20720 37868 20772 37874
rect 20720 37810 20772 37816
rect 20732 37466 20760 37810
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 20824 37274 20852 39510
rect 20916 38418 20944 40054
rect 21468 39030 21496 40394
rect 21916 40384 21968 40390
rect 21916 40326 21968 40332
rect 21456 39024 21508 39030
rect 21456 38966 21508 38972
rect 21088 38888 21140 38894
rect 21088 38830 21140 38836
rect 20904 38412 20956 38418
rect 20904 38354 20956 38360
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20732 37246 20852 37274
rect 20536 37120 20588 37126
rect 20536 37062 20588 37068
rect 20444 36780 20496 36786
rect 20444 36722 20496 36728
rect 20352 36644 20404 36650
rect 20352 36586 20404 36592
rect 20168 36576 20220 36582
rect 20168 36518 20220 36524
rect 20180 36378 20208 36518
rect 20258 36408 20314 36417
rect 20168 36372 20220 36378
rect 20258 36343 20314 36352
rect 20168 36314 20220 36320
rect 20272 35873 20300 36343
rect 20364 36310 20392 36586
rect 20456 36378 20484 36722
rect 20444 36372 20496 36378
rect 20444 36314 20496 36320
rect 20352 36304 20404 36310
rect 20352 36246 20404 36252
rect 20456 36174 20484 36314
rect 20548 36174 20576 37062
rect 20628 36712 20680 36718
rect 20628 36654 20680 36660
rect 20640 36378 20668 36654
rect 20628 36372 20680 36378
rect 20628 36314 20680 36320
rect 20444 36168 20496 36174
rect 20444 36110 20496 36116
rect 20536 36168 20588 36174
rect 20536 36110 20588 36116
rect 20628 36100 20680 36106
rect 20628 36042 20680 36048
rect 20258 35864 20314 35873
rect 20258 35799 20314 35808
rect 20534 35864 20590 35873
rect 20640 35850 20668 36042
rect 20590 35822 20668 35850
rect 20534 35799 20590 35808
rect 20732 35714 20760 37246
rect 20996 37188 21048 37194
rect 20996 37130 21048 37136
rect 21008 36854 21036 37130
rect 20812 36848 20864 36854
rect 20810 36816 20812 36825
rect 20996 36848 21048 36854
rect 20864 36816 20866 36825
rect 20996 36790 21048 36796
rect 20810 36751 20866 36760
rect 20996 36712 21048 36718
rect 20810 36680 20866 36689
rect 20996 36654 21048 36660
rect 20810 36615 20866 36624
rect 20824 36174 20852 36615
rect 20812 36168 20864 36174
rect 20812 36110 20864 36116
rect 20548 35686 20760 35714
rect 20260 35080 20312 35086
rect 20260 35022 20312 35028
rect 20076 34400 20128 34406
rect 20076 34342 20128 34348
rect 20074 34232 20130 34241
rect 20074 34167 20130 34176
rect 19616 33992 19668 33998
rect 19616 33934 19668 33940
rect 19444 33816 19564 33844
rect 19984 33856 20036 33862
rect 19444 33538 19472 33816
rect 19984 33798 20036 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 33658 20024 33798
rect 19984 33652 20036 33658
rect 19984 33594 20036 33600
rect 19444 33510 19564 33538
rect 19536 32910 19564 33510
rect 19524 32904 19576 32910
rect 19524 32846 19576 32852
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19444 32065 19472 32370
rect 19616 32360 19668 32366
rect 20088 32348 20116 34167
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 20180 33862 20208 33934
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 20168 33584 20220 33590
rect 20168 33526 20220 33532
rect 19616 32302 19668 32308
rect 19996 32320 20116 32348
rect 19430 32056 19486 32065
rect 19430 31991 19486 32000
rect 19628 31686 19656 32302
rect 19892 32292 19944 32298
rect 19892 32234 19944 32240
rect 19708 32224 19760 32230
rect 19706 32192 19708 32201
rect 19760 32192 19762 32201
rect 19706 32127 19762 32136
rect 19720 31929 19748 32127
rect 19904 31958 19932 32234
rect 19892 31952 19944 31958
rect 19706 31920 19762 31929
rect 19892 31894 19944 31900
rect 19706 31855 19762 31864
rect 19996 31793 20024 32320
rect 19982 31784 20038 31793
rect 19982 31719 20038 31728
rect 19616 31680 19668 31686
rect 19616 31622 19668 31628
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19798 31376 19854 31385
rect 19996 31346 20024 31719
rect 20074 31648 20130 31657
rect 20074 31583 20130 31592
rect 19798 31311 19854 31320
rect 19984 31340 20036 31346
rect 19338 31240 19394 31249
rect 19338 31175 19394 31184
rect 19248 31136 19300 31142
rect 19248 31078 19300 31084
rect 19260 30938 19288 31078
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19352 30410 19380 31175
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19260 30382 19380 30410
rect 19156 30116 19208 30122
rect 19156 30058 19208 30064
rect 19156 29776 19208 29782
rect 19156 29718 19208 29724
rect 19168 29594 19196 29718
rect 19260 29594 19288 30382
rect 19444 30326 19472 30670
rect 19812 30666 19840 31311
rect 19984 31282 20036 31288
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19800 30660 19852 30666
rect 19800 30602 19852 30608
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19996 30258 20024 30670
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 19352 29850 19380 30194
rect 19800 30116 19852 30122
rect 19800 30058 19852 30064
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 19432 29776 19484 29782
rect 19432 29718 19484 29724
rect 19340 29640 19392 29646
rect 19168 29588 19340 29594
rect 19168 29582 19392 29588
rect 19168 29566 19380 29582
rect 19168 29209 19196 29566
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19154 29200 19210 29209
rect 19154 29135 19210 29144
rect 19260 28490 19288 29242
rect 19340 29232 19392 29238
rect 19338 29200 19340 29209
rect 19392 29200 19394 29209
rect 19338 29135 19394 29144
rect 19444 29050 19472 29718
rect 19812 29492 19840 30058
rect 20088 30002 20116 31583
rect 20180 30258 20208 33526
rect 20272 33046 20300 35022
rect 20352 33924 20404 33930
rect 20352 33866 20404 33872
rect 20364 33590 20392 33866
rect 20352 33584 20404 33590
rect 20352 33526 20404 33532
rect 20548 33522 20576 35686
rect 20628 35624 20680 35630
rect 20628 35566 20680 35572
rect 20536 33516 20588 33522
rect 20536 33458 20588 33464
rect 20260 33040 20312 33046
rect 20260 32982 20312 32988
rect 20258 32872 20314 32881
rect 20258 32807 20314 32816
rect 20272 30870 20300 32807
rect 20548 32416 20576 33458
rect 20456 32388 20576 32416
rect 20260 30864 20312 30870
rect 20260 30806 20312 30812
rect 20260 30660 20312 30666
rect 20260 30602 20312 30608
rect 20272 30569 20300 30602
rect 20258 30560 20314 30569
rect 20258 30495 20314 30504
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 20260 30116 20312 30122
rect 20260 30058 20312 30064
rect 19904 29974 20208 30002
rect 19904 29646 19932 29974
rect 19892 29640 19944 29646
rect 19892 29582 19944 29588
rect 20076 29504 20128 29510
rect 19812 29464 20024 29492
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19996 29170 20024 29464
rect 20076 29446 20128 29452
rect 19524 29164 19576 29170
rect 19524 29106 19576 29112
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19352 29022 19472 29050
rect 19352 28626 19380 29022
rect 19432 28756 19484 28762
rect 19536 28744 19564 29106
rect 19484 28716 19564 28744
rect 19432 28698 19484 28704
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 19996 28558 20024 29106
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19064 28212 19116 28218
rect 19064 28154 19116 28160
rect 19168 28082 19196 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19246 28248 19302 28257
rect 19574 28251 19882 28260
rect 19246 28183 19302 28192
rect 19524 28212 19576 28218
rect 19260 28150 19288 28183
rect 19524 28154 19576 28160
rect 19248 28144 19300 28150
rect 19248 28086 19300 28092
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19294 27872 19346 27878
rect 18984 27798 19104 27826
rect 19294 27814 19346 27820
rect 18972 27668 19024 27674
rect 18892 27628 18972 27656
rect 18972 27610 19024 27616
rect 18972 27396 19024 27402
rect 18892 27356 18972 27384
rect 18892 27305 18920 27356
rect 18972 27338 19024 27344
rect 18878 27296 18934 27305
rect 18878 27231 18934 27240
rect 18800 27084 18920 27112
rect 18604 27066 18656 27072
rect 18786 27024 18842 27033
rect 18786 26959 18788 26968
rect 18840 26959 18842 26968
rect 18788 26930 18840 26936
rect 18604 26852 18656 26858
rect 18604 26794 18656 26800
rect 18616 26450 18644 26794
rect 18788 26784 18840 26790
rect 18788 26726 18840 26732
rect 18604 26444 18656 26450
rect 18604 26386 18656 26392
rect 18510 26208 18566 26217
rect 18510 26143 18566 26152
rect 18524 25537 18552 26143
rect 18800 26081 18828 26726
rect 18602 26072 18658 26081
rect 18602 26007 18658 26016
rect 18786 26072 18842 26081
rect 18786 26007 18842 26016
rect 18510 25528 18566 25537
rect 18510 25463 18566 25472
rect 18512 25288 18564 25294
rect 18616 25276 18644 26007
rect 18892 25974 18920 27084
rect 19076 26874 19104 27798
rect 19306 27690 19334 27814
rect 19536 27713 19564 28154
rect 19168 27662 19334 27690
rect 19522 27704 19578 27713
rect 19168 27614 19196 27662
rect 19522 27639 19578 27648
rect 19168 27586 19288 27614
rect 18984 26846 19104 26874
rect 18880 25968 18932 25974
rect 18880 25910 18932 25916
rect 18564 25248 18644 25276
rect 18892 25242 18920 25910
rect 18512 25230 18564 25236
rect 18800 25214 18920 25242
rect 18432 25078 18644 25106
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18234 24848 18290 24857
rect 18234 24783 18236 24792
rect 18288 24783 18290 24792
rect 18236 24754 18288 24760
rect 18234 24712 18290 24721
rect 18234 24647 18290 24656
rect 18064 24364 18184 24392
rect 17958 22264 18014 22273
rect 17958 22199 18014 22208
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17788 21146 17816 21354
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17972 20942 18000 21286
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17696 20097 17724 20266
rect 17682 20088 17738 20097
rect 17682 20023 17738 20032
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17696 19378 17724 19722
rect 17788 19718 17816 20402
rect 17880 19854 17908 20742
rect 17960 20392 18012 20398
rect 17958 20360 17960 20369
rect 18012 20360 18014 20369
rect 17958 20295 18014 20304
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17774 19544 17830 19553
rect 17830 19502 17908 19530
rect 17774 19479 17830 19488
rect 17880 19446 17908 19502
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17696 18290 17724 18906
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17788 18290 17816 18566
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17880 18136 17908 18838
rect 17788 18108 17908 18136
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17512 17190 17724 17218
rect 17592 17128 17644 17134
rect 17420 17088 17540 17116
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17236 16250 17264 16594
rect 17512 16590 17540 17088
rect 17592 17070 17644 17076
rect 17604 16658 17632 17070
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17328 16046 17356 16458
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17224 15904 17276 15910
rect 17276 15864 17356 15892
rect 17224 15846 17276 15852
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17236 14414 17264 15370
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17236 14249 17264 14350
rect 17222 14240 17278 14249
rect 17222 14175 17278 14184
rect 17052 14028 17264 14056
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16960 13376 16988 13942
rect 17052 13938 17080 14028
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17144 13394 17172 13874
rect 17236 13394 17264 14028
rect 17132 13388 17184 13394
rect 16960 13348 17080 13376
rect 16762 13288 16818 13297
rect 16762 13223 16818 13232
rect 16948 13252 17000 13258
rect 16776 13190 16804 13223
rect 16948 13194 17000 13200
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16960 12850 16988 13194
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17052 11898 17080 13348
rect 17132 13330 17184 13336
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17052 11354 17080 11834
rect 17144 11558 17172 12922
rect 17236 11694 17264 13330
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17040 11348 17092 11354
rect 16960 11308 17040 11336
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16868 10674 16896 10950
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16776 9042 16804 9522
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16868 8974 16896 10610
rect 16960 10538 16988 11308
rect 17040 11290 17092 11296
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 17052 10985 17080 11018
rect 17038 10976 17094 10985
rect 17038 10911 17094 10920
rect 17144 10742 17172 11494
rect 17236 11014 17264 11630
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 17328 10418 17356 15864
rect 17420 15570 17448 16186
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17420 14278 17448 14962
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17406 14104 17462 14113
rect 17406 14039 17462 14048
rect 17420 13938 17448 14039
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17420 13394 17448 13874
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 16960 10390 17356 10418
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16776 7886 16804 8774
rect 16868 8090 16896 8910
rect 16960 8362 16988 10390
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17052 8974 17080 9522
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8537 17080 8910
rect 17144 8906 17172 9522
rect 17512 9178 17540 14554
rect 17604 9450 17632 15642
rect 17696 12986 17724 17190
rect 17788 16794 17816 18108
rect 17972 18034 18000 19654
rect 18064 19174 18092 24364
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 18156 22642 18184 22918
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 18248 22438 18276 24647
rect 18432 24585 18460 24890
rect 18512 24608 18564 24614
rect 18418 24576 18474 24585
rect 18512 24550 18564 24556
rect 18616 24562 18644 25078
rect 18694 24576 18750 24585
rect 18418 24511 18474 24520
rect 18328 24336 18380 24342
rect 18328 24278 18380 24284
rect 18340 22778 18368 24278
rect 18432 23610 18460 24511
rect 18524 24041 18552 24550
rect 18616 24534 18694 24562
rect 18694 24511 18750 24520
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18510 24032 18566 24041
rect 18510 23967 18566 23976
rect 18616 23866 18644 24210
rect 18708 24206 18736 24511
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18800 24052 18828 25214
rect 18880 25152 18932 25158
rect 18880 25094 18932 25100
rect 18708 24024 18828 24052
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18708 23644 18736 24024
rect 18892 23730 18920 25094
rect 18984 24070 19012 26846
rect 19064 26784 19116 26790
rect 19064 26726 19116 26732
rect 19076 26518 19104 26726
rect 19064 26512 19116 26518
rect 19064 26454 19116 26460
rect 19156 26308 19208 26314
rect 19260 26296 19288 27586
rect 19890 27568 19946 27577
rect 19946 27526 20024 27554
rect 19890 27503 19946 27512
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19208 26268 19288 26296
rect 19156 26250 19208 26256
rect 19352 26246 19380 26930
rect 19444 26874 19472 27338
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27062 20024 27526
rect 19984 27056 20036 27062
rect 19984 26998 20036 27004
rect 19444 26846 19564 26874
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19064 26240 19116 26246
rect 19064 26182 19116 26188
rect 19340 26240 19392 26246
rect 19340 26182 19392 26188
rect 18972 24064 19024 24070
rect 18972 24006 19024 24012
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 18616 23616 18736 23644
rect 18432 23594 18552 23610
rect 18432 23588 18564 23594
rect 18432 23582 18512 23588
rect 18512 23530 18564 23536
rect 18420 23520 18472 23526
rect 18616 23508 18644 23616
rect 18984 23594 19012 24006
rect 19076 23769 19104 26182
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 19352 25514 19380 25774
rect 19168 25486 19380 25514
rect 19062 23760 19118 23769
rect 19062 23695 19118 23704
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 18972 23588 19024 23594
rect 18972 23530 19024 23536
rect 18880 23520 18932 23526
rect 18616 23480 18828 23508
rect 18420 23462 18472 23468
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18432 22658 18460 23462
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18432 22642 18552 22658
rect 18616 22642 18644 23054
rect 18800 22982 18828 23480
rect 18880 23462 18932 23468
rect 18788 22976 18840 22982
rect 18694 22944 18750 22953
rect 18788 22918 18840 22924
rect 18694 22879 18750 22888
rect 18432 22636 18564 22642
rect 18432 22630 18512 22636
rect 18512 22578 18564 22584
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18156 21622 18184 22170
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 18156 21185 18184 21422
rect 18142 21176 18198 21185
rect 18248 21146 18276 22374
rect 18340 22030 18368 22510
rect 18604 22432 18656 22438
rect 18524 22392 18604 22420
rect 18418 22264 18474 22273
rect 18418 22199 18474 22208
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18432 21554 18460 22199
rect 18524 22098 18552 22392
rect 18604 22374 18656 22380
rect 18602 22264 18658 22273
rect 18602 22199 18658 22208
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 18616 21554 18644 22199
rect 18420 21548 18472 21554
rect 18420 21490 18472 21496
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18142 21111 18198 21120
rect 18236 21140 18288 21146
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18156 18970 18184 21111
rect 18236 21082 18288 21088
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18340 19922 18368 20742
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18340 19378 18368 19858
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18142 18864 18198 18873
rect 18142 18799 18198 18808
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17880 18006 18000 18034
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17788 16114 17816 16730
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17774 15736 17830 15745
rect 17774 15671 17830 15680
rect 17788 14550 17816 15671
rect 17776 14544 17828 14550
rect 17774 14512 17776 14521
rect 17828 14512 17830 14521
rect 17774 14447 17830 14456
rect 17774 14376 17830 14385
rect 17774 14311 17830 14320
rect 17788 13938 17816 14311
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17774 13832 17830 13841
rect 17774 13767 17776 13776
rect 17828 13767 17830 13776
rect 17776 13738 17828 13744
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17880 12850 17908 18006
rect 17960 17604 18012 17610
rect 17960 17546 18012 17552
rect 17972 15162 18000 17546
rect 18064 17202 18092 18566
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18064 16590 18092 17138
rect 18156 17066 18184 18799
rect 18234 18728 18290 18737
rect 18234 18663 18290 18672
rect 18248 18290 18276 18663
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 18156 16250 18184 17002
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 18156 15706 18184 16050
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18142 15600 18198 15609
rect 18142 15535 18198 15544
rect 18156 15502 18184 15535
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18052 15428 18104 15434
rect 18052 15370 18104 15376
rect 18064 15162 18092 15370
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17960 14952 18012 14958
rect 17958 14920 17960 14929
rect 18012 14920 18014 14929
rect 17958 14855 18014 14864
rect 18156 14482 18184 15302
rect 18248 14958 18276 15846
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18144 14476 18196 14482
rect 18064 14436 18144 14464
rect 18064 13938 18092 14436
rect 18144 14418 18196 14424
rect 18142 14240 18198 14249
rect 18142 14175 18198 14184
rect 18052 13932 18104 13938
rect 18156 13936 18184 14175
rect 18052 13874 18104 13880
rect 18144 13930 18196 13936
rect 18064 13841 18092 13874
rect 18144 13872 18196 13878
rect 18050 13832 18106 13841
rect 18050 13767 18106 13776
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 17960 13728 18012 13734
rect 18144 13728 18196 13734
rect 18012 13676 18144 13682
rect 18248 13705 18276 13738
rect 17960 13670 18196 13676
rect 18234 13696 18290 13705
rect 17972 13654 18184 13670
rect 18234 13631 18290 13640
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17972 11626 18000 12718
rect 18064 11626 18092 13330
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18248 12850 18276 13262
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18156 11762 18184 12310
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 18052 11620 18104 11626
rect 18052 11562 18104 11568
rect 18064 11286 18092 11562
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17972 9042 18000 11086
rect 18064 10742 18092 11222
rect 18156 11150 18184 11698
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18248 10810 18276 11290
rect 18340 11082 18368 18090
rect 18432 17626 18460 21082
rect 18524 19334 18552 21286
rect 18616 21146 18644 21286
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18524 19306 18644 19334
rect 18432 17598 18552 17626
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17338 18460 17478
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18432 15706 18460 15982
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18418 15600 18474 15609
rect 18418 15535 18474 15544
rect 18432 15502 18460 15535
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18418 15056 18474 15065
rect 18418 14991 18474 15000
rect 18432 14890 18460 14991
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18418 14648 18474 14657
rect 18418 14583 18474 14592
rect 18432 13802 18460 14583
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18524 12900 18552 17598
rect 18616 14113 18644 19306
rect 18708 18970 18736 22879
rect 18786 22808 18842 22817
rect 18786 22743 18842 22752
rect 18800 22642 18828 22743
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18788 22160 18840 22166
rect 18788 22102 18840 22108
rect 18800 21078 18828 22102
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18800 18170 18828 19110
rect 18892 18834 18920 23462
rect 19076 23118 19104 23598
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18984 20942 19012 22578
rect 19076 22030 19104 22918
rect 19168 22681 19196 25486
rect 19248 25424 19300 25430
rect 19248 25366 19300 25372
rect 19260 24070 19288 25366
rect 19444 25362 19472 26726
rect 19536 26382 19564 26846
rect 19996 26382 20024 26998
rect 19524 26376 19576 26382
rect 19524 26318 19576 26324
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 19984 26240 20036 26246
rect 19984 26182 20036 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19892 26036 19944 26042
rect 19892 25978 19944 25984
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19904 25226 19932 25978
rect 19996 25906 20024 26182
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19892 25220 19944 25226
rect 19892 25162 19944 25168
rect 19340 24948 19392 24954
rect 19444 24936 19472 25162
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19444 24908 19564 24936
rect 19340 24890 19392 24896
rect 19352 24818 19380 24890
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19352 24342 19380 24754
rect 19536 24750 19564 24908
rect 19628 24818 19840 24834
rect 20088 24818 20116 29446
rect 20180 29034 20208 29974
rect 20168 29028 20220 29034
rect 20168 28970 20220 28976
rect 20168 28552 20220 28558
rect 20168 28494 20220 28500
rect 20180 28393 20208 28494
rect 20166 28384 20222 28393
rect 20166 28319 20222 28328
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20180 24818 20208 26726
rect 19628 24812 19852 24818
rect 19628 24806 19800 24812
rect 19524 24744 19576 24750
rect 19524 24686 19576 24692
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19536 24206 19564 24686
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19340 24064 19392 24070
rect 19628 24052 19656 24806
rect 19800 24754 19852 24760
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 19708 24744 19760 24750
rect 19708 24686 19760 24692
rect 19720 24070 19748 24686
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 20088 24206 20116 24618
rect 19800 24200 19852 24206
rect 20076 24200 20128 24206
rect 20074 24168 20076 24177
rect 20128 24168 20130 24177
rect 19852 24148 20024 24154
rect 19800 24142 20024 24148
rect 19812 24126 20024 24142
rect 19340 24006 19392 24012
rect 19444 24024 19656 24052
rect 19708 24064 19760 24070
rect 19260 23866 19288 24006
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19246 22944 19302 22953
rect 19246 22879 19302 22888
rect 19154 22672 19210 22681
rect 19154 22607 19210 22616
rect 19260 22030 19288 22879
rect 19352 22710 19380 24006
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19352 22030 19380 22646
rect 19444 22438 19472 24024
rect 19708 24006 19760 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23848 20024 24126
rect 20074 24103 20130 24112
rect 20272 23848 20300 30058
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20364 29170 20392 29786
rect 20456 29170 20484 32388
rect 20536 32292 20588 32298
rect 20536 32234 20588 32240
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20444 29164 20496 29170
rect 20444 29106 20496 29112
rect 20456 28744 20484 29106
rect 20364 28716 20484 28744
rect 20364 28218 20392 28716
rect 20442 28656 20498 28665
rect 20442 28591 20498 28600
rect 20456 28558 20484 28591
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 20352 28212 20404 28218
rect 20352 28154 20404 28160
rect 20456 28082 20484 28494
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20548 26994 20576 32234
rect 20640 29238 20668 35566
rect 20904 34944 20956 34950
rect 20904 34886 20956 34892
rect 20812 34536 20864 34542
rect 20812 34478 20864 34484
rect 20718 34232 20774 34241
rect 20718 34167 20774 34176
rect 20732 34066 20760 34167
rect 20720 34060 20772 34066
rect 20720 34002 20772 34008
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20732 33522 20760 33798
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20824 33318 20852 34478
rect 20916 33522 20944 34886
rect 20904 33516 20956 33522
rect 20904 33458 20956 33464
rect 20812 33312 20864 33318
rect 20812 33254 20864 33260
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20732 31385 20760 32778
rect 20824 32586 20852 33254
rect 20916 32745 20944 33458
rect 20902 32736 20958 32745
rect 20902 32671 20958 32680
rect 20902 32600 20958 32609
rect 20824 32558 20902 32586
rect 20902 32535 20958 32544
rect 20904 32224 20956 32230
rect 20810 32192 20866 32201
rect 20904 32166 20956 32172
rect 20810 32127 20866 32136
rect 20824 32026 20852 32127
rect 20812 32020 20864 32026
rect 20812 31962 20864 31968
rect 20812 31884 20864 31890
rect 20812 31826 20864 31832
rect 20718 31376 20774 31385
rect 20718 31311 20774 31320
rect 20720 30116 20772 30122
rect 20720 30058 20772 30064
rect 20732 29646 20760 30058
rect 20824 30054 20852 31826
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20824 29646 20852 29990
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20824 29016 20852 29582
rect 20640 28988 20852 29016
rect 20640 28762 20668 28988
rect 20810 28792 20866 28801
rect 20628 28756 20680 28762
rect 20810 28727 20866 28736
rect 20628 28698 20680 28704
rect 20640 28558 20668 28698
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20732 28257 20760 28426
rect 20718 28248 20774 28257
rect 20718 28183 20774 28192
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 20640 27606 20668 27950
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20640 27130 20668 27338
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 20732 26994 20760 28018
rect 20824 27614 20852 28727
rect 20916 28014 20944 32166
rect 21008 31958 21036 36654
rect 21100 33522 21128 38830
rect 21180 38752 21232 38758
rect 21180 38694 21232 38700
rect 21192 38418 21220 38694
rect 21468 38654 21496 38966
rect 21732 38956 21784 38962
rect 21732 38898 21784 38904
rect 21548 38888 21600 38894
rect 21548 38830 21600 38836
rect 21640 38888 21692 38894
rect 21640 38830 21692 38836
rect 21560 38729 21588 38830
rect 21546 38720 21602 38729
rect 21546 38655 21602 38664
rect 21284 38626 21496 38654
rect 21180 38412 21232 38418
rect 21180 38354 21232 38360
rect 21180 38276 21232 38282
rect 21180 38218 21232 38224
rect 21192 37505 21220 38218
rect 21178 37496 21234 37505
rect 21178 37431 21234 37440
rect 21284 36786 21312 38626
rect 21560 38350 21588 38655
rect 21548 38344 21600 38350
rect 21548 38286 21600 38292
rect 21548 38208 21600 38214
rect 21548 38150 21600 38156
rect 21560 37942 21588 38150
rect 21548 37936 21600 37942
rect 21548 37878 21600 37884
rect 21364 37460 21416 37466
rect 21364 37402 21416 37408
rect 21376 37097 21404 37402
rect 21548 37392 21600 37398
rect 21548 37334 21600 37340
rect 21362 37088 21418 37097
rect 21362 37023 21418 37032
rect 21376 36786 21404 37023
rect 21560 36802 21588 37334
rect 21272 36780 21324 36786
rect 21272 36722 21324 36728
rect 21364 36780 21416 36786
rect 21364 36722 21416 36728
rect 21468 36774 21588 36802
rect 21270 36272 21326 36281
rect 21270 36207 21326 36216
rect 21284 35698 21312 36207
rect 21468 36122 21496 36774
rect 21548 36712 21600 36718
rect 21546 36680 21548 36689
rect 21600 36680 21602 36689
rect 21546 36615 21602 36624
rect 21560 36281 21588 36615
rect 21546 36272 21602 36281
rect 21546 36207 21602 36216
rect 21468 36094 21588 36122
rect 21560 35766 21588 36094
rect 21548 35760 21600 35766
rect 21548 35702 21600 35708
rect 21272 35692 21324 35698
rect 21272 35634 21324 35640
rect 21456 35012 21508 35018
rect 21456 34954 21508 34960
rect 21468 34746 21496 34954
rect 21456 34740 21508 34746
rect 21456 34682 21508 34688
rect 21180 34400 21232 34406
rect 21180 34342 21232 34348
rect 21192 34082 21220 34342
rect 21456 34128 21508 34134
rect 21192 34054 21312 34082
rect 21456 34070 21508 34076
rect 21560 34082 21588 35702
rect 21652 34610 21680 38830
rect 21744 37942 21772 38898
rect 21822 38584 21878 38593
rect 21822 38519 21878 38528
rect 21732 37936 21784 37942
rect 21732 37878 21784 37884
rect 21732 37800 21784 37806
rect 21732 37742 21784 37748
rect 21744 35698 21772 37742
rect 21732 35692 21784 35698
rect 21732 35634 21784 35640
rect 21640 34604 21692 34610
rect 21640 34546 21692 34552
rect 21652 34202 21680 34546
rect 21640 34196 21692 34202
rect 21640 34138 21692 34144
rect 21180 33992 21232 33998
rect 21180 33934 21232 33940
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 21088 33312 21140 33318
rect 21088 33254 21140 33260
rect 21100 32026 21128 33254
rect 21192 33114 21220 33934
rect 21284 33386 21312 34054
rect 21362 33688 21418 33697
rect 21362 33623 21364 33632
rect 21416 33623 21418 33632
rect 21364 33594 21416 33600
rect 21272 33380 21324 33386
rect 21272 33322 21324 33328
rect 21180 33108 21232 33114
rect 21180 33050 21232 33056
rect 21180 32428 21232 32434
rect 21180 32370 21232 32376
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 20996 31952 21048 31958
rect 21192 31906 21220 32370
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 21284 32026 21312 32302
rect 21376 32178 21404 33594
rect 21468 32910 21496 34070
rect 21560 34054 21680 34082
rect 21546 33552 21602 33561
rect 21546 33487 21602 33496
rect 21560 33454 21588 33487
rect 21548 33448 21600 33454
rect 21548 33390 21600 33396
rect 21652 33386 21680 34054
rect 21732 33584 21784 33590
rect 21732 33526 21784 33532
rect 21640 33380 21692 33386
rect 21640 33322 21692 33328
rect 21546 33280 21602 33289
rect 21546 33215 21602 33224
rect 21456 32904 21508 32910
rect 21456 32846 21508 32852
rect 21560 32502 21588 33215
rect 21640 33108 21692 33114
rect 21640 33050 21692 33056
rect 21548 32496 21600 32502
rect 21548 32438 21600 32444
rect 21652 32434 21680 33050
rect 21744 32910 21772 33526
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21732 32768 21784 32774
rect 21732 32710 21784 32716
rect 21640 32428 21692 32434
rect 21640 32370 21692 32376
rect 21376 32150 21680 32178
rect 21454 32056 21510 32065
rect 21272 32020 21324 32026
rect 21272 31962 21324 31968
rect 21364 32020 21416 32026
rect 21454 31991 21510 32000
rect 21364 31962 21416 31968
rect 21376 31906 21404 31962
rect 20996 31894 21048 31900
rect 21100 31878 21220 31906
rect 21284 31878 21404 31906
rect 21100 31804 21128 31878
rect 21284 31822 21312 31878
rect 21008 31776 21128 31804
rect 21272 31816 21324 31822
rect 20904 28008 20956 28014
rect 20904 27950 20956 27956
rect 20824 27586 20944 27614
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20364 25752 20392 26250
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20456 25974 20484 26182
rect 20548 25974 20576 26930
rect 20628 26784 20680 26790
rect 20628 26726 20680 26732
rect 20444 25968 20496 25974
rect 20444 25910 20496 25916
rect 20536 25968 20588 25974
rect 20536 25910 20588 25916
rect 20640 25906 20668 26726
rect 20732 26024 20760 26930
rect 20824 26450 20852 27474
rect 20812 26444 20864 26450
rect 20812 26386 20864 26392
rect 20732 25996 20852 26024
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20444 25764 20496 25770
rect 20364 25724 20444 25752
rect 20364 24614 20392 25724
rect 20444 25706 20496 25712
rect 20732 25498 20760 25842
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20628 25424 20680 25430
rect 20628 25366 20680 25372
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20352 24608 20404 24614
rect 20352 24550 20404 24556
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20364 24177 20392 24346
rect 20350 24168 20406 24177
rect 20350 24103 20406 24112
rect 19904 23820 20024 23848
rect 20088 23820 20300 23848
rect 19904 23633 19932 23820
rect 20088 23780 20116 23820
rect 19996 23752 20116 23780
rect 19890 23624 19946 23633
rect 19890 23559 19892 23568
rect 19944 23559 19946 23568
rect 19892 23530 19944 23536
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19524 22092 19576 22098
rect 19444 22052 19524 22080
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19076 21729 19104 21966
rect 19062 21720 19118 21729
rect 19062 21655 19118 21664
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 19076 20584 19104 21490
rect 19260 21418 19288 21966
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 18984 20556 19104 20584
rect 18984 20466 19012 20556
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 18970 20360 19026 20369
rect 18970 20295 19026 20304
rect 18984 19922 19012 20295
rect 19076 20058 19104 20402
rect 19352 20262 19380 21830
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19168 20058 19196 20198
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19444 19922 19472 22052
rect 19524 22034 19576 22040
rect 19616 22024 19668 22030
rect 19614 21992 19616 22001
rect 19668 21992 19670 22001
rect 19614 21927 19670 21936
rect 19904 21894 19932 22510
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19890 20904 19946 20913
rect 19890 20839 19946 20848
rect 19904 20806 19932 20839
rect 19996 20806 20024 23752
rect 20168 23724 20220 23730
rect 20088 23684 20168 23712
rect 20088 23118 20116 23684
rect 20168 23666 20220 23672
rect 20260 23588 20312 23594
rect 20260 23530 20312 23536
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 20168 23044 20220 23050
rect 20168 22986 20220 22992
rect 20074 22944 20130 22953
rect 20074 22879 20130 22888
rect 20088 22545 20116 22879
rect 20180 22710 20208 22986
rect 20168 22704 20220 22710
rect 20168 22646 20220 22652
rect 20272 22624 20300 23530
rect 20364 23254 20392 24103
rect 20456 24070 20484 24754
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20548 24188 20576 24346
rect 20640 24313 20668 25366
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20732 24721 20760 24754
rect 20718 24712 20774 24721
rect 20718 24647 20774 24656
rect 20824 24596 20852 25996
rect 20916 25906 20944 27586
rect 21008 27538 21036 31776
rect 21272 31758 21324 31764
rect 21364 31816 21416 31822
rect 21364 31758 21416 31764
rect 21180 31748 21232 31754
rect 21180 31690 21232 31696
rect 21192 31346 21220 31690
rect 21088 31340 21140 31346
rect 21088 31282 21140 31288
rect 21180 31340 21232 31346
rect 21180 31282 21232 31288
rect 21100 30977 21128 31282
rect 21086 30968 21142 30977
rect 21086 30903 21142 30912
rect 21088 29572 21140 29578
rect 21088 29514 21140 29520
rect 21100 27577 21128 29514
rect 21192 29238 21220 31282
rect 21376 31210 21404 31758
rect 21364 31204 21416 31210
rect 21364 31146 21416 31152
rect 21272 30864 21324 30870
rect 21272 30806 21324 30812
rect 21284 29238 21312 30806
rect 21364 30592 21416 30598
rect 21362 30560 21364 30569
rect 21416 30560 21418 30569
rect 21362 30495 21418 30504
rect 21180 29232 21232 29238
rect 21180 29174 21232 29180
rect 21272 29232 21324 29238
rect 21272 29174 21324 29180
rect 21376 29034 21404 30495
rect 21364 29028 21416 29034
rect 21192 28988 21364 29016
rect 21086 27568 21142 27577
rect 20996 27532 21048 27538
rect 21086 27503 21142 27512
rect 20996 27474 21048 27480
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20994 27296 21050 27305
rect 20994 27231 21050 27240
rect 21008 26790 21036 27231
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 21100 26217 21128 27406
rect 21192 26382 21220 28988
rect 21364 28970 21416 28976
rect 21362 28520 21418 28529
rect 21362 28455 21364 28464
rect 21416 28455 21418 28464
rect 21364 28426 21416 28432
rect 21376 27713 21404 28426
rect 21468 28014 21496 31991
rect 21652 31822 21680 32150
rect 21744 31890 21772 32710
rect 21732 31884 21784 31890
rect 21732 31826 21784 31832
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 21560 30734 21588 31282
rect 21548 30728 21600 30734
rect 21548 30670 21600 30676
rect 21548 29776 21600 29782
rect 21548 29718 21600 29724
rect 21638 29744 21694 29753
rect 21560 29646 21588 29718
rect 21638 29679 21694 29688
rect 21548 29640 21600 29646
rect 21548 29582 21600 29588
rect 21560 29481 21588 29582
rect 21546 29472 21602 29481
rect 21546 29407 21602 29416
rect 21652 29102 21680 29679
rect 21640 29096 21692 29102
rect 21640 29038 21692 29044
rect 21638 28792 21694 28801
rect 21638 28727 21694 28736
rect 21652 28558 21680 28727
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21548 28484 21600 28490
rect 21548 28426 21600 28432
rect 21456 28008 21508 28014
rect 21456 27950 21508 27956
rect 21362 27704 21418 27713
rect 21362 27639 21418 27648
rect 21364 27600 21416 27606
rect 21362 27568 21364 27577
rect 21416 27568 21418 27577
rect 21362 27503 21418 27512
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21364 27464 21416 27470
rect 21560 27418 21588 28426
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21652 27878 21680 28358
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21744 27418 21772 31826
rect 21364 27406 21416 27412
rect 21284 27130 21312 27406
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21272 26988 21324 26994
rect 21376 26976 21404 27406
rect 21324 26948 21404 26976
rect 21272 26930 21324 26936
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 21180 26376 21232 26382
rect 21284 26364 21312 26726
rect 21376 26518 21404 26948
rect 21468 27390 21588 27418
rect 21652 27390 21772 27418
rect 21364 26512 21416 26518
rect 21364 26454 21416 26460
rect 21284 26336 21404 26364
rect 21180 26318 21232 26324
rect 21086 26208 21142 26217
rect 21008 26166 21086 26194
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20916 25294 20944 25638
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20916 24750 20944 25230
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20732 24568 20852 24596
rect 20626 24304 20682 24313
rect 20626 24239 20682 24248
rect 20548 24160 20668 24188
rect 20444 24064 20496 24070
rect 20496 24024 20576 24052
rect 20444 24006 20496 24012
rect 20442 23896 20498 23905
rect 20442 23831 20498 23840
rect 20456 23730 20484 23831
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20352 23248 20404 23254
rect 20352 23190 20404 23196
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20364 22817 20392 22918
rect 20350 22808 20406 22817
rect 20350 22743 20406 22752
rect 20352 22636 20404 22642
rect 20272 22596 20352 22624
rect 20352 22578 20404 22584
rect 20074 22536 20130 22545
rect 20074 22471 20130 22480
rect 20350 22536 20406 22545
rect 20350 22471 20406 22480
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20088 22234 20116 22374
rect 20364 22250 20392 22471
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 20272 22222 20392 22250
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20088 21690 20116 21966
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 20180 21486 20208 21898
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20272 20942 20300 22222
rect 20456 21842 20484 23462
rect 20364 21814 20484 21842
rect 20364 21554 20392 21814
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 19892 20800 19944 20806
rect 19892 20742 19944 20748
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19522 20496 19578 20505
rect 19522 20431 19524 20440
rect 19576 20431 19578 20440
rect 19524 20402 19576 20408
rect 19996 20398 20024 20742
rect 20456 20602 20484 21626
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 19984 20392 20036 20398
rect 20036 20352 20116 20380
rect 19984 20334 20036 20340
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 20233 19656 20266
rect 19800 20256 19852 20262
rect 19614 20224 19670 20233
rect 19800 20198 19852 20204
rect 19614 20159 19670 20168
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 18984 19334 19012 19858
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19156 19372 19208 19378
rect 18984 19320 19156 19334
rect 18984 19314 19208 19320
rect 18984 19306 19196 19314
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18892 18290 18920 18770
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 19076 18290 19104 18566
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18800 18142 18920 18170
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18800 17746 18828 18022
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18788 17604 18840 17610
rect 18708 17564 18788 17592
rect 18708 17202 18736 17564
rect 18788 17546 18840 17552
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18892 15502 18920 18142
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 17678 19012 18022
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17377 19012 17478
rect 18970 17368 19026 17377
rect 18970 17303 19026 17312
rect 18984 17270 19012 17303
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18602 14104 18658 14113
rect 18602 14039 18658 14048
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18616 13841 18644 13874
rect 18602 13832 18658 13841
rect 18602 13767 18658 13776
rect 18604 12912 18656 12918
rect 18524 12872 18604 12900
rect 18604 12854 18656 12860
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11898 18552 12038
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 18432 10470 18460 11834
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18524 11150 18552 11630
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18524 10810 18552 11086
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18616 10606 18644 10950
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18616 10062 18644 10542
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17144 8634 17172 8842
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17316 8560 17368 8566
rect 17038 8528 17094 8537
rect 17316 8502 17368 8508
rect 17038 8463 17094 8472
rect 17052 8430 17080 8463
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 17328 7886 17356 8502
rect 17972 8498 18000 8978
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18432 8634 18460 8774
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7886 17448 8230
rect 15936 7822 15988 7828
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 5778 15056 6054
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 15580 4282 15608 7822
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15764 7410 15792 7754
rect 15856 7546 15884 7822
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15948 7410 15976 7822
rect 16040 7806 16160 7834
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 16040 6866 16068 7806
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16132 7546 16160 7686
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15856 6458 15884 6598
rect 15948 6458 15976 6734
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16040 6254 16068 6802
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16592 5914 16620 6802
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 15016 4276 15068 4282
rect 15016 4218 15068 4224
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14844 2854 14872 3470
rect 15028 3466 15056 4218
rect 15750 4040 15806 4049
rect 15750 3975 15806 3984
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15120 3670 15148 3878
rect 15672 3738 15700 3878
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15304 3126 15332 3334
rect 15488 3126 15516 3674
rect 15764 3534 15792 3975
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 16500 2922 16528 4218
rect 16592 4214 16620 4558
rect 16776 4282 16804 7822
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17236 7410 17264 7686
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17052 6866 17080 7346
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 17052 5914 17080 6190
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17328 5370 17356 7822
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16868 4282 16896 4490
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16592 3466 16620 4150
rect 17328 4146 17356 4218
rect 17696 4146 17724 6734
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17880 5778 17908 6598
rect 17972 6458 18000 8434
rect 18708 8430 18736 14486
rect 18800 14414 18828 15098
rect 18878 14920 18934 14929
rect 18878 14855 18934 14864
rect 18892 14414 18920 14855
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18800 14074 18828 14214
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 19076 13190 19104 18226
rect 19168 17610 19196 19306
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19260 16726 19288 18226
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19352 15026 19380 19654
rect 19444 19378 19472 19858
rect 19812 19854 19840 20198
rect 20088 19854 20116 20352
rect 20548 19922 20576 24024
rect 20640 23497 20668 24160
rect 20626 23488 20682 23497
rect 20626 23423 20682 23432
rect 20628 23112 20680 23118
rect 20626 23080 20628 23089
rect 20680 23080 20682 23089
rect 20626 23015 20682 23024
rect 20732 22642 20760 24568
rect 21008 24274 21036 26166
rect 21086 26143 21142 26152
rect 21086 25800 21142 25809
rect 21086 25735 21142 25744
rect 20996 24268 21048 24274
rect 20996 24210 21048 24216
rect 20902 24168 20958 24177
rect 20902 24103 20904 24112
rect 20956 24103 20958 24112
rect 20904 24074 20956 24080
rect 20810 24032 20866 24041
rect 20810 23967 20866 23976
rect 20824 23798 20852 23967
rect 20812 23792 20864 23798
rect 20812 23734 20864 23740
rect 21008 23730 21036 24210
rect 21100 24177 21128 25735
rect 21192 25498 21220 26318
rect 21270 26072 21326 26081
rect 21270 26007 21326 26016
rect 21284 25673 21312 26007
rect 21376 25838 21404 26336
rect 21364 25832 21416 25838
rect 21364 25774 21416 25780
rect 21270 25664 21326 25673
rect 21270 25599 21326 25608
rect 21180 25492 21232 25498
rect 21180 25434 21232 25440
rect 21468 25362 21496 27390
rect 21548 26988 21600 26994
rect 21548 26930 21600 26936
rect 21560 26042 21588 26930
rect 21548 26036 21600 26042
rect 21548 25978 21600 25984
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21376 24857 21404 25230
rect 21548 25152 21600 25158
rect 21548 25094 21600 25100
rect 21362 24848 21418 24857
rect 21272 24812 21324 24818
rect 21418 24806 21496 24834
rect 21362 24783 21418 24792
rect 21272 24754 21324 24760
rect 21180 24336 21232 24342
rect 21178 24304 21180 24313
rect 21232 24304 21234 24313
rect 21178 24239 21234 24248
rect 21284 24206 21312 24754
rect 21468 24274 21496 24806
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21272 24200 21324 24206
rect 21086 24168 21142 24177
rect 21272 24142 21324 24148
rect 21086 24103 21142 24112
rect 21456 24132 21508 24138
rect 21456 24074 21508 24080
rect 21178 23760 21234 23769
rect 20996 23724 21048 23730
rect 21234 23730 21312 23746
rect 21234 23724 21324 23730
rect 21234 23718 21272 23724
rect 21178 23695 21234 23704
rect 20996 23666 21048 23672
rect 21272 23666 21324 23672
rect 21088 23656 21140 23662
rect 21086 23624 21088 23633
rect 21180 23656 21232 23662
rect 21140 23624 21142 23633
rect 21180 23598 21232 23604
rect 21086 23559 21142 23568
rect 20810 23488 20866 23497
rect 20810 23423 20866 23432
rect 20824 23118 20852 23423
rect 21192 23254 21220 23598
rect 21180 23248 21232 23254
rect 20994 23216 21050 23225
rect 21180 23190 21232 23196
rect 20994 23151 21050 23160
rect 21008 23118 21036 23151
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20996 23112 21048 23118
rect 21088 23112 21140 23118
rect 20996 23054 21048 23060
rect 21086 23080 21088 23089
rect 21180 23112 21232 23118
rect 21140 23080 21142 23089
rect 21180 23054 21232 23060
rect 21086 23015 21142 23024
rect 20720 22636 20772 22642
rect 21192 22624 21220 23054
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 20720 22578 20772 22584
rect 21008 22596 21220 22624
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20640 22030 20668 22170
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20628 21616 20680 21622
rect 20626 21584 20628 21593
rect 20680 21584 20682 21593
rect 20626 21519 20682 21528
rect 20640 20466 20668 21519
rect 20732 20602 20760 22102
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 21008 20534 21036 22596
rect 21088 22160 21140 22166
rect 21086 22128 21088 22137
rect 21140 22128 21142 22137
rect 21086 22063 21142 22072
rect 21086 21992 21142 22001
rect 21376 21962 21404 22986
rect 21468 22234 21496 24074
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21086 21927 21142 21936
rect 21364 21956 21416 21962
rect 21100 21321 21128 21927
rect 21364 21898 21416 21904
rect 21560 21554 21588 25094
rect 21652 24954 21680 27390
rect 21732 25900 21784 25906
rect 21732 25842 21784 25848
rect 21744 25809 21772 25842
rect 21730 25800 21786 25809
rect 21730 25735 21786 25744
rect 21640 24948 21692 24954
rect 21640 24890 21692 24896
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21652 24206 21680 24550
rect 21744 24342 21772 25735
rect 21732 24336 21784 24342
rect 21732 24278 21784 24284
rect 21640 24200 21692 24206
rect 21640 24142 21692 24148
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21652 21486 21680 21626
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21086 21312 21142 21321
rect 21086 21247 21142 21256
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 20996 20528 21048 20534
rect 20996 20470 21048 20476
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 21008 20262 21036 20470
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 19800 19848 19852 19854
rect 19984 19848 20036 19854
rect 19852 19808 19984 19836
rect 19800 19790 19852 19796
rect 19984 19790 20036 19796
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19890 19272 19946 19281
rect 19890 19207 19946 19216
rect 19904 18970 19932 19207
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19444 18290 19472 18702
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20088 18290 20116 19382
rect 20180 19378 20208 19858
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20272 19378 20300 19722
rect 21376 19718 21404 20402
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 20640 19514 20668 19654
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20168 18760 20220 18766
rect 20166 18728 20168 18737
rect 20220 18728 20222 18737
rect 20166 18663 20222 18672
rect 20272 18290 20300 18906
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 19996 18086 20024 18226
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 17746 20024 18022
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 20088 17610 20116 18226
rect 20364 18170 20392 18226
rect 20180 18142 20392 18170
rect 20180 18086 20208 18142
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20180 17202 20208 17478
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19432 17060 19484 17066
rect 19432 17002 19484 17008
rect 19444 16153 19472 17002
rect 19996 16969 20024 17070
rect 20168 17060 20220 17066
rect 20168 17002 20220 17008
rect 20076 16992 20128 16998
rect 19982 16960 20038 16969
rect 20076 16934 20128 16940
rect 19982 16895 20038 16904
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19430 16144 19486 16153
rect 19430 16079 19486 16088
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19340 15020 19392 15026
rect 19444 15008 19472 15438
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19524 15020 19576 15026
rect 19444 14980 19524 15008
rect 19340 14962 19392 14968
rect 19524 14962 19576 14968
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19260 12850 19288 13126
rect 19352 12918 19380 13466
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 18800 11218 18828 12786
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18892 12238 18920 12582
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 11354 18920 11630
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 19076 11218 19104 12650
rect 19168 12170 19196 12650
rect 19352 12442 19380 12854
rect 19444 12481 19472 14826
rect 19812 14414 19840 15098
rect 20088 14958 20116 16934
rect 20180 16590 20208 17002
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20272 16590 20300 16934
rect 20364 16590 20392 18022
rect 20534 17368 20590 17377
rect 20534 17303 20590 17312
rect 20548 17270 20576 17303
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20456 16726 20484 17138
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20180 15910 20208 16526
rect 20364 16250 20392 16526
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20548 16114 20576 16458
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20534 15872 20590 15881
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20180 15026 20208 15506
rect 20272 15026 20300 15846
rect 20534 15807 20590 15816
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19812 14260 19840 14350
rect 19812 14232 20024 14260
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14074 20024 14232
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19536 13569 19564 13806
rect 19720 13569 19748 13942
rect 20088 13938 20116 14894
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19522 13560 19578 13569
rect 19522 13495 19578 13504
rect 19706 13560 19762 13569
rect 19706 13495 19762 13504
rect 20180 13394 20208 14962
rect 20444 14544 20496 14550
rect 20442 14512 20444 14521
rect 20496 14512 20498 14521
rect 20442 14447 20498 14456
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20456 13938 20484 14350
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19536 12889 19564 12922
rect 19522 12880 19578 12889
rect 20272 12850 20300 13738
rect 19522 12815 19578 12824
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 19430 12472 19486 12481
rect 19340 12436 19392 12442
rect 19430 12407 19486 12416
rect 19340 12378 19392 12384
rect 19444 12322 19472 12407
rect 19352 12294 19472 12322
rect 19996 12306 20024 12786
rect 19616 12300 19668 12306
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 18788 11212 18840 11218
rect 19064 11212 19116 11218
rect 18840 11172 18920 11200
rect 18788 11154 18840 11160
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18800 10810 18828 11018
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18892 10266 18920 11172
rect 19064 11154 19116 11160
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18892 10062 18920 10202
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18984 8974 19012 9318
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 19260 7834 19288 9930
rect 19352 9518 19380 12294
rect 19616 12242 19668 12248
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19628 12186 19656 12242
rect 20180 12238 20208 12786
rect 19444 12158 19656 12186
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 19444 11354 19472 12158
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19892 11620 19944 11626
rect 19892 11562 19944 11568
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19628 11218 19656 11494
rect 19904 11218 19932 11562
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19444 10742 19472 11086
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 8498 19380 9318
rect 19536 9178 19564 9590
rect 19996 9194 20024 10746
rect 20088 9654 20116 11086
rect 20180 11082 20208 12174
rect 20272 11830 20300 12786
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20272 10606 20300 11766
rect 20364 11393 20392 11834
rect 20456 11762 20484 13874
rect 20548 12073 20576 15807
rect 20534 12064 20590 12073
rect 20534 11999 20590 12008
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20350 11384 20406 11393
rect 20350 11319 20406 11328
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19524 9172 19576 9178
rect 19996 9166 20116 9194
rect 19524 9114 19576 9120
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19444 8430 19472 8910
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19720 7886 19748 8230
rect 19432 7880 19484 7886
rect 19260 7828 19432 7834
rect 19260 7822 19484 7828
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 19260 7806 19472 7822
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17960 5568 18012 5574
rect 18064 5556 18092 6258
rect 18012 5528 18092 5556
rect 17960 5510 18012 5516
rect 17774 4856 17830 4865
rect 17774 4791 17830 4800
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16592 3194 16620 3402
rect 16776 3194 16804 3878
rect 16960 3738 16988 4082
rect 17696 3738 17724 4082
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17788 3602 17816 4791
rect 17972 4622 18000 5510
rect 18340 4826 18368 7414
rect 18616 7410 18644 7754
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18616 6186 18644 7346
rect 19076 7206 19104 7686
rect 19260 7410 19288 7806
rect 19904 7732 19932 8298
rect 19996 7886 20024 9046
rect 20088 8498 20116 9166
rect 20180 8650 20208 10542
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20180 8634 20300 8650
rect 20168 8628 20300 8634
rect 20220 8622 20300 8628
rect 20168 8570 20220 8576
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19904 7704 20024 7732
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19168 6730 19196 7142
rect 19260 7002 19288 7346
rect 19890 7304 19946 7313
rect 19890 7239 19946 7248
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19904 6866 19932 7239
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 6254 18920 6598
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6322 20024 7704
rect 20180 6866 20208 8434
rect 20272 7410 20300 8622
rect 20364 8498 20392 10406
rect 20442 9616 20498 9625
rect 20442 9551 20498 9560
rect 20456 9518 20484 9551
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20456 6934 20484 9454
rect 20444 6928 20496 6934
rect 20496 6888 20576 6916
rect 20444 6870 20496 6876
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20180 6458 20208 6802
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 17866 3904 17922 3913
rect 17866 3839 17922 3848
rect 17880 3602 17908 3839
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 17696 2854 17724 3538
rect 17972 3126 18000 4558
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18432 4282 18460 4422
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18328 4140 18380 4146
rect 18380 4100 18460 4128
rect 18328 4082 18380 4088
rect 18432 3942 18460 4100
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18708 3738 18736 4218
rect 19076 4214 19104 4558
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 20088 4078 20116 5714
rect 20168 5636 20220 5642
rect 20168 5578 20220 5584
rect 20180 5370 20208 5578
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 20088 3602 20116 4014
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20088 3194 20116 3538
rect 20364 3534 20392 4422
rect 20456 4146 20484 6734
rect 20548 5370 20576 6888
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 20180 2990 20208 3334
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 17696 2446 17724 2790
rect 19522 2680 19578 2689
rect 19522 2615 19578 2624
rect 19536 2446 19564 2615
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 20640 2378 20668 19450
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20732 17066 20760 19246
rect 21376 18630 21404 19654
rect 21652 19378 21680 20878
rect 21744 20466 21772 24006
rect 21836 22710 21864 38519
rect 21928 38049 21956 40326
rect 22112 39914 22140 40870
rect 22204 40730 22232 41534
rect 22468 41482 22520 41488
rect 22664 41274 22692 41550
rect 23202 41511 23258 41520
rect 23216 41478 23244 41511
rect 22836 41472 22888 41478
rect 22836 41414 22888 41420
rect 23204 41472 23256 41478
rect 23204 41414 23256 41420
rect 22652 41268 22704 41274
rect 22652 41210 22704 41216
rect 22664 41070 22692 41210
rect 22376 41064 22428 41070
rect 22376 41006 22428 41012
rect 22652 41064 22704 41070
rect 22652 41006 22704 41012
rect 22192 40724 22244 40730
rect 22192 40666 22244 40672
rect 22388 40662 22416 41006
rect 22744 40928 22796 40934
rect 22744 40870 22796 40876
rect 22376 40656 22428 40662
rect 22376 40598 22428 40604
rect 22388 40458 22416 40598
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22376 40452 22428 40458
rect 22376 40394 22428 40400
rect 22284 40384 22336 40390
rect 22480 40361 22508 40462
rect 22652 40452 22704 40458
rect 22652 40394 22704 40400
rect 22284 40326 22336 40332
rect 22466 40352 22522 40361
rect 22100 39908 22152 39914
rect 22100 39850 22152 39856
rect 22190 39128 22246 39137
rect 22112 39086 22190 39114
rect 22008 38820 22060 38826
rect 22008 38762 22060 38768
rect 21914 38040 21970 38049
rect 21914 37975 21970 37984
rect 21916 36712 21968 36718
rect 21916 36654 21968 36660
rect 21928 36417 21956 36654
rect 21914 36408 21970 36417
rect 21914 36343 21970 36352
rect 21914 34776 21970 34785
rect 21914 34711 21970 34720
rect 21928 34474 21956 34711
rect 21916 34468 21968 34474
rect 21916 34410 21968 34416
rect 22020 33946 22048 38762
rect 22112 38758 22140 39086
rect 22190 39063 22246 39072
rect 22192 38956 22244 38962
rect 22192 38898 22244 38904
rect 22100 38752 22152 38758
rect 22100 38694 22152 38700
rect 22098 38448 22154 38457
rect 22098 38383 22154 38392
rect 22112 37233 22140 38383
rect 22204 37806 22232 38898
rect 22296 38894 22324 40326
rect 22466 40287 22522 40296
rect 22664 40186 22692 40394
rect 22652 40180 22704 40186
rect 22652 40122 22704 40128
rect 22466 39400 22522 39409
rect 22388 39358 22466 39386
rect 22388 39098 22416 39358
rect 22466 39335 22522 39344
rect 22376 39092 22428 39098
rect 22376 39034 22428 39040
rect 22284 38888 22336 38894
rect 22284 38830 22336 38836
rect 22388 38758 22416 39034
rect 22376 38752 22428 38758
rect 22560 38752 22612 38758
rect 22376 38694 22428 38700
rect 22480 38712 22560 38740
rect 22284 38208 22336 38214
rect 22284 38150 22336 38156
rect 22192 37800 22244 37806
rect 22192 37742 22244 37748
rect 22296 37652 22324 38150
rect 22376 37868 22428 37874
rect 22376 37810 22428 37816
rect 22204 37624 22324 37652
rect 22204 37330 22232 37624
rect 22284 37460 22336 37466
rect 22284 37402 22336 37408
rect 22192 37324 22244 37330
rect 22192 37266 22244 37272
rect 22098 37224 22154 37233
rect 22098 37159 22154 37168
rect 22112 36718 22140 37159
rect 22100 36712 22152 36718
rect 22100 36654 22152 36660
rect 22192 36712 22244 36718
rect 22192 36654 22244 36660
rect 22204 36378 22232 36654
rect 22192 36372 22244 36378
rect 22192 36314 22244 36320
rect 22192 36168 22244 36174
rect 22296 36122 22324 37402
rect 22388 36961 22416 37810
rect 22374 36952 22430 36961
rect 22374 36887 22430 36896
rect 22244 36116 22324 36122
rect 22192 36110 22324 36116
rect 22204 36094 22324 36110
rect 22296 35698 22324 36094
rect 22374 35864 22430 35873
rect 22374 35799 22430 35808
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 22388 35630 22416 35799
rect 22376 35624 22428 35630
rect 22376 35566 22428 35572
rect 22376 34740 22428 34746
rect 22480 34728 22508 38712
rect 22560 38694 22612 38700
rect 22560 38276 22612 38282
rect 22560 38218 22612 38224
rect 22572 36922 22600 38218
rect 22664 37942 22692 40122
rect 22756 39846 22784 40870
rect 22744 39840 22796 39846
rect 22744 39782 22796 39788
rect 22756 38350 22784 39782
rect 22848 38729 22876 41414
rect 23020 40996 23072 41002
rect 23020 40938 23072 40944
rect 22928 40452 22980 40458
rect 22928 40394 22980 40400
rect 22940 40361 22968 40394
rect 22926 40352 22982 40361
rect 22926 40287 22982 40296
rect 23032 40066 23060 40938
rect 23110 40624 23166 40633
rect 23110 40559 23166 40568
rect 23124 40526 23152 40559
rect 23112 40520 23164 40526
rect 23112 40462 23164 40468
rect 23204 40520 23256 40526
rect 23204 40462 23256 40468
rect 22940 40038 23060 40066
rect 22834 38720 22890 38729
rect 22834 38655 22890 38664
rect 22836 38480 22888 38486
rect 22836 38422 22888 38428
rect 22744 38344 22796 38350
rect 22744 38286 22796 38292
rect 22652 37936 22704 37942
rect 22652 37878 22704 37884
rect 22848 37874 22876 38422
rect 22836 37868 22888 37874
rect 22836 37810 22888 37816
rect 22744 37800 22796 37806
rect 22744 37742 22796 37748
rect 22650 37360 22706 37369
rect 22650 37295 22706 37304
rect 22560 36916 22612 36922
rect 22560 36858 22612 36864
rect 22560 36576 22612 36582
rect 22560 36518 22612 36524
rect 22572 36174 22600 36518
rect 22664 36174 22692 37295
rect 22756 37194 22784 37742
rect 22744 37188 22796 37194
rect 22744 37130 22796 37136
rect 22940 37074 22968 40038
rect 23216 39574 23244 40462
rect 23308 40458 23336 41618
rect 23492 41614 23520 42026
rect 24308 41676 24360 41682
rect 24308 41618 24360 41624
rect 23480 41608 23532 41614
rect 23478 41576 23480 41585
rect 24124 41608 24176 41614
rect 23532 41576 23534 41585
rect 24124 41550 24176 41556
rect 23478 41511 23534 41520
rect 24032 41540 24084 41546
rect 24032 41482 24084 41488
rect 23938 41304 23994 41313
rect 23938 41239 23994 41248
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 23400 40730 23428 41074
rect 23952 41070 23980 41239
rect 23940 41064 23992 41070
rect 23940 41006 23992 41012
rect 24044 40905 24072 41482
rect 24136 41070 24164 41550
rect 24124 41064 24176 41070
rect 24124 41006 24176 41012
rect 24030 40896 24086 40905
rect 24030 40831 24086 40840
rect 23754 40760 23810 40769
rect 23388 40724 23440 40730
rect 23754 40695 23810 40704
rect 23388 40666 23440 40672
rect 23768 40662 23796 40695
rect 24044 40662 24072 40831
rect 24136 40730 24164 41006
rect 24124 40724 24176 40730
rect 24124 40666 24176 40672
rect 23756 40656 23808 40662
rect 23676 40616 23756 40644
rect 23480 40588 23532 40594
rect 23480 40530 23532 40536
rect 23296 40452 23348 40458
rect 23296 40394 23348 40400
rect 23204 39568 23256 39574
rect 23204 39510 23256 39516
rect 23020 39500 23072 39506
rect 23020 39442 23072 39448
rect 23032 39030 23060 39442
rect 23020 39024 23072 39030
rect 23020 38966 23072 38972
rect 23308 38962 23336 40394
rect 23492 39930 23520 40530
rect 23676 40050 23704 40616
rect 23756 40598 23808 40604
rect 24032 40656 24084 40662
rect 24032 40598 24084 40604
rect 24122 40624 24178 40633
rect 24122 40559 24178 40568
rect 23754 40352 23810 40361
rect 23810 40310 23888 40338
rect 23754 40287 23810 40296
rect 23664 40044 23716 40050
rect 23664 39986 23716 39992
rect 23388 39908 23440 39914
rect 23492 39902 23704 39930
rect 23388 39850 23440 39856
rect 23204 38956 23256 38962
rect 23204 38898 23256 38904
rect 23296 38956 23348 38962
rect 23296 38898 23348 38904
rect 23020 38888 23072 38894
rect 23020 38830 23072 38836
rect 23032 37262 23060 38830
rect 23216 38350 23244 38898
rect 23308 38457 23336 38898
rect 23400 38894 23428 39850
rect 23572 39296 23624 39302
rect 23572 39238 23624 39244
rect 23480 38956 23532 38962
rect 23480 38898 23532 38904
rect 23388 38888 23440 38894
rect 23388 38830 23440 38836
rect 23294 38448 23350 38457
rect 23294 38383 23350 38392
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 23296 38344 23348 38350
rect 23400 38332 23428 38830
rect 23492 38418 23520 38898
rect 23480 38412 23532 38418
rect 23480 38354 23532 38360
rect 23348 38304 23428 38332
rect 23296 38286 23348 38292
rect 23308 38214 23336 38286
rect 23296 38208 23348 38214
rect 23296 38150 23348 38156
rect 23296 38004 23348 38010
rect 23296 37946 23348 37952
rect 23112 37936 23164 37942
rect 23112 37878 23164 37884
rect 23124 37262 23152 37878
rect 23308 37874 23336 37946
rect 23296 37868 23348 37874
rect 23296 37810 23348 37816
rect 23202 37768 23258 37777
rect 23202 37703 23258 37712
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 23112 37256 23164 37262
rect 23112 37198 23164 37204
rect 22756 37046 22968 37074
rect 22756 36786 22784 37046
rect 22834 36952 22890 36961
rect 22834 36887 22890 36896
rect 22848 36786 22876 36887
rect 23216 36854 23244 37703
rect 23388 37664 23440 37670
rect 23388 37606 23440 37612
rect 23480 37664 23532 37670
rect 23480 37606 23532 37612
rect 23400 37466 23428 37606
rect 23492 37466 23520 37606
rect 23388 37460 23440 37466
rect 23388 37402 23440 37408
rect 23480 37460 23532 37466
rect 23480 37402 23532 37408
rect 23308 37318 23520 37346
rect 23308 37233 23336 37318
rect 23492 37262 23520 37318
rect 23388 37256 23440 37262
rect 23294 37224 23350 37233
rect 23388 37198 23440 37204
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 23294 37159 23350 37168
rect 23400 37126 23428 37198
rect 23388 37120 23440 37126
rect 23386 37088 23388 37097
rect 23440 37088 23442 37097
rect 23386 37023 23442 37032
rect 23478 36952 23534 36961
rect 23478 36887 23534 36896
rect 23204 36848 23256 36854
rect 23204 36790 23256 36796
rect 23492 36786 23520 36887
rect 22744 36780 22796 36786
rect 22744 36722 22796 36728
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23018 36680 23074 36689
rect 23018 36615 23074 36624
rect 22928 36304 22980 36310
rect 22928 36246 22980 36252
rect 22560 36168 22612 36174
rect 22560 36110 22612 36116
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22664 35601 22692 36110
rect 22756 35834 22784 36110
rect 22744 35828 22796 35834
rect 22744 35770 22796 35776
rect 22940 35698 22968 36246
rect 23032 35834 23060 36615
rect 23296 36304 23348 36310
rect 23584 36258 23612 39238
rect 23676 37369 23704 39902
rect 23756 39568 23808 39574
rect 23756 39510 23808 39516
rect 23768 38758 23796 39510
rect 23860 38962 23888 40310
rect 24032 40112 24084 40118
rect 24032 40054 24084 40060
rect 24044 39302 24072 40054
rect 24136 40050 24164 40559
rect 24216 40520 24268 40526
rect 24216 40462 24268 40468
rect 24124 40044 24176 40050
rect 24124 39986 24176 39992
rect 24032 39296 24084 39302
rect 24032 39238 24084 39244
rect 23848 38956 23900 38962
rect 23848 38898 23900 38904
rect 23940 38956 23992 38962
rect 23940 38898 23992 38904
rect 23756 38752 23808 38758
rect 23756 38694 23808 38700
rect 23754 38448 23810 38457
rect 23754 38383 23810 38392
rect 23662 37360 23718 37369
rect 23662 37295 23718 37304
rect 23664 37188 23716 37194
rect 23664 37130 23716 37136
rect 23676 36310 23704 37130
rect 23296 36246 23348 36252
rect 23020 35828 23072 35834
rect 23020 35770 23072 35776
rect 23308 35698 23336 36246
rect 23492 36230 23612 36258
rect 23664 36304 23716 36310
rect 23664 36246 23716 36252
rect 22928 35692 22980 35698
rect 22928 35634 22980 35640
rect 23296 35692 23348 35698
rect 23296 35634 23348 35640
rect 23388 35692 23440 35698
rect 23388 35634 23440 35640
rect 22650 35592 22706 35601
rect 22650 35527 22706 35536
rect 22560 35012 22612 35018
rect 22560 34954 22612 34960
rect 22428 34700 22508 34728
rect 22376 34682 22428 34688
rect 22572 34678 22600 34954
rect 22560 34672 22612 34678
rect 22560 34614 22612 34620
rect 22664 34610 22692 35527
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22756 35290 22784 35430
rect 22940 35290 22968 35634
rect 22744 35284 22796 35290
rect 22744 35226 22796 35232
rect 22928 35284 22980 35290
rect 22928 35226 22980 35232
rect 23204 35080 23256 35086
rect 23204 35022 23256 35028
rect 22100 34604 22152 34610
rect 22652 34604 22704 34610
rect 22152 34564 22232 34592
rect 22100 34546 22152 34552
rect 21928 33918 22048 33946
rect 22100 33992 22152 33998
rect 22100 33934 22152 33940
rect 21928 32230 21956 33918
rect 22112 33522 22140 33934
rect 22100 33516 22152 33522
rect 22100 33458 22152 33464
rect 22008 32904 22060 32910
rect 22008 32846 22060 32852
rect 22020 32570 22048 32846
rect 22112 32570 22140 33458
rect 22008 32564 22060 32570
rect 22008 32506 22060 32512
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22100 32292 22152 32298
rect 22100 32234 22152 32240
rect 21916 32224 21968 32230
rect 21916 32166 21968 32172
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21928 30734 21956 31758
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22020 31124 22048 31622
rect 22112 31278 22140 32234
rect 22204 32042 22232 34564
rect 22652 34546 22704 34552
rect 22284 34468 22336 34474
rect 22284 34410 22336 34416
rect 22296 33998 22324 34410
rect 22928 34196 22980 34202
rect 22928 34138 22980 34144
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22836 33992 22888 33998
rect 22836 33934 22888 33940
rect 22652 33924 22704 33930
rect 22652 33866 22704 33872
rect 22560 33516 22612 33522
rect 22560 33458 22612 33464
rect 22284 33448 22336 33454
rect 22336 33408 22416 33436
rect 22284 33390 22336 33396
rect 22284 32224 22336 32230
rect 22282 32192 22284 32201
rect 22336 32192 22338 32201
rect 22282 32127 22338 32136
rect 22204 32014 22324 32042
rect 22190 31376 22246 31385
rect 22190 31311 22246 31320
rect 22100 31272 22152 31278
rect 22204 31260 22232 31311
rect 22152 31232 22232 31260
rect 22100 31214 22152 31220
rect 22020 31096 22232 31124
rect 22204 30938 22232 31096
rect 22192 30932 22244 30938
rect 22192 30874 22244 30880
rect 22296 30870 22324 32014
rect 22388 31754 22416 33408
rect 22572 32910 22600 33458
rect 22560 32904 22612 32910
rect 22480 32864 22560 32892
rect 22480 31958 22508 32864
rect 22560 32846 22612 32852
rect 22558 32600 22614 32609
rect 22558 32535 22614 32544
rect 22468 31952 22520 31958
rect 22468 31894 22520 31900
rect 22376 31748 22428 31754
rect 22572 31736 22600 32535
rect 22664 31958 22692 33866
rect 22848 33833 22876 33934
rect 22834 33824 22890 33833
rect 22834 33759 22890 33768
rect 22744 33652 22796 33658
rect 22744 33594 22796 33600
rect 22652 31952 22704 31958
rect 22652 31894 22704 31900
rect 22572 31708 22692 31736
rect 22376 31690 22428 31696
rect 22468 31476 22520 31482
rect 22468 31418 22520 31424
rect 22376 31340 22428 31346
rect 22376 31282 22428 31288
rect 22284 30864 22336 30870
rect 22284 30806 22336 30812
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 22100 30388 22152 30394
rect 22100 30330 22152 30336
rect 22112 29714 22140 30330
rect 22284 30184 22336 30190
rect 22284 30126 22336 30132
rect 22296 30025 22324 30126
rect 22282 30016 22338 30025
rect 22282 29951 22338 29960
rect 22190 29880 22246 29889
rect 22190 29815 22246 29824
rect 22100 29708 22152 29714
rect 22100 29650 22152 29656
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21928 29034 21956 29582
rect 22204 29345 22232 29815
rect 22284 29776 22336 29782
rect 22284 29718 22336 29724
rect 22296 29578 22324 29718
rect 22284 29572 22336 29578
rect 22284 29514 22336 29520
rect 22190 29336 22246 29345
rect 22190 29271 22246 29280
rect 21916 29028 21968 29034
rect 21916 28970 21968 28976
rect 22008 29028 22060 29034
rect 22008 28970 22060 28976
rect 21916 28416 21968 28422
rect 21916 28358 21968 28364
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21928 22098 21956 28358
rect 22020 26790 22048 28970
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 22204 25294 22232 29271
rect 22388 29152 22416 31282
rect 22480 30938 22508 31418
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22572 30938 22600 31214
rect 22468 30932 22520 30938
rect 22468 30874 22520 30880
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22664 30716 22692 31708
rect 22756 30734 22784 33594
rect 22940 33425 22968 34138
rect 23020 33856 23072 33862
rect 23020 33798 23072 33804
rect 23032 33590 23060 33798
rect 23216 33590 23244 35022
rect 23296 34944 23348 34950
rect 23296 34886 23348 34892
rect 23308 34066 23336 34886
rect 23400 34202 23428 35634
rect 23492 34728 23520 36230
rect 23572 36168 23624 36174
rect 23572 36110 23624 36116
rect 23664 36168 23716 36174
rect 23664 36110 23716 36116
rect 23584 35834 23612 36110
rect 23572 35828 23624 35834
rect 23572 35770 23624 35776
rect 23676 35698 23704 36110
rect 23664 35692 23716 35698
rect 23664 35634 23716 35640
rect 23492 34700 23612 34728
rect 23478 34232 23534 34241
rect 23388 34196 23440 34202
rect 23478 34167 23534 34176
rect 23388 34138 23440 34144
rect 23296 34060 23348 34066
rect 23296 34002 23348 34008
rect 23020 33584 23072 33590
rect 23020 33526 23072 33532
rect 23204 33584 23256 33590
rect 23204 33526 23256 33532
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 22926 33416 22982 33425
rect 22926 33351 22982 33360
rect 23020 33380 23072 33386
rect 23020 33322 23072 33328
rect 22928 33312 22980 33318
rect 22928 33254 22980 33260
rect 22940 33114 22968 33254
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 22836 32768 22888 32774
rect 23032 32722 23060 33322
rect 22836 32710 22888 32716
rect 22848 32230 22876 32710
rect 22940 32694 23060 32722
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22836 31952 22888 31958
rect 22836 31894 22888 31900
rect 22572 30688 22692 30716
rect 22744 30728 22796 30734
rect 22466 29744 22522 29753
rect 22466 29679 22468 29688
rect 22520 29679 22522 29688
rect 22468 29650 22520 29656
rect 22468 29504 22520 29510
rect 22572 29492 22600 30688
rect 22744 30670 22796 30676
rect 22744 30592 22796 30598
rect 22744 30534 22796 30540
rect 22756 30433 22784 30534
rect 22742 30424 22798 30433
rect 22848 30394 22876 31894
rect 22742 30359 22798 30368
rect 22836 30388 22888 30394
rect 22836 30330 22888 30336
rect 22834 30288 22890 30297
rect 22834 30223 22890 30232
rect 22652 30184 22704 30190
rect 22652 30126 22704 30132
rect 22664 29646 22692 30126
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22572 29464 22692 29492
rect 22468 29446 22520 29452
rect 22480 29322 22508 29446
rect 22480 29294 22600 29322
rect 22468 29164 22520 29170
rect 22388 29124 22468 29152
rect 22468 29106 22520 29112
rect 22480 29073 22508 29106
rect 22466 29064 22522 29073
rect 22284 29028 22336 29034
rect 22572 29034 22600 29294
rect 22466 28999 22522 29008
rect 22560 29028 22612 29034
rect 22284 28970 22336 28976
rect 22560 28970 22612 28976
rect 22296 27334 22324 28970
rect 22468 28960 22520 28966
rect 22466 28928 22468 28937
rect 22520 28928 22522 28937
rect 22466 28863 22522 28872
rect 22572 28608 22600 28970
rect 22480 28580 22600 28608
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22296 26382 22324 27270
rect 22388 27169 22416 27338
rect 22374 27160 22430 27169
rect 22374 27095 22430 27104
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22204 24818 22232 25094
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22112 24206 22140 24686
rect 22190 24440 22246 24449
rect 22190 24375 22246 24384
rect 22204 24342 22232 24375
rect 22192 24336 22244 24342
rect 22192 24278 22244 24284
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 22008 24064 22060 24070
rect 22008 24006 22060 24012
rect 22020 23361 22048 24006
rect 22006 23352 22062 23361
rect 22006 23287 22062 23296
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21928 21554 21956 22034
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 22020 21350 22048 22714
rect 22296 22642 22324 24686
rect 22374 24304 22430 24313
rect 22374 24239 22430 24248
rect 22388 24138 22416 24239
rect 22376 24132 22428 24138
rect 22376 24074 22428 24080
rect 22480 23118 22508 28580
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22572 27470 22600 28426
rect 22664 27946 22692 29464
rect 22756 29170 22784 29786
rect 22848 29714 22876 30223
rect 22940 29889 22968 32694
rect 23020 32564 23072 32570
rect 23020 32506 23072 32512
rect 23032 31822 23060 32506
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23124 31686 23152 33458
rect 23308 33386 23336 34002
rect 23388 33992 23440 33998
rect 23388 33934 23440 33940
rect 23400 33454 23428 33934
rect 23492 33658 23520 34167
rect 23584 34105 23612 34700
rect 23570 34096 23626 34105
rect 23570 34031 23572 34040
rect 23624 34031 23626 34040
rect 23572 34002 23624 34008
rect 23768 33810 23796 38383
rect 23860 36242 23888 38898
rect 23952 38554 23980 38898
rect 24032 38888 24084 38894
rect 24032 38830 24084 38836
rect 23940 38548 23992 38554
rect 23940 38490 23992 38496
rect 23848 36236 23900 36242
rect 23848 36178 23900 36184
rect 23952 36174 23980 38490
rect 23940 36168 23992 36174
rect 23940 36110 23992 36116
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 23676 33782 23796 33810
rect 23480 33652 23532 33658
rect 23480 33594 23532 33600
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 23296 33380 23348 33386
rect 23296 33322 23348 33328
rect 23204 32224 23256 32230
rect 23204 32166 23256 32172
rect 23112 31680 23164 31686
rect 23112 31622 23164 31628
rect 23124 31210 23152 31622
rect 23112 31204 23164 31210
rect 23112 31146 23164 31152
rect 23112 30932 23164 30938
rect 23112 30874 23164 30880
rect 23020 30660 23072 30666
rect 23020 30602 23072 30608
rect 23032 30394 23060 30602
rect 23124 30433 23152 30874
rect 23110 30424 23166 30433
rect 23020 30388 23072 30394
rect 23110 30359 23166 30368
rect 23020 30330 23072 30336
rect 22926 29880 22982 29889
rect 23216 29866 23244 32166
rect 23400 31328 23428 33390
rect 23492 31346 23520 33594
rect 23676 33114 23704 33782
rect 23756 33380 23808 33386
rect 23860 33368 23888 36042
rect 23952 35766 23980 36110
rect 23940 35760 23992 35766
rect 23940 35702 23992 35708
rect 23940 35624 23992 35630
rect 23940 35566 23992 35572
rect 23952 35290 23980 35566
rect 23940 35284 23992 35290
rect 23940 35226 23992 35232
rect 23940 33924 23992 33930
rect 23940 33866 23992 33872
rect 23952 33522 23980 33866
rect 24044 33658 24072 38830
rect 24136 38654 24164 39986
rect 24228 38865 24256 40462
rect 24320 40032 24348 41618
rect 24412 41478 24440 42026
rect 24492 41744 24544 41750
rect 24492 41686 24544 41692
rect 24400 41472 24452 41478
rect 24400 41414 24452 41420
rect 24412 41070 24440 41414
rect 24400 41064 24452 41070
rect 24400 41006 24452 41012
rect 24504 40712 24532 41686
rect 25596 41540 25648 41546
rect 25596 41482 25648 41488
rect 25872 41540 25924 41546
rect 25872 41482 25924 41488
rect 26240 41540 26292 41546
rect 26240 41482 26292 41488
rect 25320 41268 25372 41274
rect 25240 41228 25320 41256
rect 25042 41168 25098 41177
rect 25042 41103 25044 41112
rect 25096 41103 25098 41112
rect 25044 41074 25096 41080
rect 24768 40928 24820 40934
rect 24768 40870 24820 40876
rect 24504 40684 24624 40712
rect 24596 40594 24624 40684
rect 24584 40588 24636 40594
rect 24584 40530 24636 40536
rect 24596 40050 24624 40530
rect 24676 40520 24728 40526
rect 24676 40462 24728 40468
rect 24584 40044 24636 40050
rect 24320 40004 24532 40032
rect 24504 39817 24532 40004
rect 24584 39986 24636 39992
rect 24490 39808 24546 39817
rect 24490 39743 24546 39752
rect 24308 39500 24360 39506
rect 24308 39442 24360 39448
rect 24320 39302 24348 39442
rect 24308 39296 24360 39302
rect 24308 39238 24360 39244
rect 24320 38962 24348 39238
rect 24308 38956 24360 38962
rect 24308 38898 24360 38904
rect 24214 38856 24270 38865
rect 24214 38791 24270 38800
rect 24136 38626 24440 38654
rect 24412 37913 24440 38626
rect 24122 37904 24178 37913
rect 24122 37839 24124 37848
rect 24176 37839 24178 37848
rect 24398 37904 24454 37913
rect 24504 37874 24532 39743
rect 24398 37839 24454 37848
rect 24492 37868 24544 37874
rect 24124 37810 24176 37816
rect 24492 37810 24544 37816
rect 24122 37768 24178 37777
rect 24122 37703 24178 37712
rect 24136 34513 24164 37703
rect 24306 37496 24362 37505
rect 24306 37431 24362 37440
rect 24214 36952 24270 36961
rect 24214 36887 24270 36896
rect 24228 36854 24256 36887
rect 24216 36848 24268 36854
rect 24320 36825 24348 37431
rect 24492 37392 24544 37398
rect 24492 37334 24544 37340
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24216 36790 24268 36796
rect 24306 36816 24362 36825
rect 24306 36751 24308 36760
rect 24360 36751 24362 36760
rect 24308 36744 24360 36750
rect 24216 36712 24268 36718
rect 24268 36672 24348 36700
rect 24216 36654 24268 36660
rect 24122 34504 24178 34513
rect 24122 34439 24178 34448
rect 24216 34468 24268 34474
rect 24216 34410 24268 34416
rect 24124 33924 24176 33930
rect 24124 33866 24176 33872
rect 24032 33652 24084 33658
rect 24032 33594 24084 33600
rect 24044 33561 24072 33594
rect 24030 33552 24086 33561
rect 23940 33516 23992 33522
rect 24030 33487 24086 33496
rect 23940 33458 23992 33464
rect 23808 33340 23888 33368
rect 23940 33380 23992 33386
rect 23756 33322 23808 33328
rect 23940 33322 23992 33328
rect 23664 33108 23716 33114
rect 23664 33050 23716 33056
rect 23572 32496 23624 32502
rect 23572 32438 23624 32444
rect 22926 29815 22982 29824
rect 23124 29838 23244 29866
rect 23308 31300 23428 31328
rect 23480 31340 23532 31346
rect 22836 29708 22888 29714
rect 22836 29650 22888 29656
rect 22834 29608 22890 29617
rect 22834 29543 22890 29552
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22744 29028 22796 29034
rect 22744 28970 22796 28976
rect 22756 28762 22784 28970
rect 22744 28756 22796 28762
rect 22744 28698 22796 28704
rect 22744 28144 22796 28150
rect 22744 28086 22796 28092
rect 22652 27940 22704 27946
rect 22652 27882 22704 27888
rect 22560 27464 22612 27470
rect 22560 27406 22612 27412
rect 22652 27328 22704 27334
rect 22756 27316 22784 28086
rect 22704 27288 22784 27316
rect 22652 27270 22704 27276
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22756 26625 22784 26930
rect 22742 26616 22798 26625
rect 22652 26580 22704 26586
rect 22742 26551 22798 26560
rect 22652 26522 22704 26528
rect 22664 24206 22692 26522
rect 22744 26512 22796 26518
rect 22744 26454 22796 26460
rect 22756 25770 22784 26454
rect 22744 25764 22796 25770
rect 22744 25706 22796 25712
rect 22756 24750 22784 25706
rect 22848 24818 22876 29446
rect 22940 27606 22968 29815
rect 23124 29306 23152 29838
rect 23308 29730 23336 31300
rect 23480 31282 23532 31288
rect 23584 31226 23612 32438
rect 23676 32065 23704 33050
rect 23662 32056 23718 32065
rect 23662 31991 23718 32000
rect 23662 31920 23718 31929
rect 23662 31855 23718 31864
rect 23388 31204 23440 31210
rect 23388 31146 23440 31152
rect 23492 31198 23612 31226
rect 23676 31210 23704 31855
rect 23754 31512 23810 31521
rect 23754 31447 23810 31456
rect 23664 31204 23716 31210
rect 23216 29702 23336 29730
rect 23216 29646 23244 29702
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23296 29640 23348 29646
rect 23400 29594 23428 31146
rect 23492 30258 23520 31198
rect 23664 31146 23716 31152
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23492 30054 23520 30194
rect 23480 30048 23532 30054
rect 23480 29990 23532 29996
rect 23584 29782 23612 30194
rect 23572 29776 23624 29782
rect 23570 29744 23572 29753
rect 23624 29744 23626 29753
rect 23570 29679 23626 29688
rect 23348 29588 23428 29594
rect 23296 29582 23428 29588
rect 23308 29566 23428 29582
rect 23570 29608 23626 29617
rect 23570 29543 23572 29552
rect 23624 29543 23626 29552
rect 23572 29514 23624 29520
rect 23020 29300 23072 29306
rect 23020 29242 23072 29248
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 23032 28994 23060 29242
rect 23204 29096 23256 29102
rect 23124 29056 23204 29084
rect 23124 28994 23152 29056
rect 23204 29038 23256 29044
rect 23032 28966 23152 28994
rect 23020 28416 23072 28422
rect 23020 28358 23072 28364
rect 22928 27600 22980 27606
rect 22928 27542 22980 27548
rect 22926 27160 22982 27169
rect 22926 27095 22982 27104
rect 22940 26994 22968 27095
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 22928 26512 22980 26518
rect 22928 26454 22980 26460
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22742 24576 22798 24585
rect 22742 24511 22798 24520
rect 22756 24206 22784 24511
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22112 21962 22140 22442
rect 22296 22166 22324 22578
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 22756 22030 22784 23122
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 22652 21412 22704 21418
rect 22652 21354 22704 21360
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 21732 20460 21784 20466
rect 21732 20402 21784 20408
rect 21744 19922 21772 20402
rect 21732 19916 21784 19922
rect 21732 19858 21784 19864
rect 21744 19378 21772 19858
rect 21836 19378 21864 20470
rect 21928 19854 21956 20538
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22112 19854 22140 20334
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 21928 19378 21956 19790
rect 22296 19378 22324 19994
rect 22572 19854 22600 20470
rect 22664 20398 22692 21354
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22664 20262 22692 20334
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 21732 19236 21784 19242
rect 21732 19178 21784 19184
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21560 18290 21588 18838
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 21456 18216 21508 18222
rect 21456 18158 21508 18164
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20718 16688 20774 16697
rect 20718 16623 20774 16632
rect 20732 16046 20760 16623
rect 20824 16590 20852 17002
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16726 20944 16934
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 20916 16250 20944 16458
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20902 16144 20958 16153
rect 20812 16108 20864 16114
rect 20902 16079 20904 16088
rect 20812 16050 20864 16056
rect 20956 16079 20958 16088
rect 20904 16050 20956 16056
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20732 12986 20760 14962
rect 20824 14414 20852 16050
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20916 15706 20944 15914
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 21008 14482 21036 17206
rect 21100 16114 21128 17478
rect 21272 17264 21324 17270
rect 21272 17206 21324 17212
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21192 16046 21220 16526
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 21192 14278 21220 14894
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21180 14000 21232 14006
rect 21180 13942 21232 13948
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20916 13705 20944 13874
rect 20902 13696 20958 13705
rect 20902 13631 20958 13640
rect 21192 13546 21220 13942
rect 21284 13938 21312 17206
rect 21468 16794 21496 18158
rect 21744 17270 21772 19178
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21456 16788 21508 16794
rect 21508 16748 21588 16776
rect 21456 16730 21508 16736
rect 21364 16652 21416 16658
rect 21416 16612 21496 16640
rect 21364 16594 21416 16600
rect 21364 16516 21416 16522
rect 21364 16458 21416 16464
rect 21376 16182 21404 16458
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 21468 15502 21496 16612
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 20916 13518 21220 13546
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 11880 20760 12582
rect 20824 12374 20852 12718
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 20916 12050 20944 13518
rect 20996 13456 21048 13462
rect 20996 13398 21048 13404
rect 21008 12170 21036 13398
rect 21086 12880 21142 12889
rect 21086 12815 21088 12824
rect 21140 12815 21142 12824
rect 21088 12786 21140 12792
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 20916 12022 21036 12050
rect 20904 11892 20956 11898
rect 20732 11852 20852 11880
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20732 10266 20760 11562
rect 20824 11354 20852 11852
rect 20904 11834 20956 11840
rect 20916 11762 20944 11834
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20916 11082 20944 11698
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20824 10742 20852 11018
rect 20812 10736 20864 10742
rect 20812 10678 20864 10684
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20732 9586 20760 10202
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20916 8090 20944 11018
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 21008 7392 21036 12022
rect 21100 10538 21128 12786
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21192 11898 21220 12174
rect 21376 12170 21404 15302
rect 21560 15042 21588 16748
rect 21652 16658 21680 17002
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21468 15014 21588 15042
rect 21468 14074 21496 15014
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21560 14482 21588 14894
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21652 13954 21680 16594
rect 21744 15706 21772 16934
rect 21836 16726 21864 17138
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21928 15978 21956 18770
rect 22204 18766 22232 19314
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22296 18290 22324 19178
rect 22388 18970 22416 19246
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22374 18728 22430 18737
rect 22374 18663 22430 18672
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22100 17264 22152 17270
rect 22020 17224 22100 17252
rect 22020 16969 22048 17224
rect 22100 17206 22152 17212
rect 22006 16960 22062 16969
rect 22006 16895 22062 16904
rect 22020 16590 22048 16895
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21744 15502 21772 15642
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21560 13926 21680 13954
rect 21468 13258 21496 13874
rect 21456 13252 21508 13258
rect 21456 13194 21508 13200
rect 21560 12481 21588 13926
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21546 12472 21602 12481
rect 21546 12407 21602 12416
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21284 11830 21312 12106
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21192 11665 21220 11698
rect 21272 11688 21324 11694
rect 21178 11656 21234 11665
rect 21376 11676 21404 12106
rect 21468 11830 21496 12310
rect 21560 12238 21588 12407
rect 21652 12306 21680 13806
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21456 11824 21508 11830
rect 21456 11766 21508 11772
rect 21376 11648 21496 11676
rect 21272 11630 21324 11636
rect 21178 11591 21234 11600
rect 21284 11082 21312 11630
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11218 21404 11494
rect 21468 11218 21496 11648
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21560 11150 21588 12174
rect 21638 12064 21694 12073
rect 21638 11999 21694 12008
rect 21652 11665 21680 11999
rect 21638 11656 21694 11665
rect 21638 11591 21694 11600
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21652 11150 21680 11290
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21744 10996 21772 13670
rect 21836 13462 21864 15370
rect 21914 14648 21970 14657
rect 21914 14583 21916 14592
rect 21968 14583 21970 14592
rect 21916 14554 21968 14560
rect 21824 13456 21876 13462
rect 21824 13398 21876 13404
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21836 12102 21864 13262
rect 21914 12200 21970 12209
rect 21914 12135 21970 12144
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 11937 21864 12038
rect 21822 11928 21878 11937
rect 21928 11898 21956 12135
rect 21822 11863 21878 11872
rect 21916 11892 21968 11898
rect 21836 11558 21864 11863
rect 21916 11834 21968 11840
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21652 10968 21772 10996
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21468 9518 21496 10066
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21468 9042 21496 9318
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 21100 7886 21128 8026
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21192 7750 21220 8366
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21192 7426 21220 7686
rect 21284 7546 21312 7822
rect 21376 7546 21404 7822
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21192 7410 21312 7426
rect 21560 7410 21588 8434
rect 21652 7886 21680 10968
rect 21730 10840 21786 10849
rect 21730 10775 21786 10784
rect 21744 10062 21772 10775
rect 21824 10736 21876 10742
rect 21824 10678 21876 10684
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21088 7404 21140 7410
rect 21008 7364 21088 7392
rect 21192 7404 21324 7410
rect 21192 7398 21272 7404
rect 21088 7346 21140 7352
rect 21272 7346 21324 7352
rect 21364 7404 21416 7410
rect 21548 7404 21600 7410
rect 21416 7364 21496 7392
rect 21364 7346 21416 7352
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20916 4690 20944 5170
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20824 3738 20852 3878
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 20732 2650 20760 3402
rect 20916 3346 20944 3878
rect 21008 3466 21036 4558
rect 21100 4282 21128 7346
rect 21284 7002 21312 7346
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21376 6458 21404 6598
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21192 5710 21220 6258
rect 21468 5914 21496 7364
rect 21548 7346 21600 7352
rect 21560 6866 21588 7346
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21652 6730 21680 6938
rect 21744 6848 21772 9658
rect 21836 8090 21864 10678
rect 21928 9722 21956 11834
rect 22020 11830 22048 15642
rect 22098 15464 22154 15473
rect 22098 15399 22154 15408
rect 22112 15366 22140 15399
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 22098 14648 22154 14657
rect 22098 14583 22154 14592
rect 22112 14278 22140 14583
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22112 13274 22140 14214
rect 22204 13394 22232 18022
rect 22296 15502 22324 18022
rect 22388 17746 22416 18663
rect 22480 18154 22508 18906
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22572 17678 22600 19654
rect 22664 19378 22692 20198
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22848 19310 22876 20198
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22664 18170 22692 18566
rect 22744 18216 22796 18222
rect 22664 18164 22744 18170
rect 22664 18158 22796 18164
rect 22664 18142 22784 18158
rect 22664 17678 22692 18142
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22756 17882 22784 18022
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22848 17678 22876 19246
rect 22940 18902 22968 26454
rect 23032 25294 23060 28358
rect 23020 25288 23072 25294
rect 23020 25230 23072 25236
rect 23020 24404 23072 24410
rect 23020 24346 23072 24352
rect 23032 23769 23060 24346
rect 23124 24206 23152 28966
rect 23204 28756 23256 28762
rect 23204 28698 23256 28704
rect 23216 27674 23244 28698
rect 23570 28520 23626 28529
rect 23570 28455 23572 28464
rect 23624 28455 23626 28464
rect 23572 28426 23624 28432
rect 23480 28416 23532 28422
rect 23480 28358 23532 28364
rect 23204 27668 23256 27674
rect 23204 27610 23256 27616
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23216 26790 23244 26930
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 23308 26586 23336 27406
rect 23388 27396 23440 27402
rect 23388 27338 23440 27344
rect 23400 26858 23428 27338
rect 23388 26852 23440 26858
rect 23388 26794 23440 26800
rect 23296 26580 23348 26586
rect 23296 26522 23348 26528
rect 23492 25752 23520 28358
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23584 26450 23612 27406
rect 23572 26444 23624 26450
rect 23572 26386 23624 26392
rect 23308 25724 23520 25752
rect 23308 24410 23336 25724
rect 23386 25664 23442 25673
rect 23386 25599 23442 25608
rect 23296 24404 23348 24410
rect 23296 24346 23348 24352
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 23018 23760 23074 23769
rect 23018 23695 23074 23704
rect 23124 23526 23152 24142
rect 23308 23662 23336 24346
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 23308 22982 23336 23598
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23400 22817 23428 25599
rect 23676 25294 23704 31146
rect 23768 30841 23796 31447
rect 23848 31340 23900 31346
rect 23952 31328 23980 33322
rect 24136 32881 24164 33866
rect 24228 33522 24256 34410
rect 24320 34354 24348 36672
rect 24412 36378 24440 37062
rect 24400 36372 24452 36378
rect 24400 36314 24452 36320
rect 24504 35698 24532 37334
rect 24492 35692 24544 35698
rect 24492 35634 24544 35640
rect 24504 35086 24532 35634
rect 24596 35630 24624 39986
rect 24688 38418 24716 40462
rect 24780 39574 24808 40870
rect 25240 40633 25268 41228
rect 25320 41210 25372 41216
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25412 41132 25464 41138
rect 25412 41074 25464 41080
rect 25332 40905 25360 41074
rect 25318 40896 25374 40905
rect 25318 40831 25374 40840
rect 25320 40724 25372 40730
rect 25320 40666 25372 40672
rect 25226 40624 25282 40633
rect 25226 40559 25282 40568
rect 24860 40452 24912 40458
rect 24860 40394 24912 40400
rect 24768 39568 24820 39574
rect 24768 39510 24820 39516
rect 24872 39302 24900 40394
rect 25134 40080 25190 40089
rect 25134 40015 25190 40024
rect 24950 39400 25006 39409
rect 24950 39335 24952 39344
rect 25004 39335 25006 39344
rect 24952 39306 25004 39312
rect 24860 39296 24912 39302
rect 24860 39238 24912 39244
rect 25042 39264 25098 39273
rect 24768 38820 24820 38826
rect 24768 38762 24820 38768
rect 24780 38729 24808 38762
rect 24766 38720 24822 38729
rect 24766 38655 24822 38664
rect 24872 38418 24900 39238
rect 25042 39199 25098 39208
rect 25056 39030 25084 39199
rect 25148 39080 25176 40015
rect 25240 39642 25268 40559
rect 25332 40372 25360 40666
rect 25424 40526 25452 41074
rect 25412 40520 25464 40526
rect 25412 40462 25464 40468
rect 25412 40384 25464 40390
rect 25332 40344 25412 40372
rect 25412 40326 25464 40332
rect 25228 39636 25280 39642
rect 25228 39578 25280 39584
rect 25320 39636 25372 39642
rect 25320 39578 25372 39584
rect 25332 39545 25360 39578
rect 25318 39536 25374 39545
rect 25318 39471 25374 39480
rect 25318 39400 25374 39409
rect 25424 39386 25452 40326
rect 25504 39976 25556 39982
rect 25504 39918 25556 39924
rect 25374 39358 25452 39386
rect 25318 39335 25374 39344
rect 25318 39264 25374 39273
rect 25318 39199 25374 39208
rect 25148 39052 25268 39080
rect 25044 39024 25096 39030
rect 25044 38966 25096 38972
rect 25240 38962 25268 39052
rect 24952 38956 25004 38962
rect 24952 38898 25004 38904
rect 25228 38956 25280 38962
rect 25228 38898 25280 38904
rect 24676 38412 24728 38418
rect 24676 38354 24728 38360
rect 24860 38412 24912 38418
rect 24860 38354 24912 38360
rect 24676 37868 24728 37874
rect 24676 37810 24728 37816
rect 24688 36854 24716 37810
rect 24676 36848 24728 36854
rect 24676 36790 24728 36796
rect 24676 36644 24728 36650
rect 24676 36586 24728 36592
rect 24688 36174 24716 36586
rect 24872 36242 24900 38354
rect 24964 38214 24992 38898
rect 25044 38820 25096 38826
rect 25044 38762 25096 38768
rect 25056 38457 25084 38762
rect 25134 38720 25190 38729
rect 25134 38655 25190 38664
rect 25148 38554 25176 38655
rect 25332 38654 25360 39199
rect 25516 39098 25544 39918
rect 25608 39794 25636 41482
rect 25688 41200 25740 41206
rect 25688 41142 25740 41148
rect 25700 40594 25728 41142
rect 25688 40588 25740 40594
rect 25688 40530 25740 40536
rect 25780 40520 25832 40526
rect 25780 40462 25832 40468
rect 25792 39846 25820 40462
rect 25780 39840 25832 39846
rect 25608 39766 25728 39794
rect 25780 39782 25832 39788
rect 25700 39642 25728 39766
rect 25596 39636 25648 39642
rect 25596 39578 25648 39584
rect 25688 39636 25740 39642
rect 25688 39578 25740 39584
rect 25504 39092 25556 39098
rect 25504 39034 25556 39040
rect 25516 38962 25544 39034
rect 25504 38956 25556 38962
rect 25504 38898 25556 38904
rect 25410 38720 25466 38729
rect 25410 38655 25466 38664
rect 25240 38626 25360 38654
rect 25136 38548 25188 38554
rect 25136 38490 25188 38496
rect 25042 38448 25098 38457
rect 25042 38383 25098 38392
rect 25044 38344 25096 38350
rect 25044 38286 25096 38292
rect 24952 38208 25004 38214
rect 24952 38150 25004 38156
rect 24964 37806 24992 38150
rect 24952 37800 25004 37806
rect 24952 37742 25004 37748
rect 25056 37262 25084 38286
rect 25148 38282 25176 38490
rect 25136 38276 25188 38282
rect 25136 38218 25188 38224
rect 25136 37800 25188 37806
rect 25136 37742 25188 37748
rect 25044 37256 25096 37262
rect 25044 37198 25096 37204
rect 24952 36780 25004 36786
rect 24952 36722 25004 36728
rect 24860 36236 24912 36242
rect 24860 36178 24912 36184
rect 24676 36168 24728 36174
rect 24676 36110 24728 36116
rect 24964 36106 24992 36722
rect 25056 36378 25084 37198
rect 25148 36394 25176 37742
rect 25240 37398 25268 38626
rect 25320 38276 25372 38282
rect 25320 38218 25372 38224
rect 25228 37392 25280 37398
rect 25228 37334 25280 37340
rect 25240 36650 25268 37334
rect 25228 36644 25280 36650
rect 25228 36586 25280 36592
rect 25332 36530 25360 38218
rect 25424 37126 25452 38655
rect 25516 37398 25544 38898
rect 25608 38486 25636 39578
rect 25884 39438 25912 41482
rect 26252 41206 26280 41482
rect 26332 41268 26384 41274
rect 26332 41210 26384 41216
rect 26240 41200 26292 41206
rect 26240 41142 26292 41148
rect 26252 40934 26280 41142
rect 26240 40928 26292 40934
rect 26240 40870 26292 40876
rect 26056 40520 26108 40526
rect 26056 40462 26108 40468
rect 26068 40225 26096 40462
rect 26054 40216 26110 40225
rect 26054 40151 26110 40160
rect 26344 40050 26372 41210
rect 26056 40044 26108 40050
rect 26056 39986 26108 39992
rect 26332 40044 26384 40050
rect 26332 39986 26384 39992
rect 25964 39840 26016 39846
rect 25964 39782 26016 39788
rect 25872 39432 25924 39438
rect 25872 39374 25924 39380
rect 25688 39296 25740 39302
rect 25688 39238 25740 39244
rect 25780 39296 25832 39302
rect 25780 39238 25832 39244
rect 25596 38480 25648 38486
rect 25596 38422 25648 38428
rect 25700 38418 25728 39238
rect 25792 38554 25820 39238
rect 25884 38554 25912 39374
rect 25976 38894 26004 39782
rect 26068 39273 26096 39986
rect 26240 39568 26292 39574
rect 26240 39510 26292 39516
rect 26148 39432 26200 39438
rect 26148 39374 26200 39380
rect 26054 39264 26110 39273
rect 26054 39199 26110 39208
rect 26160 38962 26188 39374
rect 26056 38956 26108 38962
rect 26056 38898 26108 38904
rect 26148 38956 26200 38962
rect 26148 38898 26200 38904
rect 25964 38888 26016 38894
rect 25964 38830 26016 38836
rect 25976 38554 26004 38830
rect 25780 38548 25832 38554
rect 25780 38490 25832 38496
rect 25872 38548 25924 38554
rect 25872 38490 25924 38496
rect 25964 38548 26016 38554
rect 25964 38490 26016 38496
rect 25688 38412 25740 38418
rect 25688 38354 25740 38360
rect 25780 38344 25832 38350
rect 25780 38286 25832 38292
rect 25596 38004 25648 38010
rect 25596 37946 25648 37952
rect 25504 37392 25556 37398
rect 25504 37334 25556 37340
rect 25412 37120 25464 37126
rect 25412 37062 25464 37068
rect 25424 36786 25452 37062
rect 25516 36786 25544 37334
rect 25608 37262 25636 37946
rect 25792 37262 25820 38286
rect 25872 38276 25924 38282
rect 25872 38218 25924 38224
rect 25596 37256 25648 37262
rect 25596 37198 25648 37204
rect 25688 37256 25740 37262
rect 25688 37198 25740 37204
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 25608 36854 25636 37198
rect 25596 36848 25648 36854
rect 25596 36790 25648 36796
rect 25412 36780 25464 36786
rect 25412 36722 25464 36728
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 25332 36502 25544 36530
rect 25044 36372 25096 36378
rect 25148 36366 25360 36394
rect 25044 36314 25096 36320
rect 24952 36100 25004 36106
rect 24952 36042 25004 36048
rect 25056 35698 25084 36314
rect 25136 36100 25188 36106
rect 25136 36042 25188 36048
rect 25228 36100 25280 36106
rect 25228 36042 25280 36048
rect 25148 35698 25176 36042
rect 24676 35692 24728 35698
rect 24676 35634 24728 35640
rect 25044 35692 25096 35698
rect 25044 35634 25096 35640
rect 25136 35692 25188 35698
rect 25136 35634 25188 35640
rect 24584 35624 24636 35630
rect 24584 35566 24636 35572
rect 24596 35222 24624 35566
rect 24584 35216 24636 35222
rect 24584 35158 24636 35164
rect 24492 35080 24544 35086
rect 24492 35022 24544 35028
rect 24320 34326 24532 34354
rect 24308 34196 24360 34202
rect 24308 34138 24360 34144
rect 24320 33590 24348 34138
rect 24308 33584 24360 33590
rect 24308 33526 24360 33532
rect 24398 33552 24454 33561
rect 24216 33516 24268 33522
rect 24398 33487 24400 33496
rect 24216 33458 24268 33464
rect 24452 33487 24454 33496
rect 24400 33458 24452 33464
rect 24122 32872 24178 32881
rect 24122 32807 24178 32816
rect 24228 32570 24256 33458
rect 24412 33318 24440 33458
rect 24504 33318 24532 34326
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24596 33454 24624 33798
rect 24584 33448 24636 33454
rect 24584 33390 24636 33396
rect 24400 33312 24452 33318
rect 24306 33280 24362 33289
rect 24400 33254 24452 33260
rect 24492 33312 24544 33318
rect 24492 33254 24544 33260
rect 24306 33215 24362 33224
rect 24320 32910 24348 33215
rect 24308 32904 24360 32910
rect 24308 32846 24360 32852
rect 24216 32564 24268 32570
rect 24216 32506 24268 32512
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24228 31346 24256 32370
rect 24308 32292 24360 32298
rect 24308 32234 24360 32240
rect 23900 31300 23980 31328
rect 24032 31340 24084 31346
rect 23848 31282 23900 31288
rect 24032 31282 24084 31288
rect 24216 31340 24268 31346
rect 24216 31282 24268 31288
rect 23754 30832 23810 30841
rect 23754 30767 23810 30776
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23768 27606 23796 29990
rect 23756 27600 23808 27606
rect 23756 27542 23808 27548
rect 23768 26926 23796 27542
rect 23756 26920 23808 26926
rect 23756 26862 23808 26868
rect 23860 26518 23888 31282
rect 24044 30734 24072 31282
rect 24032 30728 24084 30734
rect 24032 30670 24084 30676
rect 24122 30696 24178 30705
rect 24044 30054 24072 30670
rect 24122 30631 24178 30640
rect 24032 30048 24084 30054
rect 24032 29990 24084 29996
rect 23940 29844 23992 29850
rect 23940 29786 23992 29792
rect 23952 29102 23980 29786
rect 24044 29714 24072 29990
rect 24032 29708 24084 29714
rect 24032 29650 24084 29656
rect 24030 29608 24086 29617
rect 24030 29543 24086 29552
rect 23940 29096 23992 29102
rect 23940 29038 23992 29044
rect 24044 27334 24072 29543
rect 24032 27328 24084 27334
rect 24032 27270 24084 27276
rect 24136 27146 24164 30631
rect 24228 28994 24256 31282
rect 24320 30938 24348 32234
rect 24400 31952 24452 31958
rect 24400 31894 24452 31900
rect 24308 30932 24360 30938
rect 24308 30874 24360 30880
rect 24412 30258 24440 31894
rect 24504 31226 24532 33254
rect 24596 33046 24624 33390
rect 24584 33040 24636 33046
rect 24584 32982 24636 32988
rect 24584 32904 24636 32910
rect 24584 32846 24636 32852
rect 24596 31958 24624 32846
rect 24688 31958 24716 35634
rect 25056 35086 25084 35634
rect 25044 35080 25096 35086
rect 25044 35022 25096 35028
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 25044 34944 25096 34950
rect 25044 34886 25096 34892
rect 24860 33516 24912 33522
rect 24780 33476 24860 33504
rect 24780 32434 24808 33476
rect 24860 33458 24912 33464
rect 24964 33318 24992 34886
rect 25056 34202 25084 34886
rect 25148 34202 25176 35634
rect 25240 34785 25268 36042
rect 25332 35193 25360 36366
rect 25412 36372 25464 36378
rect 25412 36314 25464 36320
rect 25424 36174 25452 36314
rect 25412 36168 25464 36174
rect 25412 36110 25464 36116
rect 25318 35184 25374 35193
rect 25318 35119 25374 35128
rect 25332 35068 25360 35119
rect 25412 35080 25464 35086
rect 25332 35040 25412 35068
rect 25412 35022 25464 35028
rect 25226 34776 25282 34785
rect 25226 34711 25282 34720
rect 25228 34536 25280 34542
rect 25228 34478 25280 34484
rect 25044 34196 25096 34202
rect 25044 34138 25096 34144
rect 25136 34196 25188 34202
rect 25136 34138 25188 34144
rect 25134 33552 25190 33561
rect 25134 33487 25136 33496
rect 25188 33487 25190 33496
rect 25136 33458 25188 33464
rect 24860 33312 24912 33318
rect 24860 33254 24912 33260
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 24768 32428 24820 32434
rect 24768 32370 24820 32376
rect 24584 31952 24636 31958
rect 24584 31894 24636 31900
rect 24676 31952 24728 31958
rect 24676 31894 24728 31900
rect 24872 31498 24900 33254
rect 24952 32904 25004 32910
rect 24952 32846 25004 32852
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 24964 32366 24992 32846
rect 24952 32360 25004 32366
rect 24952 32302 25004 32308
rect 25056 32298 25084 32846
rect 25148 32609 25176 33458
rect 25134 32600 25190 32609
rect 25134 32535 25190 32544
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 25044 32292 25096 32298
rect 25044 32234 25096 32240
rect 25042 31920 25098 31929
rect 24964 31878 25042 31906
rect 24964 31822 24992 31878
rect 25042 31855 25098 31864
rect 24952 31816 25004 31822
rect 25044 31816 25096 31822
rect 24952 31758 25004 31764
rect 25042 31784 25044 31793
rect 25096 31784 25098 31793
rect 24688 31470 24900 31498
rect 24688 31414 24716 31470
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24676 31272 24728 31278
rect 24504 31198 24624 31226
rect 24676 31214 24728 31220
rect 24492 31136 24544 31142
rect 24492 31078 24544 31084
rect 24504 30870 24532 31078
rect 24492 30864 24544 30870
rect 24492 30806 24544 30812
rect 24596 30274 24624 31198
rect 24688 30841 24716 31214
rect 24674 30832 24730 30841
rect 24674 30767 24730 30776
rect 24688 30666 24716 30767
rect 24676 30660 24728 30666
rect 24676 30602 24728 30608
rect 24780 30569 24808 31282
rect 24964 31142 24992 31758
rect 25042 31719 25098 31728
rect 25148 31385 25176 32438
rect 25240 32065 25268 34478
rect 25516 34082 25544 36502
rect 25608 36174 25636 36790
rect 25596 36168 25648 36174
rect 25596 36110 25648 36116
rect 25596 35760 25648 35766
rect 25596 35702 25648 35708
rect 25608 35086 25636 35702
rect 25596 35080 25648 35086
rect 25596 35022 25648 35028
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 25608 34542 25636 34886
rect 25596 34536 25648 34542
rect 25596 34478 25648 34484
rect 25424 34054 25544 34082
rect 25320 33516 25372 33522
rect 25320 33458 25372 33464
rect 25332 33318 25360 33458
rect 25320 33312 25372 33318
rect 25320 33254 25372 33260
rect 25320 32904 25372 32910
rect 25424 32892 25452 34054
rect 25504 33992 25556 33998
rect 25504 33934 25556 33940
rect 25516 33289 25544 33934
rect 25596 33516 25648 33522
rect 25596 33458 25648 33464
rect 25502 33280 25558 33289
rect 25502 33215 25558 33224
rect 25372 32864 25452 32892
rect 25608 32858 25636 33458
rect 25700 33454 25728 37198
rect 25780 36780 25832 36786
rect 25780 36722 25832 36728
rect 25792 33522 25820 36722
rect 25884 35834 25912 38218
rect 25976 37806 26004 38490
rect 25964 37800 26016 37806
rect 25964 37742 26016 37748
rect 25962 37496 26018 37505
rect 25962 37431 25964 37440
rect 26016 37431 26018 37440
rect 25964 37402 26016 37408
rect 25964 37324 26016 37330
rect 25964 37266 26016 37272
rect 25976 36854 26004 37266
rect 25964 36848 26016 36854
rect 25964 36790 26016 36796
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25976 36174 26004 36518
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 25976 35834 26004 36110
rect 25872 35828 25924 35834
rect 25872 35770 25924 35776
rect 25964 35828 26016 35834
rect 25964 35770 26016 35776
rect 25872 35080 25924 35086
rect 25870 35048 25872 35057
rect 25924 35048 25926 35057
rect 25870 34983 25926 34992
rect 26068 34746 26096 38898
rect 26148 38820 26200 38826
rect 26148 38762 26200 38768
rect 26160 38350 26188 38762
rect 26252 38758 26280 39510
rect 26240 38752 26292 38758
rect 26240 38694 26292 38700
rect 26148 38344 26200 38350
rect 26148 38286 26200 38292
rect 26344 37262 26372 39986
rect 26436 38593 26464 43864
rect 30300 42378 30328 43864
rect 34440 42378 34468 43982
rect 38014 43982 38332 44010
rect 38014 43864 38070 43982
rect 30300 42362 30420 42378
rect 29092 42356 29144 42362
rect 30300 42356 30432 42362
rect 30300 42350 30380 42356
rect 29092 42298 29144 42304
rect 30380 42298 30432 42304
rect 32956 42356 33008 42362
rect 34440 42350 34560 42378
rect 38304 42362 38332 43982
rect 41878 43864 41934 44664
rect 41892 42362 41920 43864
rect 32956 42298 33008 42304
rect 29104 41818 29132 42298
rect 30472 42220 30524 42226
rect 30472 42162 30524 42168
rect 30484 41857 30512 42162
rect 31668 42152 31720 42158
rect 31668 42094 31720 42100
rect 32680 42152 32732 42158
rect 32680 42094 32732 42100
rect 30470 41848 30526 41857
rect 29000 41812 29052 41818
rect 29000 41754 29052 41760
rect 29092 41812 29144 41818
rect 30470 41783 30526 41792
rect 29092 41754 29144 41760
rect 28540 41676 28592 41682
rect 28540 41618 28592 41624
rect 26608 41540 26660 41546
rect 26608 41482 26660 41488
rect 27436 41540 27488 41546
rect 27436 41482 27488 41488
rect 26620 41274 26648 41482
rect 27252 41472 27304 41478
rect 27252 41414 27304 41420
rect 27264 41274 27292 41414
rect 26608 41268 26660 41274
rect 26608 41210 26660 41216
rect 26792 41268 26844 41274
rect 26792 41210 26844 41216
rect 27252 41268 27304 41274
rect 27252 41210 27304 41216
rect 26608 41132 26660 41138
rect 26608 41074 26660 41080
rect 26516 41064 26568 41070
rect 26516 41006 26568 41012
rect 26528 40526 26556 41006
rect 26516 40520 26568 40526
rect 26516 40462 26568 40468
rect 26528 39846 26556 40462
rect 26516 39840 26568 39846
rect 26516 39782 26568 39788
rect 26516 39636 26568 39642
rect 26516 39578 26568 39584
rect 26528 38962 26556 39578
rect 26620 39574 26648 41074
rect 26804 41070 26832 41210
rect 26882 41168 26938 41177
rect 27160 41132 27212 41138
rect 26938 41112 27016 41120
rect 26882 41103 26884 41112
rect 26936 41092 27016 41112
rect 26884 41074 26936 41080
rect 26792 41064 26844 41070
rect 26792 41006 26844 41012
rect 26792 40928 26844 40934
rect 26792 40870 26844 40876
rect 26884 40928 26936 40934
rect 26884 40870 26936 40876
rect 26700 40452 26752 40458
rect 26700 40394 26752 40400
rect 26608 39568 26660 39574
rect 26608 39510 26660 39516
rect 26516 38956 26568 38962
rect 26568 38916 26648 38944
rect 26516 38898 26568 38904
rect 26516 38820 26568 38826
rect 26516 38762 26568 38768
rect 26422 38584 26478 38593
rect 26422 38519 26478 38528
rect 26528 38010 26556 38762
rect 26516 38004 26568 38010
rect 26516 37946 26568 37952
rect 26424 37800 26476 37806
rect 26620 37788 26648 38916
rect 26712 38894 26740 40394
rect 26804 39846 26832 40870
rect 26896 40050 26924 40870
rect 26988 40730 27016 41092
rect 27160 41074 27212 41080
rect 27252 41132 27304 41138
rect 27252 41074 27304 41080
rect 27172 40934 27200 41074
rect 27160 40928 27212 40934
rect 27160 40870 27212 40876
rect 26976 40724 27028 40730
rect 26976 40666 27028 40672
rect 26974 40624 27030 40633
rect 26974 40559 27030 40568
rect 26988 40526 27016 40559
rect 26976 40520 27028 40526
rect 26976 40462 27028 40468
rect 27160 40452 27212 40458
rect 27160 40394 27212 40400
rect 26976 40384 27028 40390
rect 26976 40326 27028 40332
rect 26884 40044 26936 40050
rect 26884 39986 26936 39992
rect 26792 39840 26844 39846
rect 26792 39782 26844 39788
rect 26700 38888 26752 38894
rect 26700 38830 26752 38836
rect 26988 38654 27016 40326
rect 27068 39976 27120 39982
rect 27068 39918 27120 39924
rect 27080 39098 27108 39918
rect 27068 39092 27120 39098
rect 27068 39034 27120 39040
rect 26988 38626 27108 38654
rect 26882 38584 26938 38593
rect 27080 38554 27108 38626
rect 26882 38519 26938 38528
rect 27068 38548 27120 38554
rect 26896 38486 26924 38519
rect 27068 38490 27120 38496
rect 26884 38480 26936 38486
rect 26884 38422 26936 38428
rect 26884 38208 26936 38214
rect 26884 38150 26936 38156
rect 26896 38010 26924 38150
rect 26884 38004 26936 38010
rect 26884 37946 26936 37952
rect 26700 37868 26752 37874
rect 26700 37810 26752 37816
rect 26976 37868 27028 37874
rect 26976 37810 27028 37816
rect 26476 37760 26648 37788
rect 26424 37742 26476 37748
rect 26332 37256 26384 37262
rect 26332 37198 26384 37204
rect 26344 36961 26372 37198
rect 26436 37194 26464 37742
rect 26712 37448 26740 37810
rect 26884 37460 26936 37466
rect 26712 37420 26884 37448
rect 26424 37188 26476 37194
rect 26424 37130 26476 37136
rect 26516 37188 26568 37194
rect 26516 37130 26568 37136
rect 26330 36952 26386 36961
rect 26330 36887 26386 36896
rect 26146 36272 26202 36281
rect 26146 36207 26202 36216
rect 26160 36038 26188 36207
rect 26148 36032 26200 36038
rect 26148 35974 26200 35980
rect 26240 35692 26292 35698
rect 26160 35652 26240 35680
rect 26056 34740 26108 34746
rect 26056 34682 26108 34688
rect 26056 34604 26108 34610
rect 26056 34546 26108 34552
rect 26068 34513 26096 34546
rect 26054 34504 26110 34513
rect 26054 34439 26110 34448
rect 26054 34232 26110 34241
rect 26054 34167 26110 34176
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25964 33516 26016 33522
rect 25964 33458 26016 33464
rect 25688 33448 25740 33454
rect 25688 33390 25740 33396
rect 25320 32846 25372 32852
rect 25516 32830 25636 32858
rect 25412 32496 25464 32502
rect 25412 32438 25464 32444
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25226 32056 25282 32065
rect 25226 31991 25282 32000
rect 25228 31952 25280 31958
rect 25228 31894 25280 31900
rect 25134 31376 25190 31385
rect 25044 31340 25096 31346
rect 25134 31311 25136 31320
rect 25044 31282 25096 31288
rect 25188 31311 25190 31320
rect 25136 31282 25188 31288
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 24964 30734 24992 30874
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24766 30560 24822 30569
rect 24766 30495 24822 30504
rect 24400 30252 24452 30258
rect 24596 30246 24808 30274
rect 24452 30212 24532 30240
rect 24400 30194 24452 30200
rect 24398 30016 24454 30025
rect 24398 29951 24454 29960
rect 24308 29708 24360 29714
rect 24308 29650 24360 29656
rect 24320 29170 24348 29650
rect 24308 29164 24360 29170
rect 24308 29106 24360 29112
rect 24228 28966 24348 28994
rect 24320 28665 24348 28966
rect 24306 28656 24362 28665
rect 24306 28591 24362 28600
rect 24320 28558 24348 28591
rect 24308 28552 24360 28558
rect 24308 28494 24360 28500
rect 24216 27328 24268 27334
rect 24216 27270 24268 27276
rect 23952 27118 24164 27146
rect 23848 26512 23900 26518
rect 23848 26454 23900 26460
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23676 24818 23704 25230
rect 23664 24812 23716 24818
rect 23664 24754 23716 24760
rect 23754 24712 23810 24721
rect 23480 24676 23532 24682
rect 23480 24618 23532 24624
rect 23676 24670 23754 24698
rect 23492 24206 23520 24618
rect 23676 24342 23704 24670
rect 23754 24647 23810 24656
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23846 24576 23902 24585
rect 23664 24336 23716 24342
rect 23664 24278 23716 24284
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23676 23526 23704 24278
rect 23664 23520 23716 23526
rect 23492 23468 23664 23474
rect 23492 23462 23716 23468
rect 23492 23446 23704 23462
rect 23386 22808 23442 22817
rect 23386 22743 23442 22752
rect 23296 22500 23348 22506
rect 23296 22442 23348 22448
rect 23110 22264 23166 22273
rect 23110 22199 23112 22208
rect 23164 22199 23166 22208
rect 23112 22170 23164 22176
rect 23308 22094 23336 22442
rect 23400 22098 23428 22743
rect 23492 22273 23520 23446
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23478 22264 23534 22273
rect 23478 22199 23534 22208
rect 23124 22066 23336 22094
rect 23388 22092 23440 22098
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 23032 21690 23060 21966
rect 23020 21684 23072 21690
rect 23020 21626 23072 21632
rect 22928 18896 22980 18902
rect 22928 18838 22980 18844
rect 23124 18358 23152 22066
rect 23388 22034 23440 22040
rect 23492 21978 23520 22199
rect 23308 21950 23520 21978
rect 23308 19961 23336 21950
rect 23584 21842 23612 22918
rect 23676 22710 23704 22986
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 23676 22030 23704 22646
rect 23768 22098 23796 24550
rect 23846 24511 23902 24520
rect 23860 23186 23888 24511
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23846 22672 23902 22681
rect 23846 22607 23902 22616
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23492 21814 23612 21842
rect 23492 21622 23520 21814
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23676 21536 23704 21966
rect 23768 21672 23796 22034
rect 23860 22030 23888 22607
rect 23952 22522 23980 27118
rect 24124 26852 24176 26858
rect 24124 26794 24176 26800
rect 24030 25528 24086 25537
rect 24030 25463 24086 25472
rect 24044 24818 24072 25463
rect 24136 25294 24164 26794
rect 24228 26217 24256 27270
rect 24320 26246 24348 28494
rect 24412 26994 24440 29951
rect 24504 29481 24532 30212
rect 24676 30184 24728 30190
rect 24676 30126 24728 30132
rect 24584 29776 24636 29782
rect 24584 29718 24636 29724
rect 24490 29472 24546 29481
rect 24490 29407 24546 29416
rect 24504 29170 24532 29407
rect 24492 29164 24544 29170
rect 24492 29106 24544 29112
rect 24596 29102 24624 29718
rect 24584 29096 24636 29102
rect 24584 29038 24636 29044
rect 24596 28694 24624 29038
rect 24584 28688 24636 28694
rect 24584 28630 24636 28636
rect 24688 28558 24716 30126
rect 24780 29510 24808 30246
rect 24964 29714 24992 30670
rect 25056 30569 25084 31282
rect 25136 31136 25188 31142
rect 25136 31078 25188 31084
rect 25042 30560 25098 30569
rect 25042 30495 25098 30504
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 25056 30258 25084 30330
rect 25044 30252 25096 30258
rect 25044 30194 25096 30200
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 24768 29504 24820 29510
rect 25044 29504 25096 29510
rect 24820 29464 24992 29492
rect 24768 29446 24820 29452
rect 24964 29220 24992 29464
rect 25042 29472 25044 29481
rect 25096 29472 25098 29481
rect 25042 29407 25098 29416
rect 24780 29192 24992 29220
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24490 27976 24546 27985
rect 24490 27911 24546 27920
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 24504 26897 24532 27911
rect 24676 27464 24728 27470
rect 24676 27406 24728 27412
rect 24490 26888 24546 26897
rect 24688 26858 24716 27406
rect 24490 26823 24546 26832
rect 24584 26852 24636 26858
rect 24584 26794 24636 26800
rect 24676 26852 24728 26858
rect 24676 26794 24728 26800
rect 24308 26240 24360 26246
rect 24214 26208 24270 26217
rect 24308 26182 24360 26188
rect 24492 26240 24544 26246
rect 24492 26182 24544 26188
rect 24214 26143 24270 26152
rect 24124 25288 24176 25294
rect 24124 25230 24176 25236
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24044 24206 24072 24754
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 24044 23254 24072 24142
rect 24032 23248 24084 23254
rect 24032 23190 24084 23196
rect 24044 22710 24072 23190
rect 24032 22704 24084 22710
rect 24032 22646 24084 22652
rect 23952 22494 24072 22522
rect 24044 22438 24072 22494
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 24136 22098 24164 25230
rect 24228 23730 24256 26143
rect 24398 25256 24454 25265
rect 24398 25191 24454 25200
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 24320 24410 24348 24550
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 24412 24290 24440 25191
rect 24504 24614 24532 26182
rect 24596 25906 24624 26794
rect 24688 26518 24716 26794
rect 24676 26512 24728 26518
rect 24676 26454 24728 26460
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24584 25696 24636 25702
rect 24584 25638 24636 25644
rect 24492 24608 24544 24614
rect 24492 24550 24544 24556
rect 24320 24262 24440 24290
rect 24320 24206 24348 24262
rect 24308 24200 24360 24206
rect 24504 24154 24532 24550
rect 24308 24142 24360 24148
rect 24412 24126 24532 24154
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 24308 22636 24360 22642
rect 24308 22578 24360 22584
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 24320 22030 24348 22578
rect 24412 22098 24440 24126
rect 24492 23656 24544 23662
rect 24596 23633 24624 25638
rect 24674 24848 24730 24857
rect 24674 24783 24730 24792
rect 24688 24342 24716 24783
rect 24780 24750 24808 29192
rect 24952 28960 25004 28966
rect 24952 28902 25004 28908
rect 24964 28801 24992 28902
rect 24950 28792 25006 28801
rect 24950 28727 25006 28736
rect 25044 28756 25096 28762
rect 25044 28698 25096 28704
rect 25056 28082 25084 28698
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24950 27296 25006 27305
rect 24950 27231 25006 27240
rect 24964 26994 24992 27231
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24872 26761 24900 26862
rect 24964 26790 24992 26930
rect 24952 26784 25004 26790
rect 24858 26752 24914 26761
rect 24952 26726 25004 26732
rect 24858 26687 24914 26696
rect 24964 26382 24992 26726
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 25056 25974 25084 28018
rect 25148 27130 25176 31078
rect 25240 29617 25268 31894
rect 25332 31822 25360 32166
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 25320 31136 25372 31142
rect 25320 31078 25372 31084
rect 25332 30705 25360 31078
rect 25318 30696 25374 30705
rect 25318 30631 25374 30640
rect 25320 30388 25372 30394
rect 25320 30330 25372 30336
rect 25332 30104 25360 30330
rect 25424 30172 25452 32438
rect 25516 30394 25544 32830
rect 25596 32768 25648 32774
rect 25596 32710 25648 32716
rect 25608 31686 25636 32710
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25608 31346 25636 31622
rect 25700 31414 25728 33390
rect 25780 33312 25832 33318
rect 25778 33280 25780 33289
rect 25832 33280 25834 33289
rect 25778 33215 25834 33224
rect 25976 32774 26004 33458
rect 26068 32910 26096 34167
rect 26160 33561 26188 35652
rect 26240 35634 26292 35640
rect 26332 35692 26384 35698
rect 26332 35634 26384 35640
rect 26240 35556 26292 35562
rect 26240 35498 26292 35504
rect 26252 35086 26280 35498
rect 26344 35329 26372 35634
rect 26436 35562 26464 37130
rect 26424 35556 26476 35562
rect 26424 35498 26476 35504
rect 26330 35320 26386 35329
rect 26330 35255 26386 35264
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 26240 34468 26292 34474
rect 26240 34410 26292 34416
rect 26252 33930 26280 34410
rect 26332 34400 26384 34406
rect 26332 34342 26384 34348
rect 26424 34400 26476 34406
rect 26424 34342 26476 34348
rect 26344 33998 26372 34342
rect 26332 33992 26384 33998
rect 26332 33934 26384 33940
rect 26240 33924 26292 33930
rect 26240 33866 26292 33872
rect 26238 33824 26294 33833
rect 26238 33759 26294 33768
rect 26252 33590 26280 33759
rect 26240 33584 26292 33590
rect 26146 33552 26202 33561
rect 26240 33526 26292 33532
rect 26146 33487 26202 33496
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 25964 32768 26016 32774
rect 25964 32710 26016 32716
rect 25976 32502 26004 32710
rect 25964 32496 26016 32502
rect 25964 32438 26016 32444
rect 26068 32230 26096 32846
rect 26056 32224 26108 32230
rect 26056 32166 26108 32172
rect 25780 31952 25832 31958
rect 25780 31894 25832 31900
rect 25792 31793 25820 31894
rect 26068 31822 26096 32166
rect 26252 31958 26280 32846
rect 26344 31958 26372 33934
rect 26436 33522 26464 34342
rect 26424 33516 26476 33522
rect 26424 33458 26476 33464
rect 26424 32428 26476 32434
rect 26424 32370 26476 32376
rect 26240 31952 26292 31958
rect 26240 31894 26292 31900
rect 26332 31952 26384 31958
rect 26332 31894 26384 31900
rect 25964 31816 26016 31822
rect 25778 31784 25834 31793
rect 25964 31758 26016 31764
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 25778 31719 25834 31728
rect 25976 31414 26004 31758
rect 26148 31680 26200 31686
rect 26148 31622 26200 31628
rect 25688 31408 25740 31414
rect 25688 31350 25740 31356
rect 25964 31408 26016 31414
rect 25964 31350 26016 31356
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 25596 31136 25648 31142
rect 25596 31078 25648 31084
rect 25608 30938 25636 31078
rect 25596 30932 25648 30938
rect 25596 30874 25648 30880
rect 25596 30660 25648 30666
rect 25596 30602 25648 30608
rect 25504 30388 25556 30394
rect 25504 30330 25556 30336
rect 25516 30297 25544 30330
rect 25502 30288 25558 30297
rect 25502 30223 25558 30232
rect 25504 30184 25556 30190
rect 25424 30144 25504 30172
rect 25504 30126 25556 30132
rect 25332 30076 25452 30104
rect 25226 29608 25282 29617
rect 25226 29543 25282 29552
rect 25226 29472 25282 29481
rect 25226 29407 25282 29416
rect 25240 29170 25268 29407
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25226 29064 25282 29073
rect 25282 29034 25360 29050
rect 25282 29028 25372 29034
rect 25282 29022 25320 29028
rect 25226 28999 25282 29008
rect 25320 28970 25372 28976
rect 25228 28960 25280 28966
rect 25228 28902 25280 28908
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25148 26994 25176 27066
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25044 25968 25096 25974
rect 25044 25910 25096 25916
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24860 24608 24912 24614
rect 24860 24550 24912 24556
rect 24872 24342 24900 24550
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 24860 24336 24912 24342
rect 24912 24296 24992 24324
rect 24860 24278 24912 24284
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24492 23598 24544 23604
rect 24582 23624 24638 23633
rect 24504 22642 24532 23598
rect 24688 23594 24716 23802
rect 24860 23724 24912 23730
rect 24860 23666 24912 23672
rect 24582 23559 24638 23568
rect 24676 23588 24728 23594
rect 24676 23530 24728 23536
rect 24768 23520 24820 23526
rect 24768 23462 24820 23468
rect 24584 23044 24636 23050
rect 24584 22986 24636 22992
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24596 22522 24624 22986
rect 24504 22494 24624 22522
rect 24400 22092 24452 22098
rect 24400 22034 24452 22040
rect 23848 22024 23900 22030
rect 24216 22024 24268 22030
rect 23900 21984 23980 22012
rect 23848 21966 23900 21972
rect 23768 21644 23888 21672
rect 23756 21548 23808 21554
rect 23676 21508 23756 21536
rect 23756 21490 23808 21496
rect 23860 21418 23888 21644
rect 23848 21412 23900 21418
rect 23848 21354 23900 21360
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23492 21146 23520 21286
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23388 21072 23440 21078
rect 23440 21020 23520 21026
rect 23388 21014 23520 21020
rect 23400 20998 23520 21014
rect 23952 21010 23980 21984
rect 24216 21966 24268 21972
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24122 21720 24178 21729
rect 24122 21655 24178 21664
rect 23294 19952 23350 19961
rect 23294 19887 23350 19896
rect 23492 19854 23520 20998
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 24030 20496 24086 20505
rect 24030 20431 24086 20440
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23768 19990 23796 20198
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 23756 19984 23808 19990
rect 23756 19926 23808 19932
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23492 18986 23520 19246
rect 23308 18970 23520 18986
rect 23296 18964 23520 18970
rect 23348 18958 23520 18964
rect 23296 18906 23348 18912
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 23112 18352 23164 18358
rect 23110 18320 23112 18329
rect 23164 18320 23166 18329
rect 23020 18284 23072 18290
rect 23308 18290 23336 18566
rect 23400 18426 23428 18770
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23110 18255 23166 18264
rect 23296 18284 23348 18290
rect 23020 18226 23072 18232
rect 23296 18226 23348 18232
rect 23032 17882 23060 18226
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23032 16998 23060 17614
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22388 15910 22416 16050
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22296 14414 22324 15302
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22296 14074 22324 14350
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22388 13938 22416 15846
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22296 13326 22324 13398
rect 22284 13320 22336 13326
rect 22112 13246 22232 13274
rect 22284 13262 22336 13268
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22112 11898 22140 13126
rect 22204 12186 22232 13246
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22296 12345 22324 12378
rect 22282 12336 22338 12345
rect 22282 12271 22338 12280
rect 22388 12238 22416 13874
rect 22376 12232 22428 12238
rect 22204 12158 22324 12186
rect 22376 12174 22428 12180
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 22112 11762 22140 11834
rect 22296 11801 22324 12158
rect 22282 11792 22338 11801
rect 22100 11756 22152 11762
rect 22282 11727 22338 11736
rect 22100 11698 22152 11704
rect 22190 11248 22246 11257
rect 22190 11183 22246 11192
rect 22204 11150 22232 11183
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22296 10826 22324 11727
rect 22388 11354 22416 12174
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22388 11121 22416 11290
rect 22374 11112 22430 11121
rect 22374 11047 22430 11056
rect 22388 11014 22416 11047
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22296 10798 22416 10826
rect 22388 10130 22416 10798
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22480 10062 22508 16934
rect 23124 16794 23152 17138
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22836 16448 22888 16454
rect 22756 16396 22836 16402
rect 22756 16390 22888 16396
rect 22756 16374 22876 16390
rect 22756 16114 22784 16374
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22756 15910 22784 16050
rect 22940 16046 22968 16526
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 22928 16040 22980 16046
rect 22980 16000 23060 16028
rect 22928 15982 22980 15988
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22926 15872 22982 15881
rect 22572 13802 22600 15846
rect 22926 15807 22982 15816
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 22652 15632 22704 15638
rect 22652 15574 22704 15580
rect 22664 15502 22692 15574
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22664 14414 22692 15438
rect 22848 15366 22876 15642
rect 22940 15502 22968 15807
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22756 14278 22784 14486
rect 22940 14482 22968 14962
rect 23032 14906 23060 16000
rect 23124 15026 23152 16050
rect 23216 15434 23244 18022
rect 23296 17740 23348 17746
rect 23296 17682 23348 17688
rect 23308 15552 23336 17682
rect 23492 17354 23520 18770
rect 23584 18766 23612 19654
rect 23676 18902 23704 19722
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23664 18896 23716 18902
rect 23664 18838 23716 18844
rect 23676 18766 23704 18838
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23584 18290 23612 18566
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23768 18170 23796 19654
rect 23584 18154 23796 18170
rect 23572 18148 23796 18154
rect 23624 18142 23796 18148
rect 23572 18090 23624 18096
rect 23860 18034 23888 19994
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23400 17326 23520 17354
rect 23584 18006 23888 18034
rect 23400 16833 23428 17326
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23386 16824 23442 16833
rect 23386 16759 23442 16768
rect 23400 16590 23428 16759
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23492 16454 23520 16934
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23386 16280 23442 16289
rect 23386 16215 23442 16224
rect 23400 16114 23428 16215
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23308 15524 23520 15552
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 23400 15162 23428 15370
rect 23492 15162 23520 15524
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23112 15020 23164 15026
rect 23164 14980 23244 15008
rect 23112 14962 23164 14968
rect 23032 14878 23152 14906
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22742 14104 22798 14113
rect 22742 14039 22798 14048
rect 22756 13938 22784 14039
rect 22834 13968 22890 13977
rect 22744 13932 22796 13938
rect 22834 13903 22836 13912
rect 22744 13874 22796 13880
rect 22888 13903 22890 13912
rect 22836 13874 22888 13880
rect 22560 13796 22612 13802
rect 22560 13738 22612 13744
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22664 11370 22692 13126
rect 22756 13002 22784 13194
rect 22940 13190 22968 14418
rect 23032 13938 23060 14418
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 23018 13696 23074 13705
rect 23124 13682 23152 14878
rect 23074 13654 23152 13682
rect 23018 13631 23074 13640
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22756 12974 23060 13002
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22756 12102 22784 12242
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22572 11342 22692 11370
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22008 9988 22060 9994
rect 22008 9930 22060 9936
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22020 9586 22048 9930
rect 22008 9580 22060 9586
rect 21928 9540 22008 9568
rect 21928 9058 21956 9540
rect 22008 9522 22060 9528
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22020 9178 22048 9318
rect 22480 9178 22508 9998
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 21928 9042 22048 9058
rect 21928 9036 22060 9042
rect 21928 9030 22008 9036
rect 22008 8978 22060 8984
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22204 8090 22232 8434
rect 22284 8356 22336 8362
rect 22284 8298 22336 8304
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 21836 7410 21864 8026
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 21744 6820 21956 6848
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21088 4276 21140 4282
rect 21088 4218 21140 4224
rect 21100 3738 21128 4218
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 20824 3318 20944 3346
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20824 2446 20852 3318
rect 21192 3126 21220 5646
rect 21364 5092 21416 5098
rect 21364 5034 21416 5040
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21284 3194 21312 4626
rect 21376 4282 21404 5034
rect 21744 4690 21772 6666
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21836 6186 21864 6598
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 21928 5098 21956 6820
rect 21916 5092 21968 5098
rect 21916 5034 21968 5040
rect 22020 4690 22048 7822
rect 22192 6860 22244 6866
rect 22112 6820 22192 6848
rect 22112 6186 22140 6820
rect 22192 6802 22244 6808
rect 22296 6254 22324 8298
rect 22572 7528 22600 11342
rect 22836 11280 22888 11286
rect 22836 11222 22888 11228
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22664 7834 22692 11018
rect 22848 10674 22876 11222
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22756 7954 22784 9862
rect 23032 9654 23060 12974
rect 23216 12442 23244 14980
rect 23492 14074 23520 15098
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23400 13326 23428 13670
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23492 13258 23520 13874
rect 23584 13530 23612 18006
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 23676 16182 23704 17002
rect 23860 16776 23888 17478
rect 23952 17202 23980 19722
rect 24044 19310 24072 20431
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24044 18426 24072 19246
rect 24032 18420 24084 18426
rect 24032 18362 24084 18368
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24044 17882 24072 18226
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24044 17678 24072 17818
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 24044 17320 24072 17614
rect 24136 17542 24164 21655
rect 24228 20369 24256 21966
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21690 24440 21830
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24214 20360 24270 20369
rect 24214 20295 24270 20304
rect 24504 20233 24532 22494
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 24490 20224 24546 20233
rect 24490 20159 24546 20168
rect 24492 19984 24544 19990
rect 24492 19926 24544 19932
rect 24400 18896 24452 18902
rect 24400 18838 24452 18844
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24044 17292 24164 17320
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 23860 16748 23980 16776
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23664 16176 23716 16182
rect 23664 16118 23716 16124
rect 23664 15904 23716 15910
rect 23662 15872 23664 15881
rect 23716 15872 23718 15881
rect 23662 15807 23718 15816
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23662 15192 23718 15201
rect 23662 15127 23718 15136
rect 23676 15094 23704 15127
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23768 15026 23796 15506
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 13938 23704 14214
rect 23860 14074 23888 16594
rect 23952 15570 23980 16748
rect 24044 16658 24072 17138
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 24044 15416 24072 15982
rect 24136 15502 24164 17292
rect 24228 16522 24256 18702
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24320 18290 24348 18566
rect 24412 18290 24440 18838
rect 24504 18698 24532 19926
rect 24492 18692 24544 18698
rect 24492 18634 24544 18640
rect 24504 18465 24532 18634
rect 24490 18456 24546 18465
rect 24596 18426 24624 22374
rect 24780 21672 24808 23462
rect 24872 22982 24900 23666
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24872 22681 24900 22918
rect 24858 22672 24914 22681
rect 24858 22607 24914 22616
rect 24858 22264 24914 22273
rect 24858 22199 24914 22208
rect 24872 22098 24900 22199
rect 24964 22166 24992 24296
rect 25056 23254 25084 25910
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25148 24954 25176 25230
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25134 24440 25190 24449
rect 25134 24375 25190 24384
rect 25044 23248 25096 23254
rect 25044 23190 25096 23196
rect 25148 23100 25176 24375
rect 25240 23254 25268 28902
rect 25320 28076 25372 28082
rect 25320 28018 25372 28024
rect 25332 25906 25360 28018
rect 25424 27674 25452 30076
rect 25412 27668 25464 27674
rect 25412 27610 25464 27616
rect 25424 27470 25452 27610
rect 25516 27470 25544 30126
rect 25608 29714 25636 30602
rect 25596 29708 25648 29714
rect 25596 29650 25648 29656
rect 25594 29608 25650 29617
rect 25650 29566 25728 29594
rect 25594 29543 25650 29552
rect 25596 29504 25648 29510
rect 25596 29446 25648 29452
rect 25608 29306 25636 29446
rect 25596 29300 25648 29306
rect 25596 29242 25648 29248
rect 25700 29170 25728 29566
rect 25792 29170 25820 31282
rect 26068 30938 26096 31282
rect 26056 30932 26108 30938
rect 26056 30874 26108 30880
rect 25964 30796 26016 30802
rect 25964 30738 26016 30744
rect 25872 30728 25924 30734
rect 25872 30670 25924 30676
rect 25688 29164 25740 29170
rect 25688 29106 25740 29112
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25516 27130 25544 27406
rect 25504 27124 25556 27130
rect 25504 27066 25556 27072
rect 25608 26466 25636 29038
rect 25792 28778 25820 29106
rect 25884 28966 25912 30670
rect 25976 30258 26004 30738
rect 26160 30682 26188 31622
rect 26252 31346 26280 31894
rect 26330 31784 26386 31793
rect 26330 31719 26386 31728
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 26240 31204 26292 31210
rect 26240 31146 26292 31152
rect 26252 30938 26280 31146
rect 26240 30932 26292 30938
rect 26240 30874 26292 30880
rect 26160 30654 26280 30682
rect 26146 30560 26202 30569
rect 26146 30495 26202 30504
rect 26160 30410 26188 30495
rect 26068 30382 26188 30410
rect 25964 30252 26016 30258
rect 25964 30194 26016 30200
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25976 29170 26004 29582
rect 25964 29164 26016 29170
rect 25964 29106 26016 29112
rect 25964 29028 26016 29034
rect 25964 28970 26016 28976
rect 25872 28960 25924 28966
rect 25872 28902 25924 28908
rect 25792 28750 25912 28778
rect 25884 28694 25912 28750
rect 25780 28688 25832 28694
rect 25780 28630 25832 28636
rect 25872 28688 25924 28694
rect 25872 28630 25924 28636
rect 25792 28540 25820 28630
rect 25976 28540 26004 28970
rect 25792 28512 26004 28540
rect 25964 27464 26016 27470
rect 25964 27406 26016 27412
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 25688 27124 25740 27130
rect 25688 27066 25740 27072
rect 25700 26994 25728 27066
rect 25688 26988 25740 26994
rect 25688 26930 25740 26936
rect 25700 26586 25728 26930
rect 25792 26790 25820 27270
rect 25976 26926 26004 27406
rect 25964 26920 26016 26926
rect 25964 26862 26016 26868
rect 25872 26852 25924 26858
rect 25872 26794 25924 26800
rect 25780 26784 25832 26790
rect 25780 26726 25832 26732
rect 25778 26616 25834 26625
rect 25688 26580 25740 26586
rect 25884 26586 25912 26794
rect 25778 26551 25834 26560
rect 25872 26580 25924 26586
rect 25688 26522 25740 26528
rect 25792 26466 25820 26551
rect 25872 26522 25924 26528
rect 25504 26444 25556 26450
rect 25608 26438 25820 26466
rect 25964 26512 26016 26518
rect 25964 26454 26016 26460
rect 25504 26386 25556 26392
rect 25320 25900 25372 25906
rect 25516 25888 25544 26386
rect 25792 26382 25820 26438
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 25872 26376 25924 26382
rect 25872 26318 25924 26324
rect 25884 25906 25912 26318
rect 25872 25900 25924 25906
rect 25372 25860 25452 25888
rect 25516 25860 25636 25888
rect 25320 25842 25372 25848
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25332 23644 25360 25094
rect 25424 24585 25452 25860
rect 25504 25764 25556 25770
rect 25504 25706 25556 25712
rect 25516 25498 25544 25706
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25608 25294 25636 25860
rect 25872 25842 25924 25848
rect 25688 25832 25740 25838
rect 25688 25774 25740 25780
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25410 24576 25466 24585
rect 25410 24511 25466 24520
rect 25502 24032 25558 24041
rect 25502 23967 25558 23976
rect 25516 23712 25544 23967
rect 25596 23724 25648 23730
rect 25516 23684 25596 23712
rect 25596 23666 25648 23672
rect 25332 23616 25544 23644
rect 25516 23576 25544 23616
rect 25596 23588 25648 23594
rect 25516 23548 25596 23576
rect 25596 23530 25648 23536
rect 25228 23248 25280 23254
rect 25228 23190 25280 23196
rect 25228 23112 25280 23118
rect 25148 23072 25228 23100
rect 25228 23054 25280 23060
rect 25228 22228 25280 22234
rect 25228 22170 25280 22176
rect 24952 22160 25004 22166
rect 24952 22102 25004 22108
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24780 21644 24992 21672
rect 24858 21584 24914 21593
rect 24858 21519 24914 21528
rect 24768 21072 24820 21078
rect 24768 21014 24820 21020
rect 24780 19786 24808 21014
rect 24872 20942 24900 21519
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24964 20262 24992 21644
rect 25240 21622 25268 22170
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25228 21616 25280 21622
rect 25228 21558 25280 21564
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 25056 20534 25084 20742
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25044 20528 25096 20534
rect 25044 20470 25096 20476
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24768 19780 24820 19786
rect 24768 19722 24820 19728
rect 24688 19174 24716 19722
rect 24964 19514 24992 20198
rect 25148 19854 25176 20334
rect 25240 19990 25268 20538
rect 25412 20256 25464 20262
rect 25412 20198 25464 20204
rect 25228 19984 25280 19990
rect 25228 19926 25280 19932
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 25148 19417 25176 19790
rect 25134 19408 25190 19417
rect 24952 19372 25004 19378
rect 25134 19343 25190 19352
rect 24952 19314 25004 19320
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24688 18766 24716 19110
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24490 18391 24546 18400
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24308 18284 24360 18290
rect 24308 18226 24360 18232
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24584 18284 24636 18290
rect 24584 18226 24636 18232
rect 24400 17060 24452 17066
rect 24400 17002 24452 17008
rect 24412 16658 24440 17002
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24308 16584 24360 16590
rect 24308 16526 24360 16532
rect 24216 16516 24268 16522
rect 24216 16458 24268 16464
rect 24320 16046 24348 16526
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24124 15496 24176 15502
rect 24124 15438 24176 15444
rect 23952 15388 24072 15416
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23480 13252 23532 13258
rect 23480 13194 23532 13200
rect 23676 12850 23704 13874
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23768 13734 23796 13806
rect 23756 13728 23808 13734
rect 23754 13696 23756 13705
rect 23808 13696 23810 13705
rect 23754 13631 23810 13640
rect 23952 12918 23980 15388
rect 24228 15366 24256 15574
rect 24216 15360 24268 15366
rect 24030 15328 24086 15337
rect 24216 15302 24268 15308
rect 24030 15263 24086 15272
rect 24044 13870 24072 15263
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23940 12912 23992 12918
rect 23992 12872 24072 12900
rect 23940 12854 23992 12860
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23492 12714 23520 12786
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 22928 9648 22980 9654
rect 22928 9590 22980 9596
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22940 7954 22968 9590
rect 23124 9178 23152 12038
rect 23216 11762 23244 12378
rect 23952 12306 23980 12582
rect 23940 12300 23992 12306
rect 23940 12242 23992 12248
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23204 11756 23256 11762
rect 23256 11716 23336 11744
rect 23204 11698 23256 11704
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23216 11150 23244 11494
rect 23308 11354 23336 11716
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23492 11150 23520 11766
rect 23676 11762 23704 12106
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23676 11150 23704 11698
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23768 11218 23796 11494
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23860 11150 23888 11698
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23204 11008 23256 11014
rect 23202 10976 23204 10985
rect 23256 10976 23258 10985
rect 23202 10911 23258 10920
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23204 10668 23256 10674
rect 23204 10610 23256 10616
rect 23216 10062 23244 10610
rect 23492 10198 23520 10678
rect 23860 10266 23888 11086
rect 24044 10674 24072 12872
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 24044 10266 24072 10610
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 23480 10192 23532 10198
rect 23480 10134 23532 10140
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23308 8294 23336 8570
rect 23296 8288 23348 8294
rect 23296 8230 23348 8236
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 22664 7806 22784 7834
rect 22756 7750 22784 7806
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22480 7500 22600 7528
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22388 6458 22416 7346
rect 22480 7274 22508 7500
rect 22664 7478 22692 7686
rect 22652 7472 22704 7478
rect 22652 7414 22704 7420
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22572 7002 22600 7346
rect 22756 7313 22784 7686
rect 22742 7304 22798 7313
rect 22742 7239 22798 7248
rect 22940 7002 22968 7890
rect 23308 7886 23336 8230
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22560 6248 22612 6254
rect 22940 6202 22968 6938
rect 23388 6860 23440 6866
rect 23492 6848 23520 8774
rect 23768 8498 23796 8910
rect 24136 8634 24164 14962
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24228 11898 24256 12854
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24320 11830 24348 15846
rect 24596 15609 24624 18226
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24674 16008 24730 16017
rect 24674 15943 24730 15952
rect 24582 15600 24638 15609
rect 24582 15535 24638 15544
rect 24596 15502 24624 15535
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24412 15162 24440 15438
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24596 14618 24624 15302
rect 24688 15065 24716 15943
rect 24780 15910 24808 16050
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24872 15502 24900 18090
rect 24964 17241 24992 19314
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 25056 18766 25084 19246
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 25042 18184 25098 18193
rect 25042 18119 25098 18128
rect 24950 17232 25006 17241
rect 25056 17202 25084 18119
rect 24950 17167 25006 17176
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25148 16250 25176 16390
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24768 15428 24820 15434
rect 24768 15370 24820 15376
rect 24780 15337 24808 15370
rect 24766 15328 24822 15337
rect 24766 15263 24822 15272
rect 24872 15094 24900 15438
rect 25136 15428 25188 15434
rect 25136 15370 25188 15376
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24860 15088 24912 15094
rect 24674 15056 24730 15065
rect 24860 15030 24912 15036
rect 24674 14991 24730 15000
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24504 14056 24532 14554
rect 24872 14482 24900 15030
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24504 14028 24808 14056
rect 24398 13968 24454 13977
rect 24398 13903 24400 13912
rect 24452 13903 24454 13912
rect 24584 13932 24636 13938
rect 24400 13874 24452 13880
rect 24584 13874 24636 13880
rect 24676 13898 24728 13904
rect 24596 13530 24624 13874
rect 24676 13840 24728 13846
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24584 13320 24636 13326
rect 24582 13288 24584 13297
rect 24636 13288 24638 13297
rect 24582 13223 24638 13232
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24412 12832 24440 13126
rect 24584 12844 24636 12850
rect 24412 12804 24532 12832
rect 24308 11824 24360 11830
rect 24308 11766 24360 11772
rect 24504 11626 24532 12804
rect 24584 12786 24636 12792
rect 24596 12102 24624 12786
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24492 11620 24544 11626
rect 24492 11562 24544 11568
rect 24504 11150 24532 11562
rect 24688 11286 24716 13840
rect 24780 13394 24808 14028
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24964 13326 24992 15302
rect 25148 15201 25176 15370
rect 25134 15192 25190 15201
rect 25134 15127 25190 15136
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 25056 13938 25084 14758
rect 25134 13968 25190 13977
rect 25044 13932 25096 13938
rect 25134 13903 25136 13912
rect 25044 13874 25096 13880
rect 25188 13903 25190 13912
rect 25136 13874 25188 13880
rect 25044 13796 25096 13802
rect 25044 13738 25096 13744
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 25056 13190 25084 13738
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 25148 13394 25176 13670
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 24858 12472 24914 12481
rect 24858 12407 24914 12416
rect 24768 12368 24820 12374
rect 24766 12336 24768 12345
rect 24820 12336 24822 12345
rect 24766 12271 24822 12280
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24780 11694 24808 12038
rect 24872 11830 24900 12407
rect 24860 11824 24912 11830
rect 24858 11792 24860 11801
rect 24912 11792 24914 11801
rect 24858 11727 24914 11736
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24596 10985 24624 11018
rect 24582 10976 24638 10985
rect 24582 10911 24638 10920
rect 24688 10742 24716 11222
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 24492 8356 24544 8362
rect 24492 8298 24544 8304
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24228 7410 24256 7686
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24412 6934 24440 7346
rect 24400 6928 24452 6934
rect 24400 6870 24452 6876
rect 23440 6820 23520 6848
rect 23388 6802 23440 6808
rect 24412 6662 24440 6870
rect 24504 6798 24532 8298
rect 24780 8090 24808 11630
rect 24872 11150 24900 11727
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24964 10266 24992 12922
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25056 11898 25084 12718
rect 25240 12434 25268 18634
rect 25320 14340 25372 14346
rect 25320 14282 25372 14288
rect 25332 13938 25360 14282
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25424 13784 25452 20198
rect 25516 20058 25544 21626
rect 25608 21554 25636 21830
rect 25700 21672 25728 25774
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 25792 23050 25820 25434
rect 25976 25242 26004 26454
rect 26068 25974 26096 30382
rect 26252 30274 26280 30654
rect 26160 30246 26280 30274
rect 26160 28082 26188 30246
rect 26240 29776 26292 29782
rect 26240 29718 26292 29724
rect 26252 29510 26280 29718
rect 26240 29504 26292 29510
rect 26240 29446 26292 29452
rect 26240 29028 26292 29034
rect 26240 28970 26292 28976
rect 26252 28937 26280 28970
rect 26238 28928 26294 28937
rect 26238 28863 26294 28872
rect 26148 28076 26200 28082
rect 26148 28018 26200 28024
rect 26148 27328 26200 27334
rect 26148 27270 26200 27276
rect 26160 27033 26188 27270
rect 26146 27024 26202 27033
rect 26146 26959 26202 26968
rect 26240 26852 26292 26858
rect 26240 26794 26292 26800
rect 26148 26784 26200 26790
rect 26148 26726 26200 26732
rect 26160 26382 26188 26726
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26056 25968 26108 25974
rect 26056 25910 26108 25916
rect 26148 25832 26200 25838
rect 26148 25774 26200 25780
rect 26054 25392 26110 25401
rect 26054 25327 26110 25336
rect 25884 25214 26004 25242
rect 25884 24070 25912 25214
rect 25964 25152 26016 25158
rect 25964 25094 26016 25100
rect 25872 24064 25924 24070
rect 25872 24006 25924 24012
rect 25780 23044 25832 23050
rect 25780 22986 25832 22992
rect 25884 22234 25912 24006
rect 25872 22228 25924 22234
rect 25872 22170 25924 22176
rect 25700 21644 25820 21672
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25700 21457 25728 21490
rect 25686 21448 25742 21457
rect 25686 21383 25742 21392
rect 25792 21332 25820 21644
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25700 21304 25820 21332
rect 25504 20052 25556 20058
rect 25504 19994 25556 20000
rect 25504 19848 25556 19854
rect 25504 19790 25556 19796
rect 25516 19514 25544 19790
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25516 16794 25544 16934
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25608 16454 25636 16730
rect 25596 16448 25648 16454
rect 25700 16425 25728 21304
rect 25884 21078 25912 21490
rect 25872 21072 25924 21078
rect 25872 21014 25924 21020
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25596 16390 25648 16396
rect 25686 16416 25742 16425
rect 25608 16096 25636 16390
rect 25686 16351 25742 16360
rect 25688 16108 25740 16114
rect 25608 16068 25688 16096
rect 25688 16050 25740 16056
rect 25700 14634 25728 16050
rect 25608 14606 25728 14634
rect 25424 13756 25482 13784
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25332 12918 25360 13670
rect 25454 13546 25482 13756
rect 25424 13518 25482 13546
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 25148 12406 25268 12434
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 24952 10260 25004 10266
rect 24952 10202 25004 10208
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24766 7848 24822 7857
rect 24766 7783 24822 7792
rect 24780 7478 24808 7783
rect 24964 7546 24992 8434
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24768 7472 24820 7478
rect 24768 7414 24820 7420
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24596 6322 24624 7346
rect 24952 7268 25004 7274
rect 24952 7210 25004 7216
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24688 6322 24716 6598
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 22560 6190 22612 6196
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 22020 4010 22048 4626
rect 22112 4282 22140 6122
rect 22572 5914 22600 6190
rect 22848 6174 22968 6202
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22296 5370 22324 5510
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22848 4146 22876 6174
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 22940 5234 22968 6054
rect 23112 5772 23164 5778
rect 23112 5714 23164 5720
rect 23124 5302 23152 5714
rect 23768 5574 23796 6054
rect 24584 5772 24636 5778
rect 24584 5714 24636 5720
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 23860 5370 23888 5510
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23296 5160 23348 5166
rect 23296 5102 23348 5108
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3194 21864 3878
rect 23308 3602 23336 5102
rect 24032 4276 24084 4282
rect 24032 4218 24084 4224
rect 23848 3936 23900 3942
rect 23848 3878 23900 3884
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 22572 3194 22600 3402
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 21180 3120 21232 3126
rect 21180 3062 21232 3068
rect 23308 3058 23336 3538
rect 23860 3126 23888 3878
rect 24044 3738 24072 4218
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 24136 3738 24164 4082
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24596 3602 24624 5714
rect 24688 5302 24716 6258
rect 24872 6254 24900 6734
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 24688 4078 24716 5238
rect 24872 5166 24900 6190
rect 24964 5370 24992 7210
rect 25056 5642 25084 10950
rect 25148 8838 25176 12406
rect 25320 12232 25372 12238
rect 25320 12174 25372 12180
rect 25226 11928 25282 11937
rect 25226 11863 25282 11872
rect 25240 10742 25268 11863
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 25332 10062 25360 12174
rect 25424 11098 25452 13518
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25516 12238 25544 13126
rect 25608 12986 25636 14606
rect 25792 14498 25820 19110
rect 25700 14470 25820 14498
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25700 12918 25728 14470
rect 25778 13968 25834 13977
rect 25778 13903 25834 13912
rect 25792 13802 25820 13903
rect 25780 13796 25832 13802
rect 25780 13738 25832 13744
rect 25792 13462 25820 13738
rect 25780 13456 25832 13462
rect 25780 13398 25832 13404
rect 25688 12912 25740 12918
rect 25688 12854 25740 12860
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25686 11928 25742 11937
rect 25596 11892 25648 11898
rect 25686 11863 25742 11872
rect 25596 11834 25648 11840
rect 25608 11218 25636 11834
rect 25700 11762 25728 11863
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25688 11144 25740 11150
rect 25686 11112 25688 11121
rect 25740 11112 25742 11121
rect 25424 11070 25636 11098
rect 25410 10704 25466 10713
rect 25410 10639 25466 10648
rect 25424 10606 25452 10639
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25240 9586 25268 9998
rect 25424 9722 25452 10542
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25240 8430 25268 9522
rect 25332 8974 25360 9522
rect 25320 8968 25372 8974
rect 25320 8910 25372 8916
rect 25516 8566 25544 10202
rect 25608 9625 25636 11070
rect 25884 11098 25912 20742
rect 25976 19310 26004 25094
rect 26068 24410 26096 25327
rect 26056 24404 26108 24410
rect 26056 24346 26108 24352
rect 26160 23730 26188 25774
rect 26252 23866 26280 26794
rect 26344 25906 26372 31719
rect 26436 29170 26464 32370
rect 26528 32026 26556 37130
rect 26608 36916 26660 36922
rect 26608 36858 26660 36864
rect 26620 33658 26648 36858
rect 26712 36378 26740 37420
rect 26884 37402 26936 37408
rect 26988 37398 27016 37810
rect 26976 37392 27028 37398
rect 26976 37334 27028 37340
rect 26976 37256 27028 37262
rect 26896 37216 26976 37244
rect 26792 36712 26844 36718
rect 26792 36654 26844 36660
rect 26700 36372 26752 36378
rect 26700 36314 26752 36320
rect 26700 36236 26752 36242
rect 26700 36178 26752 36184
rect 26712 35222 26740 36178
rect 26804 36174 26832 36654
rect 26792 36168 26844 36174
rect 26790 36136 26792 36145
rect 26844 36136 26846 36145
rect 26790 36071 26846 36080
rect 26790 35728 26846 35737
rect 26896 35698 26924 37216
rect 26976 37198 27028 37204
rect 26974 36680 27030 36689
rect 26974 36615 27030 36624
rect 26988 36310 27016 36615
rect 26976 36304 27028 36310
rect 26976 36246 27028 36252
rect 26976 36100 27028 36106
rect 26976 36042 27028 36048
rect 26790 35663 26792 35672
rect 26844 35663 26846 35672
rect 26884 35692 26936 35698
rect 26792 35634 26844 35640
rect 26884 35634 26936 35640
rect 26804 35290 26832 35634
rect 26792 35284 26844 35290
rect 26792 35226 26844 35232
rect 26700 35216 26752 35222
rect 26700 35158 26752 35164
rect 26896 35154 26924 35634
rect 26884 35148 26936 35154
rect 26884 35090 26936 35096
rect 26896 34746 26924 35090
rect 26884 34740 26936 34746
rect 26884 34682 26936 34688
rect 26700 33924 26752 33930
rect 26700 33866 26752 33872
rect 26608 33652 26660 33658
rect 26608 33594 26660 33600
rect 26620 33318 26648 33594
rect 26608 33312 26660 33318
rect 26608 33254 26660 33260
rect 26606 32736 26662 32745
rect 26606 32671 26662 32680
rect 26620 32201 26648 32671
rect 26606 32192 26662 32201
rect 26606 32127 26662 32136
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 26608 31748 26660 31754
rect 26608 31690 26660 31696
rect 26516 31680 26568 31686
rect 26514 31648 26516 31657
rect 26568 31648 26570 31657
rect 26514 31583 26570 31592
rect 26528 31346 26556 31583
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26620 30938 26648 31690
rect 26712 31142 26740 33866
rect 26882 33688 26938 33697
rect 26792 33652 26844 33658
rect 26882 33623 26938 33632
rect 26792 33594 26844 33600
rect 26700 31136 26752 31142
rect 26700 31078 26752 31084
rect 26608 30932 26660 30938
rect 26608 30874 26660 30880
rect 26712 30734 26740 31078
rect 26516 30728 26568 30734
rect 26516 30670 26568 30676
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26700 30728 26752 30734
rect 26700 30670 26752 30676
rect 26528 30122 26556 30670
rect 26620 30598 26648 30670
rect 26608 30592 26660 30598
rect 26608 30534 26660 30540
rect 26620 30258 26648 30534
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 26516 30116 26568 30122
rect 26516 30058 26568 30064
rect 26608 30048 26660 30054
rect 26608 29990 26660 29996
rect 26514 29336 26570 29345
rect 26514 29271 26516 29280
rect 26568 29271 26570 29280
rect 26516 29242 26568 29248
rect 26620 29170 26648 29990
rect 26700 29300 26752 29306
rect 26700 29242 26752 29248
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 26516 29164 26568 29170
rect 26516 29106 26568 29112
rect 26608 29164 26660 29170
rect 26608 29106 26660 29112
rect 26436 27470 26464 29106
rect 26528 28082 26556 29106
rect 26620 28558 26648 29106
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26608 28144 26660 28150
rect 26608 28086 26660 28092
rect 26516 28076 26568 28082
rect 26516 28018 26568 28024
rect 26620 27946 26648 28086
rect 26516 27940 26568 27946
rect 26516 27882 26568 27888
rect 26608 27940 26660 27946
rect 26608 27882 26660 27888
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26436 27033 26464 27406
rect 26528 27130 26556 27882
rect 26608 27464 26660 27470
rect 26608 27406 26660 27412
rect 26516 27124 26568 27130
rect 26516 27066 26568 27072
rect 26422 27024 26478 27033
rect 26422 26959 26478 26968
rect 26528 26518 26556 27066
rect 26516 26512 26568 26518
rect 26516 26454 26568 26460
rect 26516 26376 26568 26382
rect 26516 26318 26568 26324
rect 26424 26240 26476 26246
rect 26528 26217 26556 26318
rect 26620 26246 26648 27406
rect 26608 26240 26660 26246
rect 26424 26182 26476 26188
rect 26514 26208 26570 26217
rect 26436 25906 26464 26182
rect 26608 26182 26660 26188
rect 26514 26143 26570 26152
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 26424 25900 26476 25906
rect 26424 25842 26476 25848
rect 26528 25498 26556 26143
rect 26516 25492 26568 25498
rect 26516 25434 26568 25440
rect 26332 25356 26384 25362
rect 26332 25298 26384 25304
rect 26344 23905 26372 25298
rect 26424 24064 26476 24070
rect 26476 24024 26556 24052
rect 26424 24006 26476 24012
rect 26330 23896 26386 23905
rect 26240 23860 26292 23866
rect 26386 23840 26464 23848
rect 26330 23831 26464 23840
rect 26344 23820 26464 23831
rect 26240 23802 26292 23808
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 26332 23724 26384 23730
rect 26332 23666 26384 23672
rect 26344 23633 26372 23666
rect 26330 23624 26386 23633
rect 26330 23559 26386 23568
rect 26436 23526 26464 23820
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26424 23520 26476 23526
rect 26424 23462 26476 23468
rect 26344 23118 26372 23462
rect 26332 23112 26384 23118
rect 26332 23054 26384 23060
rect 26424 23044 26476 23050
rect 26424 22986 26476 22992
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26160 21554 26188 22170
rect 26332 21888 26384 21894
rect 26332 21830 26384 21836
rect 26344 21554 26372 21830
rect 26148 21548 26200 21554
rect 26148 21490 26200 21496
rect 26332 21548 26384 21554
rect 26332 21490 26384 21496
rect 26160 20602 26188 21490
rect 26344 20913 26372 21490
rect 26330 20904 26386 20913
rect 26330 20839 26386 20848
rect 26436 20806 26464 22986
rect 26424 20800 26476 20806
rect 26330 20768 26386 20777
rect 26424 20742 26476 20748
rect 26330 20703 26386 20712
rect 26344 20618 26372 20703
rect 26148 20596 26200 20602
rect 26344 20590 26464 20618
rect 26148 20538 26200 20544
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 26068 17610 26096 17818
rect 26056 17604 26108 17610
rect 26056 17546 26108 17552
rect 26068 16454 26096 17546
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26344 17377 26372 17478
rect 26330 17368 26386 17377
rect 26330 17303 26386 17312
rect 26240 16720 26292 16726
rect 26240 16662 26292 16668
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 26252 16250 26280 16662
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26344 16250 26372 16526
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 25964 15020 26016 15026
rect 25964 14962 26016 14968
rect 25976 14929 26004 14962
rect 26252 14958 26280 15098
rect 26056 14952 26108 14958
rect 25962 14920 26018 14929
rect 26056 14894 26108 14900
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 25962 14855 26018 14864
rect 25976 14074 26004 14855
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 25964 13456 26016 13462
rect 26068 13444 26096 14894
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26016 13416 26096 13444
rect 25964 13398 26016 13404
rect 25976 13326 26004 13398
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 26160 12238 26188 14418
rect 26252 13954 26280 14894
rect 26332 14408 26384 14414
rect 26436 14396 26464 20590
rect 26528 19378 26556 24024
rect 26620 22642 26648 26182
rect 26712 25906 26740 29242
rect 26700 25900 26752 25906
rect 26700 25842 26752 25848
rect 26804 24614 26832 33594
rect 26896 33590 26924 33623
rect 26884 33584 26936 33590
rect 26884 33526 26936 33532
rect 26882 32872 26938 32881
rect 26882 32807 26938 32816
rect 26896 30666 26924 32807
rect 26988 31686 27016 36042
rect 27080 35698 27108 38490
rect 27068 35692 27120 35698
rect 27068 35634 27120 35640
rect 27068 34536 27120 34542
rect 27068 34478 27120 34484
rect 27080 33862 27108 34478
rect 27068 33856 27120 33862
rect 27068 33798 27120 33804
rect 27080 33522 27108 33798
rect 27172 33658 27200 40394
rect 27264 40225 27292 41074
rect 27448 40712 27476 41482
rect 27712 41472 27764 41478
rect 27712 41414 27764 41420
rect 27448 40684 27660 40712
rect 27526 40624 27582 40633
rect 27448 40582 27526 40610
rect 27250 40216 27306 40225
rect 27250 40151 27306 40160
rect 27344 40180 27396 40186
rect 27344 40122 27396 40128
rect 27356 40089 27384 40122
rect 27342 40080 27398 40089
rect 27342 40015 27398 40024
rect 27252 38344 27304 38350
rect 27252 38286 27304 38292
rect 27264 36038 27292 38286
rect 27344 37120 27396 37126
rect 27344 37062 27396 37068
rect 27356 36922 27384 37062
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27448 36530 27476 40582
rect 27526 40559 27582 40568
rect 27632 40508 27660 40684
rect 27724 40662 27752 41414
rect 28080 41132 28132 41138
rect 28080 41074 28132 41080
rect 28172 41132 28224 41138
rect 28172 41074 28224 41080
rect 28356 41132 28408 41138
rect 28356 41074 28408 41080
rect 28448 41132 28500 41138
rect 28448 41074 28500 41080
rect 28092 41041 28120 41074
rect 28078 41032 28134 41041
rect 28078 40967 28134 40976
rect 27712 40656 27764 40662
rect 28184 40633 28212 41074
rect 27712 40598 27764 40604
rect 28170 40624 28226 40633
rect 27540 40480 27660 40508
rect 27540 40390 27568 40480
rect 27724 40458 27752 40598
rect 28170 40559 28226 40568
rect 27712 40452 27764 40458
rect 27712 40394 27764 40400
rect 28080 40452 28132 40458
rect 28080 40394 28132 40400
rect 27528 40384 27580 40390
rect 27724 40361 27752 40394
rect 27528 40326 27580 40332
rect 27710 40352 27766 40361
rect 27710 40287 27766 40296
rect 27896 39976 27948 39982
rect 27816 39936 27896 39964
rect 27712 39432 27764 39438
rect 27712 39374 27764 39380
rect 27620 39296 27672 39302
rect 27620 39238 27672 39244
rect 27632 39098 27660 39238
rect 27620 39092 27672 39098
rect 27620 39034 27672 39040
rect 27618 38992 27674 39001
rect 27724 38978 27752 39374
rect 27674 38962 27752 38978
rect 27674 38956 27764 38962
rect 27674 38950 27712 38956
rect 27618 38927 27674 38936
rect 27712 38898 27764 38904
rect 27620 38888 27672 38894
rect 27620 38830 27672 38836
rect 27632 38654 27660 38830
rect 27540 38626 27660 38654
rect 27540 38010 27568 38626
rect 27618 38584 27674 38593
rect 27816 38554 27844 39936
rect 27896 39918 27948 39924
rect 27896 39840 27948 39846
rect 27896 39782 27948 39788
rect 27908 38962 27936 39782
rect 28092 39438 28120 40394
rect 28368 40089 28396 41074
rect 28460 40916 28488 41074
rect 28552 41070 28580 41618
rect 28724 41132 28776 41138
rect 28644 41092 28724 41120
rect 28540 41064 28592 41070
rect 28540 41006 28592 41012
rect 28540 40928 28592 40934
rect 28460 40888 28540 40916
rect 28540 40870 28592 40876
rect 28552 40526 28580 40870
rect 28540 40520 28592 40526
rect 28540 40462 28592 40468
rect 28448 40112 28500 40118
rect 28354 40080 28410 40089
rect 28448 40054 28500 40060
rect 28354 40015 28410 40024
rect 28356 39636 28408 39642
rect 28356 39578 28408 39584
rect 28080 39432 28132 39438
rect 28080 39374 28132 39380
rect 28264 39432 28316 39438
rect 28264 39374 28316 39380
rect 27896 38956 27948 38962
rect 27896 38898 27948 38904
rect 27988 38956 28040 38962
rect 27988 38898 28040 38904
rect 27618 38519 27674 38528
rect 27804 38548 27856 38554
rect 27632 38486 27660 38519
rect 27804 38490 27856 38496
rect 27620 38480 27672 38486
rect 27620 38422 27672 38428
rect 27620 38344 27672 38350
rect 27620 38286 27672 38292
rect 27632 38010 27660 38286
rect 27712 38276 27764 38282
rect 27712 38218 27764 38224
rect 27528 38004 27580 38010
rect 27528 37946 27580 37952
rect 27620 38004 27672 38010
rect 27620 37946 27672 37952
rect 27724 37874 27752 38218
rect 27816 37874 27844 38490
rect 27908 38434 27936 38898
rect 28000 38729 28028 38898
rect 27986 38720 28042 38729
rect 27986 38655 28042 38664
rect 28092 38486 28120 39374
rect 28080 38480 28132 38486
rect 27908 38406 28028 38434
rect 28080 38422 28132 38428
rect 27896 38344 27948 38350
rect 27896 38286 27948 38292
rect 27712 37868 27764 37874
rect 27712 37810 27764 37816
rect 27804 37868 27856 37874
rect 27804 37810 27856 37816
rect 27528 37800 27580 37806
rect 27580 37748 27844 37754
rect 27528 37742 27844 37748
rect 27540 37738 27844 37742
rect 27540 37732 27856 37738
rect 27540 37726 27804 37732
rect 27804 37674 27856 37680
rect 27618 37496 27674 37505
rect 27618 37431 27674 37440
rect 27632 37330 27660 37431
rect 27620 37324 27672 37330
rect 27620 37266 27672 37272
rect 27528 37256 27580 37262
rect 27528 37198 27580 37204
rect 27356 36502 27476 36530
rect 27252 36032 27304 36038
rect 27252 35974 27304 35980
rect 27356 35834 27384 36502
rect 27344 35828 27396 35834
rect 27344 35770 27396 35776
rect 27356 35601 27384 35770
rect 27540 35698 27568 37198
rect 27620 36372 27672 36378
rect 27620 36314 27672 36320
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27528 35692 27580 35698
rect 27528 35634 27580 35640
rect 27342 35592 27398 35601
rect 27342 35527 27398 35536
rect 27448 34649 27476 35634
rect 27540 35086 27568 35634
rect 27632 35494 27660 36314
rect 27908 36310 27936 38286
rect 28000 37194 28028 38406
rect 28276 38162 28304 39374
rect 28368 39370 28396 39578
rect 28356 39364 28408 39370
rect 28356 39306 28408 39312
rect 28092 38134 28304 38162
rect 27988 37188 28040 37194
rect 27988 37130 28040 37136
rect 27988 36712 28040 36718
rect 27988 36654 28040 36660
rect 27896 36304 27948 36310
rect 27896 36246 27948 36252
rect 27712 36168 27764 36174
rect 27712 36110 27764 36116
rect 27896 36168 27948 36174
rect 28000 36156 28028 36654
rect 27948 36128 28028 36156
rect 27896 36110 27948 36116
rect 27620 35488 27672 35494
rect 27618 35456 27620 35465
rect 27672 35456 27674 35465
rect 27618 35391 27674 35400
rect 27724 35290 27752 36110
rect 27908 35494 27936 36110
rect 28092 35986 28120 38134
rect 28356 37936 28408 37942
rect 28000 35958 28120 35986
rect 28184 37896 28356 37924
rect 27896 35488 27948 35494
rect 27896 35430 27948 35436
rect 27712 35284 27764 35290
rect 27712 35226 27764 35232
rect 27620 35216 27672 35222
rect 27620 35158 27672 35164
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 27632 34921 27660 35158
rect 27804 35148 27856 35154
rect 27856 35108 27936 35136
rect 27804 35090 27856 35096
rect 27618 34912 27674 34921
rect 27618 34847 27674 34856
rect 27632 34678 27660 34847
rect 27620 34672 27672 34678
rect 27434 34640 27490 34649
rect 27620 34614 27672 34620
rect 27434 34575 27490 34584
rect 27712 34604 27764 34610
rect 27712 34546 27764 34552
rect 27250 34096 27306 34105
rect 27306 34054 27384 34082
rect 27250 34031 27306 34040
rect 27160 33652 27212 33658
rect 27160 33594 27212 33600
rect 27068 33516 27120 33522
rect 27068 33458 27120 33464
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 27172 33386 27200 33458
rect 27160 33380 27212 33386
rect 27160 33322 27212 33328
rect 27172 32774 27200 33322
rect 27356 32978 27384 34054
rect 27620 34060 27672 34066
rect 27620 34002 27672 34008
rect 27528 33924 27580 33930
rect 27528 33866 27580 33872
rect 27540 33522 27568 33866
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27434 33416 27490 33425
rect 27434 33351 27490 33360
rect 27448 33318 27476 33351
rect 27436 33312 27488 33318
rect 27436 33254 27488 33260
rect 27540 33114 27568 33458
rect 27528 33108 27580 33114
rect 27528 33050 27580 33056
rect 27526 33008 27582 33017
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27344 32972 27396 32978
rect 27632 32978 27660 34002
rect 27724 33153 27752 34546
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 27710 33144 27766 33153
rect 27710 33079 27766 33088
rect 27712 33040 27764 33046
rect 27712 32982 27764 32988
rect 27526 32943 27582 32952
rect 27620 32972 27672 32978
rect 27344 32914 27396 32920
rect 27160 32768 27212 32774
rect 27160 32710 27212 32716
rect 27068 32496 27120 32502
rect 27068 32438 27120 32444
rect 26976 31680 27028 31686
rect 26976 31622 27028 31628
rect 27080 31328 27108 32438
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 27172 31414 27200 32370
rect 27264 32337 27292 32914
rect 27356 32570 27384 32914
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 27250 32328 27306 32337
rect 27250 32263 27306 32272
rect 27436 32292 27488 32298
rect 27436 32234 27488 32240
rect 27344 32224 27396 32230
rect 27344 32166 27396 32172
rect 27250 32056 27306 32065
rect 27250 31991 27306 32000
rect 27264 31822 27292 31991
rect 27252 31816 27304 31822
rect 27252 31758 27304 31764
rect 27252 31680 27304 31686
rect 27252 31622 27304 31628
rect 27160 31408 27212 31414
rect 27160 31350 27212 31356
rect 26988 31300 27108 31328
rect 26884 30660 26936 30666
rect 26884 30602 26936 30608
rect 26896 28994 26924 30602
rect 26988 30598 27016 31300
rect 27264 31260 27292 31622
rect 27080 31232 27292 31260
rect 26976 30592 27028 30598
rect 26976 30534 27028 30540
rect 26896 28966 27016 28994
rect 26882 27568 26938 27577
rect 26882 27503 26884 27512
rect 26936 27503 26938 27512
rect 26884 27474 26936 27480
rect 26896 24818 26924 27474
rect 26988 27305 27016 28966
rect 26974 27296 27030 27305
rect 26974 27231 27030 27240
rect 26988 26926 27016 27231
rect 26976 26920 27028 26926
rect 26976 26862 27028 26868
rect 27080 26382 27108 31232
rect 27158 31104 27214 31113
rect 27158 31039 27214 31048
rect 27172 30938 27200 31039
rect 27160 30932 27212 30938
rect 27160 30874 27212 30880
rect 27356 30870 27384 32166
rect 27448 31929 27476 32234
rect 27540 32230 27568 32943
rect 27620 32914 27672 32920
rect 27724 32434 27752 32982
rect 27712 32428 27764 32434
rect 27712 32370 27764 32376
rect 27528 32224 27580 32230
rect 27528 32166 27580 32172
rect 27526 32056 27582 32065
rect 27526 31991 27582 32000
rect 27434 31920 27490 31929
rect 27434 31855 27490 31864
rect 27344 30864 27396 30870
rect 27344 30806 27396 30812
rect 27448 30666 27476 31855
rect 27540 31686 27568 31991
rect 27528 31680 27580 31686
rect 27528 31622 27580 31628
rect 27620 31408 27672 31414
rect 27620 31350 27672 31356
rect 27528 31204 27580 31210
rect 27528 31146 27580 31152
rect 27436 30660 27488 30666
rect 27436 30602 27488 30608
rect 27342 30560 27398 30569
rect 27342 30495 27398 30504
rect 27160 30184 27212 30190
rect 27160 30126 27212 30132
rect 27172 28801 27200 30126
rect 27356 29322 27384 30495
rect 27434 30016 27490 30025
rect 27540 30002 27568 31146
rect 27632 30734 27660 31350
rect 27816 30802 27844 33390
rect 27804 30796 27856 30802
rect 27804 30738 27856 30744
rect 27620 30728 27672 30734
rect 27620 30670 27672 30676
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 27620 30592 27672 30598
rect 27620 30534 27672 30540
rect 27490 29974 27568 30002
rect 27434 29951 27490 29960
rect 27528 29844 27580 29850
rect 27264 29306 27384 29322
rect 27448 29804 27528 29832
rect 27264 29300 27396 29306
rect 27264 29294 27344 29300
rect 27158 28792 27214 28801
rect 27158 28727 27214 28736
rect 27158 28656 27214 28665
rect 27158 28591 27214 28600
rect 27172 28558 27200 28591
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27160 28212 27212 28218
rect 27160 28154 27212 28160
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 26988 25974 27016 26318
rect 26976 25968 27028 25974
rect 26976 25910 27028 25916
rect 26976 25832 27028 25838
rect 26974 25800 26976 25809
rect 27028 25800 27030 25809
rect 27172 25786 27200 28154
rect 27264 27169 27292 29294
rect 27344 29242 27396 29248
rect 27344 29164 27396 29170
rect 27448 29152 27476 29804
rect 27528 29786 27580 29792
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27540 29510 27568 29650
rect 27632 29646 27660 30534
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27528 29504 27580 29510
rect 27528 29446 27580 29452
rect 27396 29124 27476 29152
rect 27344 29106 27396 29112
rect 27632 28966 27660 29582
rect 27724 29102 27752 30670
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27816 29646 27844 30194
rect 27804 29640 27856 29646
rect 27804 29582 27856 29588
rect 27712 29096 27764 29102
rect 27712 29038 27764 29044
rect 27620 28960 27672 28966
rect 27620 28902 27672 28908
rect 27632 28558 27660 28902
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27712 28416 27764 28422
rect 27712 28358 27764 28364
rect 27344 28212 27396 28218
rect 27344 28154 27396 28160
rect 27356 27470 27384 28154
rect 27724 28082 27752 28358
rect 27816 28218 27844 29582
rect 27908 29306 27936 35108
rect 28000 35018 28028 35958
rect 28080 35692 28132 35698
rect 28080 35634 28132 35640
rect 27988 35012 28040 35018
rect 27988 34954 28040 34960
rect 27988 33516 28040 33522
rect 27988 33458 28040 33464
rect 28000 32609 28028 33458
rect 27986 32600 28042 32609
rect 27986 32535 28042 32544
rect 28000 32434 28028 32535
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 28092 31890 28120 35634
rect 28184 33658 28212 37896
rect 28356 37878 28408 37884
rect 28264 37800 28316 37806
rect 28264 37742 28316 37748
rect 28276 37262 28304 37742
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 28264 36916 28316 36922
rect 28264 36858 28316 36864
rect 28276 36582 28304 36858
rect 28354 36816 28410 36825
rect 28460 36786 28488 40054
rect 28552 39438 28580 40462
rect 28644 39982 28672 41092
rect 28724 41074 28776 41080
rect 29012 40916 29040 41754
rect 29276 41608 29328 41614
rect 29276 41550 29328 41556
rect 29288 41206 29316 41550
rect 31576 41472 31628 41478
rect 31576 41414 31628 41420
rect 29460 41268 29512 41274
rect 29460 41210 29512 41216
rect 29276 41200 29328 41206
rect 29276 41142 29328 41148
rect 29276 40928 29328 40934
rect 29012 40888 29276 40916
rect 29276 40870 29328 40876
rect 28724 40452 28776 40458
rect 28724 40394 28776 40400
rect 28632 39976 28684 39982
rect 28632 39918 28684 39924
rect 28540 39432 28592 39438
rect 28736 39409 28764 40394
rect 29184 40384 29236 40390
rect 29184 40326 29236 40332
rect 29092 40112 29144 40118
rect 29092 40054 29144 40060
rect 29000 39432 29052 39438
rect 28540 39374 28592 39380
rect 28722 39400 28778 39409
rect 28552 39098 28580 39374
rect 29000 39374 29052 39380
rect 28722 39335 28778 39344
rect 28816 39296 28868 39302
rect 28816 39238 28868 39244
rect 28908 39296 28960 39302
rect 28908 39238 28960 39244
rect 28540 39092 28592 39098
rect 28540 39034 28592 39040
rect 28828 39030 28856 39238
rect 28632 39024 28684 39030
rect 28538 38992 28594 39001
rect 28816 39024 28868 39030
rect 28632 38966 28684 38972
rect 28814 38992 28816 39001
rect 28868 38992 28870 39001
rect 28538 38927 28594 38936
rect 28552 38758 28580 38927
rect 28540 38752 28592 38758
rect 28540 38694 28592 38700
rect 28540 38480 28592 38486
rect 28540 38422 28592 38428
rect 28552 37262 28580 38422
rect 28644 38010 28672 38966
rect 28814 38927 28870 38936
rect 28920 38876 28948 39238
rect 28828 38865 28948 38876
rect 28814 38856 28948 38865
rect 28870 38848 28948 38856
rect 28814 38791 28870 38800
rect 28724 38752 28776 38758
rect 28724 38694 28776 38700
rect 28816 38752 28868 38758
rect 28816 38694 28868 38700
rect 28906 38720 28962 38729
rect 28736 38593 28764 38694
rect 28722 38584 28778 38593
rect 28722 38519 28778 38528
rect 28724 38276 28776 38282
rect 28724 38218 28776 38224
rect 28632 38004 28684 38010
rect 28632 37946 28684 37952
rect 28630 37904 28686 37913
rect 28630 37839 28686 37848
rect 28644 37806 28672 37839
rect 28632 37800 28684 37806
rect 28632 37742 28684 37748
rect 28736 37330 28764 38218
rect 28724 37324 28776 37330
rect 28724 37266 28776 37272
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 28354 36751 28410 36760
rect 28448 36780 28500 36786
rect 28368 36666 28396 36751
rect 28448 36722 28500 36728
rect 28368 36638 28488 36666
rect 28264 36576 28316 36582
rect 28264 36518 28316 36524
rect 28356 36576 28408 36582
rect 28356 36518 28408 36524
rect 28276 34746 28304 36518
rect 28368 36310 28396 36518
rect 28460 36310 28488 36638
rect 28356 36304 28408 36310
rect 28356 36246 28408 36252
rect 28448 36304 28500 36310
rect 28448 36246 28500 36252
rect 28354 36136 28410 36145
rect 28410 36094 28488 36122
rect 28354 36071 28410 36080
rect 28460 35698 28488 36094
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 28354 35320 28410 35329
rect 28354 35255 28410 35264
rect 28368 35154 28396 35255
rect 28356 35148 28408 35154
rect 28356 35090 28408 35096
rect 28356 35012 28408 35018
rect 28356 34954 28408 34960
rect 28264 34740 28316 34746
rect 28264 34682 28316 34688
rect 28264 33924 28316 33930
rect 28264 33866 28316 33872
rect 28172 33652 28224 33658
rect 28172 33594 28224 33600
rect 28184 33114 28212 33594
rect 28276 33522 28304 33866
rect 28264 33516 28316 33522
rect 28264 33458 28316 33464
rect 28172 33108 28224 33114
rect 28172 33050 28224 33056
rect 28172 32972 28224 32978
rect 28172 32914 28224 32920
rect 28080 31884 28132 31890
rect 28080 31826 28132 31832
rect 27988 31816 28040 31822
rect 27988 31758 28040 31764
rect 28000 30394 28028 31758
rect 28080 31272 28132 31278
rect 28080 31214 28132 31220
rect 28092 30977 28120 31214
rect 28078 30968 28134 30977
rect 28078 30903 28134 30912
rect 27988 30388 28040 30394
rect 27988 30330 28040 30336
rect 27986 30016 28042 30025
rect 27986 29951 28042 29960
rect 28000 29510 28028 29951
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 27896 29300 27948 29306
rect 27896 29242 27948 29248
rect 27908 29034 27936 29242
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 27896 29028 27948 29034
rect 27896 28970 27948 28976
rect 27804 28212 27856 28218
rect 27804 28154 27856 28160
rect 27436 28076 27488 28082
rect 27436 28018 27488 28024
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27344 27464 27396 27470
rect 27344 27406 27396 27412
rect 27250 27160 27306 27169
rect 27250 27095 27306 27104
rect 27356 26994 27384 27406
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27264 25922 27292 26930
rect 27356 26586 27384 26930
rect 27448 26926 27476 28018
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27448 26586 27476 26862
rect 27344 26580 27396 26586
rect 27344 26522 27396 26528
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 27540 26353 27568 27406
rect 27526 26344 27582 26353
rect 27526 26279 27582 26288
rect 27344 26036 27396 26042
rect 27396 25996 27568 26024
rect 27344 25978 27396 25984
rect 27264 25894 27476 25922
rect 27540 25906 27568 25996
rect 27632 25974 27660 27950
rect 27802 27704 27858 27713
rect 27908 27674 27936 28970
rect 28000 28150 28028 29106
rect 27988 28144 28040 28150
rect 27988 28086 28040 28092
rect 27802 27639 27858 27648
rect 27896 27668 27948 27674
rect 27712 27600 27764 27606
rect 27712 27542 27764 27548
rect 27724 26994 27752 27542
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27620 25968 27672 25974
rect 27620 25910 27672 25916
rect 27344 25832 27396 25838
rect 27172 25758 27292 25786
rect 27344 25774 27396 25780
rect 26974 25735 27030 25744
rect 27160 25696 27212 25702
rect 27160 25638 27212 25644
rect 26976 25220 27028 25226
rect 26976 25162 27028 25168
rect 26884 24812 26936 24818
rect 26884 24754 26936 24760
rect 26988 24682 27016 25162
rect 27068 24812 27120 24818
rect 27068 24754 27120 24760
rect 26976 24676 27028 24682
rect 26976 24618 27028 24624
rect 26792 24608 26844 24614
rect 26792 24550 26844 24556
rect 26884 24336 26936 24342
rect 26884 24278 26936 24284
rect 26792 24268 26844 24274
rect 26792 24210 26844 24216
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 26620 20262 26648 21422
rect 26608 20256 26660 20262
rect 26608 20198 26660 20204
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26712 19242 26740 23598
rect 26804 23526 26832 24210
rect 26896 23866 26924 24278
rect 26988 24052 27016 24618
rect 27080 24206 27108 24754
rect 27068 24200 27120 24206
rect 27066 24168 27068 24177
rect 27120 24168 27122 24177
rect 27066 24103 27122 24112
rect 27068 24064 27120 24070
rect 26988 24024 27068 24052
rect 27068 24006 27120 24012
rect 26884 23860 26936 23866
rect 26884 23802 26936 23808
rect 26882 23760 26938 23769
rect 26882 23695 26938 23704
rect 26896 23662 26924 23695
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26792 23520 26844 23526
rect 26792 23462 26844 23468
rect 27172 22094 27200 25638
rect 27264 24342 27292 25758
rect 27356 25498 27384 25774
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 27448 24342 27476 25894
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27540 24954 27568 25842
rect 27724 25786 27752 26930
rect 27816 25838 27844 27639
rect 27896 27610 27948 27616
rect 28000 27606 28028 28086
rect 27988 27600 28040 27606
rect 27988 27542 28040 27548
rect 28092 27520 28120 30903
rect 28184 30734 28212 32914
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28276 31346 28304 31758
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28262 31104 28318 31113
rect 28262 31039 28318 31048
rect 28172 30728 28224 30734
rect 28172 30670 28224 30676
rect 28276 30433 28304 31039
rect 28262 30424 28318 30433
rect 28262 30359 28318 30368
rect 28172 30320 28224 30326
rect 28172 30262 28224 30268
rect 28184 29889 28212 30262
rect 28170 29880 28226 29889
rect 28170 29815 28226 29824
rect 28184 29170 28212 29815
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 28092 27492 28212 27520
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27632 25758 27752 25786
rect 27804 25832 27856 25838
rect 27804 25774 27856 25780
rect 27528 24948 27580 24954
rect 27528 24890 27580 24896
rect 27632 24834 27660 25758
rect 27540 24806 27660 24834
rect 27252 24336 27304 24342
rect 27250 24304 27252 24313
rect 27436 24336 27488 24342
rect 27304 24304 27306 24313
rect 27436 24278 27488 24284
rect 27250 24239 27306 24248
rect 27436 24200 27488 24206
rect 27540 24188 27568 24806
rect 27488 24160 27568 24188
rect 27710 24168 27766 24177
rect 27436 24142 27488 24148
rect 27620 24132 27672 24138
rect 27908 24138 27936 27338
rect 28184 27112 28212 27492
rect 28276 27130 28304 30359
rect 28368 28422 28396 34954
rect 28460 34610 28488 35634
rect 28552 34921 28580 37198
rect 28644 35714 28672 37198
rect 28724 37188 28776 37194
rect 28724 37130 28776 37136
rect 28736 36378 28764 37130
rect 28828 36922 28856 38694
rect 28906 38655 28962 38664
rect 28816 36916 28868 36922
rect 28816 36858 28868 36864
rect 28920 36854 28948 38655
rect 29012 38418 29040 39374
rect 29104 38554 29132 40054
rect 29196 40050 29224 40326
rect 29184 40044 29236 40050
rect 29184 39986 29236 39992
rect 29288 39846 29316 40870
rect 29368 40520 29420 40526
rect 29368 40462 29420 40468
rect 29276 39840 29328 39846
rect 29276 39782 29328 39788
rect 29276 39636 29328 39642
rect 29276 39578 29328 39584
rect 29184 39500 29236 39506
rect 29184 39442 29236 39448
rect 29092 38548 29144 38554
rect 29092 38490 29144 38496
rect 29000 38412 29052 38418
rect 29000 38354 29052 38360
rect 29000 38004 29052 38010
rect 29000 37946 29052 37952
rect 29012 37194 29040 37946
rect 29092 37868 29144 37874
rect 29092 37810 29144 37816
rect 29104 37466 29132 37810
rect 29092 37460 29144 37466
rect 29092 37402 29144 37408
rect 29000 37188 29052 37194
rect 29000 37130 29052 37136
rect 28998 37088 29054 37097
rect 28998 37023 29054 37032
rect 29012 36854 29040 37023
rect 28908 36848 28960 36854
rect 28908 36790 28960 36796
rect 29000 36848 29052 36854
rect 29000 36790 29052 36796
rect 28816 36780 28868 36786
rect 28816 36722 28868 36728
rect 28724 36372 28776 36378
rect 28724 36314 28776 36320
rect 28722 36272 28778 36281
rect 28722 36207 28724 36216
rect 28776 36207 28778 36216
rect 28724 36178 28776 36184
rect 28724 36100 28776 36106
rect 28724 36042 28776 36048
rect 28736 35834 28764 36042
rect 28724 35828 28776 35834
rect 28724 35770 28776 35776
rect 28644 35686 28764 35714
rect 28632 35624 28684 35630
rect 28632 35566 28684 35572
rect 28644 35465 28672 35566
rect 28630 35456 28686 35465
rect 28630 35391 28686 35400
rect 28736 35306 28764 35686
rect 28644 35278 28764 35306
rect 28828 35290 28856 36722
rect 28908 36712 28960 36718
rect 28908 36654 28960 36660
rect 29090 36680 29146 36689
rect 28920 36417 28948 36654
rect 29090 36615 29146 36624
rect 28906 36408 28962 36417
rect 28906 36343 28962 36352
rect 28816 35284 28868 35290
rect 28538 34912 28594 34921
rect 28538 34847 28594 34856
rect 28448 34604 28500 34610
rect 28448 34546 28500 34552
rect 28448 34128 28500 34134
rect 28448 34070 28500 34076
rect 28460 29170 28488 34070
rect 28538 33960 28594 33969
rect 28538 33895 28594 33904
rect 28552 33522 28580 33895
rect 28540 33516 28592 33522
rect 28540 33458 28592 33464
rect 28644 33318 28672 35278
rect 28816 35226 28868 35232
rect 29000 35284 29052 35290
rect 29000 35226 29052 35232
rect 28908 35216 28960 35222
rect 28828 35164 28908 35170
rect 28828 35158 28960 35164
rect 28828 35142 28948 35158
rect 28828 35086 28856 35142
rect 28816 35080 28868 35086
rect 28814 35048 28816 35057
rect 29012 35068 29040 35226
rect 28868 35048 28870 35057
rect 28724 35012 28776 35018
rect 28814 34983 28870 34992
rect 28920 35040 29040 35068
rect 29104 35057 29132 36615
rect 29090 35048 29146 35057
rect 28724 34954 28776 34960
rect 28736 34785 28764 34954
rect 28816 34944 28868 34950
rect 28920 34932 28948 35040
rect 29090 34983 29146 34992
rect 29104 34950 29132 34983
rect 28868 34904 28948 34932
rect 29092 34944 29144 34950
rect 28816 34886 28868 34892
rect 29092 34886 29144 34892
rect 28722 34776 28778 34785
rect 28722 34711 28778 34720
rect 29092 34604 29144 34610
rect 29092 34546 29144 34552
rect 28724 33992 28776 33998
rect 28724 33934 28776 33940
rect 28632 33312 28684 33318
rect 28632 33254 28684 33260
rect 28540 33108 28592 33114
rect 28540 33050 28592 33056
rect 28552 32881 28580 33050
rect 28538 32872 28594 32881
rect 28538 32807 28594 32816
rect 28540 32360 28592 32366
rect 28540 32302 28592 32308
rect 28632 32360 28684 32366
rect 28632 32302 28684 32308
rect 28552 31346 28580 32302
rect 28540 31340 28592 31346
rect 28540 31282 28592 31288
rect 28644 30326 28672 32302
rect 28736 32178 28764 33934
rect 28908 33516 28960 33522
rect 28908 33458 28960 33464
rect 28920 33028 28948 33458
rect 28920 33000 28994 33028
rect 28966 32892 28994 33000
rect 28966 32864 29040 32892
rect 29012 32774 29040 32864
rect 29000 32768 29052 32774
rect 29000 32710 29052 32716
rect 29104 32570 29132 34546
rect 28816 32564 28868 32570
rect 28816 32506 28868 32512
rect 29092 32564 29144 32570
rect 29092 32506 29144 32512
rect 28828 32473 28856 32506
rect 28814 32464 28870 32473
rect 28814 32399 28870 32408
rect 28908 32428 28960 32434
rect 28908 32370 28960 32376
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 28736 32150 28856 32178
rect 28724 32020 28776 32026
rect 28724 31962 28776 31968
rect 28736 31414 28764 31962
rect 28828 31890 28856 32150
rect 28816 31884 28868 31890
rect 28816 31826 28868 31832
rect 28920 31822 28948 32370
rect 29104 31958 29132 32370
rect 29196 32230 29224 39442
rect 29288 38554 29316 39578
rect 29276 38548 29328 38554
rect 29276 38490 29328 38496
rect 29276 38412 29328 38418
rect 29276 38354 29328 38360
rect 29288 37942 29316 38354
rect 29276 37936 29328 37942
rect 29276 37878 29328 37884
rect 29380 37262 29408 40462
rect 29368 37256 29420 37262
rect 29368 37198 29420 37204
rect 29368 36372 29420 36378
rect 29368 36314 29420 36320
rect 29380 35086 29408 36314
rect 29276 35080 29328 35086
rect 29276 35022 29328 35028
rect 29368 35080 29420 35086
rect 29368 35022 29420 35028
rect 29288 34785 29316 35022
rect 29274 34776 29330 34785
rect 29274 34711 29330 34720
rect 29380 34610 29408 35022
rect 29472 35000 29500 41210
rect 29736 41132 29788 41138
rect 29736 41074 29788 41080
rect 30564 41132 30616 41138
rect 30564 41074 30616 41080
rect 29748 40458 29776 41074
rect 30012 40996 30064 41002
rect 30012 40938 30064 40944
rect 30024 40730 30052 40938
rect 30380 40928 30432 40934
rect 30380 40870 30432 40876
rect 30472 40928 30524 40934
rect 30472 40870 30524 40876
rect 30286 40760 30342 40769
rect 30012 40724 30064 40730
rect 30286 40695 30288 40704
rect 30012 40666 30064 40672
rect 30340 40695 30342 40704
rect 30288 40666 30340 40672
rect 29736 40452 29788 40458
rect 29736 40394 29788 40400
rect 29828 40452 29880 40458
rect 29828 40394 29880 40400
rect 29644 39840 29696 39846
rect 29644 39782 29696 39788
rect 29552 39636 29604 39642
rect 29552 39578 29604 39584
rect 29564 39098 29592 39578
rect 29656 39506 29684 39782
rect 29748 39624 29776 40394
rect 29840 40089 29868 40394
rect 29826 40080 29882 40089
rect 29826 40015 29882 40024
rect 29748 39596 29868 39624
rect 29644 39500 29696 39506
rect 29644 39442 29696 39448
rect 29736 39500 29788 39506
rect 29736 39442 29788 39448
rect 29644 39296 29696 39302
rect 29644 39238 29696 39244
rect 29552 39092 29604 39098
rect 29552 39034 29604 39040
rect 29656 38962 29684 39238
rect 29748 39137 29776 39442
rect 29734 39128 29790 39137
rect 29734 39063 29790 39072
rect 29644 38956 29696 38962
rect 29644 38898 29696 38904
rect 29840 38706 29868 39596
rect 29920 39296 29972 39302
rect 29920 39238 29972 39244
rect 29564 38678 29868 38706
rect 29564 36689 29592 38678
rect 29644 38548 29696 38554
rect 29644 38490 29696 38496
rect 29550 36680 29606 36689
rect 29550 36615 29606 36624
rect 29656 35698 29684 38490
rect 29828 38276 29880 38282
rect 29828 38218 29880 38224
rect 29840 37466 29868 38218
rect 29828 37460 29880 37466
rect 29828 37402 29880 37408
rect 29736 37188 29788 37194
rect 29736 37130 29788 37136
rect 29748 35698 29776 37130
rect 29840 36922 29868 37402
rect 29828 36916 29880 36922
rect 29828 36858 29880 36864
rect 29932 36106 29960 39238
rect 30024 38282 30052 40666
rect 30196 40044 30248 40050
rect 30196 39986 30248 39992
rect 30104 38956 30156 38962
rect 30104 38898 30156 38904
rect 30012 38276 30064 38282
rect 30012 38218 30064 38224
rect 30116 38010 30144 38898
rect 30208 38214 30236 39986
rect 30392 39846 30420 40870
rect 30484 40730 30512 40870
rect 30472 40724 30524 40730
rect 30472 40666 30524 40672
rect 30472 40384 30524 40390
rect 30576 40372 30604 41074
rect 30656 41064 30708 41070
rect 30656 41006 30708 41012
rect 30840 41064 30892 41070
rect 30840 41006 30892 41012
rect 30524 40344 30604 40372
rect 30472 40326 30524 40332
rect 30380 39840 30432 39846
rect 30380 39782 30432 39788
rect 30484 39642 30512 40326
rect 30668 40089 30696 41006
rect 30748 40112 30800 40118
rect 30654 40080 30710 40089
rect 30748 40054 30800 40060
rect 30654 40015 30710 40024
rect 30472 39636 30524 39642
rect 30472 39578 30524 39584
rect 30656 39432 30708 39438
rect 30656 39374 30708 39380
rect 30564 39364 30616 39370
rect 30564 39306 30616 39312
rect 30472 38888 30524 38894
rect 30576 38865 30604 39306
rect 30472 38830 30524 38836
rect 30562 38856 30618 38865
rect 30288 38752 30340 38758
rect 30288 38694 30340 38700
rect 30300 38593 30328 38694
rect 30286 38584 30342 38593
rect 30286 38519 30342 38528
rect 30484 38418 30512 38830
rect 30562 38791 30618 38800
rect 30472 38412 30524 38418
rect 30472 38354 30524 38360
rect 30576 38350 30604 38791
rect 30668 38758 30696 39374
rect 30656 38752 30708 38758
rect 30656 38694 30708 38700
rect 30760 38457 30788 40054
rect 30746 38448 30802 38457
rect 30746 38383 30802 38392
rect 30564 38344 30616 38350
rect 30852 38332 30880 41006
rect 31208 40384 31260 40390
rect 31208 40326 31260 40332
rect 31484 40384 31536 40390
rect 31484 40326 31536 40332
rect 31220 39982 31248 40326
rect 31208 39976 31260 39982
rect 31208 39918 31260 39924
rect 31208 39568 31260 39574
rect 31208 39510 31260 39516
rect 30932 39364 30984 39370
rect 30932 39306 30984 39312
rect 30564 38286 30616 38292
rect 30668 38304 30880 38332
rect 30380 38276 30432 38282
rect 30380 38218 30432 38224
rect 30196 38208 30248 38214
rect 30196 38150 30248 38156
rect 30288 38208 30340 38214
rect 30288 38150 30340 38156
rect 30104 38004 30156 38010
rect 30104 37946 30156 37952
rect 30012 37868 30064 37874
rect 30012 37810 30064 37816
rect 30024 37262 30052 37810
rect 30116 37330 30144 37946
rect 30300 37466 30328 38150
rect 30288 37460 30340 37466
rect 30288 37402 30340 37408
rect 30104 37324 30156 37330
rect 30104 37266 30156 37272
rect 30012 37256 30064 37262
rect 30010 37224 30012 37233
rect 30064 37224 30066 37233
rect 30010 37159 30066 37168
rect 30104 37188 30156 37194
rect 29920 36100 29972 36106
rect 29920 36042 29972 36048
rect 30024 35698 30052 37159
rect 30104 37130 30156 37136
rect 30196 37188 30248 37194
rect 30196 37130 30248 37136
rect 29644 35692 29696 35698
rect 29644 35634 29696 35640
rect 29736 35692 29788 35698
rect 29736 35634 29788 35640
rect 29828 35692 29880 35698
rect 29828 35634 29880 35640
rect 30012 35692 30064 35698
rect 30012 35634 30064 35640
rect 29642 35592 29698 35601
rect 29748 35578 29776 35634
rect 29698 35550 29776 35578
rect 29642 35527 29698 35536
rect 29644 35488 29696 35494
rect 29644 35430 29696 35436
rect 29656 35329 29684 35430
rect 29642 35320 29698 35329
rect 29642 35255 29698 35264
rect 29656 35086 29684 35255
rect 29644 35080 29696 35086
rect 29644 35022 29696 35028
rect 29472 34972 29592 35000
rect 29368 34604 29420 34610
rect 29368 34546 29420 34552
rect 29274 33552 29330 33561
rect 29274 33487 29330 33496
rect 29288 33386 29316 33487
rect 29276 33380 29328 33386
rect 29276 33322 29328 33328
rect 29184 32224 29236 32230
rect 29184 32166 29236 32172
rect 29288 32042 29316 33322
rect 29564 33318 29592 34972
rect 29748 34542 29776 35550
rect 29736 34536 29788 34542
rect 29736 34478 29788 34484
rect 29552 33312 29604 33318
rect 29552 33254 29604 33260
rect 29368 32904 29420 32910
rect 29368 32846 29420 32852
rect 29196 32014 29316 32042
rect 29000 31952 29052 31958
rect 29000 31894 29052 31900
rect 29092 31952 29144 31958
rect 29092 31894 29144 31900
rect 28908 31816 28960 31822
rect 28908 31758 28960 31764
rect 28816 31680 28868 31686
rect 28816 31622 28868 31628
rect 28724 31408 28776 31414
rect 28724 31350 28776 31356
rect 28724 31272 28776 31278
rect 28724 31214 28776 31220
rect 28736 30938 28764 31214
rect 28724 30932 28776 30938
rect 28724 30874 28776 30880
rect 28828 30734 28856 31622
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 28816 30388 28868 30394
rect 28816 30330 28868 30336
rect 28632 30320 28684 30326
rect 28632 30262 28684 30268
rect 28448 29164 28500 29170
rect 28500 29124 28672 29152
rect 28448 29106 28500 29112
rect 28644 28558 28672 29124
rect 28828 28642 28856 30330
rect 28920 28762 28948 31758
rect 29012 30938 29040 31894
rect 29092 31816 29144 31822
rect 29092 31758 29144 31764
rect 29104 31346 29132 31758
rect 29196 31686 29224 32014
rect 29276 31952 29328 31958
rect 29276 31894 29328 31900
rect 29184 31680 29236 31686
rect 29184 31622 29236 31628
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 29000 30932 29052 30938
rect 29000 30874 29052 30880
rect 29104 30818 29132 31282
rect 29012 30790 29132 30818
rect 29012 29714 29040 30790
rect 29092 30592 29144 30598
rect 29092 30534 29144 30540
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 29012 29345 29040 29650
rect 28998 29336 29054 29345
rect 28998 29271 29054 29280
rect 29000 29096 29052 29102
rect 29000 29038 29052 29044
rect 28908 28756 28960 28762
rect 28908 28698 28960 28704
rect 28828 28614 28948 28642
rect 28632 28552 28684 28558
rect 28632 28494 28684 28500
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28552 27470 28580 28426
rect 28644 27946 28672 28494
rect 28724 28416 28776 28422
rect 28724 28358 28776 28364
rect 28632 27940 28684 27946
rect 28632 27882 28684 27888
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 28356 27396 28408 27402
rect 28356 27338 28408 27344
rect 28092 27084 28212 27112
rect 28264 27124 28316 27130
rect 28092 24818 28120 27084
rect 28264 27066 28316 27072
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 28184 26518 28212 26930
rect 28172 26512 28224 26518
rect 28172 26454 28224 26460
rect 28172 25696 28224 25702
rect 28172 25638 28224 25644
rect 28184 25430 28212 25638
rect 28172 25424 28224 25430
rect 28172 25366 28224 25372
rect 28276 25362 28304 27066
rect 28368 26994 28396 27338
rect 28552 26994 28580 27406
rect 28736 27334 28764 28358
rect 28816 27464 28868 27470
rect 28816 27406 28868 27412
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28828 27130 28856 27406
rect 28816 27124 28868 27130
rect 28816 27066 28868 27072
rect 28722 27024 28778 27033
rect 28356 26988 28408 26994
rect 28356 26930 28408 26936
rect 28540 26988 28592 26994
rect 28722 26959 28724 26968
rect 28540 26930 28592 26936
rect 28776 26959 28778 26968
rect 28724 26930 28776 26936
rect 28354 26888 28410 26897
rect 28354 26823 28356 26832
rect 28408 26823 28410 26832
rect 28356 26794 28408 26800
rect 28540 26784 28592 26790
rect 28540 26726 28592 26732
rect 28356 26240 28408 26246
rect 28356 26182 28408 26188
rect 28368 26081 28396 26182
rect 28354 26072 28410 26081
rect 28354 26007 28410 26016
rect 28368 25362 28396 26007
rect 28264 25356 28316 25362
rect 28264 25298 28316 25304
rect 28356 25356 28408 25362
rect 28356 25298 28408 25304
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28552 24342 28580 26726
rect 28724 25696 28776 25702
rect 28724 25638 28776 25644
rect 28736 25294 28764 25638
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 28736 24886 28764 25230
rect 28816 25152 28868 25158
rect 28816 25094 28868 25100
rect 28724 24880 28776 24886
rect 28724 24822 28776 24828
rect 28828 24698 28856 25094
rect 28644 24670 28856 24698
rect 28540 24336 28592 24342
rect 28540 24278 28592 24284
rect 27710 24103 27766 24112
rect 27896 24132 27948 24138
rect 27620 24074 27672 24080
rect 27528 24064 27580 24070
rect 27528 24006 27580 24012
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 27080 22066 27200 22094
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26804 20466 26832 21422
rect 26792 20460 26844 20466
rect 26792 20402 26844 20408
rect 26804 19922 26832 20402
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 26882 19816 26938 19825
rect 26882 19751 26938 19760
rect 26700 19236 26752 19242
rect 26700 19178 26752 19184
rect 26896 18290 26924 19751
rect 26976 19168 27028 19174
rect 26976 19110 27028 19116
rect 26988 18766 27016 19110
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 26884 18284 26936 18290
rect 26884 18226 26936 18232
rect 26884 18080 26936 18086
rect 26514 18048 26570 18057
rect 26884 18022 26936 18028
rect 26514 17983 26570 17992
rect 26528 16794 26556 17983
rect 26700 17536 26752 17542
rect 26700 17478 26752 17484
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26516 16788 26568 16794
rect 26516 16730 26568 16736
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26528 15858 26556 16526
rect 26620 15978 26648 16934
rect 26712 16590 26740 17478
rect 26700 16584 26752 16590
rect 26700 16526 26752 16532
rect 26712 16114 26740 16526
rect 26792 16448 26844 16454
rect 26792 16390 26844 16396
rect 26804 16250 26832 16390
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26792 16108 26844 16114
rect 26792 16050 26844 16056
rect 26712 15978 26740 16050
rect 26608 15972 26660 15978
rect 26608 15914 26660 15920
rect 26700 15972 26752 15978
rect 26700 15914 26752 15920
rect 26804 15858 26832 16050
rect 26528 15830 26832 15858
rect 26516 15088 26568 15094
rect 26516 15030 26568 15036
rect 26528 14414 26556 15030
rect 26620 14482 26648 15830
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26712 14414 26740 14894
rect 26896 14618 26924 18022
rect 26976 17672 27028 17678
rect 26976 17614 27028 17620
rect 26988 17338 27016 17614
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 26976 16992 27028 16998
rect 26976 16934 27028 16940
rect 26988 16658 27016 16934
rect 26976 16652 27028 16658
rect 26976 16594 27028 16600
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 26384 14368 26464 14396
rect 26516 14408 26568 14414
rect 26332 14350 26384 14356
rect 26516 14350 26568 14356
rect 26700 14408 26752 14414
rect 26896 14362 26924 14554
rect 27080 14414 27108 22066
rect 27160 21004 27212 21010
rect 27264 20992 27292 23802
rect 27540 23769 27568 24006
rect 27526 23760 27582 23769
rect 27526 23695 27582 23704
rect 27528 23656 27580 23662
rect 27528 23598 27580 23604
rect 27434 23488 27490 23497
rect 27434 23423 27490 23432
rect 27448 23186 27476 23423
rect 27540 23254 27568 23598
rect 27528 23248 27580 23254
rect 27528 23190 27580 23196
rect 27436 23180 27488 23186
rect 27436 23122 27488 23128
rect 27632 22409 27660 24074
rect 27724 23254 27752 24103
rect 27896 24074 27948 24080
rect 27712 23248 27764 23254
rect 27712 23190 27764 23196
rect 27618 22400 27674 22409
rect 27618 22335 27674 22344
rect 27526 21992 27582 22001
rect 27526 21927 27528 21936
rect 27580 21927 27582 21936
rect 27528 21898 27580 21904
rect 27436 21888 27488 21894
rect 27436 21830 27488 21836
rect 27212 20964 27292 20992
rect 27160 20946 27212 20952
rect 27448 20942 27476 21830
rect 27908 21729 27936 24074
rect 28264 23792 28316 23798
rect 28264 23734 28316 23740
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 28000 23322 28028 23666
rect 27988 23316 28040 23322
rect 27988 23258 28040 23264
rect 28276 23118 28304 23734
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28172 22976 28224 22982
rect 28172 22918 28224 22924
rect 28448 22976 28500 22982
rect 28448 22918 28500 22924
rect 27894 21720 27950 21729
rect 27894 21655 27950 21664
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 27160 20800 27212 20806
rect 27160 20742 27212 20748
rect 27172 20534 27200 20742
rect 27160 20528 27212 20534
rect 27160 20470 27212 20476
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27172 19854 27200 20198
rect 27540 20058 27568 20946
rect 28184 20874 28212 22918
rect 28460 22778 28488 22918
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28264 21888 28316 21894
rect 28264 21830 28316 21836
rect 28276 21146 28304 21830
rect 28552 21486 28580 24278
rect 28644 22030 28672 24670
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 28828 23118 28856 24550
rect 28920 24070 28948 28614
rect 29012 28558 29040 29038
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 29012 27674 29040 28494
rect 29000 27668 29052 27674
rect 29000 27610 29052 27616
rect 29000 27464 29052 27470
rect 29000 27406 29052 27412
rect 29012 27130 29040 27406
rect 29000 27124 29052 27130
rect 29000 27066 29052 27072
rect 29000 26852 29052 26858
rect 29000 26794 29052 26800
rect 29012 26586 29040 26794
rect 29000 26580 29052 26586
rect 29000 26522 29052 26528
rect 28998 25664 29054 25673
rect 28998 25599 29054 25608
rect 29012 25158 29040 25599
rect 29104 25401 29132 30534
rect 29196 25537 29224 31622
rect 29288 30716 29316 31894
rect 29380 31822 29408 32846
rect 29840 32774 29868 35634
rect 29920 35488 29972 35494
rect 29920 35430 29972 35436
rect 29932 34746 29960 35430
rect 29920 34740 29972 34746
rect 29920 34682 29972 34688
rect 30024 34649 30052 35634
rect 30010 34640 30066 34649
rect 29920 34604 29972 34610
rect 29972 34584 30010 34592
rect 29972 34575 30066 34584
rect 29972 34564 30052 34575
rect 29920 34546 29972 34552
rect 30116 34490 30144 37130
rect 30208 35494 30236 37130
rect 30392 35873 30420 38218
rect 30564 37800 30616 37806
rect 30564 37742 30616 37748
rect 30472 37732 30524 37738
rect 30472 37674 30524 37680
rect 30484 37398 30512 37674
rect 30576 37466 30604 37742
rect 30564 37460 30616 37466
rect 30564 37402 30616 37408
rect 30472 37392 30524 37398
rect 30668 37346 30696 38304
rect 30840 38208 30892 38214
rect 30746 38176 30802 38185
rect 30840 38150 30892 38156
rect 30746 38111 30802 38120
rect 30472 37334 30524 37340
rect 30576 37318 30696 37346
rect 30378 35864 30434 35873
rect 30378 35799 30434 35808
rect 30288 35624 30340 35630
rect 30288 35566 30340 35572
rect 30380 35624 30432 35630
rect 30380 35566 30432 35572
rect 30196 35488 30248 35494
rect 30196 35430 30248 35436
rect 30196 34944 30248 34950
rect 30196 34886 30248 34892
rect 29932 34462 30144 34490
rect 29828 32768 29880 32774
rect 29828 32710 29880 32716
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29368 31816 29420 31822
rect 29368 31758 29420 31764
rect 29380 31346 29408 31758
rect 29368 31340 29420 31346
rect 29368 31282 29420 31288
rect 29564 30870 29592 32506
rect 29734 32056 29790 32065
rect 29734 31991 29736 32000
rect 29788 31991 29790 32000
rect 29736 31962 29788 31968
rect 29932 31958 29960 34462
rect 30208 34184 30236 34886
rect 30300 34785 30328 35566
rect 30392 35290 30420 35566
rect 30470 35456 30526 35465
rect 30470 35391 30526 35400
rect 30380 35284 30432 35290
rect 30380 35226 30432 35232
rect 30392 35086 30420 35226
rect 30484 35222 30512 35391
rect 30472 35216 30524 35222
rect 30472 35158 30524 35164
rect 30380 35080 30432 35086
rect 30380 35022 30432 35028
rect 30380 34944 30432 34950
rect 30378 34912 30380 34921
rect 30472 34944 30524 34950
rect 30432 34912 30434 34921
rect 30472 34886 30524 34892
rect 30378 34847 30434 34856
rect 30286 34776 30342 34785
rect 30286 34711 30288 34720
rect 30340 34711 30342 34720
rect 30288 34682 30340 34688
rect 30288 34604 30340 34610
rect 30288 34546 30340 34552
rect 30116 34156 30236 34184
rect 30116 33998 30144 34156
rect 30196 34060 30248 34066
rect 30196 34002 30248 34008
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30012 33516 30064 33522
rect 30012 33458 30064 33464
rect 30024 33046 30052 33458
rect 30208 33114 30236 34002
rect 30300 33522 30328 34546
rect 30288 33516 30340 33522
rect 30288 33458 30340 33464
rect 30196 33108 30248 33114
rect 30196 33050 30248 33056
rect 30012 33040 30064 33046
rect 30012 32982 30064 32988
rect 30104 32972 30156 32978
rect 30104 32914 30156 32920
rect 30116 32774 30144 32914
rect 30208 32910 30236 33050
rect 30196 32904 30248 32910
rect 30196 32846 30248 32852
rect 30104 32768 30156 32774
rect 30104 32710 30156 32716
rect 30196 32768 30248 32774
rect 30196 32710 30248 32716
rect 30104 32428 30156 32434
rect 30104 32370 30156 32376
rect 30012 32224 30064 32230
rect 30012 32166 30064 32172
rect 30024 32026 30052 32166
rect 30012 32020 30064 32026
rect 30012 31962 30064 31968
rect 29920 31952 29972 31958
rect 29920 31894 29972 31900
rect 30024 31754 30052 31962
rect 29932 31726 30052 31754
rect 29828 31272 29880 31278
rect 29828 31214 29880 31220
rect 29368 30864 29420 30870
rect 29366 30832 29368 30841
rect 29552 30864 29604 30870
rect 29420 30832 29422 30841
rect 29552 30806 29604 30812
rect 29642 30832 29698 30841
rect 29366 30767 29422 30776
rect 29642 30767 29644 30776
rect 29696 30767 29698 30776
rect 29644 30738 29696 30744
rect 29368 30728 29420 30734
rect 29288 30688 29368 30716
rect 29368 30670 29420 30676
rect 29460 30592 29512 30598
rect 29460 30534 29512 30540
rect 29276 29028 29328 29034
rect 29276 28970 29328 28976
rect 29288 27878 29316 28970
rect 29368 28008 29420 28014
rect 29368 27950 29420 27956
rect 29276 27872 29328 27878
rect 29276 27814 29328 27820
rect 29276 27532 29328 27538
rect 29276 27474 29328 27480
rect 29182 25528 29238 25537
rect 29182 25463 29238 25472
rect 29288 25412 29316 27474
rect 29380 27334 29408 27950
rect 29368 27328 29420 27334
rect 29368 27270 29420 27276
rect 29090 25392 29146 25401
rect 29090 25327 29146 25336
rect 29196 25384 29316 25412
rect 29092 25288 29144 25294
rect 29196 25276 29224 25384
rect 29144 25248 29224 25276
rect 29274 25256 29330 25265
rect 29092 25230 29144 25236
rect 29274 25191 29330 25200
rect 29000 25152 29052 25158
rect 29000 25094 29052 25100
rect 29090 25120 29146 25129
rect 29090 25055 29146 25064
rect 28908 24064 28960 24070
rect 28908 24006 28960 24012
rect 29104 23576 29132 25055
rect 29288 24954 29316 25191
rect 29276 24948 29328 24954
rect 29276 24890 29328 24896
rect 29274 24848 29330 24857
rect 29274 24783 29330 24792
rect 29184 24608 29236 24614
rect 29184 24550 29236 24556
rect 29196 23662 29224 24550
rect 29288 24138 29316 24783
rect 29276 24132 29328 24138
rect 29276 24074 29328 24080
rect 29184 23656 29236 23662
rect 29184 23598 29236 23604
rect 28920 23548 29132 23576
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 28920 22166 28948 23548
rect 29000 23180 29052 23186
rect 29000 23122 29052 23128
rect 29012 22642 29040 23122
rect 29092 23112 29144 23118
rect 29092 23054 29144 23060
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 29012 22234 29040 22578
rect 29000 22228 29052 22234
rect 29000 22170 29052 22176
rect 28908 22160 28960 22166
rect 28908 22102 28960 22108
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28644 21622 28672 21966
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28264 21140 28316 21146
rect 28264 21082 28316 21088
rect 28448 21140 28500 21146
rect 28552 21128 28580 21422
rect 28632 21412 28684 21418
rect 28632 21354 28684 21360
rect 28500 21100 28580 21128
rect 28448 21082 28500 21088
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 28552 20534 28580 20742
rect 28540 20528 28592 20534
rect 28540 20470 28592 20476
rect 28540 20392 28592 20398
rect 28644 20346 28672 21354
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28920 20942 28948 21286
rect 29012 20942 29040 22170
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 28908 20800 28960 20806
rect 28908 20742 28960 20748
rect 28592 20340 28672 20346
rect 28540 20334 28672 20340
rect 28552 20318 28672 20334
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27264 18902 27292 19994
rect 28552 19786 28580 20318
rect 28540 19780 28592 19786
rect 28540 19722 28592 19728
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 27252 18896 27304 18902
rect 27252 18838 27304 18844
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 27172 18426 27200 18566
rect 27160 18420 27212 18426
rect 27160 18362 27212 18368
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27264 17678 27292 18022
rect 27252 17672 27304 17678
rect 27252 17614 27304 17620
rect 27356 17218 27384 18226
rect 27448 17882 27476 19382
rect 27712 19372 27764 19378
rect 27712 19314 27764 19320
rect 27526 18456 27582 18465
rect 27526 18391 27582 18400
rect 27540 18290 27568 18391
rect 27724 18290 27752 19314
rect 28552 18698 28580 19722
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 28540 18692 28592 18698
rect 28540 18634 28592 18640
rect 27804 18420 27856 18426
rect 27804 18362 27856 18368
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27436 17876 27488 17882
rect 27436 17818 27488 17824
rect 27356 17202 27476 17218
rect 27356 17196 27488 17202
rect 27356 17190 27436 17196
rect 27436 17138 27488 17144
rect 27158 16416 27214 16425
rect 27158 16351 27214 16360
rect 26700 14350 26752 14356
rect 26252 13926 26464 13954
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26252 11762 26280 13670
rect 26436 13326 26464 13926
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26528 13258 26556 14350
rect 26608 14340 26660 14346
rect 26608 14282 26660 14288
rect 26332 13252 26384 13258
rect 26332 13194 26384 13200
rect 26516 13252 26568 13258
rect 26516 13194 26568 13200
rect 26344 12434 26372 13194
rect 26620 12646 26648 14282
rect 26712 13326 26740 14350
rect 26804 14334 26924 14362
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 26804 13802 26832 14334
rect 26884 14272 26936 14278
rect 26884 14214 26936 14220
rect 26976 14272 27028 14278
rect 26976 14214 27028 14220
rect 26896 13938 26924 14214
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 26792 13796 26844 13802
rect 26792 13738 26844 13744
rect 26790 13560 26846 13569
rect 26790 13495 26846 13504
rect 26700 13320 26752 13326
rect 26698 13288 26700 13297
rect 26752 13288 26754 13297
rect 26698 13223 26754 13232
rect 26804 13190 26832 13495
rect 26700 13184 26752 13190
rect 26700 13126 26752 13132
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26608 12640 26660 12646
rect 26608 12582 26660 12588
rect 26344 12406 26648 12434
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26528 11898 26556 12038
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26514 11792 26570 11801
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26332 11756 26384 11762
rect 26384 11716 26464 11744
rect 26514 11727 26516 11736
rect 26332 11698 26384 11704
rect 26056 11620 26108 11626
rect 26056 11562 26108 11568
rect 25962 11384 26018 11393
rect 25962 11319 26018 11328
rect 25976 11286 26004 11319
rect 25964 11280 26016 11286
rect 25964 11222 26016 11228
rect 25964 11144 26016 11150
rect 25686 11047 25742 11056
rect 25792 11070 25912 11098
rect 25962 11112 25964 11121
rect 26016 11112 26018 11121
rect 25688 10668 25740 10674
rect 25688 10610 25740 10616
rect 25700 10130 25728 10610
rect 25688 10124 25740 10130
rect 25688 10066 25740 10072
rect 25594 9616 25650 9625
rect 25594 9551 25650 9560
rect 25688 9580 25740 9586
rect 25608 9110 25636 9551
rect 25688 9522 25740 9528
rect 25596 9104 25648 9110
rect 25596 9046 25648 9052
rect 25504 8560 25556 8566
rect 25504 8502 25556 8508
rect 25228 8424 25280 8430
rect 25148 8384 25228 8412
rect 25148 7886 25176 8384
rect 25228 8366 25280 8372
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 25240 7546 25268 7822
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25136 7268 25188 7274
rect 25136 7210 25188 7216
rect 25148 6798 25176 7210
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25044 5636 25096 5642
rect 25044 5578 25096 5584
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24964 4826 24992 5170
rect 24952 4820 25004 4826
rect 24952 4762 25004 4768
rect 25056 4690 25084 5578
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 25148 4622 25176 5306
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 25240 4146 25268 7346
rect 25332 6866 25360 7822
rect 25608 7546 25636 7890
rect 25700 7886 25728 9522
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25700 7410 25728 7822
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25504 6112 25556 6118
rect 25504 6054 25556 6060
rect 25516 5710 25544 6054
rect 25792 5778 25820 11070
rect 25962 11047 26018 11056
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25884 9994 25912 10950
rect 26068 10674 26096 11562
rect 26148 11280 26200 11286
rect 26436 11257 26464 11716
rect 26568 11727 26570 11736
rect 26516 11698 26568 11704
rect 26528 11286 26556 11698
rect 26516 11280 26568 11286
rect 26148 11222 26200 11228
rect 26422 11248 26478 11257
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 25976 10470 26004 10610
rect 25964 10464 26016 10470
rect 25964 10406 26016 10412
rect 25976 10266 26004 10406
rect 25964 10260 26016 10266
rect 25964 10202 26016 10208
rect 25872 9988 25924 9994
rect 25872 9930 25924 9936
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25870 9480 25926 9489
rect 25870 9415 25872 9424
rect 25924 9415 25926 9424
rect 25872 9386 25924 9392
rect 25976 7886 26004 9522
rect 26068 8090 26096 10610
rect 26160 9674 26188 11222
rect 26516 11222 26568 11228
rect 26422 11183 26478 11192
rect 26436 11132 26464 11183
rect 26516 11144 26568 11150
rect 26436 11104 26516 11132
rect 26516 11086 26568 11092
rect 26240 11076 26292 11082
rect 26292 11036 26464 11064
rect 26240 11018 26292 11024
rect 26238 10976 26294 10985
rect 26238 10911 26294 10920
rect 26252 10674 26280 10911
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26436 10266 26464 11036
rect 26514 10976 26570 10985
rect 26514 10911 26570 10920
rect 26528 10810 26556 10911
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26160 9646 26464 9674
rect 26436 9586 26464 9646
rect 26620 9586 26648 12406
rect 26712 11082 26740 13126
rect 26988 12238 27016 14214
rect 27068 13320 27120 13326
rect 27068 13262 27120 13268
rect 27080 12714 27108 13262
rect 27068 12708 27120 12714
rect 27068 12650 27120 12656
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26896 11898 26924 12038
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 26988 11762 27016 12174
rect 27080 11762 27108 12174
rect 27172 11778 27200 16351
rect 27252 16108 27304 16114
rect 27252 16050 27304 16056
rect 27264 15570 27292 16050
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 27252 15088 27304 15094
rect 27252 15030 27304 15036
rect 27264 14074 27292 15030
rect 27342 14512 27398 14521
rect 27342 14447 27398 14456
rect 27356 14074 27384 14447
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27344 14068 27396 14074
rect 27344 14010 27396 14016
rect 27344 13796 27396 13802
rect 27344 13738 27396 13744
rect 27252 13728 27304 13734
rect 27252 13670 27304 13676
rect 27264 12238 27292 13670
rect 27356 13258 27384 13738
rect 27344 13252 27396 13258
rect 27344 13194 27396 13200
rect 27252 12232 27304 12238
rect 27252 12174 27304 12180
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 27068 11756 27120 11762
rect 27172 11750 27292 11778
rect 27068 11698 27120 11704
rect 26792 11688 26844 11694
rect 26792 11630 26844 11636
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26712 10674 26740 11018
rect 26804 10674 26832 11630
rect 26884 11552 26936 11558
rect 26882 11520 26884 11529
rect 26936 11520 26938 11529
rect 26882 11455 26938 11464
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 26896 10810 26924 11086
rect 26884 10804 26936 10810
rect 26884 10746 26936 10752
rect 26988 10713 27016 11086
rect 26974 10704 27030 10713
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26792 10668 26844 10674
rect 26974 10639 27030 10648
rect 26792 10610 26844 10616
rect 26988 10062 27016 10639
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26424 9580 26476 9586
rect 26424 9522 26476 9528
rect 26608 9580 26660 9586
rect 26608 9522 26660 9528
rect 27160 9580 27212 9586
rect 27264 9568 27292 11750
rect 27356 11694 27384 12174
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27356 10742 27384 11630
rect 27448 10810 27476 17138
rect 27540 15026 27568 18226
rect 27712 18080 27764 18086
rect 27712 18022 27764 18028
rect 27724 17678 27752 18022
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27712 16584 27764 16590
rect 27712 16526 27764 16532
rect 27724 16289 27752 16526
rect 27710 16280 27766 16289
rect 27710 16215 27766 16224
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 27724 15026 27752 15098
rect 27816 15026 27844 18362
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27620 14884 27672 14890
rect 27620 14826 27672 14832
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27540 14618 27568 14758
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 27632 14278 27660 14826
rect 27816 14414 27844 14962
rect 27804 14408 27856 14414
rect 27710 14376 27766 14385
rect 27804 14350 27856 14356
rect 27710 14311 27766 14320
rect 27724 14278 27752 14311
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27816 13954 27844 14350
rect 27724 13938 27844 13954
rect 27712 13932 27844 13938
rect 27764 13926 27844 13932
rect 27712 13874 27764 13880
rect 27724 13462 27752 13874
rect 27712 13456 27764 13462
rect 27712 13398 27764 13404
rect 27908 12434 27936 14962
rect 27724 12406 27936 12434
rect 28000 12434 28028 18226
rect 28092 15026 28120 18226
rect 28356 18216 28408 18222
rect 28356 18158 28408 18164
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 28184 16153 28212 16458
rect 28170 16144 28226 16153
rect 28170 16079 28226 16088
rect 28170 15192 28226 15201
rect 28368 15162 28396 18158
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28552 16590 28580 17478
rect 28540 16584 28592 16590
rect 28540 16526 28592 16532
rect 28552 16114 28580 16526
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 28170 15127 28226 15136
rect 28356 15156 28408 15162
rect 28080 15020 28132 15026
rect 28080 14962 28132 14968
rect 28184 14906 28212 15127
rect 28356 15098 28408 15104
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28092 14878 28212 14906
rect 28092 13870 28120 14878
rect 28172 14816 28224 14822
rect 28172 14758 28224 14764
rect 28184 14618 28212 14758
rect 28172 14612 28224 14618
rect 28172 14554 28224 14560
rect 28172 14272 28224 14278
rect 28172 14214 28224 14220
rect 28184 14113 28212 14214
rect 28170 14104 28226 14113
rect 28170 14039 28226 14048
rect 28276 13938 28304 14962
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28264 13932 28316 13938
rect 28264 13874 28316 13880
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 28368 13802 28396 14350
rect 28448 13864 28500 13870
rect 28448 13806 28500 13812
rect 28356 13796 28408 13802
rect 28356 13738 28408 13744
rect 28368 13326 28396 13738
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 28000 12406 28120 12434
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 27344 10736 27396 10742
rect 27344 10678 27396 10684
rect 27528 9580 27580 9586
rect 27264 9540 27528 9568
rect 27160 9522 27212 9528
rect 26620 9489 26648 9522
rect 26884 9512 26936 9518
rect 26606 9480 26662 9489
rect 26884 9454 26936 9460
rect 26606 9415 26662 9424
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26160 7886 26188 9318
rect 26344 8974 26372 9318
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 26424 8832 26476 8838
rect 26424 8774 26476 8780
rect 26436 8634 26464 8774
rect 26424 8628 26476 8634
rect 26424 8570 26476 8576
rect 25964 7880 26016 7886
rect 25870 7848 25926 7857
rect 25926 7828 25964 7834
rect 25926 7822 26016 7828
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 25926 7806 26004 7822
rect 25870 7783 25926 7792
rect 25976 7410 26004 7806
rect 26056 7812 26108 7818
rect 26056 7754 26108 7760
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25780 5772 25832 5778
rect 25780 5714 25832 5720
rect 25504 5704 25556 5710
rect 25504 5646 25556 5652
rect 25962 5264 26018 5273
rect 25962 5199 26018 5208
rect 25320 5160 25372 5166
rect 25320 5102 25372 5108
rect 25228 4140 25280 4146
rect 25228 4082 25280 4088
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24688 3618 24716 4014
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24780 3738 24808 3878
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 24688 3590 24808 3618
rect 24596 3466 24624 3538
rect 24688 3534 24716 3590
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24584 3460 24636 3466
rect 24584 3402 24636 3408
rect 24780 3126 24808 3590
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 24872 2854 24900 3334
rect 25240 3194 25268 4082
rect 25332 3738 25360 5102
rect 25976 4690 26004 5199
rect 25964 4684 26016 4690
rect 25964 4626 26016 4632
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25596 4004 25648 4010
rect 25596 3946 25648 3952
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 25332 3058 25360 3674
rect 25608 3602 25636 3946
rect 25596 3596 25648 3602
rect 25596 3538 25648 3544
rect 25700 3194 25728 4082
rect 25872 3392 25924 3398
rect 25976 3346 26004 4626
rect 26068 3738 26096 7754
rect 26160 7392 26188 7822
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26344 7478 26372 7686
rect 26712 7546 26740 9114
rect 26804 8974 26832 9318
rect 26896 9042 26924 9454
rect 27172 9042 27200 9522
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 27160 9036 27212 9042
rect 27160 8978 27212 8984
rect 26792 8968 26844 8974
rect 26792 8910 26844 8916
rect 26988 7750 27016 8978
rect 26976 7744 27028 7750
rect 26976 7686 27028 7692
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 26240 7404 26292 7410
rect 26160 7364 26240 7392
rect 26160 6934 26188 7364
rect 26240 7346 26292 7352
rect 26608 7268 26660 7274
rect 26608 7210 26660 7216
rect 26620 7002 26648 7210
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 26148 6928 26200 6934
rect 26148 6870 26200 6876
rect 26332 6928 26384 6934
rect 26332 6870 26384 6876
rect 26148 6724 26200 6730
rect 26148 6666 26200 6672
rect 26160 6458 26188 6666
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26252 6458 26280 6598
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 26240 4752 26292 4758
rect 26240 4694 26292 4700
rect 26252 4282 26280 4694
rect 26344 4690 26372 6870
rect 26620 6798 26648 6938
rect 26712 6866 26740 7482
rect 27356 6866 27384 9540
rect 27528 9522 27580 9528
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27436 8900 27488 8906
rect 27632 8888 27660 9114
rect 27488 8860 27660 8888
rect 27436 8842 27488 8848
rect 27632 8634 27660 8860
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27540 7342 27568 7686
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 27436 6996 27488 7002
rect 27436 6938 27488 6944
rect 27448 6866 27476 6938
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27436 6860 27488 6866
rect 27436 6802 27488 6808
rect 26608 6792 26660 6798
rect 26608 6734 26660 6740
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 26976 6724 27028 6730
rect 26976 6666 27028 6672
rect 26988 6458 27016 6666
rect 26976 6452 27028 6458
rect 26976 6394 27028 6400
rect 27080 6118 27108 6734
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 27068 6112 27120 6118
rect 27068 6054 27120 6060
rect 26528 5778 26556 6054
rect 26516 5772 26568 5778
rect 26516 5714 26568 5720
rect 26528 5166 26556 5714
rect 26608 5228 26660 5234
rect 26608 5170 26660 5176
rect 26516 5160 26568 5166
rect 26516 5102 26568 5108
rect 26528 4826 26556 5102
rect 26516 4820 26568 4826
rect 26516 4762 26568 4768
rect 26332 4684 26384 4690
rect 26332 4626 26384 4632
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26620 4010 26648 5170
rect 26700 4548 26752 4554
rect 26700 4490 26752 4496
rect 26712 4282 26740 4490
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26608 4004 26660 4010
rect 26608 3946 26660 3952
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 25924 3340 26004 3346
rect 25872 3334 26004 3340
rect 25884 3318 26004 3334
rect 25976 3194 26004 3318
rect 26068 3194 26096 3674
rect 26620 3534 26648 3946
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 27540 2990 27568 7278
rect 27724 5370 27752 12406
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 27804 9920 27856 9926
rect 27804 9862 27856 9868
rect 27816 8906 27844 9862
rect 28000 9518 28028 9998
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 27988 9512 28040 9518
rect 27988 9454 28040 9460
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27908 8634 27936 9454
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 28092 8022 28120 12406
rect 28080 8016 28132 8022
rect 28080 7958 28132 7964
rect 27712 5364 27764 5370
rect 27712 5306 27764 5312
rect 28092 4826 28120 7958
rect 28460 7290 28488 13806
rect 28644 12782 28672 19314
rect 28816 16652 28868 16658
rect 28816 16594 28868 16600
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28632 12776 28684 12782
rect 28632 12718 28684 12724
rect 28736 12442 28764 16390
rect 28828 15910 28856 16594
rect 28816 15904 28868 15910
rect 28816 15846 28868 15852
rect 28816 12912 28868 12918
rect 28816 12854 28868 12860
rect 28724 12436 28776 12442
rect 28724 12378 28776 12384
rect 28540 12096 28592 12102
rect 28540 12038 28592 12044
rect 28552 11830 28580 12038
rect 28632 11892 28684 11898
rect 28632 11834 28684 11840
rect 28540 11824 28592 11830
rect 28540 11766 28592 11772
rect 28644 9586 28672 11834
rect 28540 9580 28592 9586
rect 28540 9522 28592 9528
rect 28632 9580 28684 9586
rect 28632 9522 28684 9528
rect 28552 9110 28580 9522
rect 28644 9178 28672 9522
rect 28632 9172 28684 9178
rect 28632 9114 28684 9120
rect 28540 9104 28592 9110
rect 28540 9046 28592 9052
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28644 8566 28672 8910
rect 28632 8560 28684 8566
rect 28684 8508 28764 8514
rect 28632 8502 28764 8508
rect 28644 8486 28764 8502
rect 28460 7262 28672 7290
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 28368 6254 28396 6666
rect 28552 6458 28580 7142
rect 28644 6798 28672 7262
rect 28632 6792 28684 6798
rect 28632 6734 28684 6740
rect 28540 6452 28592 6458
rect 28540 6394 28592 6400
rect 28736 6322 28764 8486
rect 28724 6316 28776 6322
rect 28724 6258 28776 6264
rect 28356 6248 28408 6254
rect 28356 6190 28408 6196
rect 28368 5234 28396 6190
rect 28828 5710 28856 12854
rect 28920 12442 28948 20742
rect 29000 19168 29052 19174
rect 29000 19110 29052 19116
rect 29012 17678 29040 19110
rect 29104 18222 29132 23054
rect 29184 22568 29236 22574
rect 29184 22510 29236 22516
rect 29196 19378 29224 22510
rect 29380 21570 29408 27270
rect 29288 21542 29408 21570
rect 29288 21146 29316 21542
rect 29472 21486 29500 30534
rect 29840 30394 29868 31214
rect 29828 30388 29880 30394
rect 29828 30330 29880 30336
rect 29642 30288 29698 30297
rect 29642 30223 29698 30232
rect 29552 29504 29604 29510
rect 29552 29446 29604 29452
rect 29564 28558 29592 29446
rect 29656 29102 29684 30223
rect 29932 30190 29960 31726
rect 30116 31142 30144 32370
rect 30208 32366 30236 32710
rect 30300 32570 30328 33458
rect 30380 33108 30432 33114
rect 30380 33050 30432 33056
rect 30392 32842 30420 33050
rect 30380 32836 30432 32842
rect 30380 32778 30432 32784
rect 30288 32564 30340 32570
rect 30288 32506 30340 32512
rect 30196 32360 30248 32366
rect 30196 32302 30248 32308
rect 30288 32224 30340 32230
rect 30288 32166 30340 32172
rect 30300 31822 30328 32166
rect 30392 31822 30420 32778
rect 30288 31816 30340 31822
rect 30288 31758 30340 31764
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30196 31340 30248 31346
rect 30196 31282 30248 31288
rect 30104 31136 30156 31142
rect 30104 31078 30156 31084
rect 30116 30190 30144 31078
rect 29920 30184 29972 30190
rect 29920 30126 29972 30132
rect 30104 30184 30156 30190
rect 30104 30126 30156 30132
rect 29828 29776 29880 29782
rect 29828 29718 29880 29724
rect 29840 29102 29868 29718
rect 29644 29096 29696 29102
rect 29828 29096 29880 29102
rect 29644 29038 29696 29044
rect 29826 29064 29828 29073
rect 29880 29064 29882 29073
rect 29826 28999 29882 29008
rect 29642 28928 29698 28937
rect 29642 28863 29698 28872
rect 29656 28762 29684 28863
rect 29644 28756 29696 28762
rect 29644 28698 29696 28704
rect 29552 28552 29604 28558
rect 29552 28494 29604 28500
rect 29552 27940 29604 27946
rect 29552 27882 29604 27888
rect 29564 27538 29592 27882
rect 29552 27532 29604 27538
rect 29552 27474 29604 27480
rect 29656 27470 29684 28698
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29840 27946 29868 28494
rect 29932 28490 29960 30126
rect 30208 30054 30236 31282
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30104 30048 30156 30054
rect 30104 29990 30156 29996
rect 30196 30048 30248 30054
rect 30196 29990 30248 29996
rect 30116 29646 30144 29990
rect 30208 29850 30236 29990
rect 30196 29844 30248 29850
rect 30196 29786 30248 29792
rect 30300 29646 30328 30194
rect 30104 29640 30156 29646
rect 30104 29582 30156 29588
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30012 29504 30064 29510
rect 30012 29446 30064 29452
rect 30024 29170 30052 29446
rect 30300 29238 30328 29582
rect 30104 29232 30156 29238
rect 30104 29174 30156 29180
rect 30288 29232 30340 29238
rect 30288 29174 30340 29180
rect 30012 29164 30064 29170
rect 30012 29106 30064 29112
rect 30116 28914 30144 29174
rect 30392 29102 30420 29582
rect 30380 29096 30432 29102
rect 30380 29038 30432 29044
rect 30196 28960 30248 28966
rect 30116 28908 30196 28914
rect 30116 28902 30248 28908
rect 30116 28886 30236 28902
rect 30208 28558 30236 28886
rect 30196 28552 30248 28558
rect 30196 28494 30248 28500
rect 29920 28484 29972 28490
rect 29920 28426 29972 28432
rect 30288 28416 30340 28422
rect 30288 28358 30340 28364
rect 29828 27940 29880 27946
rect 29828 27882 29880 27888
rect 29644 27464 29696 27470
rect 29644 27406 29696 27412
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 29564 26926 29592 27270
rect 29840 26994 29868 27882
rect 30196 27872 30248 27878
rect 30196 27814 30248 27820
rect 30104 27396 30156 27402
rect 30104 27338 30156 27344
rect 29828 26988 29880 26994
rect 29828 26930 29880 26936
rect 29552 26920 29604 26926
rect 29552 26862 29604 26868
rect 30116 26858 30144 27338
rect 30208 27130 30236 27814
rect 30196 27124 30248 27130
rect 30196 27066 30248 27072
rect 30104 26852 30156 26858
rect 30104 26794 30156 26800
rect 29644 26784 29696 26790
rect 29644 26726 29696 26732
rect 30012 26784 30064 26790
rect 30012 26726 30064 26732
rect 29552 25832 29604 25838
rect 29552 25774 29604 25780
rect 29564 23118 29592 25774
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29552 22432 29604 22438
rect 29552 22374 29604 22380
rect 29564 22166 29592 22374
rect 29552 22160 29604 22166
rect 29552 22102 29604 22108
rect 29368 21480 29420 21486
rect 29368 21422 29420 21428
rect 29460 21480 29512 21486
rect 29460 21422 29512 21428
rect 29380 21146 29408 21422
rect 29276 21140 29328 21146
rect 29276 21082 29328 21088
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 29550 21040 29606 21049
rect 29550 20975 29552 20984
rect 29604 20975 29606 20984
rect 29552 20946 29604 20952
rect 29656 20584 29684 26726
rect 30024 26489 30052 26726
rect 30010 26480 30066 26489
rect 30010 26415 30066 26424
rect 29734 25664 29790 25673
rect 29734 25599 29790 25608
rect 29748 25294 29776 25599
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 29736 25152 29788 25158
rect 29736 25094 29788 25100
rect 29748 22642 29776 25094
rect 30196 24336 30248 24342
rect 30196 24278 30248 24284
rect 30012 23656 30064 23662
rect 30012 23598 30064 23604
rect 30024 23322 30052 23598
rect 30012 23316 30064 23322
rect 30012 23258 30064 23264
rect 29920 23248 29972 23254
rect 29920 23190 29972 23196
rect 29932 22642 29960 23190
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 30024 21962 30052 23258
rect 30208 22094 30236 24278
rect 30300 24274 30328 28358
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 30392 27674 30420 27814
rect 30380 27668 30432 27674
rect 30380 27610 30432 27616
rect 30484 26450 30512 34886
rect 30576 34513 30604 37318
rect 30656 37256 30708 37262
rect 30656 37198 30708 37204
rect 30668 35766 30696 37198
rect 30656 35760 30708 35766
rect 30656 35702 30708 35708
rect 30668 35329 30696 35702
rect 30760 35698 30788 38111
rect 30852 38010 30880 38150
rect 30840 38004 30892 38010
rect 30840 37946 30892 37952
rect 30944 37346 30972 39306
rect 31024 39024 31076 39030
rect 31022 38992 31024 39001
rect 31076 38992 31078 39001
rect 31022 38927 31078 38936
rect 31116 38888 31168 38894
rect 31116 38830 31168 38836
rect 31024 38752 31076 38758
rect 31024 38694 31076 38700
rect 31036 38554 31064 38694
rect 31024 38548 31076 38554
rect 31024 38490 31076 38496
rect 31128 37670 31156 38830
rect 31220 38758 31248 39510
rect 31392 39364 31444 39370
rect 31392 39306 31444 39312
rect 31208 38752 31260 38758
rect 31208 38694 31260 38700
rect 31300 37868 31352 37874
rect 31300 37810 31352 37816
rect 31208 37800 31260 37806
rect 31208 37742 31260 37748
rect 31116 37664 31168 37670
rect 31116 37606 31168 37612
rect 30852 37318 30972 37346
rect 31024 37392 31076 37398
rect 31024 37334 31076 37340
rect 30852 37262 30880 37318
rect 30840 37256 30892 37262
rect 30840 37198 30892 37204
rect 30932 37256 30984 37262
rect 30932 37198 30984 37204
rect 30748 35692 30800 35698
rect 30748 35634 30800 35640
rect 30852 35494 30880 37198
rect 30944 36922 30972 37198
rect 31036 37176 31064 37334
rect 31220 37330 31248 37742
rect 31208 37324 31260 37330
rect 31208 37266 31260 37272
rect 31208 37188 31260 37194
rect 31036 37148 31208 37176
rect 30932 36916 30984 36922
rect 30932 36858 30984 36864
rect 30932 36780 30984 36786
rect 30932 36722 30984 36728
rect 30840 35488 30892 35494
rect 30944 35465 30972 36722
rect 30840 35430 30892 35436
rect 30930 35456 30986 35465
rect 30930 35391 30986 35400
rect 30654 35320 30710 35329
rect 30654 35255 30710 35264
rect 30668 35000 30696 35255
rect 30944 35222 30972 35391
rect 30932 35216 30984 35222
rect 30932 35158 30984 35164
rect 30668 34972 30788 35000
rect 30654 34912 30710 34921
rect 30654 34847 30710 34856
rect 30668 34746 30696 34847
rect 30656 34740 30708 34746
rect 30656 34682 30708 34688
rect 30760 34678 30788 34972
rect 30840 34944 30892 34950
rect 30840 34886 30892 34892
rect 30852 34746 30880 34886
rect 30840 34740 30892 34746
rect 30840 34682 30892 34688
rect 30748 34672 30800 34678
rect 30852 34649 30880 34682
rect 30748 34614 30800 34620
rect 30838 34640 30894 34649
rect 30838 34575 30894 34584
rect 30562 34504 30618 34513
rect 30562 34439 30618 34448
rect 30656 34196 30708 34202
rect 30656 34138 30708 34144
rect 30668 33454 30696 34138
rect 30656 33448 30708 33454
rect 30656 33390 30708 33396
rect 30668 32298 30696 33390
rect 30840 32836 30892 32842
rect 30840 32778 30892 32784
rect 30932 32836 30984 32842
rect 30932 32778 30984 32784
rect 30852 32502 30880 32778
rect 30840 32496 30892 32502
rect 30840 32438 30892 32444
rect 30944 32434 30972 32778
rect 30932 32428 30984 32434
rect 30932 32370 30984 32376
rect 30656 32292 30708 32298
rect 30656 32234 30708 32240
rect 30840 32224 30892 32230
rect 30840 32166 30892 32172
rect 30852 32026 30880 32166
rect 30944 32026 30972 32370
rect 30840 32020 30892 32026
rect 30840 31962 30892 31968
rect 30932 32020 30984 32026
rect 30932 31962 30984 31968
rect 30932 31680 30984 31686
rect 30930 31648 30932 31657
rect 30984 31648 30986 31657
rect 30930 31583 30986 31592
rect 31036 31482 31064 37148
rect 31208 37130 31260 37136
rect 31208 36372 31260 36378
rect 31208 36314 31260 36320
rect 31220 35834 31248 36314
rect 31312 36242 31340 37810
rect 31404 36802 31432 39306
rect 31496 39098 31524 40326
rect 31588 39438 31616 41414
rect 31680 41138 31708 42094
rect 32692 41818 32720 42094
rect 32680 41812 32732 41818
rect 32680 41754 32732 41760
rect 32588 41676 32640 41682
rect 32588 41618 32640 41624
rect 32404 41540 32456 41546
rect 32404 41482 32456 41488
rect 31668 41132 31720 41138
rect 31668 41074 31720 41080
rect 32416 41070 32444 41482
rect 32404 41064 32456 41070
rect 32404 41006 32456 41012
rect 32600 40594 32628 41618
rect 32588 40588 32640 40594
rect 32588 40530 32640 40536
rect 32220 40452 32272 40458
rect 32220 40394 32272 40400
rect 32772 40452 32824 40458
rect 32772 40394 32824 40400
rect 32232 40186 32260 40394
rect 32588 40384 32640 40390
rect 32588 40326 32640 40332
rect 32600 40186 32628 40326
rect 32220 40180 32272 40186
rect 32220 40122 32272 40128
rect 32588 40180 32640 40186
rect 32588 40122 32640 40128
rect 31668 39976 31720 39982
rect 31668 39918 31720 39924
rect 32310 39944 32366 39953
rect 31576 39432 31628 39438
rect 31576 39374 31628 39380
rect 31576 39296 31628 39302
rect 31576 39238 31628 39244
rect 31588 39098 31616 39238
rect 31484 39092 31536 39098
rect 31484 39034 31536 39040
rect 31576 39092 31628 39098
rect 31576 39034 31628 39040
rect 31576 38956 31628 38962
rect 31576 38898 31628 38904
rect 31484 38548 31536 38554
rect 31484 38490 31536 38496
rect 31496 37670 31524 38490
rect 31484 37664 31536 37670
rect 31484 37606 31536 37612
rect 31588 37448 31616 38898
rect 31680 37874 31708 39918
rect 32310 39879 32366 39888
rect 32036 39840 32088 39846
rect 32036 39782 32088 39788
rect 32048 39642 32076 39782
rect 31852 39636 31904 39642
rect 31852 39578 31904 39584
rect 32036 39636 32088 39642
rect 32036 39578 32088 39584
rect 31760 38956 31812 38962
rect 31760 38898 31812 38904
rect 31772 38865 31800 38898
rect 31758 38856 31814 38865
rect 31758 38791 31814 38800
rect 31864 38758 31892 39578
rect 31944 39296 31996 39302
rect 31944 39238 31996 39244
rect 31956 39030 31984 39238
rect 31944 39024 31996 39030
rect 31944 38966 31996 38972
rect 32128 38956 32180 38962
rect 32128 38898 32180 38904
rect 31852 38752 31904 38758
rect 31852 38694 31904 38700
rect 31668 37868 31720 37874
rect 31668 37810 31720 37816
rect 31588 37420 31708 37448
rect 31574 37224 31630 37233
rect 31574 37159 31576 37168
rect 31628 37159 31630 37168
rect 31576 37130 31628 37136
rect 31484 37120 31536 37126
rect 31484 37062 31536 37068
rect 31496 36922 31524 37062
rect 31484 36916 31536 36922
rect 31484 36858 31536 36864
rect 31680 36854 31708 37420
rect 31576 36848 31628 36854
rect 31404 36774 31524 36802
rect 31576 36790 31628 36796
rect 31668 36848 31720 36854
rect 31668 36790 31720 36796
rect 31392 36644 31444 36650
rect 31392 36586 31444 36592
rect 31404 36242 31432 36586
rect 31496 36582 31524 36774
rect 31484 36576 31536 36582
rect 31484 36518 31536 36524
rect 31300 36236 31352 36242
rect 31300 36178 31352 36184
rect 31392 36236 31444 36242
rect 31392 36178 31444 36184
rect 31208 35828 31260 35834
rect 31208 35770 31260 35776
rect 31114 35728 31170 35737
rect 31114 35663 31116 35672
rect 31168 35663 31170 35672
rect 31116 35634 31168 35640
rect 31128 35290 31156 35634
rect 31484 35556 31536 35562
rect 31484 35498 31536 35504
rect 31116 35284 31168 35290
rect 31116 35226 31168 35232
rect 31298 35184 31354 35193
rect 31298 35119 31354 35128
rect 31392 35148 31444 35154
rect 31312 35086 31340 35119
rect 31392 35090 31444 35096
rect 31116 35080 31168 35086
rect 31114 35048 31116 35057
rect 31300 35080 31352 35086
rect 31168 35048 31170 35057
rect 31300 35022 31352 35028
rect 31114 34983 31170 34992
rect 31300 34740 31352 34746
rect 31404 34728 31432 35090
rect 31352 34700 31432 34728
rect 31300 34682 31352 34688
rect 31208 34468 31260 34474
rect 31208 34410 31260 34416
rect 31220 33114 31248 34410
rect 31496 33522 31524 35498
rect 31588 35222 31616 36790
rect 31680 36258 31708 36790
rect 31680 36230 31800 36258
rect 31666 36000 31722 36009
rect 31666 35935 31722 35944
rect 31576 35216 31628 35222
rect 31576 35158 31628 35164
rect 31576 35012 31628 35018
rect 31576 34954 31628 34960
rect 31588 34202 31616 34954
rect 31576 34196 31628 34202
rect 31576 34138 31628 34144
rect 31484 33516 31536 33522
rect 31404 33476 31484 33504
rect 31208 33108 31260 33114
rect 31208 33050 31260 33056
rect 31404 32910 31432 33476
rect 31484 33458 31536 33464
rect 31576 33448 31628 33454
rect 31576 33390 31628 33396
rect 31392 32904 31444 32910
rect 31392 32846 31444 32852
rect 31208 32564 31260 32570
rect 31208 32506 31260 32512
rect 31116 32360 31168 32366
rect 31116 32302 31168 32308
rect 31128 31958 31156 32302
rect 31116 31952 31168 31958
rect 31116 31894 31168 31900
rect 31220 31482 31248 32506
rect 31588 32434 31616 33390
rect 31576 32428 31628 32434
rect 31576 32370 31628 32376
rect 31300 32020 31352 32026
rect 31300 31962 31352 31968
rect 31024 31476 31076 31482
rect 31024 31418 31076 31424
rect 31208 31476 31260 31482
rect 31208 31418 31260 31424
rect 31312 31414 31340 31962
rect 31300 31408 31352 31414
rect 31300 31350 31352 31356
rect 30840 31340 30892 31346
rect 30840 31282 30892 31288
rect 31208 31340 31260 31346
rect 31208 31282 31260 31288
rect 30748 30252 30800 30258
rect 30748 30194 30800 30200
rect 30564 29776 30616 29782
rect 30564 29718 30616 29724
rect 30576 29481 30604 29718
rect 30760 29578 30788 30194
rect 30748 29572 30800 29578
rect 30748 29514 30800 29520
rect 30656 29504 30708 29510
rect 30562 29472 30618 29481
rect 30656 29446 30708 29452
rect 30562 29407 30618 29416
rect 30564 27328 30616 27334
rect 30564 27270 30616 27276
rect 30576 26994 30604 27270
rect 30564 26988 30616 26994
rect 30564 26930 30616 26936
rect 30472 26444 30524 26450
rect 30472 26386 30524 26392
rect 30378 25936 30434 25945
rect 30378 25871 30380 25880
rect 30432 25871 30434 25880
rect 30564 25900 30616 25906
rect 30380 25842 30432 25848
rect 30564 25842 30616 25848
rect 30392 25294 30420 25842
rect 30576 25362 30604 25842
rect 30668 25498 30696 29446
rect 30760 29034 30788 29514
rect 30748 29028 30800 29034
rect 30748 28970 30800 28976
rect 30852 28150 30880 31282
rect 31220 30734 31248 31282
rect 31208 30728 31260 30734
rect 31208 30670 31260 30676
rect 31576 30592 31628 30598
rect 31576 30534 31628 30540
rect 31588 30258 31616 30534
rect 31576 30252 31628 30258
rect 31576 30194 31628 30200
rect 31300 30184 31352 30190
rect 31300 30126 31352 30132
rect 31312 29646 31340 30126
rect 31300 29640 31352 29646
rect 30930 29608 30986 29617
rect 31300 29582 31352 29588
rect 31484 29640 31536 29646
rect 31484 29582 31536 29588
rect 30930 29543 30932 29552
rect 30984 29543 30986 29552
rect 30932 29514 30984 29520
rect 31300 29164 31352 29170
rect 31496 29152 31524 29582
rect 31588 29578 31616 30194
rect 31576 29572 31628 29578
rect 31576 29514 31628 29520
rect 31352 29124 31524 29152
rect 31300 29106 31352 29112
rect 31576 28960 31628 28966
rect 31576 28902 31628 28908
rect 31022 28792 31078 28801
rect 31022 28727 31078 28736
rect 31036 28150 31064 28727
rect 31588 28529 31616 28902
rect 31574 28520 31630 28529
rect 31574 28455 31630 28464
rect 30840 28144 30892 28150
rect 30840 28086 30892 28092
rect 31024 28144 31076 28150
rect 31024 28086 31076 28092
rect 30852 27946 30880 28086
rect 30840 27940 30892 27946
rect 30840 27882 30892 27888
rect 30852 27674 30880 27882
rect 30840 27668 30892 27674
rect 30840 27610 30892 27616
rect 31036 26858 31064 28086
rect 31116 28076 31168 28082
rect 31116 28018 31168 28024
rect 31128 27674 31156 28018
rect 31116 27668 31168 27674
rect 31116 27610 31168 27616
rect 31300 27328 31352 27334
rect 31300 27270 31352 27276
rect 31312 26994 31340 27270
rect 31300 26988 31352 26994
rect 31300 26930 31352 26936
rect 31024 26852 31076 26858
rect 31024 26794 31076 26800
rect 31680 26042 31708 35935
rect 31772 34921 31800 36230
rect 31864 35086 31892 38694
rect 32140 38554 32168 38898
rect 32220 38888 32272 38894
rect 32220 38830 32272 38836
rect 32128 38548 32180 38554
rect 32128 38490 32180 38496
rect 32232 38026 32260 38830
rect 32048 37998 32260 38026
rect 31944 37800 31996 37806
rect 31944 37742 31996 37748
rect 31956 36582 31984 37742
rect 32048 36854 32076 37998
rect 32220 37868 32272 37874
rect 32220 37810 32272 37816
rect 32128 37188 32180 37194
rect 32128 37130 32180 37136
rect 32036 36848 32088 36854
rect 32036 36790 32088 36796
rect 31944 36576 31996 36582
rect 31944 36518 31996 36524
rect 32140 36378 32168 37130
rect 32232 36922 32260 37810
rect 32324 37262 32352 39879
rect 32588 39364 32640 39370
rect 32588 39306 32640 39312
rect 32496 39296 32548 39302
rect 32496 39238 32548 39244
rect 32508 39098 32536 39238
rect 32600 39098 32628 39306
rect 32680 39296 32732 39302
rect 32680 39238 32732 39244
rect 32496 39092 32548 39098
rect 32496 39034 32548 39040
rect 32588 39092 32640 39098
rect 32588 39034 32640 39040
rect 32402 38992 32458 39001
rect 32402 38927 32404 38936
rect 32456 38927 32458 38936
rect 32404 38898 32456 38904
rect 32692 38758 32720 39238
rect 32784 38962 32812 40394
rect 32772 38956 32824 38962
rect 32772 38898 32824 38904
rect 32680 38752 32732 38758
rect 32680 38694 32732 38700
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32404 37256 32456 37262
rect 32404 37198 32456 37204
rect 32416 36922 32444 37198
rect 32968 37176 32996 42298
rect 34532 42294 34560 42350
rect 38292 42356 38344 42362
rect 38292 42298 38344 42304
rect 41880 42356 41932 42362
rect 41880 42298 41932 42304
rect 34520 42288 34572 42294
rect 34520 42230 34572 42236
rect 38200 42220 38252 42226
rect 38200 42162 38252 42168
rect 33324 42016 33376 42022
rect 33324 41958 33376 41964
rect 33336 41682 33364 41958
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 33324 41676 33376 41682
rect 33324 41618 33376 41624
rect 34428 41540 34480 41546
rect 34428 41482 34480 41488
rect 33876 41472 33928 41478
rect 33876 41414 33928 41420
rect 33888 41386 34008 41414
rect 33600 40588 33652 40594
rect 33600 40530 33652 40536
rect 33048 40452 33100 40458
rect 33048 40394 33100 40400
rect 33060 40186 33088 40394
rect 33048 40180 33100 40186
rect 33048 40122 33100 40128
rect 33508 39432 33560 39438
rect 33508 39374 33560 39380
rect 33520 39098 33548 39374
rect 33508 39092 33560 39098
rect 33508 39034 33560 39040
rect 33612 38962 33640 40530
rect 33692 39296 33744 39302
rect 33692 39238 33744 39244
rect 33600 38956 33652 38962
rect 33600 38898 33652 38904
rect 33612 38010 33640 38898
rect 33600 38004 33652 38010
rect 33600 37946 33652 37952
rect 33140 37664 33192 37670
rect 33140 37606 33192 37612
rect 33152 37262 33180 37606
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 32968 37148 33088 37176
rect 32588 37120 32640 37126
rect 32588 37062 32640 37068
rect 32600 36922 32628 37062
rect 32220 36916 32272 36922
rect 32220 36858 32272 36864
rect 32404 36916 32456 36922
rect 32404 36858 32456 36864
rect 32588 36916 32640 36922
rect 32588 36858 32640 36864
rect 32586 36544 32642 36553
rect 32586 36479 32642 36488
rect 32128 36372 32180 36378
rect 32128 36314 32180 36320
rect 31944 36304 31996 36310
rect 31944 36246 31996 36252
rect 31852 35080 31904 35086
rect 31852 35022 31904 35028
rect 31758 34912 31814 34921
rect 31758 34847 31814 34856
rect 31852 34672 31904 34678
rect 31852 34614 31904 34620
rect 31758 34504 31814 34513
rect 31864 34490 31892 34614
rect 31814 34462 31892 34490
rect 31956 34490 31984 36246
rect 32496 36032 32548 36038
rect 32496 35974 32548 35980
rect 32508 35698 32536 35974
rect 32496 35692 32548 35698
rect 32496 35634 32548 35640
rect 32220 35488 32272 35494
rect 32220 35430 32272 35436
rect 32312 35488 32364 35494
rect 32312 35430 32364 35436
rect 32036 35080 32088 35086
rect 32034 35048 32036 35057
rect 32088 35048 32090 35057
rect 32034 34983 32090 34992
rect 32036 34944 32088 34950
rect 32036 34886 32088 34892
rect 32048 34610 32076 34886
rect 32232 34678 32260 35430
rect 32324 35290 32352 35430
rect 32312 35284 32364 35290
rect 32312 35226 32364 35232
rect 32404 34944 32456 34950
rect 32404 34886 32456 34892
rect 32220 34672 32272 34678
rect 32220 34614 32272 34620
rect 32036 34604 32088 34610
rect 32036 34546 32088 34552
rect 32312 34604 32364 34610
rect 32312 34546 32364 34552
rect 31956 34462 32168 34490
rect 31758 34439 31814 34448
rect 31852 33924 31904 33930
rect 31852 33866 31904 33872
rect 31864 33590 31892 33866
rect 31852 33584 31904 33590
rect 31852 33526 31904 33532
rect 31852 32904 31904 32910
rect 31852 32846 31904 32852
rect 31760 29504 31812 29510
rect 31760 29446 31812 29452
rect 31772 29170 31800 29446
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31772 29073 31800 29106
rect 31758 29064 31814 29073
rect 31758 28999 31814 29008
rect 31760 28416 31812 28422
rect 31760 28358 31812 28364
rect 31772 27878 31800 28358
rect 31760 27872 31812 27878
rect 31760 27814 31812 27820
rect 31760 27532 31812 27538
rect 31760 27474 31812 27480
rect 31772 26518 31800 27474
rect 31760 26512 31812 26518
rect 31760 26454 31812 26460
rect 31668 26036 31720 26042
rect 31668 25978 31720 25984
rect 30930 25936 30986 25945
rect 30930 25871 30932 25880
rect 30984 25871 30986 25880
rect 30932 25842 30984 25848
rect 31760 25832 31812 25838
rect 31760 25774 31812 25780
rect 30656 25492 30708 25498
rect 30656 25434 30708 25440
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 31116 25288 31168 25294
rect 31116 25230 31168 25236
rect 30392 24818 30420 25230
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 31128 24750 31156 25230
rect 31668 25220 31720 25226
rect 31772 25208 31800 25774
rect 31720 25180 31800 25208
rect 31668 25162 31720 25168
rect 30748 24744 30800 24750
rect 31116 24744 31168 24750
rect 30748 24686 30800 24692
rect 30930 24712 30986 24721
rect 30562 24304 30618 24313
rect 30288 24268 30340 24274
rect 30562 24239 30618 24248
rect 30288 24210 30340 24216
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30472 23180 30524 23186
rect 30472 23122 30524 23128
rect 30286 22944 30342 22953
rect 30392 22930 30420 23122
rect 30342 22902 30420 22930
rect 30286 22879 30342 22888
rect 30392 22710 30420 22902
rect 30484 22778 30512 23122
rect 30576 22982 30604 24239
rect 30760 24206 30788 24686
rect 31116 24686 31168 24692
rect 30930 24647 30986 24656
rect 30944 24342 30972 24647
rect 31484 24608 31536 24614
rect 31484 24550 31536 24556
rect 30932 24336 30984 24342
rect 30932 24278 30984 24284
rect 31496 24206 31524 24550
rect 30748 24200 30800 24206
rect 30748 24142 30800 24148
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 30944 23866 30972 24142
rect 31576 24132 31628 24138
rect 31576 24074 31628 24080
rect 30932 23860 30984 23866
rect 30932 23802 30984 23808
rect 30656 23656 30708 23662
rect 30656 23598 30708 23604
rect 30668 23254 30696 23598
rect 31588 23254 31616 24074
rect 30656 23248 30708 23254
rect 30656 23190 30708 23196
rect 31576 23248 31628 23254
rect 31576 23190 31628 23196
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30380 22704 30432 22710
rect 30380 22646 30432 22652
rect 31116 22704 31168 22710
rect 31116 22646 31168 22652
rect 30116 22066 30236 22094
rect 30012 21956 30064 21962
rect 30012 21898 30064 21904
rect 30024 21690 30052 21898
rect 30012 21684 30064 21690
rect 30012 21626 30064 21632
rect 29564 20556 29684 20584
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 29564 19310 29592 20556
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29552 19304 29604 19310
rect 29552 19246 29604 19252
rect 29288 18834 29316 19246
rect 29564 18970 29592 19246
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29276 18828 29328 18834
rect 29196 18788 29276 18816
rect 29092 18216 29144 18222
rect 29092 18158 29144 18164
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 29196 16946 29224 18788
rect 29276 18770 29328 18776
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29564 18426 29592 18566
rect 29552 18420 29604 18426
rect 29552 18362 29604 18368
rect 29656 17542 29684 18566
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 29644 17536 29696 17542
rect 29644 17478 29696 17484
rect 29644 17332 29696 17338
rect 29644 17274 29696 17280
rect 29104 16918 29224 16946
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29104 16640 29132 16918
rect 29472 16794 29500 16934
rect 29460 16788 29512 16794
rect 29460 16730 29512 16736
rect 29368 16720 29420 16726
rect 29368 16662 29420 16668
rect 29104 16612 29316 16640
rect 29000 16448 29052 16454
rect 29000 16390 29052 16396
rect 29012 16114 29040 16390
rect 29092 16176 29144 16182
rect 29090 16144 29092 16153
rect 29184 16176 29236 16182
rect 29144 16144 29146 16153
rect 29000 16108 29052 16114
rect 29184 16118 29236 16124
rect 29090 16079 29146 16088
rect 29000 16050 29052 16056
rect 29196 15570 29224 16118
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 29288 14482 29316 16612
rect 29380 16289 29408 16662
rect 29472 16454 29500 16730
rect 29552 16720 29604 16726
rect 29552 16662 29604 16668
rect 29460 16448 29512 16454
rect 29460 16390 29512 16396
rect 29366 16280 29422 16289
rect 29366 16215 29422 16224
rect 29472 15745 29500 16390
rect 29458 15736 29514 15745
rect 29458 15671 29514 15680
rect 29472 15502 29500 15671
rect 29564 15586 29592 16662
rect 29656 16658 29684 17274
rect 29736 17196 29788 17202
rect 29736 17138 29788 17144
rect 29644 16652 29696 16658
rect 29644 16594 29696 16600
rect 29748 16562 29776 17138
rect 29920 16992 29972 16998
rect 29920 16934 29972 16940
rect 29656 16534 29776 16562
rect 29656 16454 29684 16534
rect 29644 16448 29696 16454
rect 29644 16390 29696 16396
rect 29656 16153 29684 16390
rect 29826 16280 29882 16289
rect 29826 16215 29882 16224
rect 29840 16182 29868 16215
rect 29828 16176 29880 16182
rect 29642 16144 29698 16153
rect 29828 16118 29880 16124
rect 29932 16114 29960 16934
rect 29736 16108 29788 16114
rect 29698 16088 29736 16096
rect 29642 16079 29736 16088
rect 29656 16068 29736 16079
rect 29736 16050 29788 16056
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 29644 15972 29696 15978
rect 29644 15914 29696 15920
rect 29656 15706 29684 15914
rect 29644 15700 29696 15706
rect 29644 15642 29696 15648
rect 29564 15558 29684 15586
rect 29460 15496 29512 15502
rect 29460 15438 29512 15444
rect 29552 14816 29604 14822
rect 29552 14758 29604 14764
rect 29656 14770 29684 15558
rect 30024 15162 30052 18022
rect 30116 17202 30144 22066
rect 30562 21856 30618 21865
rect 30562 21791 30618 21800
rect 30576 21622 30604 21791
rect 30564 21616 30616 21622
rect 30564 21558 30616 21564
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 30288 21004 30340 21010
rect 30288 20946 30340 20952
rect 30300 20534 30328 20946
rect 30288 20528 30340 20534
rect 30288 20470 30340 20476
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 30288 19304 30340 19310
rect 30288 19246 30340 19252
rect 30208 18426 30236 19246
rect 30300 19174 30328 19246
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30288 18828 30340 18834
rect 30288 18770 30340 18776
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 30300 18086 30328 18770
rect 30392 18766 30420 19110
rect 30380 18760 30432 18766
rect 30380 18702 30432 18708
rect 30656 18624 30708 18630
rect 30656 18566 30708 18572
rect 30668 18290 30696 18566
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30668 17338 30696 18226
rect 30748 17740 30800 17746
rect 30748 17682 30800 17688
rect 30760 17338 30788 17682
rect 30656 17332 30708 17338
rect 30656 17274 30708 17280
rect 30748 17332 30800 17338
rect 30748 17274 30800 17280
rect 30104 17196 30156 17202
rect 30104 17138 30156 17144
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30116 17082 30144 17138
rect 30116 17054 30236 17082
rect 30208 16658 30236 17054
rect 30104 16652 30156 16658
rect 30104 16594 30156 16600
rect 30196 16652 30248 16658
rect 30196 16594 30248 16600
rect 30116 16522 30144 16594
rect 30104 16516 30156 16522
rect 30104 16458 30156 16464
rect 30668 16182 30696 17138
rect 30656 16176 30708 16182
rect 30656 16118 30708 16124
rect 30104 15564 30156 15570
rect 30104 15506 30156 15512
rect 30116 15162 30144 15506
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 29734 14784 29790 14793
rect 29564 14618 29592 14758
rect 29656 14742 29734 14770
rect 29734 14719 29790 14728
rect 29552 14612 29604 14618
rect 29552 14554 29604 14560
rect 29276 14476 29328 14482
rect 29276 14418 29328 14424
rect 28998 13696 29054 13705
rect 28998 13631 29054 13640
rect 29012 13258 29040 13631
rect 29000 13252 29052 13258
rect 29000 13194 29052 13200
rect 29012 12918 29040 13194
rect 29288 12918 29316 14418
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 29276 12912 29328 12918
rect 29276 12854 29328 12860
rect 28908 12436 28960 12442
rect 28908 12378 28960 12384
rect 28920 12345 28948 12378
rect 28906 12336 28962 12345
rect 28906 12271 28962 12280
rect 29288 11898 29316 12854
rect 29748 12434 29776 14719
rect 30024 14113 30052 15098
rect 30852 14414 30880 20198
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 30944 16590 30972 17138
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30944 16046 30972 16526
rect 31036 16522 31064 21286
rect 31128 17649 31156 22646
rect 31588 21690 31616 23190
rect 31680 23118 31708 25162
rect 31864 24682 31892 32846
rect 31944 31272 31996 31278
rect 31944 31214 31996 31220
rect 31956 28218 31984 31214
rect 31944 28212 31996 28218
rect 31944 28154 31996 28160
rect 31956 28098 31984 28154
rect 31956 28070 32076 28098
rect 32048 28014 32076 28070
rect 31944 28008 31996 28014
rect 31942 27976 31944 27985
rect 32036 28008 32088 28014
rect 31996 27976 31998 27985
rect 32036 27950 32088 27956
rect 31942 27911 31998 27920
rect 32140 26586 32168 34462
rect 32324 33998 32352 34546
rect 32312 33992 32364 33998
rect 32312 33934 32364 33940
rect 32220 30184 32272 30190
rect 32220 30126 32272 30132
rect 32232 29714 32260 30126
rect 32220 29708 32272 29714
rect 32220 29650 32272 29656
rect 32232 29306 32260 29650
rect 32220 29300 32272 29306
rect 32220 29242 32272 29248
rect 32324 28994 32352 33934
rect 32416 32910 32444 34886
rect 32404 32904 32456 32910
rect 32404 32846 32456 32852
rect 32416 32570 32444 32846
rect 32404 32564 32456 32570
rect 32404 32506 32456 32512
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32416 30326 32444 31282
rect 32404 30320 32456 30326
rect 32404 30262 32456 30268
rect 32600 29730 32628 36479
rect 32864 32836 32916 32842
rect 32864 32778 32916 32784
rect 32956 32836 33008 32842
rect 32956 32778 33008 32784
rect 32876 32570 32904 32778
rect 32864 32564 32916 32570
rect 32864 32506 32916 32512
rect 32680 32428 32732 32434
rect 32680 32370 32732 32376
rect 32692 32026 32720 32370
rect 32864 32360 32916 32366
rect 32864 32302 32916 32308
rect 32680 32020 32732 32026
rect 32680 31962 32732 31968
rect 32772 31340 32824 31346
rect 32772 31282 32824 31288
rect 32680 30796 32732 30802
rect 32680 30738 32732 30744
rect 32692 30258 32720 30738
rect 32784 30666 32812 31282
rect 32772 30660 32824 30666
rect 32772 30602 32824 30608
rect 32680 30252 32732 30258
rect 32680 30194 32732 30200
rect 32508 29702 32628 29730
rect 32324 28966 32444 28994
rect 32416 28082 32444 28966
rect 32404 28076 32456 28082
rect 32404 28018 32456 28024
rect 32416 27538 32444 28018
rect 32404 27532 32456 27538
rect 32404 27474 32456 27480
rect 32128 26580 32180 26586
rect 32128 26522 32180 26528
rect 32508 26518 32536 29702
rect 32692 29646 32720 30194
rect 32680 29640 32732 29646
rect 32680 29582 32732 29588
rect 32586 29336 32642 29345
rect 32692 29306 32720 29582
rect 32586 29271 32642 29280
rect 32680 29300 32732 29306
rect 32600 28948 32628 29271
rect 32680 29242 32732 29248
rect 32784 29170 32812 30602
rect 32772 29164 32824 29170
rect 32772 29106 32824 29112
rect 32772 28960 32824 28966
rect 32600 28920 32772 28948
rect 32772 28902 32824 28908
rect 32680 28212 32732 28218
rect 32680 28154 32732 28160
rect 32692 27674 32720 28154
rect 32784 28082 32812 28902
rect 32876 28218 32904 32302
rect 32968 31278 32996 32778
rect 32956 31272 33008 31278
rect 32956 31214 33008 31220
rect 32956 30252 33008 30258
rect 32956 30194 33008 30200
rect 32968 29510 32996 30194
rect 32956 29504 33008 29510
rect 32956 29446 33008 29452
rect 32864 28212 32916 28218
rect 32864 28154 32916 28160
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 32680 27668 32732 27674
rect 32680 27610 32732 27616
rect 32876 27062 32904 28154
rect 32864 27056 32916 27062
rect 32864 26998 32916 27004
rect 32588 26784 32640 26790
rect 32588 26726 32640 26732
rect 32496 26512 32548 26518
rect 32496 26454 32548 26460
rect 32220 26376 32272 26382
rect 32220 26318 32272 26324
rect 31944 26308 31996 26314
rect 31944 26250 31996 26256
rect 31956 26042 31984 26250
rect 31944 26036 31996 26042
rect 31944 25978 31996 25984
rect 31944 25832 31996 25838
rect 31944 25774 31996 25780
rect 31956 25362 31984 25774
rect 32232 25498 32260 26318
rect 32404 26308 32456 26314
rect 32404 26250 32456 26256
rect 32416 25770 32444 26250
rect 32508 26042 32536 26454
rect 32496 26036 32548 26042
rect 32496 25978 32548 25984
rect 32404 25764 32456 25770
rect 32404 25706 32456 25712
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 31944 25356 31996 25362
rect 31944 25298 31996 25304
rect 32220 25356 32272 25362
rect 32220 25298 32272 25304
rect 31852 24676 31904 24682
rect 31852 24618 31904 24624
rect 31758 24304 31814 24313
rect 31814 24262 31892 24290
rect 31758 24239 31814 24248
rect 31760 24064 31812 24070
rect 31760 24006 31812 24012
rect 31772 23730 31800 24006
rect 31760 23724 31812 23730
rect 31760 23666 31812 23672
rect 31864 23594 31892 24262
rect 31852 23588 31904 23594
rect 31852 23530 31904 23536
rect 31956 23118 31984 25298
rect 31668 23112 31720 23118
rect 31668 23054 31720 23060
rect 31944 23112 31996 23118
rect 31944 23054 31996 23060
rect 32232 21690 32260 25298
rect 32416 24614 32444 25706
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32324 23118 32352 24142
rect 32416 23526 32444 24550
rect 32404 23520 32456 23526
rect 32404 23462 32456 23468
rect 32416 23118 32444 23462
rect 32312 23112 32364 23118
rect 32312 23054 32364 23060
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32324 22506 32352 23054
rect 32312 22500 32364 22506
rect 32312 22442 32364 22448
rect 32600 22094 32628 26726
rect 32680 26240 32732 26246
rect 32680 26182 32732 26188
rect 32692 25226 32720 26182
rect 32680 25220 32732 25226
rect 32680 25162 32732 25168
rect 33060 23866 33088 37148
rect 33416 37120 33468 37126
rect 33416 37062 33468 37068
rect 33428 36922 33456 37062
rect 33416 36916 33468 36922
rect 33416 36858 33468 36864
rect 33612 36786 33640 37946
rect 33704 37942 33732 39238
rect 33692 37936 33744 37942
rect 33692 37878 33744 37884
rect 33600 36780 33652 36786
rect 33600 36722 33652 36728
rect 33232 36576 33284 36582
rect 33232 36518 33284 36524
rect 33244 35766 33272 36518
rect 33612 36242 33640 36722
rect 33600 36236 33652 36242
rect 33600 36178 33652 36184
rect 33612 35834 33640 36178
rect 33600 35828 33652 35834
rect 33600 35770 33652 35776
rect 33232 35760 33284 35766
rect 33232 35702 33284 35708
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 33336 35154 33364 35634
rect 33324 35148 33376 35154
rect 33324 35090 33376 35096
rect 33416 33584 33468 33590
rect 33416 33526 33468 33532
rect 33232 30592 33284 30598
rect 33232 30534 33284 30540
rect 33244 30258 33272 30534
rect 33232 30252 33284 30258
rect 33232 30194 33284 30200
rect 33244 29646 33272 30194
rect 33232 29640 33284 29646
rect 33232 29582 33284 29588
rect 33428 28422 33456 33526
rect 33784 32836 33836 32842
rect 33784 32778 33836 32784
rect 33796 32434 33824 32778
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 33508 32224 33560 32230
rect 33508 32166 33560 32172
rect 33520 31822 33548 32166
rect 33796 32026 33824 32370
rect 33784 32020 33836 32026
rect 33784 31962 33836 31968
rect 33600 31884 33652 31890
rect 33600 31826 33652 31832
rect 33508 31816 33560 31822
rect 33508 31758 33560 31764
rect 33520 31278 33548 31758
rect 33612 31414 33640 31826
rect 33600 31408 33652 31414
rect 33600 31350 33652 31356
rect 33508 31272 33560 31278
rect 33508 31214 33560 31220
rect 33520 30734 33548 31214
rect 33508 30728 33560 30734
rect 33508 30670 33560 30676
rect 33520 30258 33548 30670
rect 33612 30258 33640 31350
rect 33796 31142 33824 31962
rect 33784 31136 33836 31142
rect 33784 31078 33836 31084
rect 33796 30258 33824 31078
rect 33876 30660 33928 30666
rect 33876 30602 33928 30608
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33600 30252 33652 30258
rect 33600 30194 33652 30200
rect 33784 30252 33836 30258
rect 33784 30194 33836 30200
rect 33612 29646 33640 30194
rect 33796 29646 33824 30194
rect 33600 29640 33652 29646
rect 33600 29582 33652 29588
rect 33784 29640 33836 29646
rect 33784 29582 33836 29588
rect 33416 28416 33468 28422
rect 33416 28358 33468 28364
rect 33428 28218 33456 28358
rect 33416 28212 33468 28218
rect 33416 28154 33468 28160
rect 33888 28082 33916 30602
rect 33980 28082 34008 41386
rect 34440 41070 34468 41482
rect 38212 41414 38240 42162
rect 40868 42016 40920 42022
rect 40868 41958 40920 41964
rect 38028 41386 38240 41414
rect 34612 41132 34664 41138
rect 34612 41074 34664 41080
rect 34428 41064 34480 41070
rect 34428 41006 34480 41012
rect 34440 40458 34468 41006
rect 34428 40452 34480 40458
rect 34428 40394 34480 40400
rect 34440 38010 34468 40394
rect 34520 40384 34572 40390
rect 34520 40326 34572 40332
rect 34428 38004 34480 38010
rect 34428 37946 34480 37952
rect 34532 35154 34560 40326
rect 34624 39030 34652 41074
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 37648 40520 37700 40526
rect 37648 40462 37700 40468
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 37660 39506 37688 40462
rect 37648 39500 37700 39506
rect 37648 39442 37700 39448
rect 34612 39024 34664 39030
rect 34612 38966 34664 38972
rect 34624 36854 34652 38966
rect 35348 38752 35400 38758
rect 35348 38694 35400 38700
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34796 37664 34848 37670
rect 34796 37606 34848 37612
rect 34612 36848 34664 36854
rect 34612 36790 34664 36796
rect 34624 35766 34652 36790
rect 34612 35760 34664 35766
rect 34612 35702 34664 35708
rect 34520 35148 34572 35154
rect 34348 35108 34520 35136
rect 34348 34202 34376 35108
rect 34520 35090 34572 35096
rect 34624 35086 34652 35702
rect 34808 35086 34836 37606
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34888 35148 34940 35154
rect 34888 35090 34940 35096
rect 34612 35080 34664 35086
rect 34612 35022 34664 35028
rect 34796 35080 34848 35086
rect 34796 35022 34848 35028
rect 34612 34944 34664 34950
rect 34612 34886 34664 34892
rect 34624 34610 34652 34886
rect 34808 34610 34836 35022
rect 34900 34610 34928 35090
rect 34520 34604 34572 34610
rect 34520 34546 34572 34552
rect 34612 34604 34664 34610
rect 34612 34546 34664 34552
rect 34704 34604 34756 34610
rect 34704 34546 34756 34552
rect 34796 34604 34848 34610
rect 34796 34546 34848 34552
rect 34888 34604 34940 34610
rect 34888 34546 34940 34552
rect 34428 34400 34480 34406
rect 34428 34342 34480 34348
rect 34244 34196 34296 34202
rect 34244 34138 34296 34144
rect 34336 34196 34388 34202
rect 34336 34138 34388 34144
rect 34256 33522 34284 34138
rect 34440 33946 34468 34342
rect 34532 34134 34560 34546
rect 34612 34468 34664 34474
rect 34612 34410 34664 34416
rect 34520 34128 34572 34134
rect 34520 34070 34572 34076
rect 34624 33998 34652 34410
rect 34716 34406 34744 34546
rect 34704 34400 34756 34406
rect 34704 34342 34756 34348
rect 34808 33998 34836 34546
rect 35360 34406 35388 38694
rect 37556 37256 37608 37262
rect 37556 37198 37608 37204
rect 35532 36576 35584 36582
rect 35532 36518 35584 36524
rect 35544 34610 35572 36518
rect 37280 36100 37332 36106
rect 37280 36042 37332 36048
rect 35532 34604 35584 34610
rect 35532 34546 35584 34552
rect 35348 34400 35400 34406
rect 35348 34342 35400 34348
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 34202 35388 34342
rect 35348 34196 35400 34202
rect 35348 34138 35400 34144
rect 34612 33992 34664 33998
rect 34440 33918 34560 33946
rect 34612 33934 34664 33940
rect 34704 33992 34756 33998
rect 34704 33934 34756 33940
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 34244 33516 34296 33522
rect 34244 33458 34296 33464
rect 34532 32978 34560 33918
rect 34612 33516 34664 33522
rect 34612 33458 34664 33464
rect 34624 33114 34652 33458
rect 34612 33108 34664 33114
rect 34612 33050 34664 33056
rect 34060 32972 34112 32978
rect 34060 32914 34112 32920
rect 34520 32972 34572 32978
rect 34520 32914 34572 32920
rect 34072 31754 34100 32914
rect 34336 32904 34388 32910
rect 34336 32846 34388 32852
rect 34348 32570 34376 32846
rect 34716 32842 34744 33934
rect 35360 33590 35388 34138
rect 35544 34066 35572 34546
rect 35532 34060 35584 34066
rect 35532 34002 35584 34008
rect 35348 33584 35400 33590
rect 35348 33526 35400 33532
rect 35544 33522 35572 34002
rect 35532 33516 35584 33522
rect 35532 33458 35584 33464
rect 34796 33312 34848 33318
rect 34796 33254 34848 33260
rect 35624 33312 35676 33318
rect 35624 33254 35676 33260
rect 34808 32978 34836 33254
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35636 33114 35664 33254
rect 35624 33108 35676 33114
rect 35624 33050 35676 33056
rect 34796 32972 34848 32978
rect 34796 32914 34848 32920
rect 34704 32836 34756 32842
rect 34704 32778 34756 32784
rect 34336 32564 34388 32570
rect 34336 32506 34388 32512
rect 34440 32524 34744 32552
rect 34440 32434 34468 32524
rect 34428 32428 34480 32434
rect 34428 32370 34480 32376
rect 34520 32428 34572 32434
rect 34520 32370 34572 32376
rect 34440 31890 34468 32370
rect 34428 31884 34480 31890
rect 34428 31826 34480 31832
rect 34532 31822 34560 32370
rect 34716 32298 34744 32524
rect 34808 32366 34836 32914
rect 34888 32904 34940 32910
rect 34888 32846 34940 32852
rect 34900 32570 34928 32846
rect 34980 32768 35032 32774
rect 34980 32710 35032 32716
rect 34888 32564 34940 32570
rect 34888 32506 34940 32512
rect 34796 32360 34848 32366
rect 34796 32302 34848 32308
rect 34704 32292 34756 32298
rect 34704 32234 34756 32240
rect 34900 32230 34928 32506
rect 34992 32434 35020 32710
rect 34980 32428 35032 32434
rect 34980 32370 35032 32376
rect 35636 32366 35664 33050
rect 37292 32502 37320 36042
rect 37280 32496 37332 32502
rect 37280 32438 37332 32444
rect 35532 32360 35584 32366
rect 35532 32302 35584 32308
rect 35624 32360 35676 32366
rect 35624 32302 35676 32308
rect 34888 32224 34940 32230
rect 34888 32166 34940 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34520 31816 34572 31822
rect 34520 31758 34572 31764
rect 34072 31726 34284 31754
rect 34060 30796 34112 30802
rect 34060 30738 34112 30744
rect 34072 28558 34100 30738
rect 34152 30592 34204 30598
rect 34152 30534 34204 30540
rect 34164 30258 34192 30534
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 34152 29504 34204 29510
rect 34152 29446 34204 29452
rect 34164 29170 34192 29446
rect 34152 29164 34204 29170
rect 34152 29106 34204 29112
rect 34256 28694 34284 31726
rect 34532 30682 34560 31758
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35440 30728 35492 30734
rect 34532 30654 34652 30682
rect 35440 30670 35492 30676
rect 34624 30598 34652 30654
rect 34612 30592 34664 30598
rect 34612 30534 34664 30540
rect 34520 30252 34572 30258
rect 34520 30194 34572 30200
rect 34532 29646 34560 30194
rect 34624 30122 34652 30534
rect 35256 30184 35308 30190
rect 35308 30144 35388 30172
rect 35256 30126 35308 30132
rect 34612 30116 34664 30122
rect 34612 30058 34664 30064
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34532 29170 34560 29582
rect 34624 29578 34652 30058
rect 34796 30048 34848 30054
rect 34796 29990 34848 29996
rect 34808 29646 34836 29990
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29850 35388 30144
rect 35452 29850 35480 30670
rect 35544 30054 35572 32302
rect 35624 32224 35676 32230
rect 35624 32166 35676 32172
rect 35636 32026 35664 32166
rect 35624 32020 35676 32026
rect 35624 31962 35676 31968
rect 35900 30592 35952 30598
rect 35900 30534 35952 30540
rect 35912 30394 35940 30534
rect 35900 30388 35952 30394
rect 35900 30330 35952 30336
rect 35532 30048 35584 30054
rect 35532 29990 35584 29996
rect 37568 29850 37596 37198
rect 37660 32502 37688 39442
rect 37648 32496 37700 32502
rect 37648 32438 37700 32444
rect 37740 32428 37792 32434
rect 37740 32370 37792 32376
rect 37648 32360 37700 32366
rect 37648 32302 37700 32308
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 37556 29844 37608 29850
rect 37556 29786 37608 29792
rect 35808 29708 35860 29714
rect 35808 29650 35860 29656
rect 34796 29640 34848 29646
rect 34796 29582 34848 29588
rect 35716 29640 35768 29646
rect 35716 29582 35768 29588
rect 34612 29572 34664 29578
rect 34612 29514 34664 29520
rect 35728 29306 35756 29582
rect 35716 29300 35768 29306
rect 35716 29242 35768 29248
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34244 28688 34296 28694
rect 34244 28630 34296 28636
rect 34060 28552 34112 28558
rect 34060 28494 34112 28500
rect 34072 28218 34100 28494
rect 34256 28218 34284 28630
rect 34060 28212 34112 28218
rect 34060 28154 34112 28160
rect 34244 28212 34296 28218
rect 34244 28154 34296 28160
rect 34428 28144 34480 28150
rect 34428 28086 34480 28092
rect 35162 28112 35218 28121
rect 33876 28076 33928 28082
rect 33876 28018 33928 28024
rect 33968 28076 34020 28082
rect 33968 28018 34020 28024
rect 33600 28008 33652 28014
rect 33600 27950 33652 27956
rect 33508 27328 33560 27334
rect 33508 27270 33560 27276
rect 33520 27130 33548 27270
rect 33508 27124 33560 27130
rect 33508 27066 33560 27072
rect 33612 27062 33640 27950
rect 34336 27872 34388 27878
rect 34336 27814 34388 27820
rect 34348 27470 34376 27814
rect 34336 27464 34388 27470
rect 34336 27406 34388 27412
rect 33324 27056 33376 27062
rect 33324 26998 33376 27004
rect 33600 27056 33652 27062
rect 33600 26998 33652 27004
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 33152 26586 33180 26930
rect 33140 26580 33192 26586
rect 33140 26522 33192 26528
rect 33232 26512 33284 26518
rect 33232 26454 33284 26460
rect 33244 25906 33272 26454
rect 33336 26246 33364 26998
rect 33508 26988 33560 26994
rect 33508 26930 33560 26936
rect 33324 26240 33376 26246
rect 33324 26182 33376 26188
rect 33232 25900 33284 25906
rect 33232 25842 33284 25848
rect 33336 25770 33364 26182
rect 33520 25906 33548 26930
rect 34348 26926 34376 27406
rect 34336 26920 34388 26926
rect 34336 26862 34388 26868
rect 34440 26790 34468 28086
rect 35162 28047 35164 28056
rect 35216 28047 35218 28056
rect 35716 28076 35768 28082
rect 35164 28018 35216 28024
rect 35716 28018 35768 28024
rect 35440 28008 35492 28014
rect 35440 27950 35492 27956
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35452 27554 35480 27950
rect 35532 27872 35584 27878
rect 35532 27814 35584 27820
rect 35544 27674 35572 27814
rect 35532 27668 35584 27674
rect 35532 27610 35584 27616
rect 34796 27532 34848 27538
rect 35452 27526 35572 27554
rect 34796 27474 34848 27480
rect 34808 27130 34836 27474
rect 35440 27328 35492 27334
rect 35440 27270 35492 27276
rect 34796 27124 34848 27130
rect 34796 27066 34848 27072
rect 35452 27062 35480 27270
rect 35440 27056 35492 27062
rect 35440 26998 35492 27004
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34612 26376 34664 26382
rect 34612 26318 34664 26324
rect 34336 26240 34388 26246
rect 34336 26182 34388 26188
rect 33508 25900 33560 25906
rect 33508 25842 33560 25848
rect 33324 25764 33376 25770
rect 33324 25706 33376 25712
rect 33520 25158 33548 25842
rect 34060 25220 34112 25226
rect 34060 25162 34112 25168
rect 33508 25152 33560 25158
rect 33508 25094 33560 25100
rect 33048 23860 33100 23866
rect 33048 23802 33100 23808
rect 34072 23798 34100 25162
rect 34060 23792 34112 23798
rect 34060 23734 34112 23740
rect 32680 23656 32732 23662
rect 32680 23598 32732 23604
rect 32692 23322 32720 23598
rect 32680 23316 32732 23322
rect 32680 23258 32732 23264
rect 32692 23118 32720 23258
rect 34072 23118 34100 23734
rect 32680 23112 32732 23118
rect 32680 23054 32732 23060
rect 34060 23112 34112 23118
rect 34060 23054 34112 23060
rect 32324 22066 32628 22094
rect 32692 22094 32720 23054
rect 34348 22982 34376 26182
rect 34428 25832 34480 25838
rect 34428 25774 34480 25780
rect 34440 25294 34468 25774
rect 34624 25702 34652 26318
rect 34888 26036 34940 26042
rect 34888 25978 34940 25984
rect 34900 25770 34928 25978
rect 35544 25945 35572 27526
rect 35530 25936 35586 25945
rect 35530 25871 35532 25880
rect 35584 25871 35586 25880
rect 35532 25842 35584 25848
rect 34888 25764 34940 25770
rect 34888 25706 34940 25712
rect 34612 25696 34664 25702
rect 34612 25638 34664 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34428 25288 34480 25294
rect 34428 25230 34480 25236
rect 34796 25288 34848 25294
rect 34796 25230 34848 25236
rect 34808 24274 34836 25230
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 24268 34848 24274
rect 34796 24210 34848 24216
rect 34704 23860 34756 23866
rect 34704 23802 34756 23808
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 34336 22976 34388 22982
rect 34336 22918 34388 22924
rect 34532 22778 34560 23598
rect 34716 23118 34744 23802
rect 34808 23798 34836 24210
rect 34796 23792 34848 23798
rect 34796 23734 34848 23740
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35728 23186 35756 28018
rect 35820 27538 35848 29650
rect 36268 29504 36320 29510
rect 36268 29446 36320 29452
rect 35808 27532 35860 27538
rect 35808 27474 35860 27480
rect 35808 26376 35860 26382
rect 35808 26318 35860 26324
rect 35820 25770 35848 26318
rect 36084 26240 36136 26246
rect 36084 26182 36136 26188
rect 36096 26042 36124 26182
rect 36084 26036 36136 26042
rect 36084 25978 36136 25984
rect 36280 25974 36308 29446
rect 37568 29306 37596 29786
rect 37660 29578 37688 32302
rect 37648 29572 37700 29578
rect 37648 29514 37700 29520
rect 37556 29300 37608 29306
rect 37556 29242 37608 29248
rect 36542 29200 36598 29209
rect 36542 29135 36598 29144
rect 36556 29102 36584 29135
rect 36452 29096 36504 29102
rect 36452 29038 36504 29044
rect 36544 29096 36596 29102
rect 36596 29056 36768 29084
rect 36544 29038 36596 29044
rect 36268 25968 36320 25974
rect 36268 25910 36320 25916
rect 35808 25764 35860 25770
rect 35808 25706 35860 25712
rect 36084 25696 36136 25702
rect 36084 25638 36136 25644
rect 36096 25498 36124 25638
rect 36084 25492 36136 25498
rect 36084 25434 36136 25440
rect 36280 25362 36308 25910
rect 36268 25356 36320 25362
rect 36268 25298 36320 25304
rect 35808 25152 35860 25158
rect 35808 25094 35860 25100
rect 35820 24070 35848 25094
rect 35808 24064 35860 24070
rect 35808 24006 35860 24012
rect 35820 23798 35848 24006
rect 35808 23792 35860 23798
rect 35808 23734 35860 23740
rect 35716 23180 35768 23186
rect 35716 23122 35768 23128
rect 34704 23112 34756 23118
rect 34704 23054 34756 23060
rect 34704 22976 34756 22982
rect 34704 22918 34756 22924
rect 34716 22778 34744 22918
rect 34520 22772 34572 22778
rect 34520 22714 34572 22720
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 32692 22066 32812 22094
rect 31484 21684 31536 21690
rect 31484 21626 31536 21632
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 32220 21684 32272 21690
rect 32220 21626 32272 21632
rect 31496 21554 31524 21626
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31588 21486 31616 21626
rect 31576 21480 31628 21486
rect 31576 21422 31628 21428
rect 31208 21344 31260 21350
rect 31392 21344 31444 21350
rect 31208 21286 31260 21292
rect 31312 21304 31392 21332
rect 31220 20942 31248 21286
rect 31312 21010 31340 21304
rect 31392 21286 31444 21292
rect 32220 21344 32272 21350
rect 32220 21286 32272 21292
rect 31300 21004 31352 21010
rect 31300 20946 31352 20952
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31484 20936 31536 20942
rect 31484 20878 31536 20884
rect 31300 20868 31352 20874
rect 31300 20810 31352 20816
rect 31312 17762 31340 20810
rect 31390 20088 31446 20097
rect 31496 20058 31524 20878
rect 32232 20505 32260 21286
rect 32218 20496 32274 20505
rect 32128 20460 32180 20466
rect 32218 20431 32220 20440
rect 32128 20402 32180 20408
rect 32272 20431 32274 20440
rect 32220 20402 32272 20408
rect 31760 20256 31812 20262
rect 31760 20198 31812 20204
rect 31772 20058 31800 20198
rect 31390 20023 31446 20032
rect 31484 20052 31536 20058
rect 31404 19802 31432 20023
rect 31484 19994 31536 20000
rect 31760 20052 31812 20058
rect 31760 19994 31812 20000
rect 31404 19774 31524 19802
rect 31392 19712 31444 19718
rect 31392 19654 31444 19660
rect 31404 19174 31432 19654
rect 31496 19378 31524 19774
rect 31668 19508 31720 19514
rect 31668 19450 31720 19456
rect 31484 19372 31536 19378
rect 31484 19314 31536 19320
rect 31392 19168 31444 19174
rect 31392 19110 31444 19116
rect 31496 18766 31524 19314
rect 31484 18760 31536 18766
rect 31484 18702 31536 18708
rect 31484 18284 31536 18290
rect 31484 18226 31536 18232
rect 31496 17882 31524 18226
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 31312 17734 31524 17762
rect 31300 17672 31352 17678
rect 31114 17640 31170 17649
rect 31300 17614 31352 17620
rect 31114 17575 31170 17584
rect 31024 16516 31076 16522
rect 31024 16458 31076 16464
rect 30932 16040 30984 16046
rect 30932 15982 30984 15988
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 30010 14104 30066 14113
rect 30010 14039 30066 14048
rect 30838 14104 30894 14113
rect 31036 14074 31064 16458
rect 31128 15552 31156 17575
rect 31312 17066 31340 17614
rect 31300 17060 31352 17066
rect 31300 17002 31352 17008
rect 31208 16992 31260 16998
rect 31208 16934 31260 16940
rect 31220 16590 31248 16934
rect 31312 16658 31340 17002
rect 31300 16652 31352 16658
rect 31300 16594 31352 16600
rect 31208 16584 31260 16590
rect 31208 16526 31260 16532
rect 31300 16448 31352 16454
rect 31300 16390 31352 16396
rect 31128 15524 31248 15552
rect 31116 14816 31168 14822
rect 31116 14758 31168 14764
rect 31128 14346 31156 14758
rect 31116 14340 31168 14346
rect 31116 14282 31168 14288
rect 30838 14039 30894 14048
rect 31024 14068 31076 14074
rect 30196 13932 30248 13938
rect 30196 13874 30248 13880
rect 30104 13524 30156 13530
rect 30104 13466 30156 13472
rect 29564 12406 29776 12434
rect 30012 12436 30064 12442
rect 29564 12238 29592 12406
rect 30012 12378 30064 12384
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 29276 11892 29328 11898
rect 29276 11834 29328 11840
rect 29184 9920 29236 9926
rect 29184 9862 29236 9868
rect 29196 9654 29224 9862
rect 29184 9648 29236 9654
rect 29184 9590 29236 9596
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 29104 6458 29132 7278
rect 29564 6866 29592 12174
rect 30024 11898 30052 12378
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 29644 11756 29696 11762
rect 29644 11698 29696 11704
rect 29656 9654 29684 11698
rect 29736 10464 29788 10470
rect 29736 10406 29788 10412
rect 29748 10266 29776 10406
rect 29736 10260 29788 10266
rect 29736 10202 29788 10208
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 29656 8974 29684 9590
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 30116 8566 30144 13466
rect 30208 12306 30236 13874
rect 30748 12912 30800 12918
rect 30748 12854 30800 12860
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 30300 12306 30328 12378
rect 30196 12300 30248 12306
rect 30196 12242 30248 12248
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30208 11830 30236 12242
rect 30196 11824 30248 11830
rect 30196 11766 30248 11772
rect 30300 10606 30328 12242
rect 30656 12232 30708 12238
rect 30656 12174 30708 12180
rect 30668 12050 30696 12174
rect 30760 12170 30788 12854
rect 30852 12170 30880 14039
rect 31024 14010 31076 14016
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 31036 13462 31064 13874
rect 31024 13456 31076 13462
rect 31024 13398 31076 13404
rect 31116 12232 31168 12238
rect 30944 12192 31116 12220
rect 30748 12164 30800 12170
rect 30748 12106 30800 12112
rect 30840 12164 30892 12170
rect 30840 12106 30892 12112
rect 30944 12050 30972 12192
rect 31116 12174 31168 12180
rect 30668 12022 30972 12050
rect 30472 11892 30524 11898
rect 30472 11834 30524 11840
rect 30484 11558 30512 11834
rect 30472 11552 30524 11558
rect 30472 11494 30524 11500
rect 30656 11008 30708 11014
rect 30656 10950 30708 10956
rect 30380 10736 30432 10742
rect 30380 10678 30432 10684
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 30392 9722 30420 10678
rect 30668 10062 30696 10950
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 30472 9988 30524 9994
rect 30472 9930 30524 9936
rect 30380 9716 30432 9722
rect 30380 9658 30432 9664
rect 30288 8968 30340 8974
rect 30288 8910 30340 8916
rect 30104 8560 30156 8566
rect 30104 8502 30156 8508
rect 30300 8498 30328 8910
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 29184 6656 29236 6662
rect 29184 6598 29236 6604
rect 29196 6458 29224 6598
rect 29092 6452 29144 6458
rect 29092 6394 29144 6400
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 29288 6186 29316 6258
rect 29276 6180 29328 6186
rect 29276 6122 29328 6128
rect 29288 5846 29316 6122
rect 29276 5840 29328 5846
rect 29276 5782 29328 5788
rect 30484 5778 30512 9930
rect 31128 9722 31156 10066
rect 31116 9716 31168 9722
rect 31116 9658 31168 9664
rect 30656 9512 30708 9518
rect 30656 9454 30708 9460
rect 30668 8634 30696 9454
rect 31116 8832 31168 8838
rect 31116 8774 31168 8780
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 31128 8566 31156 8774
rect 31116 8560 31168 8566
rect 31116 8502 31168 8508
rect 30564 8424 30616 8430
rect 30564 8366 30616 8372
rect 30576 7954 30604 8366
rect 31116 8288 31168 8294
rect 31116 8230 31168 8236
rect 31128 7954 31156 8230
rect 30564 7948 30616 7954
rect 30564 7890 30616 7896
rect 31116 7948 31168 7954
rect 31116 7890 31168 7896
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31128 6118 31156 6734
rect 31116 6112 31168 6118
rect 31116 6054 31168 6060
rect 30472 5772 30524 5778
rect 30472 5714 30524 5720
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 28356 5228 28408 5234
rect 28356 5170 28408 5176
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 28092 4554 28120 4762
rect 28368 4622 28396 5170
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28080 4548 28132 4554
rect 28080 4490 28132 4496
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 31128 2446 31156 6054
rect 31220 5760 31248 15524
rect 31312 14958 31340 16390
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31300 14952 31352 14958
rect 31300 14894 31352 14900
rect 31300 14816 31352 14822
rect 31300 14758 31352 14764
rect 31312 14618 31340 14758
rect 31404 14618 31432 14962
rect 31300 14612 31352 14618
rect 31300 14554 31352 14560
rect 31392 14612 31444 14618
rect 31392 14554 31444 14560
rect 31312 14414 31340 14554
rect 31496 14414 31524 17734
rect 31680 16454 31708 19450
rect 31772 19446 31800 19994
rect 32036 19848 32088 19854
rect 32036 19790 32088 19796
rect 31760 19440 31812 19446
rect 31760 19382 31812 19388
rect 31942 18728 31998 18737
rect 31942 18663 31998 18672
rect 31956 18630 31984 18663
rect 32048 18630 32076 19790
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 32036 18624 32088 18630
rect 32036 18566 32088 18572
rect 31956 18290 31984 18566
rect 31944 18284 31996 18290
rect 31944 18226 31996 18232
rect 31668 16448 31720 16454
rect 31668 16390 31720 16396
rect 31956 15434 31984 18226
rect 31944 15428 31996 15434
rect 31944 15370 31996 15376
rect 31944 15088 31996 15094
rect 31944 15030 31996 15036
rect 31576 15020 31628 15026
rect 31576 14962 31628 14968
rect 31588 14822 31616 14962
rect 31852 14952 31904 14958
rect 31852 14894 31904 14900
rect 31576 14816 31628 14822
rect 31576 14758 31628 14764
rect 31864 14550 31892 14894
rect 31852 14544 31904 14550
rect 31852 14486 31904 14492
rect 31300 14408 31352 14414
rect 31300 14350 31352 14356
rect 31484 14408 31536 14414
rect 31536 14368 31616 14396
rect 31484 14350 31536 14356
rect 31484 14272 31536 14278
rect 31484 14214 31536 14220
rect 31392 14000 31444 14006
rect 31496 13954 31524 14214
rect 31444 13948 31524 13954
rect 31392 13942 31524 13948
rect 31404 13926 31524 13942
rect 31588 13938 31616 14368
rect 31496 13326 31524 13926
rect 31576 13932 31628 13938
rect 31576 13874 31628 13880
rect 31956 13920 31984 15030
rect 32048 14822 32076 18566
rect 32140 18426 32168 20402
rect 32220 19168 32272 19174
rect 32220 19110 32272 19116
rect 32232 18766 32260 19110
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32128 18420 32180 18426
rect 32128 18362 32180 18368
rect 32232 18358 32260 18702
rect 32220 18352 32272 18358
rect 32220 18294 32272 18300
rect 32324 16538 32352 22066
rect 32496 21480 32548 21486
rect 32496 21422 32548 21428
rect 32404 20800 32456 20806
rect 32404 20742 32456 20748
rect 32416 20602 32444 20742
rect 32508 20602 32536 21422
rect 32404 20596 32456 20602
rect 32404 20538 32456 20544
rect 32496 20596 32548 20602
rect 32496 20538 32548 20544
rect 32784 20466 32812 22066
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 35348 22024 35400 22030
rect 35348 21966 35400 21972
rect 33692 21548 33744 21554
rect 33692 21490 33744 21496
rect 33140 21480 33192 21486
rect 33140 21422 33192 21428
rect 33152 20534 33180 21422
rect 33140 20528 33192 20534
rect 33140 20470 33192 20476
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32772 20460 32824 20466
rect 32772 20402 32824 20408
rect 32508 19990 32536 20402
rect 33152 20058 33180 20470
rect 33600 20392 33652 20398
rect 33600 20334 33652 20340
rect 33612 20058 33640 20334
rect 33140 20052 33192 20058
rect 33140 19994 33192 20000
rect 33600 20052 33652 20058
rect 33600 19994 33652 20000
rect 32496 19984 32548 19990
rect 32496 19926 32548 19932
rect 33704 19854 33732 21490
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34520 21004 34572 21010
rect 34520 20946 34572 20952
rect 33966 20360 34022 20369
rect 33966 20295 34022 20304
rect 33980 20262 34008 20295
rect 33968 20256 34020 20262
rect 33968 20198 34020 20204
rect 33980 19854 34008 20198
rect 34532 19990 34560 20946
rect 35256 20936 35308 20942
rect 35256 20878 35308 20884
rect 34704 20800 34756 20806
rect 34704 20742 34756 20748
rect 34796 20800 34848 20806
rect 34796 20742 34848 20748
rect 34716 20330 34744 20742
rect 34704 20324 34756 20330
rect 34704 20266 34756 20272
rect 34612 20256 34664 20262
rect 34612 20198 34664 20204
rect 34520 19984 34572 19990
rect 34520 19926 34572 19932
rect 34624 19854 34652 20198
rect 34716 20058 34744 20266
rect 34704 20052 34756 20058
rect 34704 19994 34756 20000
rect 34808 19854 34836 20742
rect 35268 20641 35296 20878
rect 35254 20632 35310 20641
rect 35360 20602 35388 21966
rect 35254 20567 35310 20576
rect 35348 20596 35400 20602
rect 35348 20538 35400 20544
rect 35348 20392 35400 20398
rect 35348 20334 35400 20340
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34980 20052 35032 20058
rect 34980 19994 35032 20000
rect 34992 19854 35020 19994
rect 35360 19854 35388 20334
rect 33692 19848 33744 19854
rect 33692 19790 33744 19796
rect 33968 19848 34020 19854
rect 33968 19790 34020 19796
rect 34612 19848 34664 19854
rect 34612 19790 34664 19796
rect 34796 19848 34848 19854
rect 34796 19790 34848 19796
rect 34980 19848 35032 19854
rect 35348 19848 35400 19854
rect 34980 19790 35032 19796
rect 35346 19816 35348 19825
rect 35400 19816 35402 19825
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 33232 19712 33284 19718
rect 33232 19654 33284 19660
rect 33324 19712 33376 19718
rect 33324 19654 33376 19660
rect 33244 19446 33272 19654
rect 33232 19440 33284 19446
rect 33232 19382 33284 19388
rect 32864 19168 32916 19174
rect 32864 19110 32916 19116
rect 32876 17218 32904 19110
rect 33138 18864 33194 18873
rect 33138 18799 33194 18808
rect 33232 18828 33284 18834
rect 33152 18766 33180 18799
rect 33232 18770 33284 18776
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 33152 18222 33180 18702
rect 33244 18426 33272 18770
rect 33336 18630 33364 19654
rect 33796 18970 33824 19722
rect 34244 19712 34296 19718
rect 34244 19654 34296 19660
rect 34256 19514 34284 19654
rect 34244 19508 34296 19514
rect 34244 19450 34296 19456
rect 34992 19334 35020 19790
rect 35346 19751 35402 19760
rect 34808 19306 35020 19334
rect 33968 19168 34020 19174
rect 33968 19110 34020 19116
rect 34152 19168 34204 19174
rect 34152 19110 34204 19116
rect 33784 18964 33836 18970
rect 33784 18906 33836 18912
rect 33876 18964 33928 18970
rect 33876 18906 33928 18912
rect 33888 18850 33916 18906
rect 33704 18822 33916 18850
rect 33324 18624 33376 18630
rect 33324 18566 33376 18572
rect 33232 18420 33284 18426
rect 33232 18362 33284 18368
rect 33336 18306 33364 18566
rect 33244 18278 33364 18306
rect 33600 18284 33652 18290
rect 33140 18216 33192 18222
rect 33140 18158 33192 18164
rect 33244 18086 33272 18278
rect 33704 18272 33732 18822
rect 33980 18766 34008 19110
rect 33784 18760 33836 18766
rect 33782 18728 33784 18737
rect 33968 18760 34020 18766
rect 33836 18728 33838 18737
rect 33968 18702 34020 18708
rect 33782 18663 33838 18672
rect 34164 18630 34192 19110
rect 34336 18760 34388 18766
rect 34336 18702 34388 18708
rect 34152 18624 34204 18630
rect 34152 18566 34204 18572
rect 33652 18244 33732 18272
rect 33784 18284 33836 18290
rect 33600 18226 33652 18232
rect 33784 18226 33836 18232
rect 33232 18080 33284 18086
rect 33232 18022 33284 18028
rect 33324 18080 33376 18086
rect 33324 18022 33376 18028
rect 33508 18080 33560 18086
rect 33508 18022 33560 18028
rect 33336 17338 33364 18022
rect 33324 17332 33376 17338
rect 33324 17274 33376 17280
rect 32876 17190 33088 17218
rect 32956 17060 33008 17066
rect 32956 17002 33008 17008
rect 32968 16590 32996 17002
rect 32956 16584 33008 16590
rect 32232 16510 32352 16538
rect 32784 16544 32956 16572
rect 32232 15706 32260 16510
rect 32312 16448 32364 16454
rect 32312 16390 32364 16396
rect 32324 16046 32352 16390
rect 32784 16114 32812 16544
rect 32956 16526 33008 16532
rect 32772 16108 32824 16114
rect 32772 16050 32824 16056
rect 32312 16040 32364 16046
rect 32784 16017 32812 16050
rect 32312 15982 32364 15988
rect 32770 16008 32826 16017
rect 32770 15943 32826 15952
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32232 15586 32260 15642
rect 32232 15558 32536 15586
rect 32220 14884 32272 14890
rect 32220 14826 32272 14832
rect 32036 14816 32088 14822
rect 32036 14758 32088 14764
rect 32232 14618 32260 14826
rect 32220 14612 32272 14618
rect 32220 14554 32272 14560
rect 32128 14544 32180 14550
rect 32128 14486 32180 14492
rect 32140 13938 32168 14486
rect 32036 13932 32088 13938
rect 31956 13892 32036 13920
rect 31588 13326 31616 13874
rect 31852 13728 31904 13734
rect 31852 13670 31904 13676
rect 31484 13320 31536 13326
rect 31484 13262 31536 13268
rect 31576 13320 31628 13326
rect 31576 13262 31628 13268
rect 31300 13184 31352 13190
rect 31300 13126 31352 13132
rect 31312 12850 31340 13126
rect 31864 12986 31892 13670
rect 31956 13444 31984 13892
rect 32036 13874 32088 13880
rect 32128 13932 32180 13938
rect 32128 13874 32180 13880
rect 32220 13932 32272 13938
rect 32220 13874 32272 13880
rect 32036 13456 32088 13462
rect 31956 13416 32036 13444
rect 32036 13398 32088 13404
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31392 12980 31444 12986
rect 31392 12922 31444 12928
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31312 12374 31340 12786
rect 31404 12782 31432 12922
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31392 12776 31444 12782
rect 31392 12718 31444 12724
rect 31668 12776 31720 12782
rect 31668 12718 31720 12724
rect 31300 12368 31352 12374
rect 31300 12310 31352 12316
rect 31404 12238 31432 12718
rect 31680 12434 31708 12718
rect 31772 12442 31800 12786
rect 31588 12406 31708 12434
rect 31760 12436 31812 12442
rect 31588 12306 31616 12406
rect 31956 12434 31984 13262
rect 32232 13190 32260 13874
rect 32220 13184 32272 13190
rect 32220 13126 32272 13132
rect 32232 12918 32260 13126
rect 32220 12912 32272 12918
rect 32220 12854 32272 12860
rect 32220 12708 32272 12714
rect 32220 12650 32272 12656
rect 32232 12434 32260 12650
rect 31956 12406 32076 12434
rect 32232 12406 32352 12434
rect 31760 12378 31812 12384
rect 31576 12300 31628 12306
rect 31576 12242 31628 12248
rect 32048 12238 32076 12406
rect 31392 12232 31444 12238
rect 31392 12174 31444 12180
rect 31668 12232 31720 12238
rect 31668 12174 31720 12180
rect 32036 12232 32088 12238
rect 32036 12174 32088 12180
rect 31300 12164 31352 12170
rect 31300 12106 31352 12112
rect 31312 10130 31340 12106
rect 31392 10600 31444 10606
rect 31392 10542 31444 10548
rect 31404 10266 31432 10542
rect 31680 10538 31708 12174
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 32140 10810 32168 11154
rect 32128 10804 32180 10810
rect 32128 10746 32180 10752
rect 31668 10532 31720 10538
rect 31668 10474 31720 10480
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31300 10124 31352 10130
rect 31300 10066 31352 10072
rect 32220 9376 32272 9382
rect 32220 9318 32272 9324
rect 31668 8968 31720 8974
rect 31668 8910 31720 8916
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 31404 8294 31432 8570
rect 31680 8498 31708 8910
rect 31760 8900 31812 8906
rect 31760 8842 31812 8848
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31392 8288 31444 8294
rect 31392 8230 31444 8236
rect 31484 8288 31536 8294
rect 31484 8230 31536 8236
rect 31496 7886 31524 8230
rect 31484 7880 31536 7886
rect 31484 7822 31536 7828
rect 31772 7546 31800 8842
rect 32232 8634 32260 9318
rect 32324 9110 32352 12406
rect 32508 11778 32536 15558
rect 32956 14068 33008 14074
rect 32956 14010 33008 14016
rect 32968 13326 32996 14010
rect 32956 13320 33008 13326
rect 32956 13262 33008 13268
rect 33060 12646 33088 17190
rect 33520 17134 33548 18022
rect 33612 17660 33640 18226
rect 33796 18086 33824 18226
rect 34164 18222 34192 18566
rect 34152 18216 34204 18222
rect 34152 18158 34204 18164
rect 33784 18080 33836 18086
rect 33784 18022 33836 18028
rect 33876 17876 33928 17882
rect 33876 17818 33928 17824
rect 33692 17672 33744 17678
rect 33612 17632 33692 17660
rect 33692 17614 33744 17620
rect 33704 17134 33732 17614
rect 33888 17202 33916 17818
rect 33876 17196 33928 17202
rect 33876 17138 33928 17144
rect 33140 17128 33192 17134
rect 33140 17070 33192 17076
rect 33508 17128 33560 17134
rect 33508 17070 33560 17076
rect 33692 17128 33744 17134
rect 33692 17070 33744 17076
rect 33784 17128 33836 17134
rect 33784 17070 33836 17076
rect 33152 16794 33180 17070
rect 33416 16992 33468 16998
rect 33416 16934 33468 16940
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 33428 16590 33456 16934
rect 33416 16584 33468 16590
rect 33520 16561 33548 17070
rect 33598 16688 33654 16697
rect 33598 16623 33600 16632
rect 33652 16623 33654 16632
rect 33600 16594 33652 16600
rect 33416 16526 33468 16532
rect 33506 16552 33562 16561
rect 33506 16487 33562 16496
rect 33520 16454 33548 16487
rect 33508 16448 33560 16454
rect 33508 16390 33560 16396
rect 33600 16108 33652 16114
rect 33520 16068 33600 16096
rect 33416 16040 33468 16046
rect 33416 15982 33468 15988
rect 33428 15706 33456 15982
rect 33416 15700 33468 15706
rect 33416 15642 33468 15648
rect 33520 15586 33548 16068
rect 33600 16050 33652 16056
rect 33600 15904 33652 15910
rect 33600 15846 33652 15852
rect 33428 15558 33548 15586
rect 33230 14376 33286 14385
rect 33286 14334 33364 14362
rect 33230 14311 33286 14320
rect 33336 14278 33364 14334
rect 33324 14272 33376 14278
rect 33324 14214 33376 14220
rect 33232 14068 33284 14074
rect 33232 14010 33284 14016
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 33152 13530 33180 13874
rect 33140 13524 33192 13530
rect 33140 13466 33192 13472
rect 33244 12918 33272 14010
rect 33336 13938 33364 14214
rect 33324 13932 33376 13938
rect 33324 13874 33376 13880
rect 33232 12912 33284 12918
rect 33232 12854 33284 12860
rect 32588 12640 32640 12646
rect 32588 12582 32640 12588
rect 33048 12640 33100 12646
rect 33048 12582 33100 12588
rect 32600 12434 32628 12582
rect 32600 12406 32812 12434
rect 32508 11750 32720 11778
rect 32496 11348 32548 11354
rect 32496 11290 32548 11296
rect 32508 10062 32536 11290
rect 32588 11280 32640 11286
rect 32588 11222 32640 11228
rect 32600 10742 32628 11222
rect 32692 11150 32720 11750
rect 32784 11218 32812 12406
rect 33060 12374 33088 12582
rect 33048 12368 33100 12374
rect 33048 12310 33100 12316
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32772 11212 32824 11218
rect 32772 11154 32824 11160
rect 32680 11144 32732 11150
rect 32680 11086 32732 11092
rect 32588 10736 32640 10742
rect 32588 10678 32640 10684
rect 32864 10600 32916 10606
rect 32864 10542 32916 10548
rect 32588 10192 32640 10198
rect 32588 10134 32640 10140
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32600 9586 32628 10134
rect 32680 9920 32732 9926
rect 32680 9862 32732 9868
rect 32772 9920 32824 9926
rect 32772 9862 32824 9868
rect 32692 9722 32720 9862
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 32588 9580 32640 9586
rect 32588 9522 32640 9528
rect 32692 9466 32720 9658
rect 32784 9654 32812 9862
rect 32876 9722 32904 10542
rect 32968 10044 32996 12174
rect 33428 11014 33456 15558
rect 33612 13938 33640 15846
rect 33704 15638 33732 17070
rect 33796 16454 33824 17070
rect 34164 16998 34192 18158
rect 34152 16992 34204 16998
rect 34152 16934 34204 16940
rect 34244 16992 34296 16998
rect 34244 16934 34296 16940
rect 33968 16584 34020 16590
rect 33968 16526 34020 16532
rect 34150 16552 34206 16561
rect 33784 16448 33836 16454
rect 33784 16390 33836 16396
rect 33876 16448 33928 16454
rect 33876 16390 33928 16396
rect 33692 15632 33744 15638
rect 33692 15574 33744 15580
rect 33796 15366 33824 16390
rect 33888 16114 33916 16390
rect 33980 16114 34008 16526
rect 34150 16487 34206 16496
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33968 16108 34020 16114
rect 33968 16050 34020 16056
rect 33980 15502 34008 16050
rect 34164 15994 34192 16487
rect 34256 16114 34284 16934
rect 34244 16108 34296 16114
rect 34244 16050 34296 16056
rect 34164 15978 34284 15994
rect 34164 15972 34296 15978
rect 34164 15966 34244 15972
rect 34244 15914 34296 15920
rect 33968 15496 34020 15502
rect 33968 15438 34020 15444
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 33784 15360 33836 15366
rect 33784 15302 33836 15308
rect 33968 15020 34020 15026
rect 33968 14962 34020 14968
rect 33980 14550 34008 14962
rect 33968 14544 34020 14550
rect 33968 14486 34020 14492
rect 33784 14476 33836 14482
rect 33784 14418 33836 14424
rect 33600 13932 33652 13938
rect 33600 13874 33652 13880
rect 33692 13728 33744 13734
rect 33692 13670 33744 13676
rect 33704 12306 33732 13670
rect 33796 12918 33824 14418
rect 33980 14074 34008 14486
rect 33968 14068 34020 14074
rect 33968 14010 34020 14016
rect 34072 13954 34100 15438
rect 34242 14104 34298 14113
rect 34242 14039 34298 14048
rect 34256 14006 34284 14039
rect 33980 13926 34100 13954
rect 34244 14000 34296 14006
rect 34244 13942 34296 13948
rect 34348 13938 34376 18702
rect 34704 18420 34756 18426
rect 34704 18362 34756 18368
rect 34612 18352 34664 18358
rect 34612 18294 34664 18300
rect 34520 18080 34572 18086
rect 34520 18022 34572 18028
rect 34532 17542 34560 18022
rect 34624 17610 34652 18294
rect 34716 17678 34744 18362
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 34612 17604 34664 17610
rect 34612 17546 34664 17552
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 34532 16794 34560 17478
rect 34520 16788 34572 16794
rect 34520 16730 34572 16736
rect 34624 16726 34652 17546
rect 34612 16720 34664 16726
rect 34612 16662 34664 16668
rect 34428 16448 34480 16454
rect 34428 16390 34480 16396
rect 34520 16448 34572 16454
rect 34520 16390 34572 16396
rect 34440 16114 34468 16390
rect 34532 16182 34560 16390
rect 34520 16176 34572 16182
rect 34520 16118 34572 16124
rect 34428 16108 34480 16114
rect 34428 16050 34480 16056
rect 34704 16108 34756 16114
rect 34704 16050 34756 16056
rect 34716 15706 34744 16050
rect 34704 15700 34756 15706
rect 34704 15642 34756 15648
rect 34612 15632 34664 15638
rect 34612 15574 34664 15580
rect 34520 14272 34572 14278
rect 34520 14214 34572 14220
rect 34152 13932 34204 13938
rect 33980 13734 34008 13926
rect 34152 13874 34204 13880
rect 34336 13932 34388 13938
rect 34336 13874 34388 13880
rect 33968 13728 34020 13734
rect 33968 13670 34020 13676
rect 34164 13326 34192 13874
rect 34532 13326 34560 14214
rect 34624 13938 34652 15574
rect 34704 15020 34756 15026
rect 34704 14962 34756 14968
rect 34716 14074 34744 14962
rect 34704 14068 34756 14074
rect 34704 14010 34756 14016
rect 34612 13932 34664 13938
rect 34612 13874 34664 13880
rect 34704 13932 34756 13938
rect 34704 13874 34756 13880
rect 34152 13320 34204 13326
rect 34428 13320 34480 13326
rect 34152 13262 34204 13268
rect 34426 13288 34428 13297
rect 34520 13320 34572 13326
rect 34480 13288 34482 13297
rect 34520 13262 34572 13268
rect 34426 13223 34482 13232
rect 33784 12912 33836 12918
rect 33784 12854 33836 12860
rect 34532 12782 34560 13262
rect 34520 12776 34572 12782
rect 34520 12718 34572 12724
rect 33692 12300 33744 12306
rect 33692 12242 33744 12248
rect 34624 12238 34652 13874
rect 34716 13462 34744 13874
rect 34808 13802 34836 19306
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35452 18426 35480 22034
rect 35532 20868 35584 20874
rect 35532 20810 35584 20816
rect 35544 20398 35572 20810
rect 35624 20596 35676 20602
rect 35624 20538 35676 20544
rect 35532 20392 35584 20398
rect 35532 20334 35584 20340
rect 35440 18420 35492 18426
rect 35440 18362 35492 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 35636 17954 35664 20538
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35544 17926 35664 17954
rect 35544 17678 35572 17926
rect 35532 17672 35584 17678
rect 35532 17614 35584 17620
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35348 15904 35400 15910
rect 35348 15846 35400 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15706 35388 15846
rect 35348 15700 35400 15706
rect 35348 15642 35400 15648
rect 35532 15360 35584 15366
rect 35532 15302 35584 15308
rect 35440 14816 35492 14822
rect 35440 14758 35492 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35256 14612 35308 14618
rect 35256 14554 35308 14560
rect 35268 14346 35296 14554
rect 35452 14482 35480 14758
rect 35348 14476 35400 14482
rect 35348 14418 35400 14424
rect 35440 14476 35492 14482
rect 35440 14418 35492 14424
rect 35256 14340 35308 14346
rect 35256 14282 35308 14288
rect 35360 14006 35388 14418
rect 35544 14414 35572 15302
rect 35624 15020 35676 15026
rect 35624 14962 35676 14968
rect 35532 14408 35584 14414
rect 35532 14350 35584 14356
rect 35348 14000 35400 14006
rect 34886 13968 34942 13977
rect 35636 13977 35664 14962
rect 35348 13942 35400 13948
rect 35622 13968 35678 13977
rect 34886 13903 34888 13912
rect 34940 13903 34942 13912
rect 35532 13932 35584 13938
rect 34888 13874 34940 13880
rect 35622 13903 35678 13912
rect 35532 13874 35584 13880
rect 34796 13796 34848 13802
rect 34796 13738 34848 13744
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35544 13546 35572 13874
rect 35452 13530 35572 13546
rect 35636 13530 35664 13903
rect 35440 13524 35572 13530
rect 35492 13518 35572 13524
rect 35624 13524 35676 13530
rect 35440 13466 35492 13472
rect 35624 13466 35676 13472
rect 34704 13456 34756 13462
rect 35728 13410 35756 23122
rect 35808 22500 35860 22506
rect 35808 22442 35860 22448
rect 35820 21078 35848 22442
rect 36464 22094 36492 29038
rect 36544 24132 36596 24138
rect 36544 24074 36596 24080
rect 36556 23866 36584 24074
rect 36544 23860 36596 23866
rect 36544 23802 36596 23808
rect 36740 23662 36768 29056
rect 37280 28552 37332 28558
rect 37280 28494 37332 28500
rect 37292 28218 37320 28494
rect 37280 28212 37332 28218
rect 37280 28154 37332 28160
rect 36820 27940 36872 27946
rect 36820 27882 36872 27888
rect 36832 27538 36860 27882
rect 36820 27532 36872 27538
rect 36820 27474 36872 27480
rect 36820 25764 36872 25770
rect 36820 25706 36872 25712
rect 36832 25294 36860 25706
rect 36820 25288 36872 25294
rect 36820 25230 36872 25236
rect 37004 24132 37056 24138
rect 37004 24074 37056 24080
rect 36636 23656 36688 23662
rect 36636 23598 36688 23604
rect 36728 23656 36780 23662
rect 36728 23598 36780 23604
rect 36280 22066 36492 22094
rect 36084 21480 36136 21486
rect 36084 21422 36136 21428
rect 35808 21072 35860 21078
rect 35808 21014 35860 21020
rect 35992 20936 36044 20942
rect 35900 20902 35952 20908
rect 35992 20878 36044 20884
rect 35900 20844 35952 20850
rect 35808 20800 35860 20806
rect 35808 20742 35860 20748
rect 35820 20505 35848 20742
rect 35806 20496 35862 20505
rect 35912 20466 35940 20844
rect 35806 20431 35862 20440
rect 35900 20460 35952 20466
rect 35820 19922 35848 20431
rect 35900 20402 35952 20408
rect 35912 20058 35940 20402
rect 35900 20052 35952 20058
rect 35900 19994 35952 20000
rect 35808 19916 35860 19922
rect 35808 19858 35860 19864
rect 36004 19802 36032 20878
rect 36096 20806 36124 21422
rect 36084 20800 36136 20806
rect 36084 20742 36136 20748
rect 36176 20800 36228 20806
rect 36176 20742 36228 20748
rect 36188 20466 36216 20742
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 36188 20058 36216 20402
rect 36176 20052 36228 20058
rect 36176 19994 36228 20000
rect 36084 19916 36136 19922
rect 36084 19858 36136 19864
rect 35820 19774 36032 19802
rect 35820 18970 35848 19774
rect 35992 19304 36044 19310
rect 35992 19246 36044 19252
rect 35808 18964 35860 18970
rect 35808 18906 35860 18912
rect 36004 18630 36032 19246
rect 36096 19242 36124 19858
rect 36084 19236 36136 19242
rect 36084 19178 36136 19184
rect 36096 18766 36124 19178
rect 36084 18760 36136 18766
rect 36084 18702 36136 18708
rect 35992 18624 36044 18630
rect 35992 18566 36044 18572
rect 35900 18216 35952 18222
rect 35900 18158 35952 18164
rect 35912 17882 35940 18158
rect 35900 17876 35952 17882
rect 35900 17818 35952 17824
rect 35900 17740 35952 17746
rect 35900 17682 35952 17688
rect 35912 16454 35940 17682
rect 36004 16590 36032 18566
rect 36280 16998 36308 22066
rect 36648 22030 36676 23598
rect 37016 22710 37044 24074
rect 37752 23798 37780 32370
rect 37924 29572 37976 29578
rect 37924 29514 37976 29520
rect 37936 28490 37964 29514
rect 37924 28484 37976 28490
rect 37924 28426 37976 28432
rect 38028 24410 38056 41386
rect 40880 41206 40908 41958
rect 40868 41200 40920 41206
rect 40868 41142 40920 41148
rect 41236 41132 41288 41138
rect 41236 41074 41288 41080
rect 40776 41064 40828 41070
rect 40776 41006 40828 41012
rect 40408 40928 40460 40934
rect 40408 40870 40460 40876
rect 40420 40730 40448 40870
rect 40408 40724 40460 40730
rect 40408 40666 40460 40672
rect 40788 40497 40816 41006
rect 41248 40905 41276 41074
rect 41234 40896 41290 40905
rect 41234 40831 41290 40840
rect 40774 40488 40830 40497
rect 38660 40452 38712 40458
rect 40774 40423 40830 40432
rect 38660 40394 38712 40400
rect 38672 39370 38700 40394
rect 39304 40384 39356 40390
rect 39304 40326 39356 40332
rect 39316 39642 39344 40326
rect 39304 39636 39356 39642
rect 39304 39578 39356 39584
rect 38660 39364 38712 39370
rect 38660 39306 38712 39312
rect 38672 38654 38700 39306
rect 39672 39296 39724 39302
rect 39672 39238 39724 39244
rect 38580 38626 38700 38654
rect 38580 37942 38608 38626
rect 38568 37936 38620 37942
rect 38568 37878 38620 37884
rect 38108 32496 38160 32502
rect 38108 32438 38160 32444
rect 38120 29646 38148 32438
rect 38580 32366 38608 37878
rect 39120 32904 39172 32910
rect 39120 32846 39172 32852
rect 38568 32360 38620 32366
rect 38568 32302 38620 32308
rect 38108 29640 38160 29646
rect 38108 29582 38160 29588
rect 38120 28626 38148 29582
rect 39132 28762 39160 32846
rect 39120 28756 39172 28762
rect 39120 28698 39172 28704
rect 38108 28620 38160 28626
rect 38108 28562 38160 28568
rect 38108 28484 38160 28490
rect 38108 28426 38160 28432
rect 38120 27334 38148 28426
rect 39132 28082 39160 28698
rect 39120 28076 39172 28082
rect 39120 28018 39172 28024
rect 38108 27328 38160 27334
rect 38108 27270 38160 27276
rect 39684 26450 39712 39238
rect 40960 37120 41012 37126
rect 40960 37062 41012 37068
rect 40972 36825 41000 37062
rect 40958 36816 41014 36825
rect 40958 36751 41014 36760
rect 40960 32768 41012 32774
rect 40958 32736 40960 32745
rect 41012 32736 41014 32745
rect 40958 32671 41014 32680
rect 40958 30152 41014 30161
rect 40958 30087 41014 30096
rect 40972 29306 41000 30087
rect 40960 29300 41012 29306
rect 40960 29242 41012 29248
rect 41328 29028 41380 29034
rect 41328 28970 41380 28976
rect 41340 28665 41368 28970
rect 41326 28656 41382 28665
rect 41326 28591 41382 28600
rect 39672 26444 39724 26450
rect 39672 26386 39724 26392
rect 41328 24676 41380 24682
rect 41328 24618 41380 24624
rect 41052 24608 41104 24614
rect 41340 24585 41368 24618
rect 41052 24550 41104 24556
rect 41326 24576 41382 24585
rect 38016 24404 38068 24410
rect 38016 24346 38068 24352
rect 38028 23866 38056 24346
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38016 23860 38068 23866
rect 38016 23802 38068 23808
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37004 22704 37056 22710
rect 37004 22646 37056 22652
rect 36636 22024 36688 22030
rect 36636 21966 36688 21972
rect 36820 21888 36872 21894
rect 36820 21830 36872 21836
rect 36832 21554 36860 21830
rect 36820 21548 36872 21554
rect 36820 21490 36872 21496
rect 37280 21548 37332 21554
rect 37280 21490 37332 21496
rect 36452 20800 36504 20806
rect 36452 20742 36504 20748
rect 37096 20800 37148 20806
rect 37096 20742 37148 20748
rect 36358 20632 36414 20641
rect 36358 20567 36414 20576
rect 36372 19854 36400 20567
rect 36464 20369 36492 20742
rect 36542 20496 36598 20505
rect 36542 20431 36544 20440
rect 36596 20431 36598 20440
rect 36728 20460 36780 20466
rect 36544 20402 36596 20408
rect 36728 20402 36780 20408
rect 36450 20360 36506 20369
rect 36450 20295 36506 20304
rect 36740 20058 36768 20402
rect 36728 20052 36780 20058
rect 36728 19994 36780 20000
rect 36360 19848 36412 19854
rect 36360 19790 36412 19796
rect 36820 18760 36872 18766
rect 36820 18702 36872 18708
rect 36728 18692 36780 18698
rect 36728 18634 36780 18640
rect 36740 18426 36768 18634
rect 36832 18426 36860 18702
rect 37108 18698 37136 20742
rect 37292 20330 37320 21490
rect 37384 20618 37412 22918
rect 37556 22568 37608 22574
rect 37556 22510 37608 22516
rect 37568 22234 37596 22510
rect 37556 22228 37608 22234
rect 37556 22170 37608 22176
rect 37752 22166 37780 23734
rect 38304 23662 38332 24142
rect 38292 23656 38344 23662
rect 38292 23598 38344 23604
rect 38304 22438 38332 23598
rect 41064 22681 41092 24550
rect 41326 24511 41382 24520
rect 41050 22672 41106 22681
rect 41050 22607 41106 22616
rect 39304 22568 39356 22574
rect 39304 22510 39356 22516
rect 38292 22432 38344 22438
rect 38292 22374 38344 22380
rect 37740 22160 37792 22166
rect 37740 22102 37792 22108
rect 37648 22092 37700 22098
rect 37648 22034 37700 22040
rect 37556 22024 37608 22030
rect 37556 21966 37608 21972
rect 37464 21888 37516 21894
rect 37464 21830 37516 21836
rect 37476 21690 37504 21830
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37384 20590 37504 20618
rect 37372 20460 37424 20466
rect 37372 20402 37424 20408
rect 37280 20324 37332 20330
rect 37280 20266 37332 20272
rect 37280 19848 37332 19854
rect 37280 19790 37332 19796
rect 37292 19310 37320 19790
rect 37384 19378 37412 20402
rect 37372 19372 37424 19378
rect 37372 19314 37424 19320
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 37384 18834 37412 19314
rect 37372 18828 37424 18834
rect 37372 18770 37424 18776
rect 37096 18692 37148 18698
rect 37148 18652 37228 18680
rect 37096 18634 37148 18640
rect 36728 18420 36780 18426
rect 36728 18362 36780 18368
rect 36820 18420 36872 18426
rect 36820 18362 36872 18368
rect 36544 18284 36596 18290
rect 36544 18226 36596 18232
rect 37096 18284 37148 18290
rect 37096 18226 37148 18232
rect 36556 17746 36584 18226
rect 36544 17740 36596 17746
rect 36544 17682 36596 17688
rect 36358 17640 36414 17649
rect 36358 17575 36360 17584
rect 36412 17575 36414 17584
rect 36360 17546 36412 17552
rect 36268 16992 36320 16998
rect 36268 16934 36320 16940
rect 35992 16584 36044 16590
rect 35992 16526 36044 16532
rect 36556 16454 36584 17682
rect 36636 17264 36688 17270
rect 36636 17206 36688 17212
rect 35900 16448 35952 16454
rect 35900 16390 35952 16396
rect 36544 16448 36596 16454
rect 36544 16390 36596 16396
rect 36556 15473 36584 16390
rect 36648 15978 36676 17206
rect 37108 16114 37136 18226
rect 36820 16108 36872 16114
rect 37096 16108 37148 16114
rect 36872 16068 37096 16096
rect 36820 16050 36872 16056
rect 37096 16050 37148 16056
rect 36636 15972 36688 15978
rect 36636 15914 36688 15920
rect 36542 15464 36598 15473
rect 36542 15399 36598 15408
rect 35808 14884 35860 14890
rect 35808 14826 35860 14832
rect 35820 14482 35848 14826
rect 35808 14476 35860 14482
rect 35808 14418 35860 14424
rect 34704 13398 34756 13404
rect 34716 13190 34744 13398
rect 35452 13382 35756 13410
rect 35072 13252 35124 13258
rect 35072 13194 35124 13200
rect 34704 13184 34756 13190
rect 34704 13126 34756 13132
rect 35084 12918 35112 13194
rect 35072 12912 35124 12918
rect 35072 12854 35124 12860
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34612 12232 34664 12238
rect 34612 12174 34664 12180
rect 34794 12064 34850 12073
rect 34794 11999 34850 12008
rect 33600 11620 33652 11626
rect 33600 11562 33652 11568
rect 33508 11212 33560 11218
rect 33508 11154 33560 11160
rect 33416 11008 33468 11014
rect 33416 10950 33468 10956
rect 33232 10804 33284 10810
rect 33232 10746 33284 10752
rect 33048 10668 33100 10674
rect 33048 10610 33100 10616
rect 33060 10266 33088 10610
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 33048 10260 33100 10266
rect 33048 10202 33100 10208
rect 33152 10062 33180 10406
rect 33048 10056 33100 10062
rect 32968 10016 33048 10044
rect 33048 9998 33100 10004
rect 33140 10056 33192 10062
rect 33140 9998 33192 10004
rect 32864 9716 32916 9722
rect 32864 9658 32916 9664
rect 32772 9648 32824 9654
rect 32772 9590 32824 9596
rect 32692 9438 32904 9466
rect 32312 9104 32364 9110
rect 32312 9046 32364 9052
rect 32220 8628 32272 8634
rect 32220 8570 32272 8576
rect 32036 8424 32088 8430
rect 32036 8366 32088 8372
rect 32048 7750 32076 8366
rect 32220 8288 32272 8294
rect 32220 8230 32272 8236
rect 32232 7818 32260 8230
rect 32220 7812 32272 7818
rect 32220 7754 32272 7760
rect 32036 7744 32088 7750
rect 32036 7686 32088 7692
rect 31760 7540 31812 7546
rect 31760 7482 31812 7488
rect 32876 5846 32904 9438
rect 33060 8838 33088 9998
rect 33140 9376 33192 9382
rect 33140 9318 33192 9324
rect 33152 9042 33180 9318
rect 33140 9036 33192 9042
rect 33140 8978 33192 8984
rect 33244 8974 33272 10746
rect 33520 10470 33548 11154
rect 33612 10810 33640 11562
rect 34808 11218 34836 11999
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11212 34848 11218
rect 34796 11154 34848 11160
rect 34808 10810 34836 11154
rect 35256 11008 35308 11014
rect 35256 10950 35308 10956
rect 35268 10810 35296 10950
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 34796 10804 34848 10810
rect 34796 10746 34848 10752
rect 35256 10804 35308 10810
rect 35256 10746 35308 10752
rect 33612 10606 33640 10746
rect 33784 10668 33836 10674
rect 33784 10610 33836 10616
rect 34612 10668 34664 10674
rect 34612 10610 34664 10616
rect 33600 10600 33652 10606
rect 33600 10542 33652 10548
rect 33508 10464 33560 10470
rect 33508 10406 33560 10412
rect 33796 9994 33824 10610
rect 34624 10062 34652 10610
rect 34796 10464 34848 10470
rect 34796 10406 34848 10412
rect 34704 10192 34756 10198
rect 34704 10134 34756 10140
rect 34612 10056 34664 10062
rect 34612 9998 34664 10004
rect 33784 9988 33836 9994
rect 33784 9930 33836 9936
rect 34624 9926 34652 9998
rect 34612 9920 34664 9926
rect 34612 9862 34664 9868
rect 34520 9172 34572 9178
rect 34520 9114 34572 9120
rect 33876 9104 33928 9110
rect 33876 9046 33928 9052
rect 33232 8968 33284 8974
rect 33232 8910 33284 8916
rect 33600 8900 33652 8906
rect 33600 8842 33652 8848
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33612 8566 33640 8842
rect 33600 8560 33652 8566
rect 33600 8502 33652 8508
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 33060 7546 33088 7822
rect 33612 7750 33640 8502
rect 33888 8498 33916 9046
rect 34532 8922 34560 9114
rect 34060 8900 34112 8906
rect 34060 8842 34112 8848
rect 34440 8894 34560 8922
rect 34612 8968 34664 8974
rect 34612 8910 34664 8916
rect 34072 8634 34100 8842
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33692 8356 33744 8362
rect 33692 8298 33744 8304
rect 33704 7886 33732 8298
rect 34072 7886 34100 8570
rect 34440 8498 34468 8894
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34532 8566 34560 8774
rect 34520 8560 34572 8566
rect 34520 8502 34572 8508
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34440 8378 34468 8434
rect 34440 8350 34560 8378
rect 34532 7886 34560 8350
rect 34624 8090 34652 8910
rect 34716 8498 34744 10134
rect 34808 10062 34836 10406
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 10056 34848 10062
rect 34796 9998 34848 10004
rect 35256 9988 35308 9994
rect 35256 9930 35308 9936
rect 34796 9920 34848 9926
rect 34796 9862 34848 9868
rect 34808 9058 34836 9862
rect 35268 9722 35296 9930
rect 35256 9716 35308 9722
rect 35256 9658 35308 9664
rect 35452 9674 35480 13382
rect 35532 13320 35584 13326
rect 35584 13268 35756 13274
rect 35532 13262 35756 13268
rect 35544 13258 35756 13262
rect 35544 13252 35768 13258
rect 35544 13246 35716 13252
rect 35716 13194 35768 13200
rect 35716 12300 35768 12306
rect 35716 12242 35768 12248
rect 35728 11830 35756 12242
rect 35716 11824 35768 11830
rect 35716 11766 35768 11772
rect 35532 11688 35584 11694
rect 35532 11630 35584 11636
rect 35544 11082 35572 11630
rect 35716 11552 35768 11558
rect 35716 11494 35768 11500
rect 35728 11354 35756 11494
rect 35716 11348 35768 11354
rect 35716 11290 35768 11296
rect 35532 11076 35584 11082
rect 35532 11018 35584 11024
rect 35452 9646 35664 9674
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34808 9030 34928 9058
rect 34900 8514 34928 9030
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34808 8486 34928 8514
rect 34612 8084 34664 8090
rect 34612 8026 34664 8032
rect 34612 7948 34664 7954
rect 34612 7890 34664 7896
rect 33692 7880 33744 7886
rect 33692 7822 33744 7828
rect 34060 7880 34112 7886
rect 34060 7822 34112 7828
rect 34520 7880 34572 7886
rect 34520 7822 34572 7828
rect 33600 7744 33652 7750
rect 33600 7686 33652 7692
rect 33048 7540 33100 7546
rect 33048 7482 33100 7488
rect 32864 5840 32916 5846
rect 32864 5782 32916 5788
rect 33060 5778 33088 7482
rect 34624 7410 34652 7890
rect 34612 7404 34664 7410
rect 34612 7346 34664 7352
rect 34624 6322 34652 7346
rect 34612 6316 34664 6322
rect 34612 6258 34664 6264
rect 31300 5772 31352 5778
rect 31220 5732 31300 5760
rect 31300 5714 31352 5720
rect 33048 5772 33100 5778
rect 33048 5714 33100 5720
rect 31760 5636 31812 5642
rect 31760 5578 31812 5584
rect 31852 5636 31904 5642
rect 31852 5578 31904 5584
rect 31772 5234 31800 5578
rect 31864 5370 31892 5578
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34532 5370 34560 5510
rect 34624 5370 34652 6258
rect 34808 5778 34836 8486
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35440 8288 35492 8294
rect 35440 8230 35492 8236
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35452 7342 35480 8230
rect 35544 8022 35572 8366
rect 35532 8016 35584 8022
rect 35532 7958 35584 7964
rect 35544 7342 35572 7958
rect 35440 7336 35492 7342
rect 35440 7278 35492 7284
rect 35532 7336 35584 7342
rect 35532 7278 35584 7284
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35636 5778 35664 9646
rect 35820 8974 35848 14418
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 35900 14340 35952 14346
rect 35900 14282 35952 14288
rect 35912 14074 35940 14282
rect 35900 14068 35952 14074
rect 35900 14010 35952 14016
rect 35900 13864 35952 13870
rect 35900 13806 35952 13812
rect 35912 13530 35940 13806
rect 35992 13728 36044 13734
rect 35992 13670 36044 13676
rect 35900 13524 35952 13530
rect 35900 13466 35952 13472
rect 36004 13394 36032 13670
rect 35992 13388 36044 13394
rect 35992 13330 36044 13336
rect 35900 13320 35952 13326
rect 35898 13288 35900 13297
rect 35952 13288 35954 13297
rect 35898 13223 35954 13232
rect 36096 12866 36124 14350
rect 36188 13240 36216 14350
rect 36268 13796 36320 13802
rect 36268 13738 36320 13744
rect 36280 13462 36308 13738
rect 36648 13682 36676 15914
rect 37200 14618 37228 18652
rect 37384 17338 37412 18770
rect 37476 18290 37504 20590
rect 37568 19922 37596 21966
rect 37660 20874 37688 22034
rect 37648 20868 37700 20874
rect 37648 20810 37700 20816
rect 37832 20392 37884 20398
rect 38304 20380 38332 22374
rect 39316 22098 39344 22510
rect 39304 22092 39356 22098
rect 39304 22034 39356 22040
rect 39120 21140 39172 21146
rect 39120 21082 39172 21088
rect 38568 20868 38620 20874
rect 38568 20810 38620 20816
rect 38844 20868 38896 20874
rect 38844 20810 38896 20816
rect 39028 20868 39080 20874
rect 39028 20810 39080 20816
rect 38384 20392 38436 20398
rect 38304 20352 38384 20380
rect 37832 20334 37884 20340
rect 38384 20334 38436 20340
rect 37556 19916 37608 19922
rect 37556 19858 37608 19864
rect 37844 19854 37872 20334
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37648 19780 37700 19786
rect 37648 19722 37700 19728
rect 37660 18970 37688 19722
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 38396 18358 38424 20334
rect 38580 18970 38608 20810
rect 38856 20602 38884 20810
rect 38844 20596 38896 20602
rect 38844 20538 38896 20544
rect 38660 20392 38712 20398
rect 38660 20334 38712 20340
rect 38672 20058 38700 20334
rect 38660 20052 38712 20058
rect 38660 19994 38712 20000
rect 38856 19854 38884 20538
rect 39040 20262 39068 20810
rect 39132 20534 39160 21082
rect 39212 20800 39264 20806
rect 39212 20742 39264 20748
rect 39120 20528 39172 20534
rect 39120 20470 39172 20476
rect 39028 20256 39080 20262
rect 39028 20198 39080 20204
rect 38936 19984 38988 19990
rect 38936 19926 38988 19932
rect 38844 19848 38896 19854
rect 38844 19790 38896 19796
rect 38568 18964 38620 18970
rect 38568 18906 38620 18912
rect 38752 18624 38804 18630
rect 38752 18566 38804 18572
rect 38384 18352 38436 18358
rect 38384 18294 38436 18300
rect 38764 18290 38792 18566
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 38752 18284 38804 18290
rect 38752 18226 38804 18232
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 38844 18216 38896 18222
rect 38844 18158 38896 18164
rect 37844 17542 37872 18158
rect 38856 17882 38884 18158
rect 38844 17876 38896 17882
rect 38844 17818 38896 17824
rect 37832 17536 37884 17542
rect 37832 17478 37884 17484
rect 37372 17332 37424 17338
rect 37372 17274 37424 17280
rect 37740 16448 37792 16454
rect 37740 16390 37792 16396
rect 37372 15972 37424 15978
rect 37372 15914 37424 15920
rect 37188 14612 37240 14618
rect 37188 14554 37240 14560
rect 36556 13654 36676 13682
rect 36268 13456 36320 13462
rect 36268 13398 36320 13404
rect 36268 13252 36320 13258
rect 36188 13212 36268 13240
rect 36188 12986 36216 13212
rect 36268 13194 36320 13200
rect 36176 12980 36228 12986
rect 36176 12922 36228 12928
rect 36096 12838 36216 12866
rect 36084 11756 36136 11762
rect 36084 11698 36136 11704
rect 35992 11552 36044 11558
rect 35992 11494 36044 11500
rect 36004 11218 36032 11494
rect 35992 11212 36044 11218
rect 35992 11154 36044 11160
rect 36096 11150 36124 11698
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 35992 10600 36044 10606
rect 35992 10542 36044 10548
rect 36004 10266 36032 10542
rect 36084 10464 36136 10470
rect 36084 10406 36136 10412
rect 35992 10260 36044 10266
rect 35992 10202 36044 10208
rect 36096 8974 36124 10406
rect 36188 9654 36216 12838
rect 36556 11558 36584 13654
rect 36636 13252 36688 13258
rect 36636 13194 36688 13200
rect 36648 12918 36676 13194
rect 37384 12968 37412 15914
rect 37384 12940 37596 12968
rect 36636 12912 36688 12918
rect 36636 12854 36688 12860
rect 36544 11552 36596 11558
rect 36544 11494 36596 11500
rect 36176 9648 36228 9654
rect 36176 9590 36228 9596
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 36084 8968 36136 8974
rect 36084 8910 36136 8916
rect 35820 8634 35848 8910
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 36188 8430 36216 9590
rect 36452 9376 36504 9382
rect 36452 9318 36504 9324
rect 36464 9042 36492 9318
rect 36452 9036 36504 9042
rect 36452 8978 36504 8984
rect 36176 8424 36228 8430
rect 36176 8366 36228 8372
rect 36648 6798 36676 12854
rect 37384 12782 37412 12940
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 37372 12776 37424 12782
rect 37372 12718 37424 12724
rect 37476 11626 37504 12786
rect 37568 11694 37596 12940
rect 37556 11688 37608 11694
rect 37556 11630 37608 11636
rect 37464 11620 37516 11626
rect 37464 11562 37516 11568
rect 36728 11552 36780 11558
rect 36728 11494 36780 11500
rect 36740 11218 36768 11494
rect 36728 11212 36780 11218
rect 36728 11154 36780 11160
rect 36820 11008 36872 11014
rect 36820 10950 36872 10956
rect 36832 10742 36860 10950
rect 36820 10736 36872 10742
rect 36820 10678 36872 10684
rect 37096 9648 37148 9654
rect 37096 9590 37148 9596
rect 37188 9648 37240 9654
rect 37188 9590 37240 9596
rect 36912 9376 36964 9382
rect 36912 9318 36964 9324
rect 36924 9042 36952 9318
rect 36912 9036 36964 9042
rect 36912 8978 36964 8984
rect 37108 8974 37136 9590
rect 37096 8968 37148 8974
rect 37096 8910 37148 8916
rect 37200 8634 37228 9590
rect 37372 9580 37424 9586
rect 37372 9522 37424 9528
rect 37384 8974 37412 9522
rect 37372 8968 37424 8974
rect 37372 8910 37424 8916
rect 37280 8832 37332 8838
rect 37280 8774 37332 8780
rect 37292 8634 37320 8774
rect 37188 8628 37240 8634
rect 37188 8570 37240 8576
rect 37280 8628 37332 8634
rect 37280 8570 37332 8576
rect 37384 8514 37412 8910
rect 37464 8832 37516 8838
rect 37464 8774 37516 8780
rect 37476 8566 37504 8774
rect 37200 8498 37412 8514
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37648 8560 37700 8566
rect 37648 8502 37700 8508
rect 37188 8492 37412 8498
rect 37240 8486 37412 8492
rect 37188 8434 37240 8440
rect 37280 8424 37332 8430
rect 37280 8366 37332 8372
rect 37384 8378 37412 8486
rect 37660 8378 37688 8502
rect 37292 7342 37320 8366
rect 37384 8350 37688 8378
rect 37280 7336 37332 7342
rect 37280 7278 37332 7284
rect 36636 6792 36688 6798
rect 36636 6734 36688 6740
rect 37292 6730 37320 7278
rect 37280 6724 37332 6730
rect 37280 6666 37332 6672
rect 37096 6316 37148 6322
rect 37096 6258 37148 6264
rect 37108 5914 37136 6258
rect 37292 6254 37320 6666
rect 37280 6248 37332 6254
rect 37280 6190 37332 6196
rect 37096 5908 37148 5914
rect 37096 5850 37148 5856
rect 34796 5772 34848 5778
rect 34796 5714 34848 5720
rect 35624 5772 35676 5778
rect 35624 5714 35676 5720
rect 34704 5704 34756 5710
rect 34704 5646 34756 5652
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 31852 5364 31904 5370
rect 31852 5306 31904 5312
rect 34520 5364 34572 5370
rect 34520 5306 34572 5312
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 34716 2774 34744 5646
rect 36280 5030 36308 5646
rect 36268 5024 36320 5030
rect 36268 4966 36320 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 36280 4826 36308 4966
rect 36268 4820 36320 4826
rect 36268 4762 36320 4768
rect 37292 4146 37320 6190
rect 37464 4752 37516 4758
rect 37464 4694 37516 4700
rect 37476 4214 37504 4694
rect 37752 4690 37780 16390
rect 37844 16114 37872 17478
rect 37924 17196 37976 17202
rect 37924 17138 37976 17144
rect 38476 17196 38528 17202
rect 38476 17138 38528 17144
rect 37936 16726 37964 17138
rect 38488 16794 38516 17138
rect 38752 17060 38804 17066
rect 38752 17002 38804 17008
rect 38476 16788 38528 16794
rect 38476 16730 38528 16736
rect 37924 16720 37976 16726
rect 38660 16720 38712 16726
rect 37924 16662 37976 16668
rect 38658 16688 38660 16697
rect 38712 16688 38714 16697
rect 38658 16623 38714 16632
rect 38660 16584 38712 16590
rect 38658 16552 38660 16561
rect 38712 16552 38714 16561
rect 38658 16487 38714 16496
rect 38476 16448 38528 16454
rect 38476 16390 38528 16396
rect 38660 16448 38712 16454
rect 38764 16436 38792 17002
rect 38948 16998 38976 19926
rect 39040 19854 39068 20198
rect 39028 19848 39080 19854
rect 39028 19790 39080 19796
rect 39132 19378 39160 20470
rect 39224 19922 39252 20742
rect 41512 20732 41564 20738
rect 41512 20674 41564 20680
rect 41524 20505 41552 20674
rect 41510 20496 41566 20505
rect 41510 20431 41566 20440
rect 39212 19916 39264 19922
rect 39212 19858 39264 19864
rect 39120 19372 39172 19378
rect 39120 19314 39172 19320
rect 40040 19372 40092 19378
rect 40040 19314 40092 19320
rect 39672 18828 39724 18834
rect 39672 18770 39724 18776
rect 39304 18692 39356 18698
rect 39304 18634 39356 18640
rect 39120 18216 39172 18222
rect 39120 18158 39172 18164
rect 38936 16992 38988 16998
rect 38936 16934 38988 16940
rect 38948 16794 38976 16934
rect 38844 16788 38896 16794
rect 38844 16730 38896 16736
rect 38936 16788 38988 16794
rect 38936 16730 38988 16736
rect 38856 16572 38884 16730
rect 38936 16584 38988 16590
rect 38856 16544 38936 16572
rect 38936 16526 38988 16532
rect 38844 16448 38896 16454
rect 38764 16408 38844 16436
rect 38660 16390 38712 16396
rect 38844 16390 38896 16396
rect 38488 16114 38516 16390
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 38476 16108 38528 16114
rect 38476 16050 38528 16056
rect 38292 14340 38344 14346
rect 38292 14282 38344 14288
rect 38304 13870 38332 14282
rect 38488 13870 38516 16050
rect 38672 15366 38700 16390
rect 39028 16040 39080 16046
rect 39028 15982 39080 15988
rect 38660 15360 38712 15366
rect 38660 15302 38712 15308
rect 38672 14822 38700 15302
rect 38660 14816 38712 14822
rect 38660 14758 38712 14764
rect 38844 14816 38896 14822
rect 38844 14758 38896 14764
rect 38856 14634 38884 14758
rect 38672 14606 38884 14634
rect 38672 14414 38700 14606
rect 38752 14544 38804 14550
rect 38804 14504 38976 14532
rect 38752 14486 38804 14492
rect 38660 14408 38712 14414
rect 38580 14368 38660 14396
rect 38292 13864 38344 13870
rect 38292 13806 38344 13812
rect 38476 13864 38528 13870
rect 38476 13806 38528 13812
rect 38384 13728 38436 13734
rect 38384 13670 38436 13676
rect 38396 13326 38424 13670
rect 38580 13394 38608 14368
rect 38660 14350 38712 14356
rect 38752 14408 38804 14414
rect 38842 14376 38898 14385
rect 38804 14356 38842 14362
rect 38752 14350 38842 14356
rect 38764 14334 38842 14350
rect 38842 14311 38898 14320
rect 38660 13932 38712 13938
rect 38660 13874 38712 13880
rect 38672 13734 38700 13874
rect 38752 13864 38804 13870
rect 38752 13806 38804 13812
rect 38660 13728 38712 13734
rect 38660 13670 38712 13676
rect 38568 13388 38620 13394
rect 38568 13330 38620 13336
rect 38384 13320 38436 13326
rect 38384 13262 38436 13268
rect 38660 13320 38712 13326
rect 38660 13262 38712 13268
rect 38396 12850 38424 13262
rect 38672 12986 38700 13262
rect 38764 13258 38792 13806
rect 38948 13530 38976 14504
rect 39040 13870 39068 15982
rect 39028 13864 39080 13870
rect 39028 13806 39080 13812
rect 38936 13524 38988 13530
rect 38936 13466 38988 13472
rect 39132 13326 39160 18158
rect 39212 17264 39264 17270
rect 39212 17206 39264 17212
rect 39224 16794 39252 17206
rect 39316 16794 39344 18634
rect 39396 17604 39448 17610
rect 39396 17546 39448 17552
rect 39408 16998 39436 17546
rect 39488 17536 39540 17542
rect 39488 17478 39540 17484
rect 39500 17066 39528 17478
rect 39488 17060 39540 17066
rect 39488 17002 39540 17008
rect 39396 16992 39448 16998
rect 39396 16934 39448 16940
rect 39212 16788 39264 16794
rect 39212 16730 39264 16736
rect 39304 16788 39356 16794
rect 39304 16730 39356 16736
rect 39316 16674 39344 16730
rect 39224 16646 39344 16674
rect 39578 16688 39634 16697
rect 39224 16250 39252 16646
rect 39578 16623 39580 16632
rect 39632 16623 39634 16632
rect 39580 16594 39632 16600
rect 39396 16584 39448 16590
rect 39394 16552 39396 16561
rect 39448 16552 39450 16561
rect 39304 16516 39356 16522
rect 39394 16487 39450 16496
rect 39304 16458 39356 16464
rect 39212 16244 39264 16250
rect 39212 16186 39264 16192
rect 39316 15910 39344 16458
rect 39488 16448 39540 16454
rect 39488 16390 39540 16396
rect 39500 16250 39528 16390
rect 39488 16244 39540 16250
rect 39488 16186 39540 16192
rect 39304 15904 39356 15910
rect 39304 15846 39356 15852
rect 39316 15026 39344 15846
rect 39488 15360 39540 15366
rect 39488 15302 39540 15308
rect 39304 15020 39356 15026
rect 39304 14962 39356 14968
rect 39316 14414 39344 14962
rect 39396 14884 39448 14890
rect 39396 14826 39448 14832
rect 39408 14414 39436 14826
rect 39500 14550 39528 15302
rect 39580 14816 39632 14822
rect 39580 14758 39632 14764
rect 39488 14544 39540 14550
rect 39488 14486 39540 14492
rect 39592 14414 39620 14758
rect 39304 14408 39356 14414
rect 39304 14350 39356 14356
rect 39396 14408 39448 14414
rect 39396 14350 39448 14356
rect 39580 14408 39632 14414
rect 39580 14350 39632 14356
rect 39304 14272 39356 14278
rect 39304 14214 39356 14220
rect 39316 14006 39344 14214
rect 39408 14074 39436 14350
rect 39396 14068 39448 14074
rect 39396 14010 39448 14016
rect 39304 14000 39356 14006
rect 39304 13942 39356 13948
rect 39120 13320 39172 13326
rect 39120 13262 39172 13268
rect 39396 13320 39448 13326
rect 39396 13262 39448 13268
rect 38752 13252 38804 13258
rect 38752 13194 38804 13200
rect 38660 12980 38712 12986
rect 38660 12922 38712 12928
rect 38384 12844 38436 12850
rect 38384 12786 38436 12792
rect 38396 11830 38424 12786
rect 39132 12434 39160 13262
rect 39132 12406 39344 12434
rect 38660 12232 38712 12238
rect 38660 12174 38712 12180
rect 38476 12096 38528 12102
rect 38476 12038 38528 12044
rect 38384 11824 38436 11830
rect 38384 11766 38436 11772
rect 38488 11694 38516 12038
rect 38476 11688 38528 11694
rect 38476 11630 38528 11636
rect 38672 11354 38700 12174
rect 38844 11824 38896 11830
rect 38844 11766 38896 11772
rect 38660 11348 38712 11354
rect 38660 11290 38712 11296
rect 38752 11212 38804 11218
rect 38752 11154 38804 11160
rect 38016 11144 38068 11150
rect 38016 11086 38068 11092
rect 37924 9580 37976 9586
rect 37924 9522 37976 9528
rect 37936 8974 37964 9522
rect 37924 8968 37976 8974
rect 37924 8910 37976 8916
rect 37832 7948 37884 7954
rect 37832 7890 37884 7896
rect 37844 5778 37872 7890
rect 38028 7886 38056 11086
rect 38660 11008 38712 11014
rect 38660 10950 38712 10956
rect 38672 10810 38700 10950
rect 38764 10810 38792 11154
rect 38660 10804 38712 10810
rect 38660 10746 38712 10752
rect 38752 10804 38804 10810
rect 38752 10746 38804 10752
rect 38660 10464 38712 10470
rect 38660 10406 38712 10412
rect 38672 9738 38700 10406
rect 38580 9722 38700 9738
rect 38568 9716 38700 9722
rect 38620 9710 38700 9716
rect 38568 9658 38620 9664
rect 38568 9512 38620 9518
rect 38568 9454 38620 9460
rect 38580 9042 38608 9454
rect 38660 9444 38712 9450
rect 38660 9386 38712 9392
rect 38672 9042 38700 9386
rect 38568 9036 38620 9042
rect 38568 8978 38620 8984
rect 38660 9036 38712 9042
rect 38660 8978 38712 8984
rect 38856 8566 38884 11766
rect 39028 11076 39080 11082
rect 39028 11018 39080 11024
rect 39040 10130 39068 11018
rect 39316 10606 39344 12406
rect 39120 10600 39172 10606
rect 39120 10542 39172 10548
rect 39304 10600 39356 10606
rect 39304 10542 39356 10548
rect 39132 10266 39160 10542
rect 39120 10260 39172 10266
rect 39120 10202 39172 10208
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 39408 10062 39436 13262
rect 39580 12776 39632 12782
rect 39580 12718 39632 12724
rect 39592 12442 39620 12718
rect 39684 12646 39712 18770
rect 39856 18624 39908 18630
rect 39856 18566 39908 18572
rect 39868 18426 39896 18566
rect 39856 18420 39908 18426
rect 39856 18362 39908 18368
rect 40052 18358 40080 19314
rect 40960 18624 41012 18630
rect 40960 18566 41012 18572
rect 40972 18426 41000 18566
rect 40960 18420 41012 18426
rect 40960 18362 41012 18368
rect 40040 18352 40092 18358
rect 40040 18294 40092 18300
rect 40052 16182 40080 18294
rect 40592 17672 40644 17678
rect 40592 17614 40644 17620
rect 40500 17604 40552 17610
rect 40500 17546 40552 17552
rect 40512 17134 40540 17546
rect 40500 17128 40552 17134
rect 40500 17070 40552 17076
rect 40512 16250 40540 17070
rect 40604 16658 40632 17614
rect 41512 17468 41564 17474
rect 41512 17410 41564 17416
rect 41052 16992 41104 16998
rect 41052 16934 41104 16940
rect 40592 16652 40644 16658
rect 40592 16594 40644 16600
rect 40500 16244 40552 16250
rect 40500 16186 40552 16192
rect 40040 16176 40092 16182
rect 40040 16118 40092 16124
rect 39764 15156 39816 15162
rect 39764 15098 39816 15104
rect 39776 14482 39804 15098
rect 39764 14476 39816 14482
rect 39764 14418 39816 14424
rect 39776 13734 39804 14418
rect 40052 14006 40080 16118
rect 40498 14376 40554 14385
rect 40498 14311 40500 14320
rect 40552 14311 40554 14320
rect 40500 14282 40552 14288
rect 40040 14000 40092 14006
rect 40040 13942 40092 13948
rect 39764 13728 39816 13734
rect 39764 13670 39816 13676
rect 39776 13326 39804 13670
rect 39764 13320 39816 13326
rect 39764 13262 39816 13268
rect 39764 13184 39816 13190
rect 39764 13126 39816 13132
rect 39856 13184 39908 13190
rect 39856 13126 39908 13132
rect 39672 12640 39724 12646
rect 39672 12582 39724 12588
rect 39580 12436 39632 12442
rect 39580 12378 39632 12384
rect 39684 11218 39712 12582
rect 39672 11212 39724 11218
rect 39672 11154 39724 11160
rect 39776 10130 39804 13126
rect 39868 12345 39896 13126
rect 40052 12918 40080 13942
rect 40040 12912 40092 12918
rect 40040 12854 40092 12860
rect 39854 12336 39910 12345
rect 40604 12306 40632 16594
rect 41064 16590 41092 16934
rect 41052 16584 41104 16590
rect 41052 16526 41104 16532
rect 41524 16425 41552 17410
rect 41510 16416 41566 16425
rect 41510 16351 41566 16360
rect 41052 13184 41104 13190
rect 41052 13126 41104 13132
rect 39854 12271 39910 12280
rect 40592 12300 40644 12306
rect 40592 12242 40644 12248
rect 41064 12238 41092 13126
rect 41052 12232 41104 12238
rect 41052 12174 41104 12180
rect 39856 11552 39908 11558
rect 39856 11494 39908 11500
rect 39868 11286 39896 11494
rect 39856 11280 39908 11286
rect 39856 11222 39908 11228
rect 39764 10124 39816 10130
rect 39764 10066 39816 10072
rect 39212 10056 39264 10062
rect 39212 9998 39264 10004
rect 39396 10056 39448 10062
rect 39396 9998 39448 10004
rect 39224 9722 39252 9998
rect 39396 9920 39448 9926
rect 39396 9862 39448 9868
rect 39580 9920 39632 9926
rect 39580 9862 39632 9868
rect 39212 9716 39264 9722
rect 39212 9658 39264 9664
rect 39408 9586 39436 9862
rect 39592 9586 39620 9862
rect 39396 9580 39448 9586
rect 39396 9522 39448 9528
rect 39580 9580 39632 9586
rect 39580 9522 39632 9528
rect 39776 9450 39804 10066
rect 39856 10056 39908 10062
rect 39856 9998 39908 10004
rect 39868 9722 39896 9998
rect 39856 9716 39908 9722
rect 39856 9658 39908 9664
rect 39764 9444 39816 9450
rect 39764 9386 39816 9392
rect 38844 8560 38896 8566
rect 38844 8502 38896 8508
rect 38016 7880 38068 7886
rect 38016 7822 38068 7828
rect 38856 7478 38884 8502
rect 40684 8492 40736 8498
rect 40684 8434 40736 8440
rect 40696 7886 40724 8434
rect 41052 8356 41104 8362
rect 41052 8298 41104 8304
rect 41064 8265 41092 8298
rect 41050 8256 41106 8265
rect 41050 8191 41106 8200
rect 40684 7880 40736 7886
rect 40684 7822 40736 7828
rect 39120 7744 39172 7750
rect 39120 7686 39172 7692
rect 38844 7472 38896 7478
rect 38844 7414 38896 7420
rect 38856 6390 38884 7414
rect 39132 7342 39160 7686
rect 40696 7546 40724 7822
rect 40684 7540 40736 7546
rect 40684 7482 40736 7488
rect 39120 7336 39172 7342
rect 39120 7278 39172 7284
rect 38844 6384 38896 6390
rect 38844 6326 38896 6332
rect 37832 5772 37884 5778
rect 37832 5714 37884 5720
rect 37844 4690 37872 5714
rect 38856 5302 38884 6326
rect 40684 6248 40736 6254
rect 40684 6190 40736 6196
rect 39764 6112 39816 6118
rect 39764 6054 39816 6060
rect 39776 5914 39804 6054
rect 39764 5908 39816 5914
rect 39764 5850 39816 5856
rect 38844 5296 38896 5302
rect 38844 5238 38896 5244
rect 37740 4684 37792 4690
rect 37740 4626 37792 4632
rect 37832 4684 37884 4690
rect 37832 4626 37884 4632
rect 38856 4214 38884 5238
rect 39028 4616 39080 4622
rect 39028 4558 39080 4564
rect 37464 4208 37516 4214
rect 37464 4150 37516 4156
rect 38844 4208 38896 4214
rect 38844 4150 38896 4156
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 39040 3942 39068 4558
rect 39028 3936 39080 3942
rect 39028 3878 39080 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34624 2746 34744 2774
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34624 2446 34652 2746
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 39040 2446 39068 3878
rect 40696 2446 40724 6190
rect 41052 4480 41104 4486
rect 41052 4422 41104 4428
rect 41064 4185 41092 4422
rect 41050 4176 41106 4185
rect 41050 4111 41106 4120
rect 20812 2440 20864 2446
rect 31116 2440 31168 2446
rect 20812 2382 20864 2388
rect 32 800 60 2314
rect 3896 800 3924 2366
rect 3988 2310 4016 2366
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 23216 2366 23336 2394
rect 31116 2382 31168 2388
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 39028 2440 39080 2446
rect 39028 2382 39080 2388
rect 40684 2440 40736 2446
rect 40684 2382 40736 2388
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 7760 800 7788 2246
rect 11624 800 11652 2246
rect 15488 800 15516 2246
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 23216 800 23244 2366
rect 23308 2310 23336 2366
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 39948 2304 40000 2310
rect 39948 2246 40000 2252
rect 27080 800 27108 2246
rect 30944 800 30972 2246
rect 34808 800 34836 2246
rect 38672 800 38700 2246
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 15474 0 15530 800
rect 19338 0 19394 800
rect 23202 0 23258 800
rect 27066 0 27122 800
rect 30930 0 30986 800
rect 34794 0 34850 800
rect 38658 0 38714 800
rect 39960 105 39988 2246
rect 39946 96 40002 105
rect 39946 31 40002 40
<< via2 >>
rect 2778 44240 2834 44296
rect 938 40160 994 40216
rect 938 36080 994 36136
rect 938 32000 994 32056
rect 938 27940 994 27976
rect 938 27920 940 27940
rect 940 27920 992 27940
rect 992 27920 994 27940
rect 938 23840 994 23896
rect 938 19780 994 19816
rect 938 19760 940 19780
rect 940 19760 992 19780
rect 992 19760 994 19780
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 14646 41792 14702 41848
rect 19430 41792 19486 41848
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 6826 34720 6882 34776
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4986 26288 5042 26344
rect 6090 32852 6092 32872
rect 6092 32852 6144 32872
rect 6144 32852 6146 32872
rect 6090 32816 6146 32852
rect 5722 31864 5778 31920
rect 10874 41384 10930 41440
rect 7378 34584 7434 34640
rect 6826 25336 6882 25392
rect 1674 19780 1730 19816
rect 1674 19760 1676 19780
rect 1676 19760 1728 19780
rect 1728 19760 1730 19780
rect 938 15680 994 15736
rect 938 11600 994 11656
rect 4526 21548 4582 21584
rect 4526 21528 4528 21548
rect 4528 21528 4580 21548
rect 4580 21528 4582 21548
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4618 19216 4674 19272
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4342 18708 4344 18728
rect 4344 18708 4396 18728
rect 4396 18708 4398 18728
rect 4342 18672 4398 18708
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 8206 33632 8262 33688
rect 7930 32020 7986 32056
rect 7930 32000 7932 32020
rect 7932 32000 7984 32020
rect 7984 32000 7986 32020
rect 8390 32952 8446 33008
rect 8942 35692 8998 35728
rect 8942 35672 8944 35692
rect 8944 35672 8996 35692
rect 8996 35672 8998 35692
rect 8298 31320 8354 31376
rect 8758 31728 8814 31784
rect 10966 40060 10968 40080
rect 10968 40060 11020 40080
rect 11020 40060 11022 40080
rect 10966 40024 11022 40060
rect 10782 37032 10838 37088
rect 9586 36760 9642 36816
rect 9586 34992 9642 35048
rect 9310 32136 9366 32192
rect 8114 26152 8170 26208
rect 9678 32272 9734 32328
rect 9586 32136 9642 32192
rect 10046 35672 10102 35728
rect 10046 34584 10102 34640
rect 9586 31728 9642 31784
rect 9402 31456 9458 31512
rect 9126 28076 9182 28112
rect 9126 28056 9128 28076
rect 9128 28056 9180 28076
rect 9180 28056 9182 28076
rect 8390 24656 8446 24712
rect 8850 27412 8852 27432
rect 8852 27412 8904 27432
rect 8904 27412 8906 27432
rect 8850 27376 8906 27412
rect 9034 26288 9090 26344
rect 9586 31356 9588 31376
rect 9588 31356 9640 31376
rect 9640 31356 9642 31376
rect 9586 31320 9642 31356
rect 9678 29028 9734 29064
rect 9678 29008 9680 29028
rect 9680 29008 9732 29028
rect 9732 29008 9734 29028
rect 9586 27412 9588 27432
rect 9588 27412 9640 27432
rect 9640 27412 9642 27432
rect 9586 27376 9642 27412
rect 10138 28872 10194 28928
rect 9402 26560 9458 26616
rect 9402 26152 9458 26208
rect 9586 25780 9588 25800
rect 9588 25780 9640 25800
rect 9640 25780 9642 25800
rect 9586 25744 9642 25780
rect 9862 25880 9918 25936
rect 10874 35672 10930 35728
rect 10690 34720 10746 34776
rect 11058 34584 11114 34640
rect 11150 32408 11206 32464
rect 10690 32000 10746 32056
rect 10782 31728 10838 31784
rect 10690 31592 10746 31648
rect 10966 30368 11022 30424
rect 11150 31320 11206 31376
rect 10506 29824 10562 29880
rect 10506 29180 10508 29200
rect 10508 29180 10560 29200
rect 10560 29180 10562 29200
rect 10506 29144 10562 29180
rect 10414 29008 10470 29064
rect 10322 27240 10378 27296
rect 10138 26868 10140 26888
rect 10140 26868 10192 26888
rect 10192 26868 10194 26888
rect 10138 26832 10194 26868
rect 9770 25744 9826 25800
rect 9034 25220 9090 25256
rect 9494 25236 9496 25256
rect 9496 25236 9548 25256
rect 9548 25236 9550 25256
rect 9034 25200 9036 25220
rect 9036 25200 9088 25220
rect 9088 25200 9090 25220
rect 9494 25200 9550 25236
rect 9218 24792 9274 24848
rect 8482 23432 8538 23488
rect 9310 24692 9312 24712
rect 9312 24692 9364 24712
rect 9364 24692 9366 24712
rect 9310 24656 9366 24692
rect 9218 23196 9220 23216
rect 9220 23196 9272 23216
rect 9272 23196 9274 23216
rect 9218 23160 9274 23196
rect 7102 21564 7104 21584
rect 7104 21564 7156 21584
rect 7156 21564 7158 21584
rect 7102 21528 7158 21564
rect 5170 20712 5226 20768
rect 5814 19236 5870 19272
rect 5814 19216 5816 19236
rect 5816 19216 5868 19236
rect 5868 19216 5870 19236
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 938 7520 994 7576
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 5262 13640 5318 13696
rect 5446 15136 5502 15192
rect 7562 21004 7618 21040
rect 7562 20984 7564 21004
rect 7564 20984 7616 21004
rect 7616 20984 7618 21004
rect 7470 18692 7526 18728
rect 7470 18672 7472 18692
rect 7472 18672 7524 18692
rect 7524 18672 7526 18692
rect 8574 22344 8630 22400
rect 8206 21956 8262 21992
rect 8206 21936 8208 21956
rect 8208 21936 8260 21956
rect 8260 21936 8262 21956
rect 8390 21548 8446 21584
rect 8390 21528 8392 21548
rect 8392 21528 8444 21548
rect 8444 21528 8446 21548
rect 11058 29416 11114 29472
rect 10874 28056 10930 28112
rect 12806 41012 12808 41032
rect 12808 41012 12860 41032
rect 12860 41012 12862 41032
rect 12806 40976 12862 41012
rect 13358 39072 13414 39128
rect 7010 11056 7066 11112
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 7838 12688 7894 12744
rect 9034 12708 9090 12744
rect 9034 12688 9036 12708
rect 9036 12688 9088 12708
rect 9088 12688 9090 12708
rect 9586 17740 9642 17776
rect 9586 17720 9588 17740
rect 9588 17720 9640 17740
rect 9640 17720 9642 17740
rect 11610 29960 11666 30016
rect 11518 28192 11574 28248
rect 11610 27920 11666 27976
rect 11426 27512 11482 27568
rect 11794 32816 11850 32872
rect 11886 32428 11942 32464
rect 11886 32408 11888 32428
rect 11888 32408 11940 32428
rect 11940 32408 11942 32428
rect 11794 32000 11850 32056
rect 10782 25608 10838 25664
rect 10598 23704 10654 23760
rect 11334 25200 11390 25256
rect 11058 24112 11114 24168
rect 11518 24384 11574 24440
rect 10782 21664 10838 21720
rect 10598 21392 10654 21448
rect 10506 18284 10562 18320
rect 10506 18264 10508 18284
rect 10508 18264 10560 18284
rect 10560 18264 10562 18284
rect 10598 18164 10600 18184
rect 10600 18164 10652 18184
rect 10652 18164 10654 18184
rect 10598 18128 10654 18164
rect 11426 22752 11482 22808
rect 9494 10004 9496 10024
rect 9496 10004 9548 10024
rect 9548 10004 9550 10024
rect 9494 9968 9550 10004
rect 9586 6704 9642 6760
rect 12530 33396 12532 33416
rect 12532 33396 12584 33416
rect 12584 33396 12586 33416
rect 12530 33360 12586 33396
rect 12530 32680 12586 32736
rect 12530 32136 12586 32192
rect 12438 29452 12440 29472
rect 12440 29452 12492 29472
rect 12492 29452 12494 29472
rect 12438 29416 12494 29452
rect 12162 28736 12218 28792
rect 15106 40180 15162 40216
rect 15106 40160 15108 40180
rect 15108 40160 15160 40180
rect 15160 40160 15162 40180
rect 15106 40044 15162 40080
rect 15106 40024 15108 40044
rect 15108 40024 15160 40044
rect 15160 40024 15162 40044
rect 14278 37984 14334 38040
rect 16210 40996 16266 41032
rect 16210 40976 16212 40996
rect 16212 40976 16264 40996
rect 16264 40976 16266 40996
rect 16578 40704 16634 40760
rect 16026 40468 16028 40488
rect 16028 40468 16080 40488
rect 16080 40468 16082 40488
rect 16026 40432 16082 40468
rect 17130 40976 17186 41032
rect 17222 40840 17278 40896
rect 16486 40296 16542 40352
rect 16762 40160 16818 40216
rect 16118 37984 16174 38040
rect 15290 37304 15346 37360
rect 16946 40060 16948 40080
rect 16948 40060 17000 40080
rect 17000 40060 17002 40080
rect 16946 40024 17002 40060
rect 18970 41656 19026 41712
rect 17682 40024 17738 40080
rect 16118 37304 16174 37360
rect 15934 37032 15990 37088
rect 15382 36624 15438 36680
rect 16762 36780 16818 36816
rect 16762 36760 16764 36780
rect 16764 36760 16816 36780
rect 16816 36760 16818 36780
rect 16578 36352 16634 36408
rect 16210 36216 16266 36272
rect 13542 35944 13598 36000
rect 13174 35012 13230 35048
rect 13174 34992 13176 35012
rect 13176 34992 13228 35012
rect 13228 34992 13230 35012
rect 12898 34584 12954 34640
rect 12990 33224 13046 33280
rect 12898 31864 12954 31920
rect 12622 29008 12678 29064
rect 12254 28328 12310 28384
rect 12162 26696 12218 26752
rect 11426 21836 11428 21856
rect 11428 21836 11480 21856
rect 11480 21836 11482 21856
rect 11426 21800 11482 21836
rect 11426 19896 11482 19952
rect 12530 28092 12532 28112
rect 12532 28092 12584 28112
rect 12584 28092 12586 28112
rect 12530 28056 12586 28092
rect 12530 24692 12532 24712
rect 12532 24692 12584 24712
rect 12584 24692 12586 24712
rect 12530 24656 12586 24692
rect 12530 23840 12586 23896
rect 12714 26424 12770 26480
rect 12714 22480 12770 22536
rect 11242 16496 11298 16552
rect 11426 16108 11482 16144
rect 11426 16088 11428 16108
rect 11428 16088 11480 16108
rect 11480 16088 11482 16108
rect 10598 12180 10600 12200
rect 10600 12180 10652 12200
rect 10652 12180 10654 12200
rect 10598 12144 10654 12180
rect 11426 10004 11428 10024
rect 11428 10004 11480 10024
rect 11480 10004 11482 10024
rect 11426 9968 11482 10004
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 938 3440 994 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 12346 20032 12402 20088
rect 13082 32272 13138 32328
rect 14094 35128 14150 35184
rect 13634 33904 13690 33960
rect 13542 33768 13598 33824
rect 13082 30232 13138 30288
rect 12990 29144 13046 29200
rect 12898 26560 12954 26616
rect 13174 29960 13230 30016
rect 14002 32952 14058 33008
rect 13542 32544 13598 32600
rect 13910 31884 13966 31920
rect 13910 31864 13912 31884
rect 13912 31864 13964 31884
rect 13964 31864 13966 31884
rect 13634 30504 13690 30560
rect 13358 29552 13414 29608
rect 14002 30232 14058 30288
rect 13266 26968 13322 27024
rect 13174 26036 13230 26072
rect 13174 26016 13176 26036
rect 13176 26016 13228 26036
rect 13228 26016 13230 26036
rect 13174 24928 13230 24984
rect 13726 27920 13782 27976
rect 14002 29280 14058 29336
rect 13634 25472 13690 25528
rect 12990 24384 13046 24440
rect 13450 23840 13506 23896
rect 13082 22208 13138 22264
rect 12530 20168 12586 20224
rect 12990 22072 13046 22128
rect 12990 21800 13046 21856
rect 12898 20576 12954 20632
rect 13910 24656 13966 24712
rect 13358 22108 13360 22128
rect 13360 22108 13412 22128
rect 13412 22108 13414 22128
rect 13358 22072 13414 22108
rect 15382 35028 15384 35048
rect 15384 35028 15436 35048
rect 15436 35028 15438 35048
rect 15382 34992 15438 35028
rect 15106 33904 15162 33960
rect 15014 32272 15070 32328
rect 14738 29280 14794 29336
rect 15106 29552 15162 29608
rect 14646 27940 14702 27976
rect 14646 27920 14648 27940
rect 14648 27920 14700 27940
rect 14700 27920 14702 27940
rect 14646 27548 14648 27568
rect 14648 27548 14700 27568
rect 14700 27548 14702 27568
rect 14646 27512 14702 27548
rect 14646 27104 14702 27160
rect 14554 25472 14610 25528
rect 14554 23568 14610 23624
rect 15382 29688 15438 29744
rect 18050 41012 18052 41032
rect 18052 41012 18104 41032
rect 18104 41012 18106 41032
rect 18050 40976 18106 41012
rect 17958 39244 17960 39264
rect 17960 39244 18012 39264
rect 18012 39244 18014 39264
rect 17958 39208 18014 39244
rect 18418 41112 18474 41168
rect 18142 40468 18144 40488
rect 18144 40468 18196 40488
rect 18196 40468 18198 40488
rect 18142 40432 18198 40468
rect 18878 40976 18934 41032
rect 18418 40024 18474 40080
rect 17222 36080 17278 36136
rect 16578 35944 16634 36000
rect 18326 39072 18382 39128
rect 18602 40568 18658 40624
rect 18602 40296 18658 40352
rect 18602 39380 18604 39400
rect 18604 39380 18656 39400
rect 18656 39380 18658 39400
rect 18602 39344 18658 39380
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 20166 41248 20222 41304
rect 19246 40840 19302 40896
rect 18970 39208 19026 39264
rect 18234 36644 18290 36680
rect 18234 36624 18236 36644
rect 18236 36624 18288 36644
rect 18288 36624 18290 36644
rect 18510 36916 18566 36952
rect 18510 36896 18512 36916
rect 18512 36896 18564 36916
rect 18564 36896 18566 36916
rect 17682 35808 17738 35864
rect 18878 36896 18934 36952
rect 19338 40296 19394 40352
rect 19982 40296 20038 40352
rect 19154 39380 19156 39400
rect 19156 39380 19208 39400
rect 19208 39380 19210 39400
rect 19154 39344 19210 39380
rect 19062 36780 19118 36816
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 20718 41656 20774 41712
rect 20166 40160 20222 40216
rect 21638 41248 21694 41304
rect 19798 39752 19854 39808
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19062 36760 19064 36780
rect 19064 36760 19116 36780
rect 19116 36760 19118 36780
rect 19246 36488 19302 36544
rect 19338 36080 19394 36136
rect 19522 36080 19578 36136
rect 18510 35944 18566 36000
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19890 35536 19946 35592
rect 16670 35164 16672 35184
rect 16672 35164 16724 35184
rect 16724 35164 16726 35184
rect 15934 34584 15990 34640
rect 16026 33088 16082 33144
rect 16210 33632 16266 33688
rect 15842 28056 15898 28112
rect 16670 35128 16726 35164
rect 16762 32816 16818 32872
rect 17038 32952 17094 33008
rect 16670 31728 16726 31784
rect 16302 30368 16358 30424
rect 16302 30232 16358 30288
rect 16026 29452 16028 29472
rect 16028 29452 16080 29472
rect 16080 29452 16082 29472
rect 16026 29416 16082 29452
rect 16026 28736 16082 28792
rect 15198 27412 15200 27432
rect 15200 27412 15252 27432
rect 15252 27412 15254 27432
rect 15198 27376 15254 27412
rect 14830 24792 14886 24848
rect 15382 26444 15438 26480
rect 15382 26424 15384 26444
rect 15384 26424 15436 26444
rect 15436 26424 15438 26444
rect 15014 24928 15070 24984
rect 14830 24520 14886 24576
rect 15382 26288 15438 26344
rect 15474 25472 15530 25528
rect 16118 28328 16174 28384
rect 15842 26444 15898 26480
rect 15842 26424 15844 26444
rect 15844 26424 15896 26444
rect 15896 26424 15898 26444
rect 16026 25472 16082 25528
rect 15658 24828 15660 24848
rect 15660 24828 15712 24848
rect 15712 24828 15714 24848
rect 15658 24792 15714 24828
rect 15198 24692 15200 24712
rect 15200 24692 15252 24712
rect 15252 24692 15254 24712
rect 15198 24656 15254 24692
rect 15198 24404 15254 24440
rect 15198 24384 15200 24404
rect 15200 24384 15252 24404
rect 15252 24384 15254 24404
rect 15658 23976 15714 24032
rect 15014 23296 15070 23352
rect 15198 23160 15254 23216
rect 15106 22616 15162 22672
rect 14002 20304 14058 20360
rect 13174 17176 13230 17232
rect 12070 16496 12126 16552
rect 11702 15156 11758 15192
rect 11702 15136 11704 15156
rect 11704 15136 11756 15156
rect 11756 15136 11758 15156
rect 12346 16108 12402 16144
rect 12346 16088 12348 16108
rect 12348 16088 12400 16108
rect 12400 16088 12402 16108
rect 12162 14456 12218 14512
rect 13082 13232 13138 13288
rect 14186 17312 14242 17368
rect 13634 11736 13690 11792
rect 14738 21256 14794 21312
rect 15658 21800 15714 21856
rect 15934 24248 15990 24304
rect 16026 23432 16082 23488
rect 16118 23024 16174 23080
rect 16118 22752 16174 22808
rect 16486 30096 16542 30152
rect 16578 29824 16634 29880
rect 17038 32272 17094 32328
rect 17130 31864 17186 31920
rect 16486 27376 16542 27432
rect 16670 27648 16726 27704
rect 16486 26324 16488 26344
rect 16488 26324 16540 26344
rect 16540 26324 16542 26344
rect 16486 26288 16542 26324
rect 17314 33224 17370 33280
rect 16946 29144 17002 29200
rect 16946 27240 17002 27296
rect 17406 31884 17462 31920
rect 17406 31864 17408 31884
rect 17408 31864 17460 31884
rect 17460 31864 17462 31884
rect 17314 28872 17370 28928
rect 17038 26696 17094 26752
rect 16670 25608 16726 25664
rect 16026 21120 16082 21176
rect 15934 19488 15990 19544
rect 16762 25472 16818 25528
rect 16670 23840 16726 23896
rect 17038 25064 17094 25120
rect 17038 24384 17094 24440
rect 17314 27104 17370 27160
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 17774 32000 17830 32056
rect 18418 32680 18474 32736
rect 18418 32544 18474 32600
rect 18142 31048 18198 31104
rect 17958 30640 18014 30696
rect 17590 30504 17646 30560
rect 17590 28736 17646 28792
rect 17314 26152 17370 26208
rect 17130 23976 17186 24032
rect 16946 22888 17002 22944
rect 16486 20304 16542 20360
rect 16578 19624 16634 19680
rect 16762 19216 16818 19272
rect 17406 23432 17462 23488
rect 17406 22616 17462 22672
rect 17774 28056 17830 28112
rect 17866 27784 17922 27840
rect 17958 26832 18014 26888
rect 17866 26152 17922 26208
rect 18234 28192 18290 28248
rect 18234 27648 18290 27704
rect 17866 25472 17922 25528
rect 17590 22752 17646 22808
rect 17590 22616 17646 22672
rect 17590 22208 17646 22264
rect 16578 18828 16634 18864
rect 16578 18808 16580 18828
rect 16580 18808 16632 18828
rect 16632 18808 16634 18828
rect 15290 16768 15346 16824
rect 14922 15136 14978 15192
rect 14922 14220 14924 14240
rect 14924 14220 14976 14240
rect 14976 14220 14978 14240
rect 14922 14184 14978 14220
rect 15106 14728 15162 14784
rect 15566 16496 15622 16552
rect 16026 17992 16082 18048
rect 15842 15544 15898 15600
rect 16118 14864 16174 14920
rect 15842 13504 15898 13560
rect 15014 8492 15070 8528
rect 15014 8472 15016 8492
rect 15016 8472 15068 8492
rect 15068 8472 15070 8492
rect 15934 12416 15990 12472
rect 16026 8472 16082 8528
rect 17222 19760 17278 19816
rect 17038 15000 17094 15056
rect 17038 14592 17094 14648
rect 18602 29824 18658 29880
rect 18602 27512 18658 27568
rect 19430 33904 19486 33960
rect 20258 37712 20314 37768
rect 20626 38936 20682 38992
rect 21730 41112 21786 41168
rect 21822 40976 21878 41032
rect 21638 40568 21694 40624
rect 22006 40588 22062 40624
rect 22006 40568 22008 40588
rect 22008 40568 22060 40588
rect 22060 40568 22062 40588
rect 20258 36352 20314 36408
rect 20258 35808 20314 35864
rect 20534 35808 20590 35864
rect 20810 36796 20812 36816
rect 20812 36796 20864 36816
rect 20864 36796 20866 36816
rect 20810 36760 20866 36796
rect 20810 36624 20866 36680
rect 20074 34176 20130 34232
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19430 32000 19486 32056
rect 19706 32172 19708 32192
rect 19708 32172 19760 32192
rect 19760 32172 19762 32192
rect 19706 32136 19762 32172
rect 19706 31864 19762 31920
rect 19982 31728 20038 31784
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19798 31320 19854 31376
rect 20074 31592 20130 31648
rect 19338 31184 19394 31240
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19154 29144 19210 29200
rect 19338 29180 19340 29200
rect 19340 29180 19392 29200
rect 19392 29180 19394 29200
rect 19338 29144 19394 29180
rect 20258 32816 20314 32872
rect 20258 30504 20314 30560
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19246 28192 19302 28248
rect 18878 27240 18934 27296
rect 18786 26988 18842 27024
rect 18786 26968 18788 26988
rect 18788 26968 18840 26988
rect 18840 26968 18842 26988
rect 18510 26152 18566 26208
rect 18602 26016 18658 26072
rect 18786 26016 18842 26072
rect 18510 25472 18566 25528
rect 19522 27648 19578 27704
rect 18234 24812 18290 24848
rect 18234 24792 18236 24812
rect 18236 24792 18288 24812
rect 18288 24792 18290 24812
rect 18234 24656 18290 24712
rect 17958 22208 18014 22264
rect 17682 20032 17738 20088
rect 17958 20340 17960 20360
rect 17960 20340 18012 20360
rect 18012 20340 18014 20360
rect 17958 20304 18014 20340
rect 17774 19488 17830 19544
rect 17222 14184 17278 14240
rect 16762 13232 16818 13288
rect 17038 10920 17094 10976
rect 17406 14048 17462 14104
rect 18418 24520 18474 24576
rect 18694 24520 18750 24576
rect 18510 23976 18566 24032
rect 19890 27512 19946 27568
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19062 23704 19118 23760
rect 18694 22888 18750 22944
rect 18142 21120 18198 21176
rect 18418 22208 18474 22264
rect 18602 22208 18658 22264
rect 18142 18808 18198 18864
rect 17774 15680 17830 15736
rect 17774 14492 17776 14512
rect 17776 14492 17828 14512
rect 17828 14492 17830 14512
rect 17774 14456 17830 14492
rect 17774 14320 17830 14376
rect 17774 13796 17830 13832
rect 17774 13776 17776 13796
rect 17776 13776 17828 13796
rect 17828 13776 17830 13796
rect 18234 18672 18290 18728
rect 18142 15544 18198 15600
rect 17958 14900 17960 14920
rect 17960 14900 18012 14920
rect 18012 14900 18014 14920
rect 17958 14864 18014 14900
rect 18142 14184 18198 14240
rect 18050 13776 18106 13832
rect 18234 13640 18290 13696
rect 18418 15544 18474 15600
rect 18418 15000 18474 15056
rect 18418 14592 18474 14648
rect 18786 22752 18842 22808
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 20166 28328 20222 28384
rect 19246 22888 19302 22944
rect 19154 22616 19210 22672
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 20074 24148 20076 24168
rect 20076 24148 20128 24168
rect 20128 24148 20130 24168
rect 20074 24112 20130 24148
rect 20442 28600 20498 28656
rect 20718 34176 20774 34232
rect 20902 32680 20958 32736
rect 20902 32544 20958 32600
rect 20810 32136 20866 32192
rect 20718 31320 20774 31376
rect 20810 28736 20866 28792
rect 20718 28192 20774 28248
rect 21546 38664 21602 38720
rect 21178 37440 21234 37496
rect 21362 37032 21418 37088
rect 21270 36216 21326 36272
rect 21546 36660 21548 36680
rect 21548 36660 21600 36680
rect 21600 36660 21602 36680
rect 21546 36624 21602 36660
rect 21546 36216 21602 36272
rect 21822 38528 21878 38584
rect 21362 33652 21418 33688
rect 21362 33632 21364 33652
rect 21364 33632 21416 33652
rect 21416 33632 21418 33652
rect 21546 33496 21602 33552
rect 21546 33224 21602 33280
rect 21454 32000 21510 32056
rect 20350 24112 20406 24168
rect 19890 23588 19946 23624
rect 19890 23568 19892 23588
rect 19892 23568 19944 23588
rect 19944 23568 19946 23588
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19062 21664 19118 21720
rect 18970 20304 19026 20360
rect 19614 21972 19616 21992
rect 19616 21972 19668 21992
rect 19668 21972 19670 21992
rect 19614 21936 19670 21972
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19890 20848 19946 20904
rect 20074 22888 20130 22944
rect 20718 24656 20774 24712
rect 21086 30912 21142 30968
rect 21362 30540 21364 30560
rect 21364 30540 21416 30560
rect 21416 30540 21418 30560
rect 21362 30504 21418 30540
rect 21086 27512 21142 27568
rect 20994 27240 21050 27296
rect 21362 28484 21418 28520
rect 21362 28464 21364 28484
rect 21364 28464 21416 28484
rect 21416 28464 21418 28484
rect 21638 29688 21694 29744
rect 21546 29416 21602 29472
rect 21638 28736 21694 28792
rect 21362 27648 21418 27704
rect 21362 27548 21364 27568
rect 21364 27548 21416 27568
rect 21416 27548 21418 27568
rect 21362 27512 21418 27548
rect 20626 24248 20682 24304
rect 20442 23840 20498 23896
rect 20350 22752 20406 22808
rect 20074 22480 20130 22536
rect 20350 22480 20406 22536
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19522 20460 19578 20496
rect 19522 20440 19524 20460
rect 19524 20440 19576 20460
rect 19576 20440 19578 20460
rect 19614 20168 19670 20224
rect 18970 17312 19026 17368
rect 18602 14048 18658 14104
rect 18602 13776 18658 13832
rect 17038 8472 17094 8528
rect 15750 3984 15806 4040
rect 18878 14864 18934 14920
rect 20626 23432 20682 23488
rect 20626 23060 20628 23080
rect 20628 23060 20680 23080
rect 20680 23060 20682 23080
rect 20626 23024 20682 23060
rect 21086 26152 21142 26208
rect 21086 25744 21142 25800
rect 20902 24132 20958 24168
rect 20902 24112 20904 24132
rect 20904 24112 20956 24132
rect 20956 24112 20958 24132
rect 20810 23976 20866 24032
rect 21270 26016 21326 26072
rect 21270 25608 21326 25664
rect 21362 24792 21418 24848
rect 21178 24284 21180 24304
rect 21180 24284 21232 24304
rect 21232 24284 21234 24304
rect 21178 24248 21234 24284
rect 21086 24112 21142 24168
rect 21178 23704 21234 23760
rect 21086 23604 21088 23624
rect 21088 23604 21140 23624
rect 21140 23604 21142 23624
rect 21086 23568 21142 23604
rect 20810 23432 20866 23488
rect 20994 23160 21050 23216
rect 21086 23060 21088 23080
rect 21088 23060 21140 23080
rect 21140 23060 21142 23080
rect 21086 23024 21142 23060
rect 20626 21564 20628 21584
rect 20628 21564 20680 21584
rect 20680 21564 20682 21584
rect 20626 21528 20682 21564
rect 21086 22108 21088 22128
rect 21088 22108 21140 22128
rect 21140 22108 21142 22128
rect 21086 22072 21142 22108
rect 21086 21936 21142 21992
rect 21730 25744 21786 25800
rect 21086 21256 21142 21312
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19890 19216 19946 19272
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20166 18708 20168 18728
rect 20168 18708 20220 18728
rect 20220 18708 20222 18728
rect 20166 18672 20222 18708
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19982 16904 20038 16960
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19430 16088 19486 16144
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20534 17312 20590 17368
rect 20534 15816 20590 15872
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19522 13504 19578 13560
rect 19706 13504 19762 13560
rect 20442 14492 20444 14512
rect 20444 14492 20496 14512
rect 20496 14492 20498 14512
rect 20442 14456 20498 14492
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19522 12824 19578 12880
rect 19430 12416 19486 12472
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 20534 12008 20590 12064
rect 20350 11328 20406 11384
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 17774 4800 17830 4856
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19890 7248 19946 7304
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20442 9560 20498 9616
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 17866 3848 17922 3904
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19522 2624 19578 2680
rect 23202 41520 23258 41576
rect 21914 37984 21970 38040
rect 21914 36352 21970 36408
rect 21914 34720 21970 34776
rect 22190 39072 22246 39128
rect 22098 38392 22154 38448
rect 22466 40296 22522 40352
rect 22466 39344 22522 39400
rect 22098 37168 22154 37224
rect 22374 36896 22430 36952
rect 22374 35808 22430 35864
rect 22926 40296 22982 40352
rect 23110 40568 23166 40624
rect 22834 38664 22890 38720
rect 22650 37304 22706 37360
rect 23478 41556 23480 41576
rect 23480 41556 23532 41576
rect 23532 41556 23534 41576
rect 23478 41520 23534 41556
rect 23938 41248 23994 41304
rect 24030 40840 24086 40896
rect 23754 40704 23810 40760
rect 24122 40568 24178 40624
rect 23754 40296 23810 40352
rect 23294 38392 23350 38448
rect 23202 37712 23258 37768
rect 22834 36896 22890 36952
rect 23294 37168 23350 37224
rect 23386 37068 23388 37088
rect 23388 37068 23440 37088
rect 23440 37068 23442 37088
rect 23386 37032 23442 37068
rect 23478 36896 23534 36952
rect 23018 36624 23074 36680
rect 23754 38392 23810 38448
rect 23662 37304 23718 37360
rect 22650 35536 22706 35592
rect 22282 32172 22284 32192
rect 22284 32172 22336 32192
rect 22336 32172 22338 32192
rect 22282 32136 22338 32172
rect 22190 31320 22246 31376
rect 22558 32544 22614 32600
rect 22834 33768 22890 33824
rect 22282 29960 22338 30016
rect 22190 29824 22246 29880
rect 22190 29280 22246 29336
rect 23478 34176 23534 34232
rect 22926 33360 22982 33416
rect 22466 29708 22522 29744
rect 22466 29688 22468 29708
rect 22468 29688 22520 29708
rect 22520 29688 22522 29708
rect 22742 30368 22798 30424
rect 22834 30232 22890 30288
rect 22466 29008 22522 29064
rect 22466 28908 22468 28928
rect 22468 28908 22520 28928
rect 22520 28908 22522 28928
rect 22466 28872 22522 28908
rect 22374 27104 22430 27160
rect 22190 24384 22246 24440
rect 22006 23296 22062 23352
rect 22374 24248 22430 24304
rect 23570 34060 23626 34096
rect 23570 34040 23572 34060
rect 23572 34040 23624 34060
rect 23624 34040 23626 34060
rect 23110 30368 23166 30424
rect 22926 29824 22982 29880
rect 25042 41132 25098 41168
rect 25042 41112 25044 41132
rect 25044 41112 25096 41132
rect 25096 41112 25098 41132
rect 24490 39752 24546 39808
rect 24214 38800 24270 38856
rect 24122 37868 24178 37904
rect 24122 37848 24124 37868
rect 24124 37848 24176 37868
rect 24176 37848 24178 37868
rect 24398 37848 24454 37904
rect 24122 37712 24178 37768
rect 24306 37440 24362 37496
rect 24214 36896 24270 36952
rect 24306 36802 24362 36816
rect 24306 36760 24308 36802
rect 24308 36760 24360 36802
rect 24360 36760 24362 36802
rect 24122 34448 24178 34504
rect 24030 33496 24086 33552
rect 22834 29606 22890 29608
rect 22834 29554 22836 29606
rect 22836 29554 22888 29606
rect 22888 29554 22890 29606
rect 22834 29552 22890 29554
rect 22742 26560 22798 26616
rect 23662 32000 23718 32056
rect 23662 31864 23718 31920
rect 23754 31456 23810 31512
rect 23570 29724 23572 29744
rect 23572 29724 23624 29744
rect 23624 29724 23626 29744
rect 23570 29688 23626 29724
rect 23570 29572 23626 29608
rect 23570 29552 23572 29572
rect 23572 29552 23624 29572
rect 23624 29552 23626 29572
rect 22926 27104 22982 27160
rect 22742 24520 22798 24576
rect 20718 16632 20774 16688
rect 20902 16108 20958 16144
rect 20902 16088 20904 16108
rect 20904 16088 20956 16108
rect 20956 16088 20958 16108
rect 20902 13640 20958 13696
rect 21086 12844 21142 12880
rect 21086 12824 21088 12844
rect 21088 12824 21140 12844
rect 21140 12824 21142 12844
rect 22374 18672 22430 18728
rect 22006 16904 22062 16960
rect 21546 12416 21602 12472
rect 21178 11600 21234 11656
rect 21638 12008 21694 12064
rect 21638 11600 21694 11656
rect 21914 14612 21970 14648
rect 21914 14592 21916 14612
rect 21916 14592 21968 14612
rect 21968 14592 21970 14612
rect 21914 12144 21970 12200
rect 21822 11872 21878 11928
rect 21730 10784 21786 10840
rect 22098 15408 22154 15464
rect 22098 14592 22154 14648
rect 23570 28484 23626 28520
rect 23570 28464 23572 28484
rect 23572 28464 23624 28484
rect 23624 28464 23626 28484
rect 23386 25608 23442 25664
rect 23018 23704 23074 23760
rect 25318 40840 25374 40896
rect 25226 40568 25282 40624
rect 25134 40024 25190 40080
rect 24950 39364 25006 39400
rect 24950 39344 24952 39364
rect 24952 39344 25004 39364
rect 25004 39344 25006 39364
rect 24766 38664 24822 38720
rect 25042 39208 25098 39264
rect 25318 39480 25374 39536
rect 25318 39344 25374 39400
rect 25318 39208 25374 39264
rect 25134 38664 25190 38720
rect 25410 38664 25466 38720
rect 25042 38392 25098 38448
rect 26054 40160 26110 40216
rect 26054 39208 26110 39264
rect 24398 33516 24454 33552
rect 24398 33496 24400 33516
rect 24400 33496 24452 33516
rect 24452 33496 24454 33516
rect 24122 32816 24178 32872
rect 24306 33224 24362 33280
rect 23754 30776 23810 30832
rect 24122 30640 24178 30696
rect 24030 29552 24086 29608
rect 25318 35128 25374 35184
rect 25226 34720 25282 34776
rect 25134 33516 25190 33552
rect 25134 33496 25136 33516
rect 25136 33496 25188 33516
rect 25188 33496 25190 33516
rect 25134 32544 25190 32600
rect 25042 31864 25098 31920
rect 25042 31764 25044 31784
rect 25044 31764 25096 31784
rect 25096 31764 25098 31784
rect 24674 30776 24730 30832
rect 25042 31728 25098 31764
rect 25502 33224 25558 33280
rect 25962 37460 26018 37496
rect 25962 37440 25964 37460
rect 25964 37440 26016 37460
rect 26016 37440 26018 37460
rect 25870 35028 25872 35048
rect 25872 35028 25924 35048
rect 25924 35028 25926 35048
rect 25870 34992 25926 35028
rect 30470 41792 30526 41848
rect 26882 41132 26938 41168
rect 26882 41112 26884 41132
rect 26884 41112 26936 41132
rect 26936 41112 26938 41132
rect 26422 38528 26478 38584
rect 26974 40568 27030 40624
rect 26882 38528 26938 38584
rect 26330 36896 26386 36952
rect 26146 36216 26202 36272
rect 26054 34448 26110 34504
rect 26054 34176 26110 34232
rect 25226 32000 25282 32056
rect 25134 31340 25190 31376
rect 25134 31320 25136 31340
rect 25136 31320 25188 31340
rect 25188 31320 25190 31340
rect 24766 30504 24822 30560
rect 24398 29960 24454 30016
rect 24306 28600 24362 28656
rect 23754 24656 23810 24712
rect 23386 22752 23442 22808
rect 23110 22228 23166 22264
rect 23110 22208 23112 22228
rect 23112 22208 23164 22228
rect 23164 22208 23166 22228
rect 23478 22208 23534 22264
rect 23846 24520 23902 24576
rect 23846 22616 23902 22672
rect 24030 25472 24086 25528
rect 24490 29416 24546 29472
rect 25042 30504 25098 30560
rect 25042 29452 25044 29472
rect 25044 29452 25096 29472
rect 25096 29452 25098 29472
rect 25042 29416 25098 29452
rect 24490 27920 24546 27976
rect 24490 26832 24546 26888
rect 24214 26152 24270 26208
rect 24398 25200 24454 25256
rect 24674 24792 24730 24848
rect 24950 28736 25006 28792
rect 24950 27240 25006 27296
rect 24858 26696 24914 26752
rect 25318 30640 25374 30696
rect 25778 33260 25780 33280
rect 25780 33260 25832 33280
rect 25832 33260 25834 33280
rect 25778 33224 25834 33260
rect 26330 35264 26386 35320
rect 26238 33768 26294 33824
rect 26146 33496 26202 33552
rect 25778 31728 25834 31784
rect 25502 30232 25558 30288
rect 25226 29552 25282 29608
rect 25226 29416 25282 29472
rect 25226 29008 25282 29064
rect 24582 23568 24638 23624
rect 24122 21664 24178 21720
rect 23294 19896 23350 19952
rect 24030 20440 24086 20496
rect 23110 18300 23112 18320
rect 23112 18300 23164 18320
rect 23164 18300 23166 18320
rect 23110 18264 23166 18300
rect 22282 12280 22338 12336
rect 22282 11736 22338 11792
rect 22190 11192 22246 11248
rect 22374 11056 22430 11112
rect 22926 15816 22982 15872
rect 23386 16768 23442 16824
rect 23386 16224 23442 16280
rect 22742 14048 22798 14104
rect 22834 13932 22890 13968
rect 22834 13912 22836 13932
rect 22836 13912 22888 13932
rect 22888 13912 22890 13932
rect 23018 13640 23074 13696
rect 24214 20304 24270 20360
rect 24490 20168 24546 20224
rect 23662 15852 23664 15872
rect 23664 15852 23716 15872
rect 23716 15852 23718 15872
rect 23662 15816 23718 15852
rect 23662 15136 23718 15192
rect 24490 18400 24546 18456
rect 24858 22616 24914 22672
rect 24858 22208 24914 22264
rect 25134 24384 25190 24440
rect 25594 29552 25650 29608
rect 26330 31728 26386 31784
rect 26146 30504 26202 30560
rect 25778 26560 25834 26616
rect 25410 24520 25466 24576
rect 25502 23976 25558 24032
rect 24858 21528 24914 21584
rect 25134 19352 25190 19408
rect 23754 13676 23756 13696
rect 23756 13676 23808 13696
rect 23808 13676 23810 13696
rect 23754 13640 23810 13676
rect 24030 15272 24086 15328
rect 23202 10956 23204 10976
rect 23204 10956 23256 10976
rect 23256 10956 23258 10976
rect 23202 10920 23258 10956
rect 22742 7248 22798 7304
rect 24674 15952 24730 16008
rect 24582 15544 24638 15600
rect 25042 18128 25098 18184
rect 24950 17176 25006 17232
rect 24766 15272 24822 15328
rect 24674 15000 24730 15056
rect 24398 13932 24454 13968
rect 24398 13912 24400 13932
rect 24400 13912 24452 13932
rect 24452 13912 24454 13932
rect 24582 13268 24584 13288
rect 24584 13268 24636 13288
rect 24636 13268 24638 13288
rect 24582 13232 24638 13268
rect 25134 15136 25190 15192
rect 25134 13932 25190 13968
rect 25134 13912 25136 13932
rect 25136 13912 25188 13932
rect 25188 13912 25190 13932
rect 24858 12416 24914 12472
rect 24766 12316 24768 12336
rect 24768 12316 24820 12336
rect 24820 12316 24822 12336
rect 24766 12280 24822 12316
rect 24858 11772 24860 11792
rect 24860 11772 24912 11792
rect 24912 11772 24914 11792
rect 24858 11736 24914 11772
rect 24582 10920 24638 10976
rect 26238 28872 26294 28928
rect 26146 26968 26202 27024
rect 26054 25336 26110 25392
rect 25686 21392 25742 21448
rect 25686 16360 25742 16416
rect 24766 7792 24822 7848
rect 25226 11872 25282 11928
rect 25778 13912 25834 13968
rect 25686 11872 25742 11928
rect 25410 10648 25466 10704
rect 25686 11092 25688 11112
rect 25688 11092 25740 11112
rect 25740 11092 25742 11112
rect 26790 36116 26792 36136
rect 26792 36116 26844 36136
rect 26844 36116 26846 36136
rect 26790 36080 26846 36116
rect 26790 35692 26846 35728
rect 26974 36624 27030 36680
rect 26790 35672 26792 35692
rect 26792 35672 26844 35692
rect 26844 35672 26846 35692
rect 26606 32680 26662 32736
rect 26606 32136 26662 32192
rect 26514 31628 26516 31648
rect 26516 31628 26568 31648
rect 26568 31628 26570 31648
rect 26514 31592 26570 31628
rect 26882 33632 26938 33688
rect 26514 29300 26570 29336
rect 26514 29280 26516 29300
rect 26516 29280 26568 29300
rect 26568 29280 26570 29300
rect 26422 26968 26478 27024
rect 26514 26152 26570 26208
rect 26330 23840 26386 23896
rect 26330 23568 26386 23624
rect 26330 20848 26386 20904
rect 26330 20712 26386 20768
rect 26330 17312 26386 17368
rect 25962 14864 26018 14920
rect 26882 32816 26938 32872
rect 27250 40160 27306 40216
rect 27342 40024 27398 40080
rect 27526 40568 27582 40624
rect 28078 40976 28134 41032
rect 28170 40568 28226 40624
rect 27710 40296 27766 40352
rect 27618 38936 27674 38992
rect 27618 38528 27674 38584
rect 28354 40024 28410 40080
rect 27986 38664 28042 38720
rect 27618 37440 27674 37496
rect 27342 35536 27398 35592
rect 27618 35436 27620 35456
rect 27620 35436 27672 35456
rect 27672 35436 27674 35456
rect 27618 35400 27674 35436
rect 27618 34856 27674 34912
rect 27434 34584 27490 34640
rect 27250 34040 27306 34096
rect 27434 33360 27490 33416
rect 27526 32952 27582 33008
rect 27710 33088 27766 33144
rect 27250 32272 27306 32328
rect 27250 32000 27306 32056
rect 26882 27532 26938 27568
rect 26882 27512 26884 27532
rect 26884 27512 26936 27532
rect 26936 27512 26938 27532
rect 26974 27240 27030 27296
rect 27158 31048 27214 31104
rect 27526 32000 27582 32056
rect 27434 31864 27490 31920
rect 27342 30504 27398 30560
rect 27434 29960 27490 30016
rect 27158 28736 27214 28792
rect 27158 28600 27214 28656
rect 26974 25780 26976 25800
rect 26976 25780 27028 25800
rect 27028 25780 27030 25800
rect 26974 25744 27030 25780
rect 27986 32544 28042 32600
rect 28354 36760 28410 36816
rect 28722 39344 28778 39400
rect 28538 38936 28594 38992
rect 28814 38972 28816 38992
rect 28816 38972 28868 38992
rect 28868 38972 28870 38992
rect 28814 38936 28870 38972
rect 28814 38800 28870 38856
rect 28722 38528 28778 38584
rect 28630 37848 28686 37904
rect 28354 36080 28410 36136
rect 28354 35264 28410 35320
rect 28078 30912 28134 30968
rect 27986 29960 28042 30016
rect 27250 27104 27306 27160
rect 27526 26288 27582 26344
rect 27802 27648 27858 27704
rect 27066 24148 27068 24168
rect 27068 24148 27120 24168
rect 27120 24148 27122 24168
rect 27066 24112 27122 24148
rect 26882 23704 26938 23760
rect 28262 31048 28318 31104
rect 28262 30368 28318 30424
rect 28170 29824 28226 29880
rect 27250 24284 27252 24304
rect 27252 24284 27304 24304
rect 27304 24284 27306 24304
rect 27250 24248 27306 24284
rect 27710 24112 27766 24168
rect 28906 38664 28962 38720
rect 28998 37032 29054 37088
rect 28722 36236 28778 36272
rect 28722 36216 28724 36236
rect 28724 36216 28776 36236
rect 28776 36216 28778 36236
rect 28630 35400 28686 35456
rect 29090 36624 29146 36680
rect 28906 36352 28962 36408
rect 28538 34856 28594 34912
rect 28538 33904 28594 33960
rect 28814 35028 28816 35048
rect 28816 35028 28868 35048
rect 28868 35028 28870 35048
rect 28814 34992 28870 35028
rect 29090 34992 29146 35048
rect 28722 34720 28778 34776
rect 28538 32816 28594 32872
rect 28814 32408 28870 32464
rect 29274 34720 29330 34776
rect 30286 40724 30342 40760
rect 30286 40704 30288 40724
rect 30288 40704 30340 40724
rect 30340 40704 30342 40724
rect 29826 40024 29882 40080
rect 29734 39072 29790 39128
rect 29550 36624 29606 36680
rect 30654 40024 30710 40080
rect 30286 38528 30342 38584
rect 30562 38800 30618 38856
rect 30746 38392 30802 38448
rect 30010 37204 30012 37224
rect 30012 37204 30064 37224
rect 30064 37204 30066 37224
rect 30010 37168 30066 37204
rect 29642 35536 29698 35592
rect 29642 35264 29698 35320
rect 29274 33496 29330 33552
rect 28998 29280 29054 29336
rect 28722 26988 28778 27024
rect 28722 26968 28724 26988
rect 28724 26968 28776 26988
rect 28776 26968 28778 26988
rect 28354 26852 28410 26888
rect 28354 26832 28356 26852
rect 28356 26832 28408 26852
rect 28408 26832 28410 26852
rect 28354 26016 28410 26072
rect 26882 19760 26938 19816
rect 26514 17992 26570 18048
rect 27526 23704 27582 23760
rect 27434 23432 27490 23488
rect 27618 22344 27674 22400
rect 27526 21956 27582 21992
rect 27526 21936 27528 21956
rect 27528 21936 27580 21956
rect 27580 21936 27582 21956
rect 27894 21664 27950 21720
rect 28998 25608 29054 25664
rect 30010 34584 30066 34640
rect 30746 38120 30802 38176
rect 30378 35808 30434 35864
rect 29734 32020 29790 32056
rect 29734 32000 29736 32020
rect 29736 32000 29788 32020
rect 29788 32000 29790 32020
rect 30470 35400 30526 35456
rect 30378 34892 30380 34912
rect 30380 34892 30432 34912
rect 30432 34892 30434 34912
rect 30378 34856 30434 34892
rect 30286 34740 30342 34776
rect 30286 34720 30288 34740
rect 30288 34720 30340 34740
rect 30340 34720 30342 34740
rect 29366 30812 29368 30832
rect 29368 30812 29420 30832
rect 29420 30812 29422 30832
rect 29366 30776 29422 30812
rect 29642 30796 29698 30832
rect 29642 30776 29644 30796
rect 29644 30776 29696 30796
rect 29696 30776 29698 30796
rect 29182 25472 29238 25528
rect 29090 25336 29146 25392
rect 29274 25200 29330 25256
rect 29090 25064 29146 25120
rect 29274 24792 29330 24848
rect 27526 18400 27582 18456
rect 27158 16360 27214 16416
rect 26790 13504 26846 13560
rect 26698 13268 26700 13288
rect 26700 13268 26752 13288
rect 26752 13268 26754 13288
rect 26698 13232 26754 13268
rect 26514 11756 26570 11792
rect 26514 11736 26516 11756
rect 26516 11736 26568 11756
rect 26568 11736 26570 11756
rect 25962 11328 26018 11384
rect 25686 11056 25742 11092
rect 25962 11092 25964 11112
rect 25964 11092 26016 11112
rect 26016 11092 26018 11112
rect 25594 9560 25650 9616
rect 25962 11056 26018 11092
rect 25870 9444 25926 9480
rect 25870 9424 25872 9444
rect 25872 9424 25924 9444
rect 25924 9424 25926 9444
rect 26422 11192 26478 11248
rect 26238 10920 26294 10976
rect 26514 10920 26570 10976
rect 27342 14456 27398 14512
rect 26882 11500 26884 11520
rect 26884 11500 26936 11520
rect 26936 11500 26938 11520
rect 26882 11464 26938 11500
rect 26974 10648 27030 10704
rect 27710 16224 27766 16280
rect 27710 14320 27766 14376
rect 28170 16088 28226 16144
rect 28170 15136 28226 15192
rect 28170 14048 28226 14104
rect 26606 9424 26662 9480
rect 25870 7792 25926 7848
rect 25962 5208 26018 5264
rect 29642 30232 29698 30288
rect 29826 29044 29828 29064
rect 29828 29044 29880 29064
rect 29880 29044 29882 29064
rect 29826 29008 29882 29044
rect 29642 28872 29698 28928
rect 29550 21004 29606 21040
rect 29550 20984 29552 21004
rect 29552 20984 29604 21004
rect 29604 20984 29606 21004
rect 30010 26424 30066 26480
rect 29734 25608 29790 25664
rect 31022 38972 31024 38992
rect 31024 38972 31076 38992
rect 31076 38972 31078 38992
rect 31022 38936 31078 38972
rect 30930 35400 30986 35456
rect 30654 35264 30710 35320
rect 30654 34856 30710 34912
rect 30838 34584 30894 34640
rect 30562 34448 30618 34504
rect 30930 31628 30932 31648
rect 30932 31628 30984 31648
rect 30984 31628 30986 31648
rect 30930 31592 30986 31628
rect 32310 39888 32366 39944
rect 31758 38800 31814 38856
rect 31574 37188 31630 37224
rect 31574 37168 31576 37188
rect 31576 37168 31628 37188
rect 31628 37168 31630 37188
rect 31114 35692 31170 35728
rect 31114 35672 31116 35692
rect 31116 35672 31168 35692
rect 31168 35672 31170 35692
rect 31298 35128 31354 35184
rect 31114 35028 31116 35048
rect 31116 35028 31168 35048
rect 31168 35028 31170 35048
rect 31114 34992 31170 35028
rect 31666 35944 31722 36000
rect 30562 29416 30618 29472
rect 30378 25900 30434 25936
rect 30378 25880 30380 25900
rect 30380 25880 30432 25900
rect 30432 25880 30434 25900
rect 30930 29572 30986 29608
rect 30930 29552 30932 29572
rect 30932 29552 30984 29572
rect 30984 29552 30986 29572
rect 31022 28736 31078 28792
rect 31574 28464 31630 28520
rect 32402 38956 32458 38992
rect 32402 38936 32404 38956
rect 32404 38936 32456 38956
rect 32456 38936 32458 38956
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 32586 36488 32642 36544
rect 31758 34856 31814 34912
rect 31758 34448 31814 34504
rect 32034 35028 32036 35048
rect 32036 35028 32088 35048
rect 32088 35028 32090 35048
rect 32034 34992 32090 35028
rect 31758 29008 31814 29064
rect 30930 25900 30986 25936
rect 30930 25880 30932 25900
rect 30932 25880 30984 25900
rect 30984 25880 30986 25900
rect 30562 24248 30618 24304
rect 30286 22888 30342 22944
rect 30930 24656 30986 24712
rect 29090 16124 29092 16144
rect 29092 16124 29144 16144
rect 29144 16124 29146 16144
rect 29090 16088 29146 16124
rect 29366 16224 29422 16280
rect 29458 15680 29514 15736
rect 29826 16224 29882 16280
rect 29642 16088 29698 16144
rect 30562 21800 30618 21856
rect 29734 14728 29790 14784
rect 28998 13640 29054 13696
rect 28906 12280 28962 12336
rect 31942 27956 31944 27976
rect 31944 27956 31996 27976
rect 31996 27956 31998 27976
rect 31942 27920 31998 27956
rect 32586 29280 32642 29336
rect 31758 24248 31814 24304
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35162 28076 35218 28112
rect 35162 28056 35164 28076
rect 35164 28056 35216 28076
rect 35216 28056 35218 28076
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35530 25900 35586 25936
rect 35530 25880 35532 25900
rect 35532 25880 35584 25900
rect 35584 25880 35586 25900
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 36542 29144 36598 29200
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 31390 20032 31446 20088
rect 32218 20460 32274 20496
rect 32218 20440 32220 20460
rect 32220 20440 32272 20460
rect 32272 20440 32274 20460
rect 31114 17584 31170 17640
rect 30010 14048 30066 14104
rect 30838 14048 30894 14104
rect 31942 18672 31998 18728
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 33966 20304 34022 20360
rect 35254 20576 35310 20632
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35346 19796 35348 19816
rect 35348 19796 35400 19816
rect 35400 19796 35402 19816
rect 33138 18808 33194 18864
rect 35346 19760 35402 19796
rect 33782 18708 33784 18728
rect 33784 18708 33836 18728
rect 33836 18708 33838 18728
rect 33782 18672 33838 18708
rect 32770 15952 32826 16008
rect 33598 16652 33654 16688
rect 33598 16632 33600 16652
rect 33600 16632 33652 16652
rect 33652 16632 33654 16652
rect 33506 16496 33562 16552
rect 33230 14320 33286 14376
rect 34150 16496 34206 16552
rect 34242 14048 34298 14104
rect 34426 13268 34428 13288
rect 34428 13268 34480 13288
rect 34480 13268 34482 13288
rect 34426 13232 34482 13268
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34886 13932 34942 13968
rect 34886 13912 34888 13932
rect 34888 13912 34940 13932
rect 34940 13912 34942 13932
rect 35622 13912 35678 13968
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35806 20440 35862 20496
rect 41234 40840 41290 40896
rect 40774 40432 40830 40488
rect 40958 36760 41014 36816
rect 40958 32716 40960 32736
rect 40960 32716 41012 32736
rect 41012 32716 41014 32736
rect 40958 32680 41014 32716
rect 40958 30096 41014 30152
rect 41326 28600 41382 28656
rect 36358 20576 36414 20632
rect 36542 20460 36598 20496
rect 36542 20440 36544 20460
rect 36544 20440 36596 20460
rect 36596 20440 36598 20460
rect 36450 20304 36506 20360
rect 41326 24520 41382 24576
rect 41050 22616 41106 22672
rect 36358 17604 36414 17640
rect 36358 17584 36360 17604
rect 36360 17584 36412 17604
rect 36412 17584 36414 17604
rect 36542 15408 36598 15464
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34794 12008 34850 12064
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35898 13268 35900 13288
rect 35900 13268 35952 13288
rect 35952 13268 35954 13288
rect 35898 13232 35954 13268
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 38658 16668 38660 16688
rect 38660 16668 38712 16688
rect 38712 16668 38714 16688
rect 38658 16632 38714 16668
rect 38658 16532 38660 16552
rect 38660 16532 38712 16552
rect 38712 16532 38714 16552
rect 38658 16496 38714 16532
rect 41510 20440 41566 20496
rect 38842 14320 38898 14376
rect 39578 16652 39634 16688
rect 39578 16632 39580 16652
rect 39580 16632 39632 16652
rect 39632 16632 39634 16652
rect 39394 16532 39396 16552
rect 39396 16532 39448 16552
rect 39448 16532 39450 16552
rect 39394 16496 39450 16532
rect 40498 14340 40554 14376
rect 40498 14320 40500 14340
rect 40500 14320 40552 14340
rect 40552 14320 40554 14340
rect 39854 12280 39910 12336
rect 41510 16360 41566 16416
rect 41050 8200 41106 8256
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 41050 4120 41106 4176
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 39946 40 40002 96
<< metal3 >>
rect 0 44298 800 44328
rect 2773 44298 2839 44301
rect 0 44296 2839 44298
rect 0 44240 2778 44296
rect 2834 44240 2839 44296
rect 0 44238 2839 44240
rect 0 44208 800 44238
rect 2773 44235 2839 44238
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 14641 41850 14707 41853
rect 19425 41852 19491 41853
rect 14774 41850 14780 41852
rect 14641 41848 14780 41850
rect 14641 41792 14646 41848
rect 14702 41792 14780 41848
rect 14641 41790 14780 41792
rect 14641 41787 14707 41790
rect 14774 41788 14780 41790
rect 14844 41788 14850 41852
rect 19374 41850 19380 41852
rect 19334 41790 19380 41850
rect 19444 41848 19491 41852
rect 19486 41792 19491 41848
rect 19374 41788 19380 41790
rect 19444 41788 19491 41792
rect 19425 41787 19491 41788
rect 30465 41850 30531 41853
rect 30598 41850 30604 41852
rect 30465 41848 30604 41850
rect 30465 41792 30470 41848
rect 30526 41792 30604 41848
rect 30465 41790 30604 41792
rect 30465 41787 30531 41790
rect 30598 41788 30604 41790
rect 30668 41788 30674 41852
rect 18965 41714 19031 41717
rect 20713 41716 20779 41717
rect 20662 41714 20668 41716
rect 18965 41712 20668 41714
rect 20732 41714 20779 41716
rect 20732 41712 20860 41714
rect 18965 41656 18970 41712
rect 19026 41656 20668 41712
rect 20774 41656 20860 41712
rect 18965 41654 20668 41656
rect 18965 41651 19031 41654
rect 20662 41652 20668 41654
rect 20732 41654 20860 41656
rect 20732 41652 20779 41654
rect 20713 41651 20779 41652
rect 23197 41578 23263 41581
rect 19290 41576 23263 41578
rect 19290 41520 23202 41576
rect 23258 41520 23263 41576
rect 19290 41518 23263 41520
rect 10542 41380 10548 41444
rect 10612 41442 10618 41444
rect 10869 41442 10935 41445
rect 10612 41440 10935 41442
rect 10612 41384 10874 41440
rect 10930 41384 10935 41440
rect 10612 41382 10935 41384
rect 10612 41380 10618 41382
rect 10869 41379 10935 41382
rect 18413 41170 18479 41173
rect 19290 41170 19350 41518
rect 23197 41515 23263 41518
rect 23473 41578 23539 41581
rect 23606 41578 23612 41580
rect 23473 41576 23612 41578
rect 23473 41520 23478 41576
rect 23534 41520 23612 41576
rect 23473 41518 23612 41520
rect 23473 41515 23539 41518
rect 23606 41516 23612 41518
rect 23676 41516 23682 41580
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 20161 41308 20227 41309
rect 20110 41306 20116 41308
rect 20070 41246 20116 41306
rect 20180 41304 20227 41308
rect 20222 41248 20227 41304
rect 20110 41244 20116 41246
rect 20180 41244 20227 41248
rect 20161 41243 20227 41244
rect 21633 41306 21699 41309
rect 23933 41306 23999 41309
rect 21633 41304 23999 41306
rect 21633 41248 21638 41304
rect 21694 41248 23938 41304
rect 23994 41248 23999 41304
rect 21633 41246 23999 41248
rect 21633 41243 21699 41246
rect 23933 41243 23999 41246
rect 18413 41168 19350 41170
rect 18413 41112 18418 41168
rect 18474 41112 19350 41168
rect 18413 41110 19350 41112
rect 21725 41170 21791 41173
rect 25037 41170 25103 41173
rect 26877 41170 26943 41173
rect 21725 41168 22248 41170
rect 21725 41112 21730 41168
rect 21786 41112 22248 41168
rect 21725 41110 22248 41112
rect 18413 41107 18479 41110
rect 21725 41107 21791 41110
rect 12801 41034 12867 41037
rect 16205 41034 16271 41037
rect 12801 41032 16271 41034
rect 12801 40976 12806 41032
rect 12862 40976 16210 41032
rect 16266 40976 16271 41032
rect 12801 40974 16271 40976
rect 12801 40971 12867 40974
rect 16205 40971 16271 40974
rect 17125 41034 17191 41037
rect 18045 41034 18111 41037
rect 18873 41034 18939 41037
rect 21817 41034 21883 41037
rect 17125 41032 21883 41034
rect 17125 40976 17130 41032
rect 17186 40976 18050 41032
rect 18106 40976 18878 41032
rect 18934 40976 21822 41032
rect 21878 40976 21883 41032
rect 17125 40974 21883 40976
rect 22188 41034 22248 41110
rect 25037 41168 26943 41170
rect 25037 41112 25042 41168
rect 25098 41112 26882 41168
rect 26938 41112 26943 41168
rect 25037 41110 26943 41112
rect 25037 41107 25103 41110
rect 26877 41107 26943 41110
rect 28073 41034 28139 41037
rect 22188 41032 28139 41034
rect 22188 40976 28078 41032
rect 28134 40976 28139 41032
rect 22188 40974 28139 40976
rect 17125 40971 17191 40974
rect 18045 40971 18111 40974
rect 18873 40971 18939 40974
rect 21817 40971 21883 40974
rect 28073 40971 28139 40974
rect 17217 40898 17283 40901
rect 19241 40898 19307 40901
rect 24025 40898 24091 40901
rect 17217 40896 24091 40898
rect 17217 40840 17222 40896
rect 17278 40840 19246 40896
rect 19302 40840 24030 40896
rect 24086 40840 24091 40896
rect 17217 40838 24091 40840
rect 17217 40835 17283 40838
rect 19241 40835 19307 40838
rect 24025 40835 24091 40838
rect 24894 40836 24900 40900
rect 24964 40898 24970 40900
rect 25313 40898 25379 40901
rect 24964 40896 25379 40898
rect 24964 40840 25318 40896
rect 25374 40840 25379 40896
rect 24964 40838 25379 40840
rect 24964 40836 24970 40838
rect 25313 40835 25379 40838
rect 41229 40898 41295 40901
rect 41720 40898 42520 40928
rect 41229 40896 42520 40898
rect 41229 40840 41234 40896
rect 41290 40840 42520 40896
rect 41229 40838 42520 40840
rect 41229 40835 41295 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 41720 40808 42520 40838
rect 34930 40767 35246 40768
rect 16573 40762 16639 40765
rect 23749 40762 23815 40765
rect 30281 40762 30347 40765
rect 16573 40760 23674 40762
rect 16573 40704 16578 40760
rect 16634 40704 23674 40760
rect 16573 40702 23674 40704
rect 16573 40699 16639 40702
rect 18597 40626 18663 40629
rect 21633 40626 21699 40629
rect 18597 40624 21699 40626
rect 18597 40568 18602 40624
rect 18658 40568 21638 40624
rect 21694 40568 21699 40624
rect 18597 40566 21699 40568
rect 18597 40563 18663 40566
rect 21633 40563 21699 40566
rect 22001 40626 22067 40629
rect 23105 40626 23171 40629
rect 22001 40624 23171 40626
rect 22001 40568 22006 40624
rect 22062 40568 23110 40624
rect 23166 40568 23171 40624
rect 22001 40566 23171 40568
rect 23614 40626 23674 40702
rect 23749 40760 30347 40762
rect 23749 40704 23754 40760
rect 23810 40704 30286 40760
rect 30342 40704 30347 40760
rect 23749 40702 30347 40704
rect 23749 40699 23815 40702
rect 30281 40699 30347 40702
rect 24117 40626 24183 40629
rect 23614 40624 24183 40626
rect 23614 40568 24122 40624
rect 24178 40568 24183 40624
rect 23614 40566 24183 40568
rect 22001 40563 22067 40566
rect 23105 40563 23171 40566
rect 24117 40563 24183 40566
rect 25221 40626 25287 40629
rect 26969 40626 27035 40629
rect 27521 40626 27587 40629
rect 28165 40626 28231 40629
rect 25221 40624 28231 40626
rect 25221 40568 25226 40624
rect 25282 40568 26974 40624
rect 27030 40568 27526 40624
rect 27582 40568 28170 40624
rect 28226 40568 28231 40624
rect 25221 40566 28231 40568
rect 25221 40563 25287 40566
rect 26969 40563 27035 40566
rect 27521 40563 27587 40566
rect 28165 40563 28231 40566
rect 16021 40490 16087 40493
rect 18137 40490 18203 40493
rect 40769 40490 40835 40493
rect 16021 40488 40835 40490
rect 16021 40432 16026 40488
rect 16082 40432 18142 40488
rect 18198 40432 40774 40488
rect 40830 40432 40835 40488
rect 16021 40430 40835 40432
rect 16021 40427 16087 40430
rect 18137 40427 18203 40430
rect 40769 40427 40835 40430
rect 16481 40354 16547 40357
rect 18597 40354 18663 40357
rect 16481 40352 18663 40354
rect 16481 40296 16486 40352
rect 16542 40296 18602 40352
rect 18658 40296 18663 40352
rect 16481 40294 18663 40296
rect 16481 40291 16547 40294
rect 18597 40291 18663 40294
rect 19333 40356 19399 40357
rect 19333 40352 19380 40356
rect 19444 40354 19450 40356
rect 19977 40354 20043 40357
rect 22461 40354 22527 40357
rect 19333 40296 19338 40352
rect 19333 40292 19380 40296
rect 19444 40294 19490 40354
rect 19977 40352 22527 40354
rect 19977 40296 19982 40352
rect 20038 40296 22466 40352
rect 22522 40296 22527 40352
rect 19977 40294 22527 40296
rect 19444 40292 19450 40294
rect 19333 40291 19399 40292
rect 19977 40291 20043 40294
rect 22461 40291 22527 40294
rect 22921 40354 22987 40357
rect 23749 40354 23815 40357
rect 27705 40354 27771 40357
rect 22921 40352 27771 40354
rect 22921 40296 22926 40352
rect 22982 40296 23754 40352
rect 23810 40296 27710 40352
rect 27766 40296 27771 40352
rect 22921 40294 27771 40296
rect 22921 40291 22987 40294
rect 23749 40291 23815 40294
rect 27705 40291 27771 40294
rect 19570 40288 19886 40289
rect 0 40218 800 40248
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 933 40218 999 40221
rect 0 40216 999 40218
rect 0 40160 938 40216
rect 994 40160 999 40216
rect 0 40158 999 40160
rect 0 40128 800 40158
rect 933 40155 999 40158
rect 15101 40218 15167 40221
rect 16757 40218 16823 40221
rect 20161 40220 20227 40221
rect 15101 40216 18706 40218
rect 15101 40160 15106 40216
rect 15162 40160 16762 40216
rect 16818 40160 18706 40216
rect 15101 40158 18706 40160
rect 15101 40155 15167 40158
rect 16757 40155 16823 40158
rect 10961 40082 11027 40085
rect 15101 40082 15167 40085
rect 10961 40080 15167 40082
rect 10961 40024 10966 40080
rect 11022 40024 15106 40080
rect 15162 40024 15167 40080
rect 10961 40022 15167 40024
rect 10961 40019 11027 40022
rect 15101 40019 15167 40022
rect 16941 40082 17007 40085
rect 17677 40082 17743 40085
rect 18413 40084 18479 40085
rect 18413 40082 18460 40084
rect 16941 40080 17743 40082
rect 16941 40024 16946 40080
rect 17002 40024 17682 40080
rect 17738 40024 17743 40080
rect 16941 40022 17743 40024
rect 18368 40080 18460 40082
rect 18368 40024 18418 40080
rect 18368 40022 18460 40024
rect 16941 40019 17007 40022
rect 17677 40019 17743 40022
rect 18413 40020 18460 40022
rect 18524 40020 18530 40084
rect 18646 40082 18706 40158
rect 20110 40156 20116 40220
rect 20180 40218 20227 40220
rect 26049 40218 26115 40221
rect 27245 40220 27311 40221
rect 26182 40218 26188 40220
rect 20180 40216 20272 40218
rect 20222 40160 20272 40216
rect 20180 40158 20272 40160
rect 26049 40216 26188 40218
rect 26049 40160 26054 40216
rect 26110 40160 26188 40216
rect 26049 40158 26188 40160
rect 20180 40156 20227 40158
rect 20161 40155 20227 40156
rect 26049 40155 26115 40158
rect 26182 40156 26188 40158
rect 26252 40156 26258 40220
rect 27245 40216 27292 40220
rect 27356 40218 27362 40220
rect 27245 40160 27250 40216
rect 27245 40156 27292 40160
rect 27356 40158 27402 40218
rect 27356 40156 27362 40158
rect 27245 40155 27311 40156
rect 25129 40082 25195 40085
rect 18646 40080 25195 40082
rect 18646 40024 25134 40080
rect 25190 40024 25195 40080
rect 18646 40022 25195 40024
rect 18413 40019 18479 40020
rect 25129 40019 25195 40022
rect 27337 40082 27403 40085
rect 28349 40084 28415 40085
rect 27337 40080 27538 40082
rect 27337 40024 27342 40080
rect 27398 40024 27538 40080
rect 27337 40022 27538 40024
rect 27337 40019 27403 40022
rect 27478 39946 27538 40022
rect 28349 40080 28396 40084
rect 28460 40082 28466 40084
rect 28349 40024 28354 40080
rect 28349 40020 28396 40024
rect 28460 40022 28506 40082
rect 28460 40020 28466 40022
rect 29678 40020 29684 40084
rect 29748 40082 29754 40084
rect 29821 40082 29887 40085
rect 29748 40080 29887 40082
rect 29748 40024 29826 40080
rect 29882 40024 29887 40080
rect 29748 40022 29887 40024
rect 29748 40020 29754 40022
rect 28349 40019 28415 40020
rect 29821 40019 29887 40022
rect 30649 40082 30715 40085
rect 31150 40082 31156 40084
rect 30649 40080 31156 40082
rect 30649 40024 30654 40080
rect 30710 40024 31156 40080
rect 30649 40022 31156 40024
rect 30649 40019 30715 40022
rect 31150 40020 31156 40022
rect 31220 40020 31226 40084
rect 32305 39946 32371 39949
rect 27478 39944 32371 39946
rect 27478 39888 32310 39944
rect 32366 39888 32371 39944
rect 27478 39886 32371 39888
rect 32305 39883 32371 39886
rect 19793 39810 19859 39813
rect 24485 39810 24551 39813
rect 19793 39808 24551 39810
rect 19793 39752 19798 39808
rect 19854 39752 24490 39808
rect 24546 39752 24551 39808
rect 19793 39750 24551 39752
rect 19793 39747 19859 39750
rect 24485 39747 24551 39750
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 25313 39540 25379 39541
rect 25262 39538 25268 39540
rect 25222 39478 25268 39538
rect 25332 39536 25379 39540
rect 25374 39480 25379 39536
rect 25262 39476 25268 39478
rect 25332 39476 25379 39480
rect 25313 39475 25379 39476
rect 18597 39402 18663 39405
rect 19149 39402 19215 39405
rect 18597 39400 19215 39402
rect 18597 39344 18602 39400
rect 18658 39344 19154 39400
rect 19210 39344 19215 39400
rect 18597 39342 19215 39344
rect 18597 39339 18663 39342
rect 19149 39339 19215 39342
rect 22461 39402 22527 39405
rect 24945 39402 25011 39405
rect 22461 39400 25011 39402
rect 22461 39344 22466 39400
rect 22522 39344 24950 39400
rect 25006 39344 25011 39400
rect 22461 39342 25011 39344
rect 22461 39339 22527 39342
rect 24945 39339 25011 39342
rect 25313 39400 25379 39405
rect 25313 39344 25318 39400
rect 25374 39344 25379 39400
rect 25313 39339 25379 39344
rect 27102 39340 27108 39404
rect 27172 39402 27178 39404
rect 28717 39402 28783 39405
rect 27172 39400 28783 39402
rect 27172 39344 28722 39400
rect 28778 39344 28783 39400
rect 27172 39342 28783 39344
rect 27172 39340 27178 39342
rect 28717 39339 28783 39342
rect 25316 39269 25376 39339
rect 17953 39266 18019 39269
rect 18965 39266 19031 39269
rect 17953 39264 19031 39266
rect 17953 39208 17958 39264
rect 18014 39208 18970 39264
rect 19026 39208 19031 39264
rect 17953 39206 19031 39208
rect 17953 39203 18019 39206
rect 18965 39203 19031 39206
rect 24342 39204 24348 39268
rect 24412 39266 24418 39268
rect 25037 39266 25103 39269
rect 24412 39264 25103 39266
rect 24412 39208 25042 39264
rect 25098 39208 25103 39264
rect 24412 39206 25103 39208
rect 24412 39204 24418 39206
rect 25037 39203 25103 39206
rect 25313 39264 25379 39269
rect 26049 39268 26115 39269
rect 25998 39266 26004 39268
rect 25313 39208 25318 39264
rect 25374 39208 25379 39264
rect 25313 39203 25379 39208
rect 25958 39206 26004 39266
rect 26068 39264 26115 39268
rect 26110 39208 26115 39264
rect 25998 39204 26004 39206
rect 26068 39204 26115 39208
rect 26049 39203 26115 39204
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 13353 39130 13419 39133
rect 18321 39130 18387 39133
rect 13353 39128 18387 39130
rect 13353 39072 13358 39128
rect 13414 39072 18326 39128
rect 18382 39072 18387 39128
rect 13353 39070 18387 39072
rect 13353 39067 13419 39070
rect 18321 39067 18387 39070
rect 22185 39130 22251 39133
rect 29729 39130 29795 39133
rect 22185 39128 29795 39130
rect 22185 39072 22190 39128
rect 22246 39072 29734 39128
rect 29790 39072 29795 39128
rect 22185 39070 29795 39072
rect 22185 39067 22251 39070
rect 29729 39067 29795 39070
rect 20621 38994 20687 38997
rect 27613 38994 27679 38997
rect 20621 38992 27679 38994
rect 20621 38936 20626 38992
rect 20682 38936 27618 38992
rect 27674 38936 27679 38992
rect 20621 38934 27679 38936
rect 20621 38931 20687 38934
rect 27613 38931 27679 38934
rect 28533 38994 28599 38997
rect 28809 38994 28875 38997
rect 28533 38992 28875 38994
rect 28533 38936 28538 38992
rect 28594 38936 28814 38992
rect 28870 38936 28875 38992
rect 28533 38934 28875 38936
rect 28533 38931 28599 38934
rect 28809 38931 28875 38934
rect 31017 38994 31083 38997
rect 32397 38994 32463 38997
rect 31017 38992 32463 38994
rect 31017 38936 31022 38992
rect 31078 38936 32402 38992
rect 32458 38936 32463 38992
rect 31017 38934 32463 38936
rect 31017 38931 31083 38934
rect 32397 38931 32463 38934
rect 23422 38796 23428 38860
rect 23492 38858 23498 38860
rect 24209 38858 24275 38861
rect 23492 38856 24275 38858
rect 23492 38800 24214 38856
rect 24270 38800 24275 38856
rect 23492 38798 24275 38800
rect 23492 38796 23498 38798
rect 24209 38795 24275 38798
rect 28809 38858 28875 38861
rect 30557 38858 30623 38861
rect 31753 38858 31819 38861
rect 28809 38856 29010 38858
rect 28809 38800 28814 38856
rect 28870 38800 29010 38856
rect 28809 38798 29010 38800
rect 28809 38795 28875 38798
rect 28950 38725 29010 38798
rect 30557 38856 31819 38858
rect 30557 38800 30562 38856
rect 30618 38800 31758 38856
rect 31814 38800 31819 38856
rect 30557 38798 31819 38800
rect 30557 38795 30623 38798
rect 31753 38795 31819 38798
rect 21541 38722 21607 38725
rect 22829 38722 22895 38725
rect 24761 38722 24827 38725
rect 25129 38722 25195 38725
rect 21541 38720 25195 38722
rect 21541 38664 21546 38720
rect 21602 38664 22834 38720
rect 22890 38664 24766 38720
rect 24822 38664 25134 38720
rect 25190 38664 25195 38720
rect 21541 38662 25195 38664
rect 21541 38659 21607 38662
rect 22829 38659 22895 38662
rect 24761 38659 24827 38662
rect 25129 38659 25195 38662
rect 25262 38660 25268 38724
rect 25332 38722 25338 38724
rect 25405 38722 25471 38725
rect 25332 38720 25471 38722
rect 25332 38664 25410 38720
rect 25466 38664 25471 38720
rect 25332 38662 25471 38664
rect 25332 38660 25338 38662
rect 25405 38659 25471 38662
rect 27981 38724 28047 38725
rect 27981 38720 28028 38724
rect 28092 38722 28098 38724
rect 27981 38664 27986 38720
rect 27981 38660 28028 38664
rect 28092 38662 28138 38722
rect 28901 38720 29010 38725
rect 28901 38664 28906 38720
rect 28962 38664 29010 38720
rect 28901 38662 29010 38664
rect 28092 38660 28098 38662
rect 27981 38659 28047 38660
rect 28901 38659 28967 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 21817 38586 21883 38589
rect 26417 38586 26483 38589
rect 21817 38584 26483 38586
rect 21817 38528 21822 38584
rect 21878 38528 26422 38584
rect 26478 38528 26483 38584
rect 21817 38526 26483 38528
rect 21817 38523 21883 38526
rect 26417 38523 26483 38526
rect 26877 38586 26943 38589
rect 27613 38586 27679 38589
rect 26877 38584 27679 38586
rect 26877 38528 26882 38584
rect 26938 38528 27618 38584
rect 27674 38528 27679 38584
rect 26877 38526 27679 38528
rect 26877 38523 26943 38526
rect 27613 38523 27679 38526
rect 28717 38586 28783 38589
rect 30281 38586 30347 38589
rect 28717 38584 30347 38586
rect 28717 38528 28722 38584
rect 28778 38528 30286 38584
rect 30342 38528 30347 38584
rect 28717 38526 30347 38528
rect 28717 38523 28783 38526
rect 30281 38523 30347 38526
rect 22093 38450 22159 38453
rect 23289 38450 23355 38453
rect 22093 38448 23355 38450
rect 22093 38392 22098 38448
rect 22154 38392 23294 38448
rect 23350 38392 23355 38448
rect 22093 38390 23355 38392
rect 22093 38387 22159 38390
rect 23289 38387 23355 38390
rect 23749 38450 23815 38453
rect 25037 38450 25103 38453
rect 23749 38448 25103 38450
rect 23749 38392 23754 38448
rect 23810 38392 25042 38448
rect 25098 38392 25103 38448
rect 23749 38390 25103 38392
rect 23749 38387 23815 38390
rect 25037 38387 25103 38390
rect 30741 38448 30807 38453
rect 30741 38392 30746 38448
rect 30802 38392 30807 38448
rect 30741 38387 30807 38392
rect 30744 38181 30804 38387
rect 30741 38176 30807 38181
rect 30741 38120 30746 38176
rect 30802 38120 30807 38176
rect 30741 38115 30807 38120
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 14273 38042 14339 38045
rect 16113 38042 16179 38045
rect 14273 38040 16179 38042
rect 14273 37984 14278 38040
rect 14334 37984 16118 38040
rect 16174 37984 16179 38040
rect 14273 37982 16179 37984
rect 14273 37979 14339 37982
rect 16113 37979 16179 37982
rect 21909 38042 21975 38045
rect 29494 38042 29500 38044
rect 21909 38040 29500 38042
rect 21909 37984 21914 38040
rect 21970 37984 29500 38040
rect 21909 37982 29500 37984
rect 21909 37979 21975 37982
rect 29494 37980 29500 37982
rect 29564 37980 29570 38044
rect 24117 37908 24183 37909
rect 24117 37904 24164 37908
rect 24228 37906 24234 37908
rect 24393 37906 24459 37909
rect 28625 37906 28691 37909
rect 24117 37848 24122 37904
rect 24117 37844 24164 37848
rect 24228 37846 24274 37906
rect 24393 37904 28691 37906
rect 24393 37848 24398 37904
rect 24454 37848 28630 37904
rect 28686 37848 28691 37904
rect 24393 37846 28691 37848
rect 24228 37844 24234 37846
rect 24117 37843 24183 37844
rect 24393 37843 24459 37846
rect 28625 37843 28691 37846
rect 20253 37770 20319 37773
rect 23197 37770 23263 37773
rect 20253 37768 23263 37770
rect 20253 37712 20258 37768
rect 20314 37712 23202 37768
rect 23258 37712 23263 37768
rect 20253 37710 23263 37712
rect 20253 37707 20319 37710
rect 23197 37707 23263 37710
rect 23606 37708 23612 37772
rect 23676 37770 23682 37772
rect 24117 37770 24183 37773
rect 23676 37768 24183 37770
rect 23676 37712 24122 37768
rect 24178 37712 24183 37768
rect 23676 37710 24183 37712
rect 23676 37708 23682 37710
rect 24117 37707 24183 37710
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 21173 37498 21239 37501
rect 24301 37498 24367 37501
rect 21173 37496 24367 37498
rect 21173 37440 21178 37496
rect 21234 37440 24306 37496
rect 24362 37440 24367 37496
rect 21173 37438 24367 37440
rect 21173 37435 21239 37438
rect 24301 37435 24367 37438
rect 25957 37498 26023 37501
rect 27613 37498 27679 37501
rect 25957 37496 27679 37498
rect 25957 37440 25962 37496
rect 26018 37440 27618 37496
rect 27674 37440 27679 37496
rect 25957 37438 27679 37440
rect 25957 37435 26023 37438
rect 27613 37435 27679 37438
rect 10910 37300 10916 37364
rect 10980 37362 10986 37364
rect 15285 37362 15351 37365
rect 16113 37362 16179 37365
rect 10980 37360 16179 37362
rect 10980 37304 15290 37360
rect 15346 37304 16118 37360
rect 16174 37304 16179 37360
rect 10980 37302 16179 37304
rect 10980 37300 10986 37302
rect 15285 37299 15351 37302
rect 16113 37299 16179 37302
rect 22645 37362 22711 37365
rect 23657 37362 23723 37365
rect 22645 37360 23723 37362
rect 22645 37304 22650 37360
rect 22706 37304 23662 37360
rect 23718 37304 23723 37360
rect 22645 37302 23723 37304
rect 22645 37299 22711 37302
rect 23657 37299 23723 37302
rect 22093 37226 22159 37229
rect 23289 37226 23355 37229
rect 22093 37224 23355 37226
rect 22093 37168 22098 37224
rect 22154 37168 23294 37224
rect 23350 37168 23355 37224
rect 22093 37166 23355 37168
rect 22093 37163 22159 37166
rect 23289 37163 23355 37166
rect 30005 37226 30071 37229
rect 31569 37226 31635 37229
rect 30005 37224 31635 37226
rect 30005 37168 30010 37224
rect 30066 37168 31574 37224
rect 31630 37168 31635 37224
rect 30005 37166 31635 37168
rect 30005 37163 30071 37166
rect 31569 37163 31635 37166
rect 10777 37090 10843 37093
rect 15929 37090 15995 37093
rect 10777 37088 15995 37090
rect 10777 37032 10782 37088
rect 10838 37032 15934 37088
rect 15990 37032 15995 37088
rect 10777 37030 15995 37032
rect 10777 37027 10843 37030
rect 15929 37027 15995 37030
rect 21357 37090 21423 37093
rect 23381 37090 23447 37093
rect 28993 37090 29059 37093
rect 21357 37088 23076 37090
rect 21357 37032 21362 37088
rect 21418 37032 23076 37088
rect 21357 37030 23076 37032
rect 21357 37027 21423 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 18505 36954 18571 36957
rect 18873 36954 18939 36957
rect 22369 36954 22435 36957
rect 22829 36954 22895 36957
rect 18505 36952 18939 36954
rect 18505 36896 18510 36952
rect 18566 36896 18878 36952
rect 18934 36896 18939 36952
rect 18505 36894 18939 36896
rect 18505 36891 18571 36894
rect 18873 36891 18939 36894
rect 22050 36952 22895 36954
rect 22050 36896 22374 36952
rect 22430 36896 22834 36952
rect 22890 36896 22895 36952
rect 22050 36894 22895 36896
rect 23016 36954 23076 37030
rect 23381 37088 29059 37090
rect 23381 37032 23386 37088
rect 23442 37032 28998 37088
rect 29054 37032 29059 37088
rect 23381 37030 29059 37032
rect 23381 37027 23447 37030
rect 28993 37027 29059 37030
rect 23473 36954 23539 36957
rect 24209 36954 24275 36957
rect 26325 36954 26391 36957
rect 23016 36952 26391 36954
rect 23016 36896 23478 36952
rect 23534 36896 24214 36952
rect 24270 36896 26330 36952
rect 26386 36896 26391 36952
rect 23016 36894 26391 36896
rect 9581 36818 9647 36821
rect 16757 36818 16823 36821
rect 9581 36816 16823 36818
rect 9581 36760 9586 36816
rect 9642 36760 16762 36816
rect 16818 36760 16823 36816
rect 9581 36758 16823 36760
rect 9581 36755 9647 36758
rect 16757 36755 16823 36758
rect 19057 36818 19123 36821
rect 19190 36818 19196 36820
rect 19057 36816 19196 36818
rect 19057 36760 19062 36816
rect 19118 36760 19196 36816
rect 19057 36758 19196 36760
rect 19057 36755 19123 36758
rect 19190 36756 19196 36758
rect 19260 36756 19266 36820
rect 20805 36818 20871 36821
rect 22050 36818 22110 36894
rect 22369 36891 22435 36894
rect 22829 36891 22895 36894
rect 23473 36891 23539 36894
rect 24209 36891 24275 36894
rect 26325 36891 26391 36894
rect 20805 36816 22110 36818
rect 20805 36760 20810 36816
rect 20866 36760 22110 36816
rect 20805 36758 22110 36760
rect 24301 36818 24367 36821
rect 28349 36818 28415 36821
rect 24301 36816 28415 36818
rect 24301 36760 24306 36816
rect 24362 36760 28354 36816
rect 28410 36760 28415 36816
rect 24301 36758 28415 36760
rect 20805 36755 20871 36758
rect 24301 36755 24367 36758
rect 28349 36755 28415 36758
rect 40953 36818 41019 36821
rect 41720 36818 42520 36848
rect 40953 36816 42520 36818
rect 40953 36760 40958 36816
rect 41014 36760 42520 36816
rect 40953 36758 42520 36760
rect 40953 36755 41019 36758
rect 41720 36728 42520 36758
rect 15142 36620 15148 36684
rect 15212 36682 15218 36684
rect 15377 36682 15443 36685
rect 15212 36680 15443 36682
rect 15212 36624 15382 36680
rect 15438 36624 15443 36680
rect 15212 36622 15443 36624
rect 15212 36620 15218 36622
rect 15377 36619 15443 36622
rect 18229 36682 18295 36685
rect 20805 36682 20871 36685
rect 21541 36682 21607 36685
rect 18229 36680 21607 36682
rect 18229 36624 18234 36680
rect 18290 36624 20810 36680
rect 20866 36624 21546 36680
rect 21602 36624 21607 36680
rect 18229 36622 21607 36624
rect 18229 36619 18295 36622
rect 20805 36619 20871 36622
rect 21541 36619 21607 36622
rect 23013 36682 23079 36685
rect 26969 36682 27035 36685
rect 29085 36682 29151 36685
rect 29545 36682 29611 36685
rect 23013 36680 29611 36682
rect 23013 36624 23018 36680
rect 23074 36624 26974 36680
rect 27030 36624 29090 36680
rect 29146 36624 29550 36680
rect 29606 36624 29611 36680
rect 23013 36622 29611 36624
rect 23013 36619 23079 36622
rect 26969 36619 27035 36622
rect 29085 36619 29151 36622
rect 29545 36619 29611 36622
rect 19241 36546 19307 36549
rect 32581 36546 32647 36549
rect 19241 36544 32647 36546
rect 19241 36488 19246 36544
rect 19302 36488 32586 36544
rect 32642 36488 32647 36544
rect 19241 36486 32647 36488
rect 19241 36483 19307 36486
rect 32581 36483 32647 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 16573 36410 16639 36413
rect 20253 36410 20319 36413
rect 16573 36408 20319 36410
rect 16573 36352 16578 36408
rect 16634 36352 20258 36408
rect 20314 36352 20319 36408
rect 16573 36350 20319 36352
rect 16573 36347 16639 36350
rect 20253 36347 20319 36350
rect 21909 36410 21975 36413
rect 28901 36410 28967 36413
rect 21909 36408 28967 36410
rect 21909 36352 21914 36408
rect 21970 36352 28906 36408
rect 28962 36352 28967 36408
rect 21909 36350 28967 36352
rect 21909 36347 21975 36350
rect 28901 36347 28967 36350
rect 16205 36274 16271 36277
rect 21265 36274 21331 36277
rect 16205 36272 21331 36274
rect 16205 36216 16210 36272
rect 16266 36216 21270 36272
rect 21326 36216 21331 36272
rect 16205 36214 21331 36216
rect 16205 36211 16271 36214
rect 21265 36211 21331 36214
rect 21541 36274 21607 36277
rect 26141 36274 26207 36277
rect 28717 36274 28783 36277
rect 21541 36272 26066 36274
rect 21541 36216 21546 36272
rect 21602 36216 26066 36272
rect 21541 36214 26066 36216
rect 21541 36211 21607 36214
rect 0 36138 800 36168
rect 933 36138 999 36141
rect 0 36136 999 36138
rect 0 36080 938 36136
rect 994 36080 999 36136
rect 0 36078 999 36080
rect 0 36048 800 36078
rect 933 36075 999 36078
rect 17217 36138 17283 36141
rect 17534 36138 17540 36140
rect 17217 36136 17540 36138
rect 17217 36080 17222 36136
rect 17278 36080 17540 36136
rect 17217 36078 17540 36080
rect 17217 36075 17283 36078
rect 17534 36076 17540 36078
rect 17604 36138 17610 36140
rect 19333 36138 19399 36141
rect 17604 36136 19399 36138
rect 17604 36080 19338 36136
rect 19394 36080 19399 36136
rect 17604 36078 19399 36080
rect 17604 36076 17610 36078
rect 19333 36075 19399 36078
rect 19517 36138 19583 36141
rect 20110 36138 20116 36140
rect 19517 36136 20116 36138
rect 19517 36080 19522 36136
rect 19578 36080 20116 36136
rect 19517 36078 20116 36080
rect 19517 36075 19583 36078
rect 20110 36076 20116 36078
rect 20180 36076 20186 36140
rect 13537 36002 13603 36005
rect 16573 36002 16639 36005
rect 13537 36000 16639 36002
rect 13537 35944 13542 36000
rect 13598 35944 16578 36000
rect 16634 35944 16639 36000
rect 13537 35942 16639 35944
rect 13537 35939 13603 35942
rect 16573 35939 16639 35942
rect 18505 36002 18571 36005
rect 18638 36002 18644 36004
rect 18505 36000 18644 36002
rect 18505 35944 18510 36000
rect 18566 35944 18644 36000
rect 18505 35942 18644 35944
rect 18505 35939 18571 35942
rect 18638 35940 18644 35942
rect 18708 35940 18714 36004
rect 26006 36002 26066 36214
rect 26141 36272 28783 36274
rect 26141 36216 26146 36272
rect 26202 36216 28722 36272
rect 28778 36216 28783 36272
rect 26141 36214 28783 36216
rect 26141 36211 26207 36214
rect 28717 36211 28783 36214
rect 26785 36138 26851 36141
rect 28349 36138 28415 36141
rect 26785 36136 28415 36138
rect 26785 36080 26790 36136
rect 26846 36080 28354 36136
rect 28410 36080 28415 36136
rect 26785 36078 28415 36080
rect 26785 36075 26851 36078
rect 28349 36075 28415 36078
rect 31661 36002 31727 36005
rect 26006 36000 31727 36002
rect 26006 35944 31666 36000
rect 31722 35944 31727 36000
rect 26006 35942 31727 35944
rect 31661 35939 31727 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 17677 35868 17743 35869
rect 17677 35866 17724 35868
rect 17632 35864 17724 35866
rect 17632 35808 17682 35864
rect 17632 35806 17724 35808
rect 17677 35804 17724 35806
rect 17788 35804 17794 35868
rect 20253 35866 20319 35869
rect 20529 35866 20595 35869
rect 20253 35864 20595 35866
rect 20253 35808 20258 35864
rect 20314 35808 20534 35864
rect 20590 35808 20595 35864
rect 20253 35806 20595 35808
rect 17677 35803 17743 35804
rect 20253 35803 20319 35806
rect 20529 35803 20595 35806
rect 22369 35866 22435 35869
rect 30373 35866 30439 35869
rect 22369 35864 30439 35866
rect 22369 35808 22374 35864
rect 22430 35808 30378 35864
rect 30434 35808 30439 35864
rect 22369 35806 30439 35808
rect 22369 35803 22435 35806
rect 30373 35803 30439 35806
rect 8937 35730 9003 35733
rect 10041 35730 10107 35733
rect 10869 35730 10935 35733
rect 8937 35728 10935 35730
rect 8937 35672 8942 35728
rect 8998 35672 10046 35728
rect 10102 35672 10874 35728
rect 10930 35672 10935 35728
rect 8937 35670 10935 35672
rect 20532 35730 20592 35803
rect 25262 35730 25268 35732
rect 20532 35670 25268 35730
rect 8937 35667 9003 35670
rect 10041 35667 10107 35670
rect 10869 35667 10935 35670
rect 25262 35668 25268 35670
rect 25332 35668 25338 35732
rect 26785 35730 26851 35733
rect 31109 35730 31175 35733
rect 26785 35728 31175 35730
rect 26785 35672 26790 35728
rect 26846 35672 31114 35728
rect 31170 35672 31175 35728
rect 26785 35670 31175 35672
rect 26785 35667 26851 35670
rect 31109 35667 31175 35670
rect 19885 35594 19951 35597
rect 22645 35594 22711 35597
rect 19885 35592 22711 35594
rect 19885 35536 19890 35592
rect 19946 35536 22650 35592
rect 22706 35536 22711 35592
rect 19885 35534 22711 35536
rect 19885 35531 19951 35534
rect 22645 35531 22711 35534
rect 27337 35594 27403 35597
rect 29637 35594 29703 35597
rect 27337 35592 29703 35594
rect 27337 35536 27342 35592
rect 27398 35536 29642 35592
rect 29698 35536 29703 35592
rect 27337 35534 29703 35536
rect 27337 35531 27403 35534
rect 29637 35531 29703 35534
rect 27613 35458 27679 35461
rect 28625 35458 28691 35461
rect 27613 35456 28691 35458
rect 27613 35400 27618 35456
rect 27674 35400 28630 35456
rect 28686 35400 28691 35456
rect 27613 35398 28691 35400
rect 27613 35395 27679 35398
rect 28625 35395 28691 35398
rect 30465 35458 30531 35461
rect 30925 35458 30991 35461
rect 30465 35456 30991 35458
rect 30465 35400 30470 35456
rect 30526 35400 30930 35456
rect 30986 35400 30991 35456
rect 30465 35398 30991 35400
rect 30465 35395 30531 35398
rect 30925 35395 30991 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 26325 35322 26391 35325
rect 28349 35322 28415 35325
rect 26325 35320 28415 35322
rect 26325 35264 26330 35320
rect 26386 35264 28354 35320
rect 28410 35264 28415 35320
rect 26325 35262 28415 35264
rect 26325 35259 26391 35262
rect 28349 35259 28415 35262
rect 29637 35322 29703 35325
rect 30649 35322 30715 35325
rect 29637 35320 30715 35322
rect 29637 35264 29642 35320
rect 29698 35264 30654 35320
rect 30710 35264 30715 35320
rect 29637 35262 30715 35264
rect 29637 35259 29703 35262
rect 30649 35259 30715 35262
rect 14089 35186 14155 35189
rect 16665 35186 16731 35189
rect 14089 35184 16731 35186
rect 14089 35128 14094 35184
rect 14150 35128 16670 35184
rect 16726 35128 16731 35184
rect 14089 35126 16731 35128
rect 14089 35123 14155 35126
rect 16665 35123 16731 35126
rect 25313 35186 25379 35189
rect 31293 35186 31359 35189
rect 25313 35184 31359 35186
rect 25313 35128 25318 35184
rect 25374 35128 31298 35184
rect 31354 35128 31359 35184
rect 25313 35126 31359 35128
rect 25313 35123 25379 35126
rect 31293 35123 31359 35126
rect 9254 34988 9260 35052
rect 9324 35050 9330 35052
rect 9581 35050 9647 35053
rect 9324 35048 9647 35050
rect 9324 34992 9586 35048
rect 9642 34992 9647 35048
rect 9324 34990 9647 34992
rect 9324 34988 9330 34990
rect 9581 34987 9647 34990
rect 13169 35050 13235 35053
rect 15377 35050 15443 35053
rect 13169 35048 15443 35050
rect 13169 34992 13174 35048
rect 13230 34992 15382 35048
rect 15438 34992 15443 35048
rect 13169 34990 15443 34992
rect 13169 34987 13235 34990
rect 15377 34987 15443 34990
rect 25865 35050 25931 35053
rect 28809 35050 28875 35053
rect 25865 35048 28875 35050
rect 25865 34992 25870 35048
rect 25926 34992 28814 35048
rect 28870 34992 28875 35048
rect 25865 34990 28875 34992
rect 25865 34987 25931 34990
rect 28809 34987 28875 34990
rect 29085 35050 29151 35053
rect 31109 35050 31175 35053
rect 32029 35050 32095 35053
rect 29085 35048 32095 35050
rect 29085 34992 29090 35048
rect 29146 34992 31114 35048
rect 31170 34992 32034 35048
rect 32090 34992 32095 35048
rect 29085 34990 32095 34992
rect 29085 34987 29151 34990
rect 31109 34987 31175 34990
rect 32029 34987 32095 34990
rect 27613 34914 27679 34917
rect 28533 34914 28599 34917
rect 30373 34914 30439 34917
rect 27613 34912 30439 34914
rect 27613 34856 27618 34912
rect 27674 34856 28538 34912
rect 28594 34856 30378 34912
rect 30434 34856 30439 34912
rect 27613 34854 30439 34856
rect 27613 34851 27679 34854
rect 28533 34851 28599 34854
rect 30373 34851 30439 34854
rect 30649 34914 30715 34917
rect 31753 34914 31819 34917
rect 30649 34912 31819 34914
rect 30649 34856 30654 34912
rect 30710 34856 31758 34912
rect 31814 34856 31819 34912
rect 30649 34854 31819 34856
rect 30649 34851 30715 34854
rect 31753 34851 31819 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 6821 34778 6887 34781
rect 10685 34778 10751 34781
rect 6821 34776 10751 34778
rect 6821 34720 6826 34776
rect 6882 34720 10690 34776
rect 10746 34720 10751 34776
rect 6821 34718 10751 34720
rect 6821 34715 6887 34718
rect 10685 34715 10751 34718
rect 21909 34778 21975 34781
rect 24894 34778 24900 34780
rect 21909 34776 24900 34778
rect 21909 34720 21914 34776
rect 21970 34720 24900 34776
rect 21909 34718 24900 34720
rect 21909 34715 21975 34718
rect 24894 34716 24900 34718
rect 24964 34716 24970 34780
rect 25221 34778 25287 34781
rect 27654 34778 27660 34780
rect 25221 34776 27660 34778
rect 25221 34720 25226 34776
rect 25282 34720 27660 34776
rect 25221 34718 27660 34720
rect 25221 34715 25287 34718
rect 27654 34716 27660 34718
rect 27724 34778 27730 34780
rect 28717 34778 28783 34781
rect 27724 34776 28783 34778
rect 27724 34720 28722 34776
rect 28778 34720 28783 34776
rect 27724 34718 28783 34720
rect 27724 34716 27730 34718
rect 28717 34715 28783 34718
rect 29269 34778 29335 34781
rect 30281 34778 30347 34781
rect 29269 34776 30347 34778
rect 29269 34720 29274 34776
rect 29330 34720 30286 34776
rect 30342 34720 30347 34776
rect 29269 34718 30347 34720
rect 29269 34715 29335 34718
rect 30281 34715 30347 34718
rect 7373 34642 7439 34645
rect 10041 34642 10107 34645
rect 7373 34640 10107 34642
rect 7373 34584 7378 34640
rect 7434 34584 10046 34640
rect 10102 34584 10107 34640
rect 7373 34582 10107 34584
rect 7373 34579 7439 34582
rect 10041 34579 10107 34582
rect 11053 34644 11119 34645
rect 11053 34640 11100 34644
rect 11164 34642 11170 34644
rect 11053 34584 11058 34640
rect 11053 34580 11100 34584
rect 11164 34582 11210 34642
rect 11164 34580 11170 34582
rect 11462 34580 11468 34644
rect 11532 34642 11538 34644
rect 12893 34642 12959 34645
rect 11532 34640 12959 34642
rect 11532 34584 12898 34640
rect 12954 34584 12959 34640
rect 11532 34582 12959 34584
rect 11532 34580 11538 34582
rect 11053 34579 11119 34580
rect 12893 34579 12959 34582
rect 15929 34642 15995 34645
rect 27429 34644 27495 34645
rect 16798 34642 16804 34644
rect 15929 34640 16804 34642
rect 15929 34584 15934 34640
rect 15990 34584 16804 34640
rect 15929 34582 16804 34584
rect 15929 34579 15995 34582
rect 16798 34580 16804 34582
rect 16868 34580 16874 34644
rect 19190 34580 19196 34644
rect 19260 34642 19266 34644
rect 21766 34642 21772 34644
rect 19260 34582 21772 34642
rect 19260 34580 19266 34582
rect 21766 34580 21772 34582
rect 21836 34580 21842 34644
rect 27429 34640 27476 34644
rect 27540 34642 27546 34644
rect 30005 34642 30071 34645
rect 30833 34642 30899 34645
rect 27429 34584 27434 34640
rect 27429 34580 27476 34584
rect 27540 34582 27586 34642
rect 30005 34640 30899 34642
rect 30005 34584 30010 34640
rect 30066 34584 30838 34640
rect 30894 34584 30899 34640
rect 30005 34582 30899 34584
rect 27540 34580 27546 34582
rect 27429 34579 27495 34580
rect 30005 34579 30071 34582
rect 30833 34579 30899 34582
rect 24117 34506 24183 34509
rect 24710 34506 24716 34508
rect 24117 34504 24716 34506
rect 24117 34448 24122 34504
rect 24178 34448 24716 34504
rect 24117 34446 24716 34448
rect 24117 34443 24183 34446
rect 24710 34444 24716 34446
rect 24780 34444 24786 34508
rect 26049 34506 26115 34509
rect 30557 34506 30623 34509
rect 31753 34506 31819 34509
rect 26049 34504 31819 34506
rect 26049 34448 26054 34504
rect 26110 34448 30562 34504
rect 30618 34448 31758 34504
rect 31814 34448 31819 34504
rect 26049 34446 31819 34448
rect 26049 34443 26115 34446
rect 30557 34443 30623 34446
rect 31753 34443 31819 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 20069 34234 20135 34237
rect 20713 34234 20779 34237
rect 20069 34232 20779 34234
rect 20069 34176 20074 34232
rect 20130 34176 20718 34232
rect 20774 34176 20779 34232
rect 20069 34174 20779 34176
rect 20069 34171 20135 34174
rect 20713 34171 20779 34174
rect 23473 34234 23539 34237
rect 24342 34234 24348 34236
rect 23473 34232 24348 34234
rect 23473 34176 23478 34232
rect 23534 34176 24348 34232
rect 23473 34174 24348 34176
rect 23473 34171 23539 34174
rect 24342 34172 24348 34174
rect 24412 34172 24418 34236
rect 26049 34234 26115 34237
rect 26182 34234 26188 34236
rect 26049 34232 26188 34234
rect 26049 34176 26054 34232
rect 26110 34176 26188 34232
rect 26049 34174 26188 34176
rect 26049 34171 26115 34174
rect 26182 34172 26188 34174
rect 26252 34172 26258 34236
rect 23565 34098 23631 34101
rect 27245 34098 27311 34101
rect 23565 34096 27311 34098
rect 23565 34040 23570 34096
rect 23626 34040 27250 34096
rect 27306 34040 27311 34096
rect 23565 34038 27311 34040
rect 23565 34035 23631 34038
rect 27245 34035 27311 34038
rect 13629 33962 13695 33965
rect 15101 33962 15167 33965
rect 13629 33960 15167 33962
rect 13629 33904 13634 33960
rect 13690 33904 15106 33960
rect 15162 33904 15167 33960
rect 13629 33902 15167 33904
rect 13629 33899 13695 33902
rect 15101 33899 15167 33902
rect 19425 33962 19491 33965
rect 28533 33962 28599 33965
rect 19425 33960 28599 33962
rect 19425 33904 19430 33960
rect 19486 33904 28538 33960
rect 28594 33904 28599 33960
rect 19425 33902 28599 33904
rect 19425 33899 19491 33902
rect 28533 33899 28599 33902
rect 9622 33764 9628 33828
rect 9692 33826 9698 33828
rect 13537 33826 13603 33829
rect 9692 33824 13603 33826
rect 9692 33768 13542 33824
rect 13598 33768 13603 33824
rect 9692 33766 13603 33768
rect 9692 33764 9698 33766
rect 13537 33763 13603 33766
rect 22829 33826 22895 33829
rect 25998 33826 26004 33828
rect 22829 33824 26004 33826
rect 22829 33768 22834 33824
rect 22890 33768 26004 33824
rect 22829 33766 26004 33768
rect 22829 33763 22895 33766
rect 25998 33764 26004 33766
rect 26068 33826 26074 33828
rect 26233 33826 26299 33829
rect 26068 33824 26299 33826
rect 26068 33768 26238 33824
rect 26294 33768 26299 33824
rect 26068 33766 26299 33768
rect 26068 33764 26074 33766
rect 26233 33763 26299 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 8201 33690 8267 33693
rect 16205 33690 16271 33693
rect 8201 33688 16271 33690
rect 8201 33632 8206 33688
rect 8262 33632 16210 33688
rect 16266 33632 16271 33688
rect 8201 33630 16271 33632
rect 8201 33627 8267 33630
rect 16205 33627 16271 33630
rect 21357 33690 21423 33693
rect 26877 33690 26943 33693
rect 21357 33688 26943 33690
rect 21357 33632 21362 33688
rect 21418 33632 26882 33688
rect 26938 33632 26943 33688
rect 21357 33630 26943 33632
rect 21357 33627 21423 33630
rect 26877 33627 26943 33630
rect 21541 33554 21607 33557
rect 24025 33554 24091 33557
rect 21541 33552 24091 33554
rect 21541 33496 21546 33552
rect 21602 33496 24030 33552
rect 24086 33496 24091 33552
rect 21541 33494 24091 33496
rect 21541 33491 21607 33494
rect 24025 33491 24091 33494
rect 24393 33554 24459 33557
rect 25129 33554 25195 33557
rect 24393 33552 25195 33554
rect 24393 33496 24398 33552
rect 24454 33496 25134 33552
rect 25190 33496 25195 33552
rect 24393 33494 25195 33496
rect 24393 33491 24459 33494
rect 25129 33491 25195 33494
rect 26141 33554 26207 33557
rect 29269 33554 29335 33557
rect 26141 33552 29335 33554
rect 26141 33496 26146 33552
rect 26202 33496 29274 33552
rect 29330 33496 29335 33552
rect 26141 33494 29335 33496
rect 26141 33491 26207 33494
rect 29269 33491 29335 33494
rect 12525 33418 12591 33421
rect 22921 33418 22987 33421
rect 27429 33418 27495 33421
rect 12525 33416 22987 33418
rect 12525 33360 12530 33416
rect 12586 33360 22926 33416
rect 22982 33360 22987 33416
rect 12525 33358 22987 33360
rect 12525 33355 12591 33358
rect 22921 33355 22987 33358
rect 24166 33416 27495 33418
rect 24166 33360 27434 33416
rect 27490 33360 27495 33416
rect 24166 33358 27495 33360
rect 12985 33282 13051 33285
rect 17309 33282 17375 33285
rect 12985 33280 17375 33282
rect 12985 33224 12990 33280
rect 13046 33224 17314 33280
rect 17370 33224 17375 33280
rect 12985 33222 17375 33224
rect 12985 33219 13051 33222
rect 17309 33219 17375 33222
rect 21541 33282 21607 33285
rect 24166 33282 24226 33358
rect 27429 33355 27495 33358
rect 21541 33280 24226 33282
rect 21541 33224 21546 33280
rect 21602 33224 24226 33280
rect 21541 33222 24226 33224
rect 24301 33282 24367 33285
rect 25497 33282 25563 33285
rect 24301 33280 25563 33282
rect 24301 33224 24306 33280
rect 24362 33224 25502 33280
rect 25558 33224 25563 33280
rect 24301 33222 25563 33224
rect 21541 33219 21607 33222
rect 24301 33219 24367 33222
rect 25497 33219 25563 33222
rect 25773 33284 25839 33285
rect 25773 33280 25820 33284
rect 25884 33282 25890 33284
rect 25773 33224 25778 33280
rect 25773 33220 25820 33224
rect 25884 33222 25930 33282
rect 25884 33220 25890 33222
rect 25773 33219 25839 33220
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 16021 33146 16087 33149
rect 26918 33146 26924 33148
rect 16021 33144 26924 33146
rect 16021 33088 16026 33144
rect 16082 33088 26924 33144
rect 16021 33086 26924 33088
rect 16021 33083 16087 33086
rect 26918 33084 26924 33086
rect 26988 33146 26994 33148
rect 27705 33146 27771 33149
rect 26988 33144 27771 33146
rect 26988 33088 27710 33144
rect 27766 33088 27771 33144
rect 26988 33086 27771 33088
rect 26988 33084 26994 33086
rect 27705 33083 27771 33086
rect 8385 33010 8451 33013
rect 13997 33010 14063 33013
rect 17033 33010 17099 33013
rect 8385 33008 12450 33010
rect 8385 32952 8390 33008
rect 8446 32952 12450 33008
rect 8385 32950 12450 32952
rect 8385 32947 8451 32950
rect 6085 32874 6151 32877
rect 11789 32874 11855 32877
rect 6085 32872 11855 32874
rect 6085 32816 6090 32872
rect 6146 32816 11794 32872
rect 11850 32816 11855 32872
rect 6085 32814 11855 32816
rect 12390 32874 12450 32950
rect 13997 33008 17099 33010
rect 13997 32952 14002 33008
rect 14058 32952 17038 33008
rect 17094 32952 17099 33008
rect 13997 32950 17099 32952
rect 13997 32947 14063 32950
rect 17033 32947 17099 32950
rect 23422 32948 23428 33012
rect 23492 33010 23498 33012
rect 27102 33010 27108 33012
rect 23492 32950 27108 33010
rect 23492 32948 23498 32950
rect 27102 32948 27108 32950
rect 27172 33010 27178 33012
rect 27521 33010 27587 33013
rect 27172 33008 27587 33010
rect 27172 32952 27526 33008
rect 27582 32952 27587 33008
rect 27172 32950 27587 32952
rect 27172 32948 27178 32950
rect 27521 32947 27587 32950
rect 16757 32874 16823 32877
rect 20253 32874 20319 32877
rect 12390 32872 20319 32874
rect 12390 32816 16762 32872
rect 16818 32816 20258 32872
rect 20314 32816 20319 32872
rect 12390 32814 20319 32816
rect 6085 32811 6151 32814
rect 11789 32811 11855 32814
rect 16757 32811 16823 32814
rect 20253 32811 20319 32814
rect 24117 32874 24183 32877
rect 26877 32874 26943 32877
rect 28533 32874 28599 32877
rect 24117 32872 28599 32874
rect 24117 32816 24122 32872
rect 24178 32816 26882 32872
rect 26938 32816 28538 32872
rect 28594 32816 28599 32872
rect 24117 32814 28599 32816
rect 24117 32811 24183 32814
rect 26877 32811 26943 32814
rect 28533 32811 28599 32814
rect 12525 32738 12591 32741
rect 18413 32738 18479 32741
rect 12525 32736 18479 32738
rect 12525 32680 12530 32736
rect 12586 32680 18418 32736
rect 18474 32680 18479 32736
rect 12525 32678 18479 32680
rect 12525 32675 12591 32678
rect 18413 32675 18479 32678
rect 20897 32738 20963 32741
rect 26601 32738 26667 32741
rect 20897 32736 26667 32738
rect 20897 32680 20902 32736
rect 20958 32680 26606 32736
rect 26662 32680 26667 32736
rect 20897 32678 26667 32680
rect 20897 32675 20963 32678
rect 26601 32675 26667 32678
rect 40953 32738 41019 32741
rect 41720 32738 42520 32768
rect 40953 32736 42520 32738
rect 40953 32680 40958 32736
rect 41014 32680 42520 32736
rect 40953 32678 42520 32680
rect 40953 32675 41019 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 41720 32648 42520 32678
rect 19570 32607 19886 32608
rect 13537 32602 13603 32605
rect 18413 32602 18479 32605
rect 13537 32600 18479 32602
rect 13537 32544 13542 32600
rect 13598 32544 18418 32600
rect 18474 32544 18479 32600
rect 13537 32542 18479 32544
rect 13537 32539 13603 32542
rect 18413 32539 18479 32542
rect 20897 32602 20963 32605
rect 22553 32602 22619 32605
rect 20897 32600 22619 32602
rect 20897 32544 20902 32600
rect 20958 32544 22558 32600
rect 22614 32544 22619 32600
rect 20897 32542 22619 32544
rect 20897 32539 20963 32542
rect 22553 32539 22619 32542
rect 25129 32602 25195 32605
rect 27981 32602 28047 32605
rect 25129 32600 28047 32602
rect 25129 32544 25134 32600
rect 25190 32544 27986 32600
rect 28042 32544 28047 32600
rect 25129 32542 28047 32544
rect 25129 32539 25195 32542
rect 27981 32539 28047 32542
rect 11145 32466 11211 32469
rect 11278 32466 11284 32468
rect 11145 32464 11284 32466
rect 11145 32408 11150 32464
rect 11206 32408 11284 32464
rect 11145 32406 11284 32408
rect 11145 32403 11211 32406
rect 11278 32404 11284 32406
rect 11348 32404 11354 32468
rect 11881 32466 11947 32469
rect 28809 32466 28875 32469
rect 11881 32464 28875 32466
rect 11881 32408 11886 32464
rect 11942 32408 28814 32464
rect 28870 32408 28875 32464
rect 11881 32406 28875 32408
rect 11881 32403 11947 32406
rect 28809 32403 28875 32406
rect 9673 32330 9739 32333
rect 13077 32330 13143 32333
rect 9673 32328 13143 32330
rect 9673 32272 9678 32328
rect 9734 32272 13082 32328
rect 13138 32272 13143 32328
rect 9673 32270 13143 32272
rect 9673 32267 9739 32270
rect 13077 32267 13143 32270
rect 15009 32330 15075 32333
rect 17033 32330 17099 32333
rect 27245 32330 27311 32333
rect 29126 32330 29132 32332
rect 15009 32328 21834 32330
rect 15009 32272 15014 32328
rect 15070 32272 17038 32328
rect 17094 32272 21834 32328
rect 15009 32270 21834 32272
rect 15009 32267 15075 32270
rect 17033 32267 17099 32270
rect 9305 32194 9371 32197
rect 9581 32194 9647 32197
rect 12525 32194 12591 32197
rect 9305 32192 9647 32194
rect 9305 32136 9310 32192
rect 9366 32136 9586 32192
rect 9642 32136 9647 32192
rect 9305 32134 9647 32136
rect 9305 32131 9371 32134
rect 9581 32131 9647 32134
rect 11654 32192 12591 32194
rect 11654 32136 12530 32192
rect 12586 32136 12591 32192
rect 11654 32134 12591 32136
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 933 32058 999 32061
rect 0 32056 999 32058
rect 0 32000 938 32056
rect 994 32000 999 32056
rect 0 31998 999 32000
rect 0 31968 800 31998
rect 933 31995 999 31998
rect 7925 32058 7991 32061
rect 10358 32058 10364 32060
rect 7925 32056 10364 32058
rect 7925 32000 7930 32056
rect 7986 32000 10364 32056
rect 7925 31998 10364 32000
rect 7925 31995 7991 31998
rect 10358 31996 10364 31998
rect 10428 32058 10434 32060
rect 10685 32058 10751 32061
rect 10428 32056 10751 32058
rect 10428 32000 10690 32056
rect 10746 32000 10751 32056
rect 10428 31998 10751 32000
rect 10428 31996 10434 31998
rect 10685 31995 10751 31998
rect 5717 31922 5783 31925
rect 11654 31922 11714 32134
rect 12525 32131 12591 32134
rect 16246 32132 16252 32196
rect 16316 32194 16322 32196
rect 19701 32194 19767 32197
rect 16316 32192 19767 32194
rect 16316 32136 19706 32192
rect 19762 32136 19767 32192
rect 16316 32134 19767 32136
rect 16316 32132 16322 32134
rect 19701 32131 19767 32134
rect 20805 32194 20871 32197
rect 21398 32194 21404 32196
rect 20805 32192 21404 32194
rect 20805 32136 20810 32192
rect 20866 32136 21404 32192
rect 20805 32134 21404 32136
rect 20805 32131 20871 32134
rect 21398 32132 21404 32134
rect 21468 32132 21474 32196
rect 11789 32058 11855 32061
rect 17769 32058 17835 32061
rect 19425 32058 19491 32061
rect 21449 32058 21515 32061
rect 11789 32056 17835 32058
rect 11789 32000 11794 32056
rect 11850 32000 17774 32056
rect 17830 32000 17835 32056
rect 11789 31998 17835 32000
rect 11789 31995 11855 31998
rect 17769 31995 17835 31998
rect 19290 32056 21515 32058
rect 19290 32000 19430 32056
rect 19486 32000 21454 32056
rect 21510 32000 21515 32056
rect 19290 31998 21515 32000
rect 21774 32058 21834 32270
rect 27245 32328 29132 32330
rect 27245 32272 27250 32328
rect 27306 32272 29132 32328
rect 27245 32270 29132 32272
rect 27245 32267 27311 32270
rect 29126 32268 29132 32270
rect 29196 32268 29202 32332
rect 22134 32132 22140 32196
rect 22204 32194 22210 32196
rect 22277 32194 22343 32197
rect 23606 32194 23612 32196
rect 22204 32192 22343 32194
rect 22204 32136 22282 32192
rect 22338 32136 22343 32192
rect 22204 32134 22343 32136
rect 22204 32132 22210 32134
rect 22277 32131 22343 32134
rect 23246 32134 23612 32194
rect 23246 32058 23306 32134
rect 23606 32132 23612 32134
rect 23676 32132 23682 32196
rect 26601 32194 26667 32197
rect 26601 32192 27538 32194
rect 26601 32136 26606 32192
rect 26662 32136 27538 32192
rect 26601 32134 27538 32136
rect 26601 32131 26667 32134
rect 27478 32061 27538 32134
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 21774 31998 23306 32058
rect 23657 32058 23723 32061
rect 25221 32058 25287 32061
rect 27245 32058 27311 32061
rect 23657 32056 23858 32058
rect 23657 32000 23662 32056
rect 23718 32000 23858 32056
rect 23657 31998 23858 32000
rect 5717 31920 11714 31922
rect 5717 31864 5722 31920
rect 5778 31864 11714 31920
rect 5717 31862 11714 31864
rect 12893 31922 12959 31925
rect 13905 31922 13971 31925
rect 17125 31922 17191 31925
rect 12893 31920 17191 31922
rect 12893 31864 12898 31920
rect 12954 31864 13910 31920
rect 13966 31864 17130 31920
rect 17186 31864 17191 31920
rect 12893 31862 17191 31864
rect 5717 31859 5783 31862
rect 12893 31859 12959 31862
rect 13905 31859 13971 31862
rect 17125 31859 17191 31862
rect 17401 31922 17467 31925
rect 19290 31922 19350 31998
rect 19425 31995 19491 31998
rect 21449 31995 21515 31998
rect 23657 31995 23723 31998
rect 17401 31920 19350 31922
rect 17401 31864 17406 31920
rect 17462 31864 19350 31920
rect 17401 31862 19350 31864
rect 19701 31922 19767 31925
rect 23657 31922 23723 31925
rect 19701 31920 23723 31922
rect 19701 31864 19706 31920
rect 19762 31864 23662 31920
rect 23718 31864 23723 31920
rect 19701 31862 23723 31864
rect 17401 31859 17467 31862
rect 19701 31859 19767 31862
rect 23657 31859 23723 31862
rect 8753 31786 8819 31789
rect 9581 31786 9647 31789
rect 10777 31786 10843 31789
rect 8753 31784 9000 31786
rect 8753 31728 8758 31784
rect 8814 31728 9000 31784
rect 8753 31726 9000 31728
rect 8753 31723 8819 31726
rect 8940 31650 9000 31726
rect 9581 31784 10843 31786
rect 9581 31728 9586 31784
rect 9642 31728 10782 31784
rect 10838 31728 10843 31784
rect 9581 31726 10843 31728
rect 9581 31723 9647 31726
rect 10777 31723 10843 31726
rect 16665 31786 16731 31789
rect 19977 31786 20043 31789
rect 23798 31786 23858 31998
rect 25221 32056 27311 32058
rect 25221 32000 25226 32056
rect 25282 32000 27250 32056
rect 27306 32000 27311 32056
rect 25221 31998 27311 32000
rect 27478 32058 27587 32061
rect 29729 32058 29795 32061
rect 27478 32056 29795 32058
rect 27478 32000 27526 32056
rect 27582 32000 29734 32056
rect 29790 32000 29795 32056
rect 27478 31998 29795 32000
rect 25221 31995 25287 31998
rect 27245 31995 27311 31998
rect 27521 31995 27587 31998
rect 29729 31995 29795 31998
rect 25037 31922 25103 31925
rect 27429 31922 27495 31925
rect 25037 31920 27495 31922
rect 25037 31864 25042 31920
rect 25098 31864 27434 31920
rect 27490 31864 27495 31920
rect 25037 31862 27495 31864
rect 25037 31859 25103 31862
rect 27429 31859 27495 31862
rect 16665 31784 20043 31786
rect 16665 31728 16670 31784
rect 16726 31728 19982 31784
rect 20038 31728 20043 31784
rect 16665 31726 20043 31728
rect 16665 31723 16731 31726
rect 19977 31723 20043 31726
rect 21544 31726 23858 31786
rect 10685 31650 10751 31653
rect 8940 31648 10751 31650
rect 8940 31592 10690 31648
rect 10746 31592 10751 31648
rect 8940 31590 10751 31592
rect 10685 31587 10751 31590
rect 20069 31650 20135 31653
rect 21544 31650 21604 31726
rect 24894 31724 24900 31788
rect 24964 31786 24970 31788
rect 25037 31786 25103 31789
rect 24964 31784 25103 31786
rect 24964 31728 25042 31784
rect 25098 31728 25103 31784
rect 24964 31726 25103 31728
rect 24964 31724 24970 31726
rect 25037 31723 25103 31726
rect 25773 31786 25839 31789
rect 26325 31786 26391 31789
rect 25773 31784 26391 31786
rect 25773 31728 25778 31784
rect 25834 31728 26330 31784
rect 26386 31728 26391 31784
rect 25773 31726 26391 31728
rect 25773 31723 25839 31726
rect 26325 31723 26391 31726
rect 26509 31650 26575 31653
rect 20069 31648 21604 31650
rect 20069 31592 20074 31648
rect 20130 31592 21604 31648
rect 20069 31590 21604 31592
rect 22050 31648 26575 31650
rect 22050 31592 26514 31648
rect 26570 31592 26575 31648
rect 22050 31590 26575 31592
rect 20069 31587 20135 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 9397 31514 9463 31517
rect 9622 31514 9628 31516
rect 9397 31512 9628 31514
rect 9397 31456 9402 31512
rect 9458 31456 9628 31512
rect 9397 31454 9628 31456
rect 9397 31451 9463 31454
rect 9622 31452 9628 31454
rect 9692 31452 9698 31516
rect 8293 31378 8359 31381
rect 9581 31378 9647 31381
rect 8293 31376 9647 31378
rect 8293 31320 8298 31376
rect 8354 31320 9586 31376
rect 9642 31320 9647 31376
rect 8293 31318 9647 31320
rect 8293 31315 8359 31318
rect 9581 31315 9647 31318
rect 11145 31378 11211 31381
rect 19793 31378 19859 31381
rect 11145 31376 19859 31378
rect 11145 31320 11150 31376
rect 11206 31320 19798 31376
rect 19854 31320 19859 31376
rect 11145 31318 19859 31320
rect 11145 31315 11211 31318
rect 19793 31315 19859 31318
rect 20713 31378 20779 31381
rect 22050 31378 22110 31590
rect 26509 31587 26575 31590
rect 27286 31588 27292 31652
rect 27356 31650 27362 31652
rect 30925 31650 30991 31653
rect 27356 31648 30991 31650
rect 27356 31592 30930 31648
rect 30986 31592 30991 31648
rect 27356 31590 30991 31592
rect 27356 31588 27362 31590
rect 23749 31514 23815 31517
rect 27102 31514 27108 31516
rect 23749 31512 27108 31514
rect 23749 31456 23754 31512
rect 23810 31456 27108 31512
rect 23749 31454 27108 31456
rect 23749 31451 23815 31454
rect 27102 31452 27108 31454
rect 27172 31452 27178 31516
rect 20713 31376 22110 31378
rect 20713 31320 20718 31376
rect 20774 31320 22110 31376
rect 20713 31318 22110 31320
rect 22185 31378 22251 31381
rect 25129 31378 25195 31381
rect 22185 31376 25195 31378
rect 22185 31320 22190 31376
rect 22246 31320 25134 31376
rect 25190 31320 25195 31376
rect 22185 31318 25195 31320
rect 20713 31315 20779 31318
rect 22185 31315 22251 31318
rect 25129 31315 25195 31318
rect 19333 31242 19399 31245
rect 27294 31242 27354 31588
rect 30925 31587 30991 31590
rect 19333 31240 27354 31242
rect 19333 31184 19338 31240
rect 19394 31184 27354 31240
rect 19333 31182 27354 31184
rect 19333 31179 19399 31182
rect 18137 31106 18203 31109
rect 27153 31106 27219 31109
rect 18137 31104 27219 31106
rect 18137 31048 18142 31104
rect 18198 31048 27158 31104
rect 27214 31048 27219 31104
rect 18137 31046 27219 31048
rect 18137 31043 18203 31046
rect 27153 31043 27219 31046
rect 28022 31044 28028 31108
rect 28092 31106 28098 31108
rect 28257 31106 28323 31109
rect 28092 31104 28323 31106
rect 28092 31048 28262 31104
rect 28318 31048 28323 31104
rect 28092 31046 28323 31048
rect 28092 31044 28098 31046
rect 28257 31043 28323 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 21081 30970 21147 30973
rect 21081 30968 22110 30970
rect 21081 30912 21086 30968
rect 21142 30912 22110 30968
rect 21081 30910 22110 30912
rect 21081 30907 21147 30910
rect 22050 30834 22110 30910
rect 23606 30908 23612 30972
rect 23676 30970 23682 30972
rect 28073 30970 28139 30973
rect 23676 30968 28139 30970
rect 23676 30912 28078 30968
rect 28134 30912 28139 30968
rect 23676 30910 28139 30912
rect 23676 30908 23682 30910
rect 28073 30907 28139 30910
rect 23749 30834 23815 30837
rect 22050 30832 23815 30834
rect 22050 30776 23754 30832
rect 23810 30776 23815 30832
rect 22050 30774 23815 30776
rect 23749 30771 23815 30774
rect 24158 30772 24164 30836
rect 24228 30834 24234 30836
rect 24669 30834 24735 30837
rect 29361 30836 29427 30837
rect 24228 30832 24735 30834
rect 24228 30776 24674 30832
rect 24730 30776 24735 30832
rect 24228 30774 24735 30776
rect 24228 30772 24234 30774
rect 24669 30771 24735 30774
rect 29310 30772 29316 30836
rect 29380 30834 29427 30836
rect 29637 30834 29703 30837
rect 29380 30832 29703 30834
rect 29422 30776 29642 30832
rect 29698 30776 29703 30832
rect 29380 30774 29703 30776
rect 29380 30772 29427 30774
rect 29361 30771 29427 30772
rect 29637 30771 29703 30774
rect 17953 30698 18019 30701
rect 21030 30698 21036 30700
rect 17953 30696 21036 30698
rect 17953 30640 17958 30696
rect 18014 30640 21036 30696
rect 17953 30638 21036 30640
rect 17953 30635 18019 30638
rect 21030 30636 21036 30638
rect 21100 30636 21106 30700
rect 21766 30636 21772 30700
rect 21836 30698 21842 30700
rect 24117 30698 24183 30701
rect 21836 30696 24183 30698
rect 21836 30640 24122 30696
rect 24178 30640 24183 30696
rect 21836 30638 24183 30640
rect 21836 30636 21842 30638
rect 24117 30635 24183 30638
rect 24526 30636 24532 30700
rect 24596 30698 24602 30700
rect 25313 30698 25379 30701
rect 24596 30696 25379 30698
rect 24596 30640 25318 30696
rect 25374 30640 25379 30696
rect 24596 30638 25379 30640
rect 24596 30636 24602 30638
rect 25313 30635 25379 30638
rect 13629 30562 13695 30565
rect 17585 30562 17651 30565
rect 13629 30560 17651 30562
rect 13629 30504 13634 30560
rect 13690 30504 17590 30560
rect 17646 30504 17651 30560
rect 13629 30502 17651 30504
rect 13629 30499 13695 30502
rect 17585 30499 17651 30502
rect 20253 30562 20319 30565
rect 20478 30562 20484 30564
rect 20253 30560 20484 30562
rect 20253 30504 20258 30560
rect 20314 30504 20484 30560
rect 20253 30502 20484 30504
rect 20253 30499 20319 30502
rect 20478 30500 20484 30502
rect 20548 30500 20554 30564
rect 21357 30562 21423 30565
rect 24761 30562 24827 30565
rect 21357 30560 24827 30562
rect 21357 30504 21362 30560
rect 21418 30504 24766 30560
rect 24822 30504 24827 30560
rect 21357 30502 24827 30504
rect 21357 30499 21423 30502
rect 24761 30499 24827 30502
rect 25037 30562 25103 30565
rect 26141 30562 26207 30565
rect 27337 30564 27403 30565
rect 25037 30560 26207 30562
rect 25037 30504 25042 30560
rect 25098 30504 26146 30560
rect 26202 30504 26207 30560
rect 25037 30502 26207 30504
rect 25037 30499 25103 30502
rect 26141 30499 26207 30502
rect 27286 30500 27292 30564
rect 27356 30562 27403 30564
rect 27356 30560 27448 30562
rect 27398 30504 27448 30560
rect 27356 30502 27448 30504
rect 27356 30500 27403 30502
rect 27337 30499 27403 30500
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 10961 30426 11027 30429
rect 10961 30424 12450 30426
rect 10961 30368 10966 30424
rect 11022 30368 12450 30424
rect 10961 30366 12450 30368
rect 10961 30363 11027 30366
rect 12390 30290 12450 30366
rect 16062 30364 16068 30428
rect 16132 30426 16138 30428
rect 16297 30426 16363 30429
rect 22737 30428 22803 30429
rect 22686 30426 22692 30428
rect 16132 30424 19488 30426
rect 16132 30368 16302 30424
rect 16358 30368 19488 30424
rect 16132 30366 19488 30368
rect 16132 30364 16138 30366
rect 16297 30363 16363 30366
rect 13077 30290 13143 30293
rect 12390 30288 13143 30290
rect 12390 30232 13082 30288
rect 13138 30232 13143 30288
rect 12390 30230 13143 30232
rect 13077 30227 13143 30230
rect 13997 30290 14063 30293
rect 16297 30290 16363 30293
rect 13997 30288 16363 30290
rect 13997 30232 14002 30288
rect 14058 30232 16302 30288
rect 16358 30232 16363 30288
rect 13997 30230 16363 30232
rect 19428 30290 19488 30366
rect 20118 30366 22692 30426
rect 22756 30426 22803 30428
rect 23105 30426 23171 30429
rect 28257 30426 28323 30429
rect 22756 30424 22848 30426
rect 22798 30368 22848 30424
rect 20118 30290 20178 30366
rect 22686 30364 22692 30366
rect 22756 30366 22848 30368
rect 23105 30424 28323 30426
rect 23105 30368 23110 30424
rect 23166 30368 28262 30424
rect 28318 30368 28323 30424
rect 23105 30366 28323 30368
rect 22756 30364 22803 30366
rect 22737 30363 22803 30364
rect 23105 30363 23171 30366
rect 28257 30363 28323 30366
rect 19428 30230 20178 30290
rect 22829 30290 22895 30293
rect 25497 30290 25563 30293
rect 22829 30288 25563 30290
rect 22829 30232 22834 30288
rect 22890 30232 25502 30288
rect 25558 30232 25563 30288
rect 22829 30230 25563 30232
rect 13997 30227 14063 30230
rect 16297 30227 16363 30230
rect 22829 30227 22895 30230
rect 25497 30227 25563 30230
rect 29494 30228 29500 30292
rect 29564 30290 29570 30292
rect 29637 30290 29703 30293
rect 29564 30288 29703 30290
rect 29564 30232 29642 30288
rect 29698 30232 29703 30288
rect 29564 30230 29703 30232
rect 29564 30228 29570 30230
rect 29637 30227 29703 30230
rect 11646 30092 11652 30156
rect 11716 30154 11722 30156
rect 16481 30154 16547 30157
rect 11716 30152 16547 30154
rect 11716 30096 16486 30152
rect 16542 30096 16547 30152
rect 11716 30094 16547 30096
rect 11716 30092 11722 30094
rect 16481 30091 16547 30094
rect 18638 30092 18644 30156
rect 18708 30154 18714 30156
rect 40953 30154 41019 30157
rect 18708 30152 41019 30154
rect 18708 30096 40958 30152
rect 41014 30096 41019 30152
rect 18708 30094 41019 30096
rect 18708 30092 18714 30094
rect 40953 30091 41019 30094
rect 11605 30018 11671 30021
rect 12566 30018 12572 30020
rect 11605 30016 12572 30018
rect 11605 29960 11610 30016
rect 11666 29960 12572 30016
rect 11605 29958 12572 29960
rect 11605 29955 11671 29958
rect 12566 29956 12572 29958
rect 12636 30018 12642 30020
rect 13169 30018 13235 30021
rect 22277 30018 22343 30021
rect 24393 30018 24459 30021
rect 12636 30016 24459 30018
rect 12636 29960 13174 30016
rect 13230 29960 22282 30016
rect 22338 29960 24398 30016
rect 24454 29960 24459 30016
rect 12636 29958 24459 29960
rect 12636 29956 12642 29958
rect 13169 29955 13235 29958
rect 22277 29955 22343 29958
rect 24393 29955 24459 29958
rect 27429 30018 27495 30021
rect 27981 30018 28047 30021
rect 27429 30016 28047 30018
rect 27429 29960 27434 30016
rect 27490 29960 27986 30016
rect 28042 29960 28047 30016
rect 27429 29958 28047 29960
rect 27429 29955 27495 29958
rect 27981 29955 28047 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 10501 29882 10567 29885
rect 16573 29882 16639 29885
rect 10501 29880 16639 29882
rect 10501 29824 10506 29880
rect 10562 29824 16578 29880
rect 16634 29824 16639 29880
rect 10501 29822 16639 29824
rect 10501 29819 10567 29822
rect 16573 29819 16639 29822
rect 18597 29882 18663 29885
rect 22185 29882 22251 29885
rect 18597 29880 22251 29882
rect 18597 29824 18602 29880
rect 18658 29824 22190 29880
rect 22246 29824 22251 29880
rect 18597 29822 22251 29824
rect 18597 29819 18663 29822
rect 22185 29819 22251 29822
rect 22921 29882 22987 29885
rect 28165 29882 28231 29885
rect 22921 29880 28231 29882
rect 22921 29824 22926 29880
rect 22982 29824 28170 29880
rect 28226 29824 28231 29880
rect 22921 29822 28231 29824
rect 22921 29819 22987 29822
rect 28165 29819 28231 29822
rect 14038 29684 14044 29748
rect 14108 29746 14114 29748
rect 15377 29746 15443 29749
rect 21633 29746 21699 29749
rect 14108 29744 15443 29746
rect 14108 29688 15382 29744
rect 15438 29688 15443 29744
rect 14108 29686 15443 29688
rect 14108 29684 14114 29686
rect 15377 29683 15443 29686
rect 15518 29744 21699 29746
rect 15518 29688 21638 29744
rect 21694 29688 21699 29744
rect 15518 29686 21699 29688
rect 13353 29610 13419 29613
rect 15101 29610 15167 29613
rect 15518 29610 15578 29686
rect 21633 29683 21699 29686
rect 22461 29746 22527 29749
rect 23565 29746 23631 29749
rect 29310 29746 29316 29748
rect 22461 29744 23631 29746
rect 22461 29688 22466 29744
rect 22522 29688 23570 29744
rect 23626 29688 23631 29744
rect 22461 29686 23631 29688
rect 22461 29683 22527 29686
rect 23565 29683 23631 29686
rect 23798 29686 29316 29746
rect 13353 29608 15578 29610
rect 13353 29552 13358 29608
rect 13414 29552 15106 29608
rect 15162 29552 15578 29608
rect 13353 29550 15578 29552
rect 13353 29547 13419 29550
rect 15101 29547 15167 29550
rect 17902 29548 17908 29612
rect 17972 29610 17978 29612
rect 22134 29610 22140 29612
rect 17972 29550 22140 29610
rect 17972 29548 17978 29550
rect 22134 29548 22140 29550
rect 22204 29548 22210 29612
rect 22829 29610 22895 29613
rect 23565 29610 23631 29613
rect 22829 29608 23631 29610
rect 22829 29552 22834 29608
rect 22890 29552 23570 29608
rect 23626 29552 23631 29608
rect 22829 29550 23631 29552
rect 22829 29547 22895 29550
rect 23565 29547 23631 29550
rect 11053 29474 11119 29477
rect 11646 29474 11652 29476
rect 11053 29472 11652 29474
rect 11053 29416 11058 29472
rect 11114 29416 11652 29472
rect 11053 29414 11652 29416
rect 11053 29411 11119 29414
rect 11646 29412 11652 29414
rect 11716 29412 11722 29476
rect 12433 29474 12499 29477
rect 16021 29474 16087 29477
rect 12433 29472 16087 29474
rect 12433 29416 12438 29472
rect 12494 29416 16026 29472
rect 16082 29416 16087 29472
rect 12433 29414 16087 29416
rect 12433 29411 12499 29414
rect 16021 29411 16087 29414
rect 21541 29474 21607 29477
rect 23798 29474 23858 29686
rect 29310 29684 29316 29686
rect 29380 29684 29386 29748
rect 24025 29610 24091 29613
rect 25221 29610 25287 29613
rect 25589 29610 25655 29613
rect 30925 29610 30991 29613
rect 24025 29608 30991 29610
rect 24025 29552 24030 29608
rect 24086 29552 25226 29608
rect 25282 29552 25594 29608
rect 25650 29552 30930 29608
rect 30986 29552 30991 29608
rect 24025 29550 30991 29552
rect 24025 29547 24091 29550
rect 25221 29547 25287 29550
rect 25589 29547 25655 29550
rect 30925 29547 30991 29550
rect 21541 29472 23858 29474
rect 21541 29416 21546 29472
rect 21602 29416 23858 29472
rect 21541 29414 23858 29416
rect 24485 29474 24551 29477
rect 25037 29474 25103 29477
rect 24485 29472 25103 29474
rect 24485 29416 24490 29472
rect 24546 29416 25042 29472
rect 25098 29416 25103 29472
rect 24485 29414 25103 29416
rect 21541 29411 21607 29414
rect 24485 29411 24551 29414
rect 25037 29411 25103 29414
rect 25221 29474 25287 29477
rect 27654 29474 27660 29476
rect 25221 29472 27660 29474
rect 25221 29416 25226 29472
rect 25282 29416 27660 29472
rect 25221 29414 27660 29416
rect 25221 29411 25287 29414
rect 27654 29412 27660 29414
rect 27724 29474 27730 29476
rect 30557 29474 30623 29477
rect 27724 29472 30623 29474
rect 27724 29416 30562 29472
rect 30618 29416 30623 29472
rect 27724 29414 30623 29416
rect 27724 29412 27730 29414
rect 30557 29411 30623 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 13997 29338 14063 29341
rect 14733 29338 14799 29341
rect 13997 29336 14799 29338
rect 13997 29280 14002 29336
rect 14058 29280 14738 29336
rect 14794 29280 14799 29336
rect 13997 29278 14799 29280
rect 13997 29275 14063 29278
rect 14733 29275 14799 29278
rect 22185 29338 22251 29341
rect 26509 29338 26575 29341
rect 22185 29336 26575 29338
rect 22185 29280 22190 29336
rect 22246 29280 26514 29336
rect 26570 29280 26575 29336
rect 22185 29278 26575 29280
rect 22185 29275 22251 29278
rect 26509 29275 26575 29278
rect 28993 29338 29059 29341
rect 32581 29338 32647 29341
rect 28993 29336 32647 29338
rect 28993 29280 28998 29336
rect 29054 29280 32586 29336
rect 32642 29280 32647 29336
rect 28993 29278 32647 29280
rect 28993 29275 29059 29278
rect 32581 29275 32647 29278
rect 9990 29140 9996 29204
rect 10060 29202 10066 29204
rect 10501 29202 10567 29205
rect 10060 29200 10567 29202
rect 10060 29144 10506 29200
rect 10562 29144 10567 29200
rect 10060 29142 10567 29144
rect 10060 29140 10066 29142
rect 10501 29139 10567 29142
rect 12985 29202 13051 29205
rect 16941 29202 17007 29205
rect 19149 29204 19215 29205
rect 19149 29202 19196 29204
rect 12985 29200 17007 29202
rect 12985 29144 12990 29200
rect 13046 29144 16946 29200
rect 17002 29144 17007 29200
rect 12985 29142 17007 29144
rect 19104 29200 19196 29202
rect 19104 29144 19154 29200
rect 19104 29142 19196 29144
rect 12985 29139 13051 29142
rect 16941 29139 17007 29142
rect 19149 29140 19196 29142
rect 19260 29140 19266 29204
rect 19333 29202 19399 29205
rect 36537 29202 36603 29205
rect 19333 29200 36603 29202
rect 19333 29144 19338 29200
rect 19394 29144 36542 29200
rect 36598 29144 36603 29200
rect 19333 29142 36603 29144
rect 19149 29139 19215 29140
rect 19333 29139 19399 29142
rect 36537 29139 36603 29142
rect 9673 29066 9739 29069
rect 10409 29066 10475 29069
rect 9673 29064 10475 29066
rect 9673 29008 9678 29064
rect 9734 29008 10414 29064
rect 10470 29008 10475 29064
rect 9673 29006 10475 29008
rect 9673 29003 9739 29006
rect 10409 29003 10475 29006
rect 12617 29066 12683 29069
rect 16246 29066 16252 29068
rect 12617 29064 16252 29066
rect 12617 29008 12622 29064
rect 12678 29008 16252 29064
rect 12617 29006 16252 29008
rect 12617 29003 12683 29006
rect 16246 29004 16252 29006
rect 16316 29004 16322 29068
rect 18454 29004 18460 29068
rect 18524 29066 18530 29068
rect 20846 29066 20852 29068
rect 18524 29006 20852 29066
rect 18524 29004 18530 29006
rect 20846 29004 20852 29006
rect 20916 29004 20922 29068
rect 22461 29066 22527 29069
rect 25221 29066 25287 29069
rect 22461 29064 25287 29066
rect 22461 29008 22466 29064
rect 22522 29008 25226 29064
rect 25282 29008 25287 29064
rect 22461 29006 25287 29008
rect 22461 29003 22527 29006
rect 25221 29003 25287 29006
rect 29821 29066 29887 29069
rect 31753 29066 31819 29069
rect 29821 29064 31819 29066
rect 29821 29008 29826 29064
rect 29882 29008 31758 29064
rect 31814 29008 31819 29064
rect 29821 29006 31819 29008
rect 29821 29003 29887 29006
rect 31753 29003 31819 29006
rect 10133 28930 10199 28933
rect 17309 28930 17375 28933
rect 10133 28928 17375 28930
rect 10133 28872 10138 28928
rect 10194 28872 17314 28928
rect 17370 28872 17375 28928
rect 10133 28870 17375 28872
rect 10133 28867 10199 28870
rect 17309 28867 17375 28870
rect 22461 28930 22527 28933
rect 26233 28930 26299 28933
rect 29637 28932 29703 28933
rect 29637 28930 29684 28932
rect 22461 28928 26299 28930
rect 22461 28872 22466 28928
rect 22522 28872 26238 28928
rect 26294 28872 26299 28928
rect 22461 28870 26299 28872
rect 29592 28928 29684 28930
rect 29592 28872 29642 28928
rect 29592 28870 29684 28872
rect 22461 28867 22527 28870
rect 26233 28867 26299 28870
rect 29637 28868 29684 28870
rect 29748 28868 29754 28932
rect 29637 28867 29703 28868
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 12157 28794 12223 28797
rect 16021 28794 16087 28797
rect 12157 28792 16087 28794
rect 12157 28736 12162 28792
rect 12218 28736 16026 28792
rect 16082 28736 16087 28792
rect 12157 28734 16087 28736
rect 12157 28731 12223 28734
rect 16021 28731 16087 28734
rect 17585 28794 17651 28797
rect 20805 28794 20871 28797
rect 21633 28794 21699 28797
rect 17585 28792 21699 28794
rect 17585 28736 17590 28792
rect 17646 28736 20810 28792
rect 20866 28736 21638 28792
rect 21694 28736 21699 28792
rect 17585 28734 21699 28736
rect 17585 28731 17651 28734
rect 20805 28731 20871 28734
rect 21633 28731 21699 28734
rect 24945 28794 25011 28797
rect 27153 28794 27219 28797
rect 24945 28792 27219 28794
rect 24945 28736 24950 28792
rect 25006 28736 27158 28792
rect 27214 28736 27219 28792
rect 24945 28734 27219 28736
rect 24945 28731 25011 28734
rect 27153 28731 27219 28734
rect 31017 28794 31083 28797
rect 31150 28794 31156 28796
rect 31017 28792 31156 28794
rect 31017 28736 31022 28792
rect 31078 28736 31156 28792
rect 31017 28734 31156 28736
rect 31017 28731 31083 28734
rect 31150 28732 31156 28734
rect 31220 28732 31226 28796
rect 20437 28658 20503 28661
rect 23422 28658 23428 28660
rect 20437 28656 23428 28658
rect 20437 28600 20442 28656
rect 20498 28600 23428 28656
rect 20437 28598 23428 28600
rect 20437 28595 20503 28598
rect 23422 28596 23428 28598
rect 23492 28596 23498 28660
rect 24301 28658 24367 28661
rect 27153 28658 27219 28661
rect 24301 28656 27219 28658
rect 24301 28600 24306 28656
rect 24362 28600 27158 28656
rect 27214 28600 27219 28656
rect 24301 28598 27219 28600
rect 24301 28595 24367 28598
rect 27153 28595 27219 28598
rect 41321 28658 41387 28661
rect 41720 28658 42520 28688
rect 41321 28656 42520 28658
rect 41321 28600 41326 28656
rect 41382 28600 42520 28656
rect 41321 28598 42520 28600
rect 41321 28595 41387 28598
rect 41720 28568 42520 28598
rect 21357 28522 21423 28525
rect 18094 28520 21423 28522
rect 18094 28464 21362 28520
rect 21418 28464 21423 28520
rect 18094 28462 21423 28464
rect 12249 28386 12315 28389
rect 16113 28386 16179 28389
rect 18094 28386 18154 28462
rect 21357 28459 21423 28462
rect 23565 28522 23631 28525
rect 31569 28522 31635 28525
rect 23565 28520 31635 28522
rect 23565 28464 23570 28520
rect 23626 28464 31574 28520
rect 31630 28464 31635 28520
rect 23565 28462 31635 28464
rect 23565 28459 23631 28462
rect 31569 28459 31635 28462
rect 12249 28384 18154 28386
rect 12249 28328 12254 28384
rect 12310 28328 16118 28384
rect 16174 28328 18154 28384
rect 12249 28326 18154 28328
rect 20161 28386 20227 28389
rect 24894 28386 24900 28388
rect 20161 28384 24900 28386
rect 20161 28328 20166 28384
rect 20222 28328 24900 28384
rect 20161 28326 24900 28328
rect 12249 28323 12315 28326
rect 16113 28323 16179 28326
rect 20161 28323 20227 28326
rect 24894 28324 24900 28326
rect 24964 28324 24970 28388
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 11513 28250 11579 28253
rect 14590 28250 14596 28252
rect 11513 28248 14596 28250
rect 11513 28192 11518 28248
rect 11574 28192 14596 28248
rect 11513 28190 14596 28192
rect 11513 28187 11579 28190
rect 14590 28188 14596 28190
rect 14660 28250 14666 28252
rect 18229 28250 18295 28253
rect 19241 28250 19307 28253
rect 14660 28190 17970 28250
rect 14660 28188 14666 28190
rect 9121 28114 9187 28117
rect 9254 28114 9260 28116
rect 9121 28112 9260 28114
rect 9121 28056 9126 28112
rect 9182 28056 9260 28112
rect 9121 28054 9260 28056
rect 9121 28051 9187 28054
rect 9254 28052 9260 28054
rect 9324 28052 9330 28116
rect 10869 28114 10935 28117
rect 12525 28114 12591 28117
rect 10869 28112 12591 28114
rect 10869 28056 10874 28112
rect 10930 28056 12530 28112
rect 12586 28056 12591 28112
rect 10869 28054 12591 28056
rect 10869 28051 10935 28054
rect 12525 28051 12591 28054
rect 15837 28116 15903 28117
rect 15837 28112 15884 28116
rect 15948 28114 15954 28116
rect 15837 28056 15842 28112
rect 15837 28052 15884 28056
rect 15948 28054 15994 28114
rect 15948 28052 15954 28054
rect 16614 28052 16620 28116
rect 16684 28114 16690 28116
rect 17769 28114 17835 28117
rect 16684 28112 17835 28114
rect 16684 28056 17774 28112
rect 17830 28056 17835 28112
rect 16684 28054 17835 28056
rect 17910 28114 17970 28190
rect 18229 28248 19307 28250
rect 18229 28192 18234 28248
rect 18290 28192 19246 28248
rect 19302 28192 19307 28248
rect 18229 28190 19307 28192
rect 18229 28187 18295 28190
rect 19241 28187 19307 28190
rect 20294 28188 20300 28252
rect 20364 28250 20370 28252
rect 20713 28250 20779 28253
rect 20364 28248 20779 28250
rect 20364 28192 20718 28248
rect 20774 28192 20779 28248
rect 20364 28190 20779 28192
rect 20364 28188 20370 28190
rect 20713 28187 20779 28190
rect 35157 28114 35223 28117
rect 17910 28112 35223 28114
rect 17910 28056 35162 28112
rect 35218 28056 35223 28112
rect 17910 28054 35223 28056
rect 16684 28052 16690 28054
rect 15837 28051 15903 28052
rect 17769 28051 17835 28054
rect 35157 28051 35223 28054
rect 0 27978 800 28008
rect 933 27978 999 27981
rect 0 27976 999 27978
rect 0 27920 938 27976
rect 994 27920 999 27976
rect 0 27918 999 27920
rect 0 27888 800 27918
rect 933 27915 999 27918
rect 11605 27978 11671 27981
rect 13721 27978 13787 27981
rect 11605 27976 13787 27978
rect 11605 27920 11610 27976
rect 11666 27920 13726 27976
rect 13782 27920 13787 27976
rect 11605 27918 13787 27920
rect 11605 27915 11671 27918
rect 13721 27915 13787 27918
rect 14641 27978 14707 27981
rect 22134 27978 22140 27980
rect 14641 27976 22140 27978
rect 14641 27920 14646 27976
rect 14702 27920 22140 27976
rect 14641 27918 22140 27920
rect 14641 27915 14707 27918
rect 22134 27916 22140 27918
rect 22204 27916 22210 27980
rect 24485 27978 24551 27981
rect 31937 27978 32003 27981
rect 24485 27976 32003 27978
rect 24485 27920 24490 27976
rect 24546 27920 31942 27976
rect 31998 27920 32003 27976
rect 24485 27918 32003 27920
rect 24485 27915 24551 27918
rect 31937 27915 32003 27918
rect 17861 27842 17927 27845
rect 23422 27842 23428 27844
rect 17861 27840 23428 27842
rect 17861 27784 17866 27840
rect 17922 27784 23428 27840
rect 17861 27782 23428 27784
rect 17861 27779 17927 27782
rect 23422 27780 23428 27782
rect 23492 27780 23498 27844
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 16246 27644 16252 27708
rect 16316 27706 16322 27708
rect 16665 27706 16731 27709
rect 16316 27704 16731 27706
rect 16316 27648 16670 27704
rect 16726 27648 16731 27704
rect 16316 27646 16731 27648
rect 16316 27644 16322 27646
rect 16665 27643 16731 27646
rect 18086 27644 18092 27708
rect 18156 27706 18162 27708
rect 18229 27706 18295 27709
rect 19517 27706 19583 27709
rect 18156 27704 18295 27706
rect 18156 27648 18234 27704
rect 18290 27648 18295 27704
rect 18156 27646 18295 27648
rect 18156 27644 18162 27646
rect 18229 27643 18295 27646
rect 19244 27704 19583 27706
rect 19244 27648 19522 27704
rect 19578 27648 19583 27704
rect 19244 27646 19583 27648
rect 11421 27570 11487 27573
rect 12750 27570 12756 27572
rect 11421 27568 12756 27570
rect 11421 27512 11426 27568
rect 11482 27512 12756 27568
rect 11421 27510 12756 27512
rect 11421 27507 11487 27510
rect 12750 27508 12756 27510
rect 12820 27508 12826 27572
rect 14641 27570 14707 27573
rect 18597 27570 18663 27573
rect 14641 27568 18663 27570
rect 14641 27512 14646 27568
rect 14702 27512 18602 27568
rect 18658 27512 18663 27568
rect 14641 27510 18663 27512
rect 19244 27570 19304 27646
rect 19517 27643 19583 27646
rect 21357 27706 21423 27709
rect 27797 27706 27863 27709
rect 21357 27704 27863 27706
rect 21357 27648 21362 27704
rect 21418 27648 27802 27704
rect 27858 27648 27863 27704
rect 21357 27646 27863 27648
rect 21357 27643 21423 27646
rect 27797 27643 27863 27646
rect 19885 27570 19951 27573
rect 19244 27568 19951 27570
rect 19244 27512 19890 27568
rect 19946 27512 19951 27568
rect 19244 27510 19951 27512
rect 14641 27507 14707 27510
rect 18597 27507 18663 27510
rect 19885 27507 19951 27510
rect 21081 27568 21147 27573
rect 21081 27512 21086 27568
rect 21142 27512 21147 27568
rect 21081 27507 21147 27512
rect 21357 27568 21423 27573
rect 26877 27572 26943 27573
rect 26877 27570 26924 27572
rect 21357 27512 21362 27568
rect 21418 27512 21423 27568
rect 21357 27507 21423 27512
rect 26832 27568 26924 27570
rect 26832 27512 26882 27568
rect 26832 27510 26924 27512
rect 26877 27508 26924 27510
rect 26988 27508 26994 27572
rect 26877 27507 26943 27508
rect 8845 27434 8911 27437
rect 9581 27434 9647 27437
rect 8845 27432 9647 27434
rect 8845 27376 8850 27432
rect 8906 27376 9586 27432
rect 9642 27376 9647 27432
rect 8845 27374 9647 27376
rect 8845 27371 8911 27374
rect 9581 27371 9647 27374
rect 15193 27434 15259 27437
rect 16481 27434 16547 27437
rect 21084 27434 21144 27507
rect 15193 27432 16547 27434
rect 15193 27376 15198 27432
rect 15254 27376 16486 27432
rect 16542 27376 16547 27432
rect 15193 27374 16547 27376
rect 15193 27371 15259 27374
rect 16481 27371 16547 27374
rect 16806 27374 21144 27434
rect 10317 27298 10383 27301
rect 16806 27298 16866 27374
rect 10317 27296 16866 27298
rect 10317 27240 10322 27296
rect 10378 27240 16866 27296
rect 10317 27238 16866 27240
rect 16941 27298 17007 27301
rect 18873 27298 18939 27301
rect 16941 27296 18939 27298
rect 16941 27240 16946 27296
rect 17002 27240 18878 27296
rect 18934 27240 18939 27296
rect 16941 27238 18939 27240
rect 10317 27235 10383 27238
rect 16941 27235 17007 27238
rect 18873 27235 18939 27238
rect 20989 27298 21055 27301
rect 21360 27298 21420 27507
rect 20989 27296 21420 27298
rect 20989 27240 20994 27296
rect 21050 27240 21420 27296
rect 20989 27238 21420 27240
rect 24945 27298 25011 27301
rect 26969 27298 27035 27301
rect 24945 27296 27035 27298
rect 24945 27240 24950 27296
rect 25006 27240 26974 27296
rect 27030 27240 27035 27296
rect 24945 27238 27035 27240
rect 20989 27235 21055 27238
rect 24945 27235 25011 27238
rect 26969 27235 27035 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 14641 27162 14707 27165
rect 17309 27162 17375 27165
rect 14641 27160 17375 27162
rect 14641 27104 14646 27160
rect 14702 27104 17314 27160
rect 17370 27104 17375 27160
rect 14641 27102 17375 27104
rect 14641 27099 14707 27102
rect 17309 27099 17375 27102
rect 22369 27162 22435 27165
rect 22921 27162 22987 27165
rect 22369 27160 26434 27162
rect 22369 27104 22374 27160
rect 22430 27104 22926 27160
rect 22982 27104 26434 27160
rect 22369 27102 26434 27104
rect 22369 27099 22435 27102
rect 22921 27099 22987 27102
rect 26374 27029 26434 27102
rect 26550 27100 26556 27164
rect 26620 27162 26626 27164
rect 27245 27162 27311 27165
rect 26620 27160 27311 27162
rect 26620 27104 27250 27160
rect 27306 27104 27311 27160
rect 26620 27102 27311 27104
rect 26620 27100 26626 27102
rect 27245 27099 27311 27102
rect 13261 27026 13327 27029
rect 18781 27026 18847 27029
rect 26141 27026 26207 27029
rect 13261 27024 26207 27026
rect 13261 26968 13266 27024
rect 13322 26968 18786 27024
rect 18842 26968 26146 27024
rect 26202 26968 26207 27024
rect 13261 26966 26207 26968
rect 26374 27026 26483 27029
rect 28717 27026 28783 27029
rect 26374 27024 28783 27026
rect 26374 26968 26422 27024
rect 26478 26968 28722 27024
rect 28778 26968 28783 27024
rect 26374 26966 28783 26968
rect 13261 26963 13327 26966
rect 18781 26963 18847 26966
rect 26141 26963 26207 26966
rect 26417 26963 26483 26966
rect 28717 26963 28783 26966
rect 10133 26890 10199 26893
rect 12566 26890 12572 26892
rect 10133 26888 12572 26890
rect 10133 26832 10138 26888
rect 10194 26832 12572 26888
rect 10133 26830 12572 26832
rect 10133 26827 10199 26830
rect 12566 26828 12572 26830
rect 12636 26828 12642 26892
rect 17953 26890 18019 26893
rect 24485 26890 24551 26893
rect 17953 26888 24551 26890
rect 17953 26832 17958 26888
rect 18014 26832 24490 26888
rect 24546 26832 24551 26888
rect 17953 26830 24551 26832
rect 17953 26827 18019 26830
rect 24485 26827 24551 26830
rect 28349 26892 28415 26893
rect 28349 26888 28396 26892
rect 28460 26890 28466 26892
rect 28349 26832 28354 26888
rect 28349 26828 28396 26832
rect 28460 26830 28506 26890
rect 28460 26828 28466 26830
rect 28349 26827 28415 26828
rect 12157 26754 12223 26757
rect 15142 26754 15148 26756
rect 12157 26752 15148 26754
rect 12157 26696 12162 26752
rect 12218 26696 15148 26752
rect 12157 26694 15148 26696
rect 12157 26691 12223 26694
rect 15142 26692 15148 26694
rect 15212 26692 15218 26756
rect 17033 26754 17099 26757
rect 24853 26754 24919 26757
rect 17033 26752 24919 26754
rect 17033 26696 17038 26752
rect 17094 26696 24858 26752
rect 24914 26696 24919 26752
rect 17033 26694 24919 26696
rect 17033 26691 17099 26694
rect 24853 26691 24919 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 9397 26618 9463 26621
rect 12893 26618 12959 26621
rect 9397 26616 12959 26618
rect 9397 26560 9402 26616
rect 9458 26560 12898 26616
rect 12954 26560 12959 26616
rect 9397 26558 12959 26560
rect 9397 26555 9463 26558
rect 12893 26555 12959 26558
rect 22737 26618 22803 26621
rect 25773 26618 25839 26621
rect 22737 26616 25839 26618
rect 22737 26560 22742 26616
rect 22798 26560 25778 26616
rect 25834 26560 25839 26616
rect 22737 26558 25839 26560
rect 22737 26555 22803 26558
rect 25773 26555 25839 26558
rect 12709 26482 12775 26485
rect 9998 26480 12775 26482
rect 9998 26424 12714 26480
rect 12770 26424 12775 26480
rect 9998 26422 12775 26424
rect 4981 26348 5047 26349
rect 4981 26344 5028 26348
rect 5092 26346 5098 26348
rect 9029 26346 9095 26349
rect 9998 26348 10058 26422
rect 12709 26419 12775 26422
rect 15377 26482 15443 26485
rect 15837 26482 15903 26485
rect 30005 26482 30071 26485
rect 15377 26480 30071 26482
rect 15377 26424 15382 26480
rect 15438 26424 15842 26480
rect 15898 26424 30010 26480
rect 30066 26424 30071 26480
rect 15377 26422 30071 26424
rect 15377 26419 15443 26422
rect 15837 26419 15903 26422
rect 30005 26419 30071 26422
rect 9990 26346 9996 26348
rect 4981 26288 4986 26344
rect 4981 26284 5028 26288
rect 5092 26286 5138 26346
rect 9029 26344 9996 26346
rect 9029 26288 9034 26344
rect 9090 26288 9996 26344
rect 9029 26286 9996 26288
rect 5092 26284 5098 26286
rect 4981 26283 5047 26284
rect 9029 26283 9095 26286
rect 9990 26284 9996 26286
rect 10060 26284 10066 26348
rect 15377 26346 15443 26349
rect 16481 26346 16547 26349
rect 27521 26346 27587 26349
rect 15377 26344 27587 26346
rect 15377 26288 15382 26344
rect 15438 26288 16486 26344
rect 16542 26288 27526 26344
rect 27582 26288 27587 26344
rect 15377 26286 27587 26288
rect 15377 26283 15443 26286
rect 16481 26283 16547 26286
rect 27521 26283 27587 26286
rect 8109 26210 8175 26213
rect 9397 26210 9463 26213
rect 8109 26208 9463 26210
rect 8109 26152 8114 26208
rect 8170 26152 9402 26208
rect 9458 26152 9463 26208
rect 8109 26150 9463 26152
rect 8109 26147 8175 26150
rect 9397 26147 9463 26150
rect 10358 26148 10364 26212
rect 10428 26210 10434 26212
rect 17309 26210 17375 26213
rect 10428 26208 17375 26210
rect 10428 26152 17314 26208
rect 17370 26152 17375 26208
rect 10428 26150 17375 26152
rect 10428 26148 10434 26150
rect 17309 26147 17375 26150
rect 17861 26210 17927 26213
rect 18505 26210 18571 26213
rect 17861 26208 18571 26210
rect 17861 26152 17866 26208
rect 17922 26152 18510 26208
rect 18566 26152 18571 26208
rect 17861 26150 18571 26152
rect 17861 26147 17927 26150
rect 18505 26147 18571 26150
rect 21081 26210 21147 26213
rect 24209 26210 24275 26213
rect 21081 26208 24275 26210
rect 21081 26152 21086 26208
rect 21142 26152 24214 26208
rect 24270 26152 24275 26208
rect 21081 26150 24275 26152
rect 21081 26147 21147 26150
rect 24209 26147 24275 26150
rect 26509 26212 26575 26213
rect 26509 26208 26556 26212
rect 26620 26210 26626 26212
rect 26509 26152 26514 26208
rect 26509 26148 26556 26152
rect 26620 26150 26666 26210
rect 26620 26148 26626 26150
rect 26509 26147 26575 26148
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 13169 26074 13235 26077
rect 18597 26074 18663 26077
rect 13169 26072 18663 26074
rect 13169 26016 13174 26072
rect 13230 26016 18602 26072
rect 18658 26016 18663 26072
rect 13169 26014 18663 26016
rect 13169 26011 13235 26014
rect 18597 26011 18663 26014
rect 18781 26076 18847 26077
rect 18781 26072 18828 26076
rect 18892 26074 18898 26076
rect 21265 26074 21331 26077
rect 28349 26074 28415 26077
rect 18781 26016 18786 26072
rect 18781 26012 18828 26016
rect 18892 26014 18938 26074
rect 21265 26072 28415 26074
rect 21265 26016 21270 26072
rect 21326 26016 28354 26072
rect 28410 26016 28415 26072
rect 21265 26014 28415 26016
rect 18892 26012 18898 26014
rect 18781 26011 18847 26012
rect 21265 26011 21331 26014
rect 28349 26011 28415 26014
rect 9857 25938 9923 25941
rect 30373 25938 30439 25941
rect 9857 25936 30439 25938
rect 9857 25880 9862 25936
rect 9918 25880 30378 25936
rect 30434 25880 30439 25936
rect 9857 25878 30439 25880
rect 9857 25875 9923 25878
rect 30373 25875 30439 25878
rect 30925 25938 30991 25941
rect 35525 25938 35591 25941
rect 30925 25936 35591 25938
rect 30925 25880 30930 25936
rect 30986 25880 35530 25936
rect 35586 25880 35591 25936
rect 30925 25878 35591 25880
rect 30925 25875 30991 25878
rect 35525 25875 35591 25878
rect 9581 25800 9647 25805
rect 9581 25744 9586 25800
rect 9642 25744 9647 25800
rect 9581 25739 9647 25744
rect 9765 25802 9831 25805
rect 21081 25802 21147 25805
rect 9765 25800 21147 25802
rect 9765 25744 9770 25800
rect 9826 25744 21086 25800
rect 21142 25744 21147 25800
rect 9765 25742 21147 25744
rect 9765 25739 9831 25742
rect 21081 25739 21147 25742
rect 21725 25802 21791 25805
rect 26969 25802 27035 25805
rect 21725 25800 27035 25802
rect 21725 25744 21730 25800
rect 21786 25744 26974 25800
rect 27030 25744 27035 25800
rect 21725 25742 27035 25744
rect 21725 25739 21791 25742
rect 26969 25739 27035 25742
rect 9584 25666 9644 25739
rect 10777 25666 10843 25669
rect 9584 25664 10843 25666
rect 9584 25608 10782 25664
rect 10838 25608 10843 25664
rect 9584 25606 10843 25608
rect 10777 25603 10843 25606
rect 16665 25666 16731 25669
rect 21265 25666 21331 25669
rect 16665 25664 21331 25666
rect 16665 25608 16670 25664
rect 16726 25608 21270 25664
rect 21326 25608 21331 25664
rect 16665 25606 21331 25608
rect 16665 25603 16731 25606
rect 21265 25603 21331 25606
rect 23381 25666 23447 25669
rect 28993 25666 29059 25669
rect 29729 25666 29795 25669
rect 23381 25664 29795 25666
rect 23381 25608 23386 25664
rect 23442 25608 28998 25664
rect 29054 25608 29734 25664
rect 29790 25608 29795 25664
rect 23381 25606 29795 25608
rect 23381 25603 23447 25606
rect 28993 25603 29059 25606
rect 29729 25603 29795 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 13629 25530 13695 25533
rect 14549 25530 14615 25533
rect 13629 25528 14615 25530
rect 13629 25472 13634 25528
rect 13690 25472 14554 25528
rect 14610 25472 14615 25528
rect 13629 25470 14615 25472
rect 13629 25467 13695 25470
rect 14549 25467 14615 25470
rect 15469 25530 15535 25533
rect 16021 25530 16087 25533
rect 15469 25528 16087 25530
rect 15469 25472 15474 25528
rect 15530 25472 16026 25528
rect 16082 25472 16087 25528
rect 15469 25470 16087 25472
rect 15469 25467 15535 25470
rect 16021 25467 16087 25470
rect 16757 25530 16823 25533
rect 17861 25530 17927 25533
rect 16757 25528 17927 25530
rect 16757 25472 16762 25528
rect 16818 25472 17866 25528
rect 17922 25472 17927 25528
rect 16757 25470 17927 25472
rect 16757 25467 16823 25470
rect 17861 25467 17927 25470
rect 18505 25530 18571 25533
rect 24025 25530 24091 25533
rect 18505 25528 24091 25530
rect 18505 25472 18510 25528
rect 18566 25472 24030 25528
rect 24086 25472 24091 25528
rect 18505 25470 24091 25472
rect 18505 25467 18571 25470
rect 24025 25467 24091 25470
rect 29177 25530 29243 25533
rect 29177 25528 29378 25530
rect 29177 25472 29182 25528
rect 29238 25472 29378 25528
rect 29177 25470 29378 25472
rect 29177 25467 29243 25470
rect 6821 25394 6887 25397
rect 26049 25394 26115 25397
rect 6821 25392 26115 25394
rect 6821 25336 6826 25392
rect 6882 25336 26054 25392
rect 26110 25336 26115 25392
rect 6821 25334 26115 25336
rect 6821 25331 6887 25334
rect 26049 25331 26115 25334
rect 29085 25394 29151 25397
rect 29085 25392 29194 25394
rect 29085 25336 29090 25392
rect 29146 25336 29194 25392
rect 29085 25331 29194 25336
rect 9029 25258 9095 25261
rect 9489 25258 9555 25261
rect 9029 25256 9555 25258
rect 9029 25200 9034 25256
rect 9090 25200 9494 25256
rect 9550 25200 9555 25256
rect 9029 25198 9555 25200
rect 9029 25195 9095 25198
rect 9489 25195 9555 25198
rect 11329 25258 11395 25261
rect 24393 25258 24459 25261
rect 11329 25256 24459 25258
rect 11329 25200 11334 25256
rect 11390 25200 24398 25256
rect 24454 25200 24459 25256
rect 11329 25198 24459 25200
rect 11329 25195 11395 25198
rect 24393 25195 24459 25198
rect 29134 25125 29194 25331
rect 29318 25261 29378 25470
rect 29269 25256 29378 25261
rect 29269 25200 29274 25256
rect 29330 25200 29378 25256
rect 29269 25198 29378 25200
rect 29269 25195 29335 25198
rect 17033 25122 17099 25125
rect 18086 25122 18092 25124
rect 17033 25120 18092 25122
rect 17033 25064 17038 25120
rect 17094 25064 18092 25120
rect 17033 25062 18092 25064
rect 17033 25059 17099 25062
rect 18086 25060 18092 25062
rect 18156 25060 18162 25124
rect 29085 25120 29194 25125
rect 29085 25064 29090 25120
rect 29146 25064 29194 25120
rect 29085 25062 29194 25064
rect 29085 25059 29151 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 13169 24986 13235 24989
rect 15009 24986 15075 24989
rect 13169 24984 15075 24986
rect 13169 24928 13174 24984
rect 13230 24928 15014 24984
rect 15070 24928 15075 24984
rect 13169 24926 15075 24928
rect 13169 24923 13235 24926
rect 15009 24923 15075 24926
rect 9213 24850 9279 24853
rect 11646 24850 11652 24852
rect 9213 24848 11652 24850
rect 9213 24792 9218 24848
rect 9274 24792 11652 24848
rect 9213 24790 11652 24792
rect 9213 24787 9279 24790
rect 11646 24788 11652 24790
rect 11716 24788 11722 24852
rect 14825 24850 14891 24853
rect 15653 24850 15719 24853
rect 14825 24848 15719 24850
rect 14825 24792 14830 24848
rect 14886 24792 15658 24848
rect 15714 24792 15719 24848
rect 14825 24790 15719 24792
rect 14825 24787 14891 24790
rect 15653 24787 15719 24790
rect 18229 24850 18295 24853
rect 21357 24850 21423 24853
rect 18229 24848 21423 24850
rect 18229 24792 18234 24848
rect 18290 24792 21362 24848
rect 21418 24792 21423 24848
rect 18229 24790 21423 24792
rect 18229 24787 18295 24790
rect 21357 24787 21423 24790
rect 24669 24850 24735 24853
rect 29269 24852 29335 24853
rect 25814 24850 25820 24852
rect 24669 24848 25820 24850
rect 24669 24792 24674 24848
rect 24730 24792 25820 24848
rect 24669 24790 25820 24792
rect 24669 24787 24735 24790
rect 25814 24788 25820 24790
rect 25884 24788 25890 24852
rect 29269 24850 29316 24852
rect 29224 24848 29316 24850
rect 29224 24792 29274 24848
rect 29224 24790 29316 24792
rect 29269 24788 29316 24790
rect 29380 24788 29386 24852
rect 29269 24787 29335 24788
rect 8385 24714 8451 24717
rect 9305 24714 9371 24717
rect 8385 24712 9371 24714
rect 8385 24656 8390 24712
rect 8446 24656 9310 24712
rect 9366 24656 9371 24712
rect 8385 24654 9371 24656
rect 8385 24651 8451 24654
rect 9305 24651 9371 24654
rect 12525 24714 12591 24717
rect 13905 24714 13971 24717
rect 15193 24714 15259 24717
rect 18229 24714 18295 24717
rect 12525 24712 18295 24714
rect 12525 24656 12530 24712
rect 12586 24656 13910 24712
rect 13966 24656 15198 24712
rect 15254 24656 18234 24712
rect 18290 24656 18295 24712
rect 12525 24654 18295 24656
rect 12525 24651 12591 24654
rect 13905 24651 13971 24654
rect 15193 24651 15259 24654
rect 18229 24651 18295 24654
rect 20713 24714 20779 24717
rect 23749 24714 23815 24717
rect 24894 24714 24900 24716
rect 20713 24712 23674 24714
rect 20713 24656 20718 24712
rect 20774 24656 23674 24712
rect 20713 24654 23674 24656
rect 20713 24651 20779 24654
rect 14825 24578 14891 24581
rect 18413 24578 18479 24581
rect 14825 24576 18479 24578
rect 14825 24520 14830 24576
rect 14886 24520 18418 24576
rect 18474 24520 18479 24576
rect 14825 24518 18479 24520
rect 14825 24515 14891 24518
rect 18413 24515 18479 24518
rect 18689 24578 18755 24581
rect 22737 24580 22803 24581
rect 22686 24578 22692 24580
rect 18689 24576 22386 24578
rect 18689 24520 18694 24576
rect 18750 24520 22386 24576
rect 18689 24518 22386 24520
rect 22646 24518 22692 24578
rect 22756 24576 22803 24580
rect 22798 24520 22803 24576
rect 18689 24515 18755 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 11513 24442 11579 24445
rect 12985 24442 13051 24445
rect 11513 24440 13051 24442
rect 11513 24384 11518 24440
rect 11574 24384 12990 24440
rect 13046 24384 13051 24440
rect 11513 24382 13051 24384
rect 11513 24379 11579 24382
rect 12985 24379 13051 24382
rect 15193 24442 15259 24445
rect 17033 24442 17099 24445
rect 22185 24442 22251 24445
rect 15193 24440 16314 24442
rect 15193 24384 15198 24440
rect 15254 24384 16314 24440
rect 15193 24382 16314 24384
rect 15193 24379 15259 24382
rect 15929 24306 15995 24309
rect 16062 24306 16068 24308
rect 15929 24304 16068 24306
rect 15929 24248 15934 24304
rect 15990 24248 16068 24304
rect 15929 24246 16068 24248
rect 15929 24243 15995 24246
rect 16062 24244 16068 24246
rect 16132 24244 16138 24308
rect 16254 24306 16314 24382
rect 17033 24440 22251 24442
rect 17033 24384 17038 24440
rect 17094 24384 22190 24440
rect 22246 24384 22251 24440
rect 17033 24382 22251 24384
rect 22326 24442 22386 24518
rect 22686 24516 22692 24518
rect 22756 24516 22803 24520
rect 23614 24578 23674 24654
rect 23749 24712 24900 24714
rect 23749 24656 23754 24712
rect 23810 24656 24900 24712
rect 23749 24654 24900 24656
rect 23749 24651 23815 24654
rect 24894 24652 24900 24654
rect 24964 24652 24970 24716
rect 25262 24652 25268 24716
rect 25332 24714 25338 24716
rect 30925 24714 30991 24717
rect 25332 24712 30991 24714
rect 25332 24656 30930 24712
rect 30986 24656 30991 24712
rect 25332 24654 30991 24656
rect 25332 24652 25338 24654
rect 30925 24651 30991 24654
rect 23841 24578 23907 24581
rect 25405 24578 25471 24581
rect 23614 24576 25471 24578
rect 23614 24520 23846 24576
rect 23902 24520 25410 24576
rect 25466 24520 25471 24576
rect 23614 24518 25471 24520
rect 22737 24515 22803 24516
rect 23841 24515 23907 24518
rect 25405 24515 25471 24518
rect 41321 24578 41387 24581
rect 41720 24578 42520 24608
rect 41321 24576 42520 24578
rect 41321 24520 41326 24576
rect 41382 24520 42520 24576
rect 41321 24518 42520 24520
rect 41321 24515 41387 24518
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 41720 24488 42520 24518
rect 34930 24447 35246 24448
rect 25129 24442 25195 24445
rect 22326 24440 25195 24442
rect 22326 24384 25134 24440
rect 25190 24384 25195 24440
rect 22326 24382 25195 24384
rect 17033 24379 17099 24382
rect 22185 24379 22251 24382
rect 25129 24379 25195 24382
rect 20621 24306 20687 24309
rect 16254 24304 20687 24306
rect 16254 24248 20626 24304
rect 20682 24248 20687 24304
rect 16254 24246 20687 24248
rect 20621 24243 20687 24246
rect 21173 24306 21239 24309
rect 22369 24306 22435 24309
rect 27245 24306 27311 24309
rect 30557 24308 30623 24309
rect 30557 24306 30604 24308
rect 21173 24304 27311 24306
rect 21173 24248 21178 24304
rect 21234 24248 22374 24304
rect 22430 24248 27250 24304
rect 27306 24248 27311 24304
rect 21173 24246 27311 24248
rect 30476 24304 30604 24306
rect 30668 24306 30674 24308
rect 31753 24306 31819 24309
rect 30668 24304 31819 24306
rect 30476 24248 30562 24304
rect 30668 24248 31758 24304
rect 31814 24248 31819 24304
rect 30476 24246 30604 24248
rect 21173 24243 21239 24246
rect 22369 24243 22435 24246
rect 27245 24243 27311 24246
rect 30557 24244 30604 24246
rect 30668 24246 31819 24248
rect 30668 24244 30674 24246
rect 30557 24243 30623 24244
rect 31753 24243 31819 24246
rect 11053 24170 11119 24173
rect 20069 24170 20135 24173
rect 20345 24172 20411 24173
rect 11053 24168 20135 24170
rect 11053 24112 11058 24168
rect 11114 24112 20074 24168
rect 20130 24112 20135 24168
rect 11053 24110 20135 24112
rect 11053 24107 11119 24110
rect 20069 24107 20135 24110
rect 20294 24108 20300 24172
rect 20364 24170 20411 24172
rect 20897 24170 20963 24173
rect 21081 24170 21147 24173
rect 20364 24168 20456 24170
rect 20406 24112 20456 24168
rect 20364 24110 20456 24112
rect 20897 24168 21147 24170
rect 20897 24112 20902 24168
rect 20958 24112 21086 24168
rect 21142 24112 21147 24168
rect 20897 24110 21147 24112
rect 20364 24108 20411 24110
rect 20345 24107 20411 24108
rect 20897 24107 20963 24110
rect 21081 24107 21147 24110
rect 27061 24170 27127 24173
rect 27705 24170 27771 24173
rect 27061 24168 27771 24170
rect 27061 24112 27066 24168
rect 27122 24112 27710 24168
rect 27766 24112 27771 24168
rect 27061 24110 27771 24112
rect 27061 24107 27127 24110
rect 27705 24107 27771 24110
rect 15653 24034 15719 24037
rect 16614 24034 16620 24036
rect 15653 24032 16620 24034
rect 15653 23976 15658 24032
rect 15714 23976 16620 24032
rect 15653 23974 16620 23976
rect 15653 23971 15719 23974
rect 16614 23972 16620 23974
rect 16684 23972 16690 24036
rect 17125 24034 17191 24037
rect 18505 24034 18571 24037
rect 17125 24032 18571 24034
rect 17125 23976 17130 24032
rect 17186 23976 18510 24032
rect 18566 23976 18571 24032
rect 17125 23974 18571 23976
rect 17125 23971 17191 23974
rect 18505 23971 18571 23974
rect 20805 24034 20871 24037
rect 25497 24034 25563 24037
rect 20805 24032 25563 24034
rect 20805 23976 20810 24032
rect 20866 23976 25502 24032
rect 25558 23976 25563 24032
rect 20805 23974 25563 23976
rect 20805 23971 20871 23974
rect 25497 23971 25563 23974
rect 19570 23968 19886 23969
rect 0 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 933 23898 999 23901
rect 0 23896 999 23898
rect 0 23840 938 23896
rect 994 23840 999 23896
rect 0 23838 999 23840
rect 0 23808 800 23838
rect 933 23835 999 23838
rect 12525 23898 12591 23901
rect 13445 23898 13511 23901
rect 16665 23898 16731 23901
rect 12525 23896 16731 23898
rect 12525 23840 12530 23896
rect 12586 23840 13450 23896
rect 13506 23840 16670 23896
rect 16726 23840 16731 23896
rect 12525 23838 16731 23840
rect 12525 23835 12591 23838
rect 13445 23835 13511 23838
rect 16665 23835 16731 23838
rect 20437 23898 20503 23901
rect 26325 23898 26391 23901
rect 20437 23896 26391 23898
rect 20437 23840 20442 23896
rect 20498 23840 26330 23896
rect 26386 23840 26391 23896
rect 20437 23838 26391 23840
rect 20437 23835 20503 23838
rect 26325 23835 26391 23838
rect 10593 23762 10659 23765
rect 18086 23762 18092 23764
rect 10593 23760 18092 23762
rect 10593 23704 10598 23760
rect 10654 23704 18092 23760
rect 10593 23702 18092 23704
rect 10593 23699 10659 23702
rect 18086 23700 18092 23702
rect 18156 23762 18162 23764
rect 19057 23762 19123 23765
rect 21173 23762 21239 23765
rect 23013 23762 23079 23765
rect 26877 23762 26943 23765
rect 27521 23762 27587 23765
rect 18156 23760 19123 23762
rect 18156 23704 19062 23760
rect 19118 23704 19123 23760
rect 18156 23702 19123 23704
rect 18156 23700 18162 23702
rect 19057 23699 19123 23702
rect 19290 23760 22938 23762
rect 19290 23704 21178 23760
rect 21234 23704 22938 23760
rect 19290 23702 22938 23704
rect 14549 23626 14615 23629
rect 19290 23626 19350 23702
rect 21173 23699 21239 23702
rect 14549 23624 19350 23626
rect 14549 23568 14554 23624
rect 14610 23568 19350 23624
rect 14549 23566 19350 23568
rect 19885 23626 19951 23629
rect 21081 23626 21147 23629
rect 19885 23624 21147 23626
rect 19885 23568 19890 23624
rect 19946 23568 21086 23624
rect 21142 23568 21147 23624
rect 19885 23566 21147 23568
rect 22878 23626 22938 23702
rect 23013 23760 27587 23762
rect 23013 23704 23018 23760
rect 23074 23704 26882 23760
rect 26938 23704 27526 23760
rect 27582 23704 27587 23760
rect 23013 23702 27587 23704
rect 23013 23699 23079 23702
rect 26877 23699 26943 23702
rect 27521 23699 27587 23702
rect 24577 23626 24643 23629
rect 26325 23626 26391 23629
rect 22878 23624 26391 23626
rect 22878 23568 24582 23624
rect 24638 23568 26330 23624
rect 26386 23568 26391 23624
rect 22878 23566 26391 23568
rect 14549 23563 14615 23566
rect 19885 23563 19951 23566
rect 21081 23563 21147 23566
rect 24577 23563 24643 23566
rect 26325 23563 26391 23566
rect 8477 23490 8543 23493
rect 12382 23490 12388 23492
rect 8477 23488 12388 23490
rect 8477 23432 8482 23488
rect 8538 23432 12388 23488
rect 8477 23430 12388 23432
rect 8477 23427 8543 23430
rect 12382 23428 12388 23430
rect 12452 23428 12458 23492
rect 16021 23490 16087 23493
rect 17401 23490 17467 23493
rect 20621 23490 20687 23493
rect 16021 23488 20687 23490
rect 16021 23432 16026 23488
rect 16082 23432 17406 23488
rect 17462 23432 20626 23488
rect 20682 23432 20687 23488
rect 16021 23430 20687 23432
rect 16021 23427 16087 23430
rect 17401 23427 17467 23430
rect 20621 23427 20687 23430
rect 20805 23490 20871 23493
rect 21398 23490 21404 23492
rect 20805 23488 21404 23490
rect 20805 23432 20810 23488
rect 20866 23432 21404 23488
rect 20805 23430 21404 23432
rect 20805 23427 20871 23430
rect 21398 23428 21404 23430
rect 21468 23428 21474 23492
rect 27429 23490 27495 23493
rect 29126 23490 29132 23492
rect 27429 23488 29132 23490
rect 27429 23432 27434 23488
rect 27490 23432 29132 23488
rect 27429 23430 29132 23432
rect 27429 23427 27495 23430
rect 29126 23428 29132 23430
rect 29196 23428 29202 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 15009 23354 15075 23357
rect 22001 23354 22067 23357
rect 15009 23352 22067 23354
rect 15009 23296 15014 23352
rect 15070 23296 22006 23352
rect 22062 23296 22067 23352
rect 15009 23294 22067 23296
rect 15009 23291 15075 23294
rect 22001 23291 22067 23294
rect 9213 23218 9279 23221
rect 9438 23218 9444 23220
rect 9213 23216 9444 23218
rect 9213 23160 9218 23216
rect 9274 23160 9444 23216
rect 9213 23158 9444 23160
rect 9213 23155 9279 23158
rect 9438 23156 9444 23158
rect 9508 23156 9514 23220
rect 15193 23218 15259 23221
rect 20989 23218 21055 23221
rect 15193 23216 21055 23218
rect 15193 23160 15198 23216
rect 15254 23160 20994 23216
rect 21050 23160 21055 23216
rect 15193 23158 21055 23160
rect 15193 23155 15259 23158
rect 20989 23155 21055 23158
rect 16113 23082 16179 23085
rect 20621 23082 20687 23085
rect 21081 23084 21147 23085
rect 16113 23080 20687 23082
rect 16113 23024 16118 23080
rect 16174 23024 20626 23080
rect 20682 23024 20687 23080
rect 16113 23022 20687 23024
rect 16113 23019 16179 23022
rect 20621 23019 20687 23022
rect 21030 23020 21036 23084
rect 21100 23082 21147 23084
rect 21100 23080 21192 23082
rect 21142 23024 21192 23080
rect 21100 23022 21192 23024
rect 21100 23020 21147 23022
rect 21081 23019 21147 23020
rect 16941 22946 17007 22949
rect 17902 22946 17908 22948
rect 16941 22944 17908 22946
rect 16941 22888 16946 22944
rect 17002 22888 17908 22944
rect 16941 22886 17908 22888
rect 16941 22883 17007 22886
rect 17902 22884 17908 22886
rect 17972 22884 17978 22948
rect 18689 22946 18755 22949
rect 19241 22948 19307 22949
rect 18822 22946 18828 22948
rect 18689 22944 18828 22946
rect 18689 22888 18694 22944
rect 18750 22888 18828 22944
rect 18689 22886 18828 22888
rect 18689 22883 18755 22886
rect 18822 22884 18828 22886
rect 18892 22884 18898 22948
rect 19190 22946 19196 22948
rect 19150 22886 19196 22946
rect 19260 22944 19307 22948
rect 19302 22888 19307 22944
rect 19190 22884 19196 22886
rect 19260 22884 19307 22888
rect 19241 22883 19307 22884
rect 20069 22946 20135 22949
rect 30281 22946 30347 22949
rect 20069 22944 30347 22946
rect 20069 22888 20074 22944
rect 20130 22888 30286 22944
rect 30342 22888 30347 22944
rect 20069 22886 30347 22888
rect 20069 22883 20135 22886
rect 30281 22883 30347 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 11421 22810 11487 22813
rect 16113 22810 16179 22813
rect 11421 22808 16179 22810
rect 11421 22752 11426 22808
rect 11482 22752 16118 22808
rect 16174 22752 16179 22808
rect 11421 22750 16179 22752
rect 11421 22747 11487 22750
rect 16113 22747 16179 22750
rect 17585 22810 17651 22813
rect 18781 22810 18847 22813
rect 17585 22808 18847 22810
rect 17585 22752 17590 22808
rect 17646 22752 18786 22808
rect 18842 22752 18847 22808
rect 17585 22750 18847 22752
rect 17585 22747 17651 22750
rect 18781 22747 18847 22750
rect 20345 22810 20411 22813
rect 23381 22810 23447 22813
rect 20345 22808 23447 22810
rect 20345 22752 20350 22808
rect 20406 22752 23386 22808
rect 23442 22752 23447 22808
rect 20345 22750 23447 22752
rect 20345 22747 20411 22750
rect 23381 22747 23447 22750
rect 15101 22674 15167 22677
rect 17401 22674 17467 22677
rect 15101 22672 17467 22674
rect 15101 22616 15106 22672
rect 15162 22616 17406 22672
rect 17462 22616 17467 22672
rect 15101 22614 17467 22616
rect 15101 22611 15167 22614
rect 17401 22611 17467 22614
rect 17585 22674 17651 22677
rect 19149 22674 19215 22677
rect 23841 22674 23907 22677
rect 24853 22674 24919 22677
rect 41045 22674 41111 22677
rect 17585 22672 24919 22674
rect 17585 22616 17590 22672
rect 17646 22616 19154 22672
rect 19210 22616 23846 22672
rect 23902 22616 24858 22672
rect 24914 22616 24919 22672
rect 17585 22614 24919 22616
rect 17585 22611 17651 22614
rect 19149 22611 19215 22614
rect 23841 22611 23907 22614
rect 24853 22611 24919 22614
rect 31710 22672 41111 22674
rect 31710 22616 41050 22672
rect 41106 22616 41111 22672
rect 31710 22614 41111 22616
rect 12709 22538 12775 22541
rect 20069 22538 20135 22541
rect 12709 22536 20135 22538
rect 12709 22480 12714 22536
rect 12770 22480 20074 22536
rect 20130 22480 20135 22536
rect 12709 22478 20135 22480
rect 12709 22475 12775 22478
rect 20069 22475 20135 22478
rect 20345 22538 20411 22541
rect 31710 22538 31770 22614
rect 41045 22611 41111 22614
rect 20345 22536 31770 22538
rect 20345 22480 20350 22536
rect 20406 22480 31770 22536
rect 20345 22478 31770 22480
rect 20345 22475 20411 22478
rect 8569 22402 8635 22405
rect 27613 22402 27679 22405
rect 8569 22400 27679 22402
rect 8569 22344 8574 22400
rect 8630 22344 27618 22400
rect 27674 22344 27679 22400
rect 8569 22342 27679 22344
rect 8569 22339 8635 22342
rect 27613 22339 27679 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 13077 22266 13143 22269
rect 17585 22266 17651 22269
rect 13077 22264 17651 22266
rect 13077 22208 13082 22264
rect 13138 22208 17590 22264
rect 17646 22208 17651 22264
rect 13077 22206 17651 22208
rect 13077 22203 13143 22206
rect 17585 22203 17651 22206
rect 17953 22266 18019 22269
rect 18413 22266 18479 22269
rect 17953 22264 18479 22266
rect 17953 22208 17958 22264
rect 18014 22208 18418 22264
rect 18474 22208 18479 22264
rect 17953 22206 18479 22208
rect 17953 22203 18019 22206
rect 18413 22203 18479 22206
rect 18597 22266 18663 22269
rect 23105 22266 23171 22269
rect 18597 22264 23171 22266
rect 18597 22208 18602 22264
rect 18658 22208 23110 22264
rect 23166 22208 23171 22264
rect 18597 22206 23171 22208
rect 18597 22203 18663 22206
rect 23105 22203 23171 22206
rect 23473 22266 23539 22269
rect 24853 22266 24919 22269
rect 23473 22264 24919 22266
rect 23473 22208 23478 22264
rect 23534 22208 24858 22264
rect 24914 22208 24919 22264
rect 23473 22206 24919 22208
rect 23473 22203 23539 22206
rect 24853 22203 24919 22206
rect 12985 22130 13051 22133
rect 13353 22130 13419 22133
rect 21081 22130 21147 22133
rect 12985 22128 13419 22130
rect 12985 22072 12990 22128
rect 13046 22072 13358 22128
rect 13414 22072 13419 22128
rect 12985 22070 13419 22072
rect 12985 22067 13051 22070
rect 13353 22067 13419 22070
rect 15150 22128 21147 22130
rect 15150 22072 21086 22128
rect 21142 22072 21147 22128
rect 15150 22070 21147 22072
rect 8201 21994 8267 21997
rect 15150 21994 15210 22070
rect 21081 22067 21147 22070
rect 19609 21994 19675 21997
rect 8201 21992 15210 21994
rect 8201 21936 8206 21992
rect 8262 21936 15210 21992
rect 8201 21934 15210 21936
rect 19382 21992 19675 21994
rect 19382 21936 19614 21992
rect 19670 21936 19675 21992
rect 19382 21934 19675 21936
rect 8201 21931 8267 21934
rect 11421 21860 11487 21861
rect 11421 21856 11468 21860
rect 11532 21858 11538 21860
rect 11421 21800 11426 21856
rect 11421 21796 11468 21800
rect 11532 21798 11578 21858
rect 11532 21796 11538 21798
rect 12382 21796 12388 21860
rect 12452 21858 12458 21860
rect 12985 21858 13051 21861
rect 12452 21856 13051 21858
rect 12452 21800 12990 21856
rect 13046 21800 13051 21856
rect 12452 21798 13051 21800
rect 12452 21796 12458 21798
rect 11421 21795 11487 21796
rect 12985 21795 13051 21798
rect 15653 21858 15719 21861
rect 19382 21858 19442 21934
rect 19609 21931 19675 21934
rect 21081 21994 21147 21997
rect 27521 21994 27587 21997
rect 21081 21992 27587 21994
rect 21081 21936 21086 21992
rect 21142 21936 27526 21992
rect 27582 21936 27587 21992
rect 21081 21934 27587 21936
rect 21081 21931 21147 21934
rect 27521 21931 27587 21934
rect 15653 21856 19442 21858
rect 15653 21800 15658 21856
rect 15714 21800 19442 21856
rect 15653 21798 19442 21800
rect 15653 21795 15719 21798
rect 22134 21796 22140 21860
rect 22204 21858 22210 21860
rect 30557 21858 30623 21861
rect 22204 21856 30623 21858
rect 22204 21800 30562 21856
rect 30618 21800 30623 21856
rect 22204 21798 30623 21800
rect 22204 21796 22210 21798
rect 30557 21795 30623 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 10777 21722 10843 21725
rect 19057 21722 19123 21725
rect 24117 21722 24183 21725
rect 27889 21722 27955 21725
rect 10777 21720 19123 21722
rect 10777 21664 10782 21720
rect 10838 21664 19062 21720
rect 19118 21664 19123 21720
rect 10777 21662 19123 21664
rect 10777 21659 10843 21662
rect 19057 21659 19123 21662
rect 20118 21720 27955 21722
rect 20118 21664 24122 21720
rect 24178 21664 27894 21720
rect 27950 21664 27955 21720
rect 20118 21662 27955 21664
rect 4521 21586 4587 21589
rect 7097 21586 7163 21589
rect 4521 21584 7163 21586
rect 4521 21528 4526 21584
rect 4582 21528 7102 21584
rect 7158 21528 7163 21584
rect 4521 21526 7163 21528
rect 4521 21523 4587 21526
rect 7097 21523 7163 21526
rect 8385 21586 8451 21589
rect 20118 21586 20178 21662
rect 24117 21659 24183 21662
rect 27889 21659 27955 21662
rect 8385 21584 20178 21586
rect 8385 21528 8390 21584
rect 8446 21528 20178 21584
rect 8385 21526 20178 21528
rect 8385 21523 8451 21526
rect 20478 21524 20484 21588
rect 20548 21586 20554 21588
rect 20621 21586 20687 21589
rect 20548 21584 20687 21586
rect 20548 21528 20626 21584
rect 20682 21528 20687 21584
rect 20548 21526 20687 21528
rect 20548 21524 20554 21526
rect 20621 21523 20687 21526
rect 24526 21524 24532 21588
rect 24596 21586 24602 21588
rect 24853 21586 24919 21589
rect 24596 21584 24919 21586
rect 24596 21528 24858 21584
rect 24914 21528 24919 21584
rect 24596 21526 24919 21528
rect 24596 21524 24602 21526
rect 24853 21523 24919 21526
rect 10593 21450 10659 21453
rect 25681 21450 25747 21453
rect 10593 21448 25747 21450
rect 10593 21392 10598 21448
rect 10654 21392 25686 21448
rect 25742 21392 25747 21448
rect 10593 21390 25747 21392
rect 10593 21387 10659 21390
rect 25681 21387 25747 21390
rect 14733 21316 14799 21317
rect 14733 21314 14780 21316
rect 14652 21312 14780 21314
rect 14844 21314 14850 21316
rect 21081 21314 21147 21317
rect 14844 21312 21147 21314
rect 14652 21256 14738 21312
rect 14844 21256 21086 21312
rect 21142 21256 21147 21312
rect 14652 21254 14780 21256
rect 14733 21252 14780 21254
rect 14844 21254 21147 21256
rect 14844 21252 14850 21254
rect 14733 21251 14799 21252
rect 21081 21251 21147 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 15878 21116 15884 21180
rect 15948 21178 15954 21180
rect 16021 21178 16087 21181
rect 18137 21180 18203 21181
rect 18086 21178 18092 21180
rect 15948 21176 16087 21178
rect 15948 21120 16026 21176
rect 16082 21120 16087 21176
rect 15948 21118 16087 21120
rect 18046 21118 18092 21178
rect 18156 21176 18203 21180
rect 18198 21120 18203 21176
rect 15948 21116 15954 21118
rect 16021 21115 16087 21118
rect 18086 21116 18092 21118
rect 18156 21116 18203 21120
rect 18137 21115 18203 21116
rect 7557 21042 7623 21045
rect 29545 21042 29611 21045
rect 7557 21040 29611 21042
rect 7557 20984 7562 21040
rect 7618 20984 29550 21040
rect 29606 20984 29611 21040
rect 7557 20982 29611 20984
rect 7557 20979 7623 20982
rect 19885 20906 19951 20909
rect 26325 20908 26391 20909
rect 20294 20906 20300 20908
rect 19885 20904 20300 20906
rect 19885 20848 19890 20904
rect 19946 20848 20300 20904
rect 19885 20846 20300 20848
rect 19885 20843 19951 20846
rect 20294 20844 20300 20846
rect 20364 20844 20370 20908
rect 26325 20906 26372 20908
rect 26280 20904 26372 20906
rect 26280 20848 26330 20904
rect 26280 20846 26372 20848
rect 26325 20844 26372 20846
rect 26436 20844 26442 20908
rect 26325 20843 26391 20844
rect 5165 20772 5231 20773
rect 5165 20770 5212 20772
rect 5120 20768 5212 20770
rect 5120 20712 5170 20768
rect 5120 20710 5212 20712
rect 5165 20708 5212 20710
rect 5276 20708 5282 20772
rect 24710 20708 24716 20772
rect 24780 20770 24786 20772
rect 26325 20770 26391 20773
rect 24780 20768 26391 20770
rect 24780 20712 26330 20768
rect 26386 20712 26391 20768
rect 24780 20710 26391 20712
rect 24780 20708 24786 20710
rect 5165 20707 5231 20708
rect 26325 20707 26391 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 12566 20572 12572 20636
rect 12636 20634 12642 20636
rect 12893 20634 12959 20637
rect 28950 20636 29010 20982
rect 29545 20979 29611 20982
rect 12636 20632 12959 20634
rect 12636 20576 12898 20632
rect 12954 20576 12959 20632
rect 12636 20574 12959 20576
rect 12636 20572 12642 20574
rect 12893 20571 12959 20574
rect 15142 20572 15148 20636
rect 15212 20572 15218 20636
rect 28942 20572 28948 20636
rect 29012 20572 29018 20636
rect 35249 20634 35315 20637
rect 36353 20634 36419 20637
rect 35249 20632 36419 20634
rect 35249 20576 35254 20632
rect 35310 20576 36358 20632
rect 36414 20576 36419 20632
rect 35249 20574 36419 20576
rect 15150 20498 15210 20572
rect 35249 20571 35315 20574
rect 36353 20571 36419 20574
rect 19517 20498 19583 20501
rect 15150 20496 19583 20498
rect 15150 20440 19522 20496
rect 19578 20440 19583 20496
rect 15150 20438 19583 20440
rect 19517 20435 19583 20438
rect 24025 20498 24091 20501
rect 32213 20498 32279 20501
rect 24025 20496 32279 20498
rect 24025 20440 24030 20496
rect 24086 20440 32218 20496
rect 32274 20440 32279 20496
rect 24025 20438 32279 20440
rect 24025 20435 24091 20438
rect 32213 20435 32279 20438
rect 35801 20498 35867 20501
rect 36537 20498 36603 20501
rect 35801 20496 36603 20498
rect 35801 20440 35806 20496
rect 35862 20440 36542 20496
rect 36598 20440 36603 20496
rect 35801 20438 36603 20440
rect 35801 20435 35867 20438
rect 36537 20435 36603 20438
rect 41505 20498 41571 20501
rect 41720 20498 42520 20528
rect 41505 20496 42520 20498
rect 41505 20440 41510 20496
rect 41566 20440 42520 20496
rect 41505 20438 42520 20440
rect 41505 20435 41571 20438
rect 41720 20408 42520 20438
rect 13997 20364 14063 20365
rect 13997 20362 14044 20364
rect 13952 20360 14044 20362
rect 13952 20304 14002 20360
rect 13952 20302 14044 20304
rect 13997 20300 14044 20302
rect 14108 20300 14114 20364
rect 16481 20362 16547 20365
rect 17953 20362 18019 20365
rect 18965 20362 19031 20365
rect 24209 20362 24275 20365
rect 16481 20360 19031 20362
rect 16481 20304 16486 20360
rect 16542 20304 17958 20360
rect 18014 20304 18970 20360
rect 19026 20304 19031 20360
rect 16481 20302 19031 20304
rect 13997 20299 14063 20300
rect 16481 20299 16547 20302
rect 17953 20299 18019 20302
rect 18965 20299 19031 20302
rect 19290 20360 24275 20362
rect 19290 20304 24214 20360
rect 24270 20304 24275 20360
rect 19290 20302 24275 20304
rect 12525 20226 12591 20229
rect 19290 20226 19350 20302
rect 24209 20299 24275 20302
rect 33961 20362 34027 20365
rect 36445 20362 36511 20365
rect 33961 20360 36511 20362
rect 33961 20304 33966 20360
rect 34022 20304 36450 20360
rect 36506 20304 36511 20360
rect 33961 20302 36511 20304
rect 33961 20299 34027 20302
rect 36445 20299 36511 20302
rect 12525 20224 19350 20226
rect 12525 20168 12530 20224
rect 12586 20168 19350 20224
rect 12525 20166 19350 20168
rect 19609 20226 19675 20229
rect 24485 20226 24551 20229
rect 19609 20224 24551 20226
rect 19609 20168 19614 20224
rect 19670 20168 24490 20224
rect 24546 20168 24551 20224
rect 19609 20166 24551 20168
rect 12525 20163 12591 20166
rect 19609 20163 19675 20166
rect 24485 20163 24551 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 12341 20090 12407 20093
rect 17677 20090 17743 20093
rect 12341 20088 17743 20090
rect 12341 20032 12346 20088
rect 12402 20032 17682 20088
rect 17738 20032 17743 20088
rect 12341 20030 17743 20032
rect 12341 20027 12407 20030
rect 17677 20027 17743 20030
rect 23422 20028 23428 20092
rect 23492 20090 23498 20092
rect 31385 20090 31451 20093
rect 23492 20088 31451 20090
rect 23492 20032 31390 20088
rect 31446 20032 31451 20088
rect 23492 20030 31451 20032
rect 23492 20028 23498 20030
rect 31385 20027 31451 20030
rect 11421 19954 11487 19957
rect 23289 19954 23355 19957
rect 11421 19952 23355 19954
rect 11421 19896 11426 19952
rect 11482 19896 23294 19952
rect 23350 19896 23355 19952
rect 11421 19894 23355 19896
rect 11421 19891 11487 19894
rect 23289 19891 23355 19894
rect 0 19818 800 19848
rect 933 19818 999 19821
rect 0 19816 999 19818
rect 0 19760 938 19816
rect 994 19760 999 19816
rect 0 19758 999 19760
rect 0 19728 800 19758
rect 933 19755 999 19758
rect 1669 19818 1735 19821
rect 17217 19818 17283 19821
rect 1669 19816 17283 19818
rect 1669 19760 1674 19816
rect 1730 19760 17222 19816
rect 17278 19760 17283 19816
rect 1669 19758 17283 19760
rect 1669 19755 1735 19758
rect 17217 19755 17283 19758
rect 26877 19818 26943 19821
rect 35341 19818 35407 19821
rect 26877 19816 35407 19818
rect 26877 19760 26882 19816
rect 26938 19760 35346 19816
rect 35402 19760 35407 19816
rect 26877 19758 35407 19760
rect 26877 19755 26943 19758
rect 35341 19755 35407 19758
rect 11278 19620 11284 19684
rect 11348 19682 11354 19684
rect 16573 19682 16639 19685
rect 11348 19680 16639 19682
rect 11348 19624 16578 19680
rect 16634 19624 16639 19680
rect 11348 19622 16639 19624
rect 11348 19620 11354 19622
rect 16573 19619 16639 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 15929 19546 15995 19549
rect 17769 19546 17835 19549
rect 15929 19544 17835 19546
rect 15929 19488 15934 19544
rect 15990 19488 17774 19544
rect 17830 19488 17835 19544
rect 15929 19486 17835 19488
rect 15929 19483 15995 19486
rect 17769 19483 17835 19486
rect 23422 19348 23428 19412
rect 23492 19410 23498 19412
rect 25129 19410 25195 19413
rect 23492 19408 25195 19410
rect 23492 19352 25134 19408
rect 25190 19352 25195 19408
rect 23492 19350 25195 19352
rect 23492 19348 23498 19350
rect 25129 19347 25195 19350
rect 4613 19274 4679 19277
rect 5809 19274 5875 19277
rect 16757 19276 16823 19277
rect 16757 19274 16804 19276
rect 4613 19272 5875 19274
rect 4613 19216 4618 19272
rect 4674 19216 5814 19272
rect 5870 19216 5875 19272
rect 4613 19214 5875 19216
rect 16712 19272 16804 19274
rect 16712 19216 16762 19272
rect 16712 19214 16804 19216
rect 4613 19211 4679 19214
rect 5809 19211 5875 19214
rect 16757 19212 16804 19214
rect 16868 19212 16874 19276
rect 19885 19274 19951 19277
rect 20110 19274 20116 19276
rect 19885 19272 20116 19274
rect 19885 19216 19890 19272
rect 19946 19216 20116 19272
rect 19885 19214 20116 19216
rect 16757 19211 16823 19212
rect 19885 19211 19951 19214
rect 20110 19212 20116 19214
rect 20180 19212 20186 19276
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 11094 18804 11100 18868
rect 11164 18866 11170 18868
rect 16573 18866 16639 18869
rect 11164 18864 16639 18866
rect 11164 18808 16578 18864
rect 16634 18808 16639 18864
rect 11164 18806 16639 18808
rect 11164 18804 11170 18806
rect 16573 18803 16639 18806
rect 18137 18866 18203 18869
rect 33133 18866 33199 18869
rect 18137 18864 33199 18866
rect 18137 18808 18142 18864
rect 18198 18808 33138 18864
rect 33194 18808 33199 18864
rect 18137 18806 33199 18808
rect 18137 18803 18203 18806
rect 33133 18803 33199 18806
rect 4337 18730 4403 18733
rect 7465 18730 7531 18733
rect 4337 18728 7531 18730
rect 4337 18672 4342 18728
rect 4398 18672 7470 18728
rect 7526 18672 7531 18728
rect 4337 18670 7531 18672
rect 4337 18667 4403 18670
rect 7465 18667 7531 18670
rect 18229 18730 18295 18733
rect 20161 18730 20227 18733
rect 20846 18730 20852 18732
rect 18229 18728 20852 18730
rect 18229 18672 18234 18728
rect 18290 18672 20166 18728
rect 20222 18672 20852 18728
rect 18229 18670 20852 18672
rect 18229 18667 18295 18670
rect 20161 18667 20227 18670
rect 20846 18668 20852 18670
rect 20916 18730 20922 18732
rect 22369 18730 22435 18733
rect 20916 18728 22435 18730
rect 20916 18672 22374 18728
rect 22430 18672 22435 18728
rect 20916 18670 22435 18672
rect 20916 18668 20922 18670
rect 22369 18667 22435 18670
rect 31937 18730 32003 18733
rect 33777 18730 33843 18733
rect 31937 18728 33843 18730
rect 31937 18672 31942 18728
rect 31998 18672 33782 18728
rect 33838 18672 33843 18728
rect 31937 18670 33843 18672
rect 31937 18667 32003 18670
rect 33777 18667 33843 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 24485 18458 24551 18461
rect 27521 18458 27587 18461
rect 24485 18456 27587 18458
rect 24485 18400 24490 18456
rect 24546 18400 27526 18456
rect 27582 18400 27587 18456
rect 24485 18398 27587 18400
rect 24485 18395 24551 18398
rect 27521 18395 27587 18398
rect 10501 18324 10567 18325
rect 10501 18320 10548 18324
rect 10612 18322 10618 18324
rect 23105 18322 23171 18325
rect 29126 18322 29132 18324
rect 10501 18264 10506 18320
rect 10501 18260 10548 18264
rect 10612 18262 10658 18322
rect 23105 18320 29132 18322
rect 23105 18264 23110 18320
rect 23166 18264 29132 18320
rect 23105 18262 29132 18264
rect 10612 18260 10618 18262
rect 10501 18259 10567 18260
rect 23105 18259 23171 18262
rect 29126 18260 29132 18262
rect 29196 18260 29202 18324
rect 10593 18186 10659 18189
rect 25037 18186 25103 18189
rect 10593 18184 25103 18186
rect 10593 18128 10598 18184
rect 10654 18128 25042 18184
rect 25098 18128 25103 18184
rect 10593 18126 25103 18128
rect 10593 18123 10659 18126
rect 25037 18123 25103 18126
rect 16021 18050 16087 18053
rect 26509 18050 26575 18053
rect 16021 18048 26575 18050
rect 16021 17992 16026 18048
rect 16082 17992 26514 18048
rect 26570 17992 26575 18048
rect 16021 17990 26575 17992
rect 16021 17987 16087 17990
rect 26509 17987 26575 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 9581 17778 9647 17781
rect 25446 17778 25452 17780
rect 9581 17776 25452 17778
rect 9581 17720 9586 17776
rect 9642 17720 25452 17776
rect 9581 17718 25452 17720
rect 9581 17715 9647 17718
rect 25446 17716 25452 17718
rect 25516 17716 25522 17780
rect 31109 17642 31175 17645
rect 36353 17642 36419 17645
rect 31109 17640 36419 17642
rect 31109 17584 31114 17640
rect 31170 17584 36358 17640
rect 36414 17584 36419 17640
rect 31109 17582 36419 17584
rect 31109 17579 31175 17582
rect 36353 17579 36419 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 14181 17370 14247 17373
rect 18965 17370 19031 17373
rect 14181 17368 19031 17370
rect 14181 17312 14186 17368
rect 14242 17312 18970 17368
rect 19026 17312 19031 17368
rect 14181 17310 19031 17312
rect 14181 17307 14247 17310
rect 18965 17307 19031 17310
rect 20529 17370 20595 17373
rect 26325 17370 26391 17373
rect 20529 17368 26391 17370
rect 20529 17312 20534 17368
rect 20590 17312 26330 17368
rect 26386 17312 26391 17368
rect 20529 17310 26391 17312
rect 20529 17307 20595 17310
rect 26325 17307 26391 17310
rect 13169 17234 13235 17237
rect 23238 17234 23244 17236
rect 13169 17232 23244 17234
rect 13169 17176 13174 17232
rect 13230 17176 23244 17232
rect 13169 17174 23244 17176
rect 13169 17171 13235 17174
rect 23238 17172 23244 17174
rect 23308 17234 23314 17236
rect 24945 17234 25011 17237
rect 23308 17232 25011 17234
rect 23308 17176 24950 17232
rect 25006 17176 25011 17232
rect 23308 17174 25011 17176
rect 23308 17172 23314 17174
rect 24945 17171 25011 17174
rect 19977 16962 20043 16965
rect 22001 16962 22067 16965
rect 19977 16960 22067 16962
rect 19977 16904 19982 16960
rect 20038 16904 22006 16960
rect 22062 16904 22067 16960
rect 19977 16902 22067 16904
rect 19977 16899 20043 16902
rect 22001 16899 22067 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 15285 16826 15351 16829
rect 17534 16826 17540 16828
rect 15285 16824 17540 16826
rect 15285 16768 15290 16824
rect 15346 16768 17540 16824
rect 15285 16766 17540 16768
rect 15285 16763 15351 16766
rect 17534 16764 17540 16766
rect 17604 16826 17610 16828
rect 23381 16826 23447 16829
rect 17604 16824 23447 16826
rect 17604 16768 23386 16824
rect 23442 16768 23447 16824
rect 17604 16766 23447 16768
rect 17604 16764 17610 16766
rect 23381 16763 23447 16766
rect 20713 16690 20779 16693
rect 33593 16690 33659 16693
rect 20713 16688 33659 16690
rect 20713 16632 20718 16688
rect 20774 16632 33598 16688
rect 33654 16632 33659 16688
rect 20713 16630 33659 16632
rect 20713 16627 20779 16630
rect 33593 16627 33659 16630
rect 38653 16690 38719 16693
rect 39573 16690 39639 16693
rect 38653 16688 39639 16690
rect 38653 16632 38658 16688
rect 38714 16632 39578 16688
rect 39634 16632 39639 16688
rect 38653 16630 39639 16632
rect 38653 16627 38719 16630
rect 39573 16627 39639 16630
rect 11237 16554 11303 16557
rect 12065 16554 12131 16557
rect 15561 16554 15627 16557
rect 33501 16554 33567 16557
rect 34145 16554 34211 16557
rect 11237 16552 34211 16554
rect 11237 16496 11242 16552
rect 11298 16496 12070 16552
rect 12126 16496 15566 16552
rect 15622 16496 33506 16552
rect 33562 16496 34150 16552
rect 34206 16496 34211 16552
rect 11237 16494 34211 16496
rect 11237 16491 11303 16494
rect 12065 16491 12131 16494
rect 15561 16491 15627 16494
rect 33501 16491 33567 16494
rect 34145 16491 34211 16494
rect 38653 16554 38719 16557
rect 39389 16554 39455 16557
rect 38653 16552 39455 16554
rect 38653 16496 38658 16552
rect 38714 16496 39394 16552
rect 39450 16496 39455 16552
rect 38653 16494 39455 16496
rect 38653 16491 38719 16494
rect 39389 16491 39455 16494
rect 25681 16418 25747 16421
rect 27153 16418 27219 16421
rect 25681 16416 27219 16418
rect 25681 16360 25686 16416
rect 25742 16360 27158 16416
rect 27214 16360 27219 16416
rect 25681 16358 27219 16360
rect 25681 16355 25747 16358
rect 27153 16355 27219 16358
rect 41505 16418 41571 16421
rect 41720 16418 42520 16448
rect 41505 16416 42520 16418
rect 41505 16360 41510 16416
rect 41566 16360 42520 16416
rect 41505 16358 42520 16360
rect 41505 16355 41571 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 41720 16328 42520 16358
rect 19570 16287 19886 16288
rect 23381 16282 23447 16285
rect 27705 16282 27771 16285
rect 23381 16280 27771 16282
rect 23381 16224 23386 16280
rect 23442 16224 27710 16280
rect 27766 16224 27771 16280
rect 23381 16222 27771 16224
rect 23381 16219 23447 16222
rect 27705 16219 27771 16222
rect 29361 16282 29427 16285
rect 29821 16282 29887 16285
rect 29361 16280 29887 16282
rect 29361 16224 29366 16280
rect 29422 16224 29826 16280
rect 29882 16224 29887 16280
rect 29361 16222 29887 16224
rect 29361 16219 29427 16222
rect 29821 16219 29887 16222
rect 11421 16146 11487 16149
rect 12341 16146 12407 16149
rect 11421 16144 12407 16146
rect 11421 16088 11426 16144
rect 11482 16088 12346 16144
rect 12402 16088 12407 16144
rect 11421 16086 12407 16088
rect 11421 16083 11487 16086
rect 12341 16083 12407 16086
rect 19425 16146 19491 16149
rect 20897 16146 20963 16149
rect 19425 16144 20963 16146
rect 19425 16088 19430 16144
rect 19486 16088 20902 16144
rect 20958 16088 20963 16144
rect 19425 16086 20963 16088
rect 19425 16083 19491 16086
rect 20897 16083 20963 16086
rect 25446 16084 25452 16148
rect 25516 16146 25522 16148
rect 25998 16146 26004 16148
rect 25516 16086 26004 16146
rect 25516 16084 25522 16086
rect 25998 16084 26004 16086
rect 26068 16146 26074 16148
rect 28165 16146 28231 16149
rect 26068 16144 28231 16146
rect 26068 16088 28170 16144
rect 28226 16088 28231 16144
rect 26068 16086 28231 16088
rect 26068 16084 26074 16086
rect 28165 16083 28231 16086
rect 29085 16146 29151 16149
rect 29637 16146 29703 16149
rect 29085 16144 29703 16146
rect 29085 16088 29090 16144
rect 29146 16088 29642 16144
rect 29698 16088 29703 16144
rect 29085 16086 29703 16088
rect 29085 16083 29151 16086
rect 29637 16083 29703 16086
rect 24669 16010 24735 16013
rect 32765 16010 32831 16013
rect 24669 16008 32831 16010
rect 24669 15952 24674 16008
rect 24730 15952 32770 16008
rect 32826 15952 32831 16008
rect 24669 15950 32831 15952
rect 24669 15947 24735 15950
rect 32765 15947 32831 15950
rect 5022 15812 5028 15876
rect 5092 15874 5098 15876
rect 20529 15874 20595 15877
rect 5092 15872 20595 15874
rect 5092 15816 20534 15872
rect 20590 15816 20595 15872
rect 5092 15814 20595 15816
rect 5092 15812 5098 15814
rect 20529 15811 20595 15814
rect 22921 15874 22987 15877
rect 23657 15874 23723 15877
rect 22921 15872 23723 15874
rect 22921 15816 22926 15872
rect 22982 15816 23662 15872
rect 23718 15816 23723 15872
rect 22921 15814 23723 15816
rect 22921 15811 22987 15814
rect 23657 15811 23723 15814
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 17769 15738 17835 15741
rect 29453 15738 29519 15741
rect 17769 15736 29519 15738
rect 17769 15680 17774 15736
rect 17830 15680 29458 15736
rect 29514 15680 29519 15736
rect 17769 15678 29519 15680
rect 17769 15675 17835 15678
rect 29453 15675 29519 15678
rect 10910 15540 10916 15604
rect 10980 15602 10986 15604
rect 15837 15602 15903 15605
rect 10980 15600 15903 15602
rect 10980 15544 15842 15600
rect 15898 15544 15903 15600
rect 10980 15542 15903 15544
rect 10980 15540 10986 15542
rect 15837 15539 15903 15542
rect 18137 15602 18203 15605
rect 18270 15602 18276 15604
rect 18137 15600 18276 15602
rect 18137 15544 18142 15600
rect 18198 15544 18276 15600
rect 18137 15542 18276 15544
rect 18137 15539 18203 15542
rect 18270 15540 18276 15542
rect 18340 15540 18346 15604
rect 18413 15602 18479 15605
rect 24577 15602 24643 15605
rect 18413 15600 24643 15602
rect 18413 15544 18418 15600
rect 18474 15544 24582 15600
rect 24638 15544 24643 15600
rect 18413 15542 24643 15544
rect 18278 15466 18338 15540
rect 18413 15539 18479 15542
rect 24577 15539 24643 15542
rect 22093 15466 22159 15469
rect 36537 15466 36603 15469
rect 18278 15406 20178 15466
rect 20118 15330 20178 15406
rect 22093 15464 36603 15466
rect 22093 15408 22098 15464
rect 22154 15408 36542 15464
rect 36598 15408 36603 15464
rect 22093 15406 36603 15408
rect 22093 15403 22159 15406
rect 36537 15403 36603 15406
rect 24025 15330 24091 15333
rect 24761 15330 24827 15333
rect 20118 15328 24827 15330
rect 20118 15272 24030 15328
rect 24086 15272 24766 15328
rect 24822 15272 24827 15328
rect 20118 15270 24827 15272
rect 24025 15267 24091 15270
rect 24761 15267 24827 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 5441 15194 5507 15197
rect 11697 15194 11763 15197
rect 14917 15196 14983 15197
rect 14917 15194 14964 15196
rect 5441 15192 11763 15194
rect 5441 15136 5446 15192
rect 5502 15136 11702 15192
rect 11758 15136 11763 15192
rect 5441 15134 11763 15136
rect 14872 15192 14964 15194
rect 14872 15136 14922 15192
rect 14872 15134 14964 15136
rect 5441 15131 5507 15134
rect 11697 15131 11763 15134
rect 14917 15132 14964 15134
rect 15028 15132 15034 15196
rect 17718 15132 17724 15196
rect 17788 15132 17794 15196
rect 23657 15194 23723 15197
rect 25129 15194 25195 15197
rect 23657 15192 25195 15194
rect 23657 15136 23662 15192
rect 23718 15136 25134 15192
rect 25190 15136 25195 15192
rect 23657 15134 25195 15136
rect 14917 15131 15026 15132
rect 14966 15058 15026 15131
rect 17033 15058 17099 15061
rect 14966 15056 17099 15058
rect 14966 15000 17038 15056
rect 17094 15000 17099 15056
rect 14966 14998 17099 15000
rect 17726 15058 17786 15132
rect 23657 15131 23723 15134
rect 25129 15131 25195 15134
rect 28165 15194 28231 15197
rect 28942 15194 28948 15196
rect 28165 15192 28948 15194
rect 28165 15136 28170 15192
rect 28226 15136 28948 15192
rect 28165 15134 28948 15136
rect 28165 15131 28231 15134
rect 28942 15132 28948 15134
rect 29012 15132 29018 15196
rect 18413 15058 18479 15061
rect 24669 15058 24735 15061
rect 17726 14998 18338 15058
rect 17033 14995 17099 14998
rect 16113 14922 16179 14925
rect 17953 14922 18019 14925
rect 16113 14920 18019 14922
rect 16113 14864 16118 14920
rect 16174 14864 17958 14920
rect 18014 14864 18019 14920
rect 16113 14862 18019 14864
rect 18278 14922 18338 14998
rect 18413 15056 24735 15058
rect 18413 15000 18418 15056
rect 18474 15000 24674 15056
rect 24730 15000 24735 15056
rect 18413 14998 24735 15000
rect 18413 14995 18479 14998
rect 24669 14995 24735 14998
rect 18873 14922 18939 14925
rect 25957 14922 26023 14925
rect 18278 14920 26023 14922
rect 18278 14864 18878 14920
rect 18934 14864 25962 14920
rect 26018 14864 26023 14920
rect 18278 14862 26023 14864
rect 16113 14859 16179 14862
rect 17953 14859 18019 14862
rect 18873 14859 18939 14862
rect 25957 14859 26023 14862
rect 15101 14786 15167 14789
rect 29729 14786 29795 14789
rect 15101 14784 29795 14786
rect 15101 14728 15106 14784
rect 15162 14728 29734 14784
rect 29790 14728 29795 14784
rect 15101 14726 29795 14728
rect 15101 14723 15167 14726
rect 29729 14723 29795 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 17033 14650 17099 14653
rect 18086 14650 18092 14652
rect 17033 14648 18092 14650
rect 17033 14592 17038 14648
rect 17094 14592 18092 14648
rect 17033 14590 18092 14592
rect 17033 14587 17099 14590
rect 18086 14588 18092 14590
rect 18156 14588 18162 14652
rect 18413 14650 18479 14653
rect 20662 14650 20668 14652
rect 18413 14648 20668 14650
rect 18413 14592 18418 14648
rect 18474 14592 20668 14648
rect 18413 14590 20668 14592
rect 18413 14587 18479 14590
rect 20662 14588 20668 14590
rect 20732 14650 20738 14652
rect 21909 14650 21975 14653
rect 20732 14648 21975 14650
rect 20732 14592 21914 14648
rect 21970 14592 21975 14648
rect 20732 14590 21975 14592
rect 20732 14588 20738 14590
rect 21909 14587 21975 14590
rect 22093 14650 22159 14653
rect 23422 14650 23428 14652
rect 22093 14648 23428 14650
rect 22093 14592 22098 14648
rect 22154 14592 23428 14648
rect 22093 14590 23428 14592
rect 22093 14587 22159 14590
rect 23422 14588 23428 14590
rect 23492 14588 23498 14652
rect 12157 14514 12223 14517
rect 17769 14514 17835 14517
rect 12157 14512 17835 14514
rect 12157 14456 12162 14512
rect 12218 14456 17774 14512
rect 17830 14456 17835 14512
rect 12157 14454 17835 14456
rect 12157 14451 12223 14454
rect 17769 14451 17835 14454
rect 20437 14514 20503 14517
rect 27337 14514 27403 14517
rect 20437 14512 27403 14514
rect 20437 14456 20442 14512
rect 20498 14456 27342 14512
rect 27398 14456 27403 14512
rect 20437 14454 27403 14456
rect 20437 14451 20503 14454
rect 27337 14451 27403 14454
rect 17769 14378 17835 14381
rect 27705 14378 27771 14381
rect 33225 14378 33291 14381
rect 17769 14376 33291 14378
rect 17769 14320 17774 14376
rect 17830 14320 27710 14376
rect 27766 14320 33230 14376
rect 33286 14320 33291 14376
rect 17769 14318 33291 14320
rect 17769 14315 17835 14318
rect 27705 14315 27771 14318
rect 33225 14315 33291 14318
rect 38837 14378 38903 14381
rect 40493 14378 40559 14381
rect 38837 14376 40559 14378
rect 38837 14320 38842 14376
rect 38898 14320 40498 14376
rect 40554 14320 40559 14376
rect 38837 14318 40559 14320
rect 38837 14315 38903 14318
rect 40493 14315 40559 14318
rect 14917 14242 14983 14245
rect 17217 14242 17283 14245
rect 18137 14242 18203 14245
rect 14917 14240 18203 14242
rect 14917 14184 14922 14240
rect 14978 14184 17222 14240
rect 17278 14184 18142 14240
rect 18198 14184 18203 14240
rect 14917 14182 18203 14184
rect 14917 14179 14983 14182
rect 17217 14179 17283 14182
rect 18137 14179 18203 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 17401 14106 17467 14109
rect 18597 14106 18663 14109
rect 17401 14104 18663 14106
rect 17401 14048 17406 14104
rect 17462 14048 18602 14104
rect 18658 14048 18663 14104
rect 17401 14046 18663 14048
rect 17401 14043 17467 14046
rect 18597 14043 18663 14046
rect 22737 14106 22803 14109
rect 28165 14106 28231 14109
rect 22737 14104 28231 14106
rect 22737 14048 22742 14104
rect 22798 14048 28170 14104
rect 28226 14048 28231 14104
rect 22737 14046 28231 14048
rect 22737 14043 22803 14046
rect 28165 14043 28231 14046
rect 30005 14106 30071 14109
rect 30833 14106 30899 14109
rect 34237 14106 34303 14109
rect 30005 14104 34303 14106
rect 30005 14048 30010 14104
rect 30066 14048 30838 14104
rect 30894 14048 34242 14104
rect 34298 14048 34303 14104
rect 30005 14046 34303 14048
rect 30005 14043 30071 14046
rect 30833 14043 30899 14046
rect 34237 14043 34303 14046
rect 22829 13970 22895 13973
rect 17772 13968 22895 13970
rect 17772 13912 22834 13968
rect 22890 13912 22895 13968
rect 17772 13910 22895 13912
rect 17772 13837 17832 13910
rect 22829 13907 22895 13910
rect 24393 13970 24459 13973
rect 25129 13970 25195 13973
rect 25773 13970 25839 13973
rect 24393 13968 25839 13970
rect 24393 13912 24398 13968
rect 24454 13912 25134 13968
rect 25190 13912 25778 13968
rect 25834 13912 25839 13968
rect 24393 13910 25839 13912
rect 24393 13907 24459 13910
rect 25129 13907 25195 13910
rect 25773 13907 25839 13910
rect 34881 13970 34947 13973
rect 35617 13970 35683 13973
rect 34881 13968 35683 13970
rect 34881 13912 34886 13968
rect 34942 13912 35622 13968
rect 35678 13912 35683 13968
rect 34881 13910 35683 13912
rect 34881 13907 34947 13910
rect 35617 13907 35683 13910
rect 17769 13832 17835 13837
rect 17769 13776 17774 13832
rect 17830 13776 17835 13832
rect 17769 13771 17835 13776
rect 18045 13834 18111 13837
rect 18597 13834 18663 13837
rect 18045 13832 18663 13834
rect 18045 13776 18050 13832
rect 18106 13776 18602 13832
rect 18658 13776 18663 13832
rect 18045 13774 18663 13776
rect 18045 13771 18111 13774
rect 18597 13771 18663 13774
rect 5257 13700 5323 13701
rect 5206 13698 5212 13700
rect 5166 13638 5212 13698
rect 5276 13696 5323 13700
rect 5318 13640 5323 13696
rect 5206 13636 5212 13638
rect 5276 13636 5323 13640
rect 18086 13636 18092 13700
rect 18156 13698 18162 13700
rect 18229 13698 18295 13701
rect 18156 13696 18295 13698
rect 18156 13640 18234 13696
rect 18290 13640 18295 13696
rect 18156 13638 18295 13640
rect 18156 13636 18162 13638
rect 5257 13635 5323 13636
rect 18229 13635 18295 13638
rect 20897 13698 20963 13701
rect 23013 13698 23079 13701
rect 23749 13698 23815 13701
rect 20897 13696 23815 13698
rect 20897 13640 20902 13696
rect 20958 13640 23018 13696
rect 23074 13640 23754 13696
rect 23810 13640 23815 13696
rect 20897 13638 23815 13640
rect 20897 13635 20963 13638
rect 23013 13635 23079 13638
rect 23749 13635 23815 13638
rect 28993 13698 29059 13701
rect 29126 13698 29132 13700
rect 28993 13696 29132 13698
rect 28993 13640 28998 13696
rect 29054 13640 29132 13696
rect 28993 13638 29132 13640
rect 28993 13635 29059 13638
rect 29126 13636 29132 13638
rect 29196 13636 29202 13700
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 15837 13562 15903 13565
rect 19517 13562 19583 13565
rect 15837 13560 19583 13562
rect 15837 13504 15842 13560
rect 15898 13504 19522 13560
rect 19578 13504 19583 13560
rect 15837 13502 19583 13504
rect 15837 13499 15903 13502
rect 19517 13499 19583 13502
rect 19701 13562 19767 13565
rect 26785 13562 26851 13565
rect 19701 13560 26851 13562
rect 19701 13504 19706 13560
rect 19762 13504 26790 13560
rect 26846 13504 26851 13560
rect 19701 13502 26851 13504
rect 19701 13499 19767 13502
rect 26785 13499 26851 13502
rect 13077 13290 13143 13293
rect 16757 13290 16823 13293
rect 13077 13288 16823 13290
rect 13077 13232 13082 13288
rect 13138 13232 16762 13288
rect 16818 13232 16823 13288
rect 13077 13230 16823 13232
rect 13077 13227 13143 13230
rect 16757 13227 16823 13230
rect 24577 13290 24643 13293
rect 26693 13290 26759 13293
rect 24577 13288 26759 13290
rect 24577 13232 24582 13288
rect 24638 13232 26698 13288
rect 26754 13232 26759 13288
rect 24577 13230 26759 13232
rect 24577 13227 24643 13230
rect 26693 13227 26759 13230
rect 34421 13290 34487 13293
rect 35893 13290 35959 13293
rect 34421 13288 35959 13290
rect 34421 13232 34426 13288
rect 34482 13232 35898 13288
rect 35954 13232 35959 13288
rect 34421 13230 35959 13232
rect 34421 13227 34487 13230
rect 35893 13227 35959 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 19517 12882 19583 12885
rect 21081 12882 21147 12885
rect 19517 12880 21147 12882
rect 19517 12824 19522 12880
rect 19578 12824 21086 12880
rect 21142 12824 21147 12880
rect 19517 12822 21147 12824
rect 19517 12819 19583 12822
rect 21081 12819 21147 12822
rect 7833 12746 7899 12749
rect 9029 12746 9095 12749
rect 7833 12744 9095 12746
rect 7833 12688 7838 12744
rect 7894 12688 9034 12744
rect 9090 12688 9095 12744
rect 7833 12686 9095 12688
rect 7833 12683 7899 12686
rect 9029 12683 9095 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 15929 12474 15995 12477
rect 19425 12474 19491 12477
rect 15929 12472 19491 12474
rect 15929 12416 15934 12472
rect 15990 12416 19430 12472
rect 19486 12416 19491 12472
rect 15929 12414 19491 12416
rect 15929 12411 15995 12414
rect 19425 12411 19491 12414
rect 21541 12474 21607 12477
rect 24853 12474 24919 12477
rect 21541 12472 24919 12474
rect 21541 12416 21546 12472
rect 21602 12416 24858 12472
rect 24914 12416 24919 12472
rect 21541 12414 24919 12416
rect 21541 12411 21607 12414
rect 24853 12411 24919 12414
rect 22277 12338 22343 12341
rect 24761 12338 24827 12341
rect 28901 12338 28967 12341
rect 22277 12336 28967 12338
rect 22277 12280 22282 12336
rect 22338 12280 24766 12336
rect 24822 12280 28906 12336
rect 28962 12280 28967 12336
rect 22277 12278 28967 12280
rect 22277 12275 22343 12278
rect 24761 12275 24827 12278
rect 28901 12275 28967 12278
rect 39849 12338 39915 12341
rect 41720 12338 42520 12368
rect 39849 12336 42520 12338
rect 39849 12280 39854 12336
rect 39910 12280 42520 12336
rect 39849 12278 42520 12280
rect 39849 12275 39915 12278
rect 41720 12248 42520 12278
rect 10593 12202 10659 12205
rect 21909 12202 21975 12205
rect 10593 12200 21975 12202
rect 10593 12144 10598 12200
rect 10654 12144 21914 12200
rect 21970 12144 21975 12200
rect 10593 12142 21975 12144
rect 10593 12139 10659 12142
rect 21909 12139 21975 12142
rect 20529 12066 20595 12069
rect 21633 12066 21699 12069
rect 34789 12066 34855 12069
rect 20529 12064 34855 12066
rect 20529 12008 20534 12064
rect 20590 12008 21638 12064
rect 21694 12008 34794 12064
rect 34850 12008 34855 12064
rect 20529 12006 34855 12008
rect 20529 12003 20595 12006
rect 21633 12003 21699 12006
rect 34789 12003 34855 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 21817 11930 21883 11933
rect 25221 11930 25287 11933
rect 25681 11930 25747 11933
rect 21817 11928 25747 11930
rect 21817 11872 21822 11928
rect 21878 11872 25226 11928
rect 25282 11872 25686 11928
rect 25742 11872 25747 11928
rect 21817 11870 25747 11872
rect 21817 11867 21883 11870
rect 25221 11867 25287 11870
rect 25681 11867 25747 11870
rect 13629 11794 13695 11797
rect 22277 11794 22343 11797
rect 13629 11792 22343 11794
rect 13629 11736 13634 11792
rect 13690 11736 22282 11792
rect 22338 11736 22343 11792
rect 13629 11734 22343 11736
rect 13629 11731 13695 11734
rect 22277 11731 22343 11734
rect 24853 11794 24919 11797
rect 26509 11794 26575 11797
rect 24853 11792 26575 11794
rect 24853 11736 24858 11792
rect 24914 11736 26514 11792
rect 26570 11736 26575 11792
rect 24853 11734 26575 11736
rect 24853 11731 24919 11734
rect 26509 11731 26575 11734
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 21173 11658 21239 11661
rect 21633 11658 21699 11661
rect 21173 11656 21699 11658
rect 21173 11600 21178 11656
rect 21234 11600 21638 11656
rect 21694 11600 21699 11656
rect 21173 11598 21699 11600
rect 21173 11595 21239 11598
rect 21633 11595 21699 11598
rect 26550 11460 26556 11524
rect 26620 11522 26626 11524
rect 26877 11522 26943 11525
rect 26620 11520 26943 11522
rect 26620 11464 26882 11520
rect 26938 11464 26943 11520
rect 26620 11462 26943 11464
rect 26620 11460 26626 11462
rect 26877 11459 26943 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 20345 11386 20411 11389
rect 25957 11386 26023 11389
rect 20345 11384 26023 11386
rect 20345 11328 20350 11384
rect 20406 11328 25962 11384
rect 26018 11328 26023 11384
rect 20345 11326 26023 11328
rect 20345 11323 20411 11326
rect 25957 11323 26023 11326
rect 22185 11250 22251 11253
rect 26417 11250 26483 11253
rect 22185 11248 26483 11250
rect 22185 11192 22190 11248
rect 22246 11192 26422 11248
rect 26478 11192 26483 11248
rect 22185 11190 26483 11192
rect 22185 11187 22251 11190
rect 26417 11187 26483 11190
rect 7005 11114 7071 11117
rect 22369 11114 22435 11117
rect 25681 11114 25747 11117
rect 7005 11112 9690 11114
rect 7005 11056 7010 11112
rect 7066 11056 9690 11112
rect 7005 11054 9690 11056
rect 7005 11051 7071 11054
rect 9630 10978 9690 11054
rect 22369 11112 25747 11114
rect 22369 11056 22374 11112
rect 22430 11056 25686 11112
rect 25742 11056 25747 11112
rect 22369 11054 25747 11056
rect 22369 11051 22435 11054
rect 25681 11051 25747 11054
rect 25957 11114 26023 11117
rect 25957 11112 26572 11114
rect 25957 11056 25962 11112
rect 26018 11056 26572 11112
rect 25957 11054 26572 11056
rect 25957 11051 26023 11054
rect 26512 10981 26572 11054
rect 15878 10978 15884 10980
rect 9630 10918 15884 10978
rect 15878 10916 15884 10918
rect 15948 10978 15954 10980
rect 17033 10978 17099 10981
rect 23197 10980 23263 10981
rect 23197 10978 23244 10980
rect 15948 10976 17099 10978
rect 15948 10920 17038 10976
rect 17094 10920 17099 10976
rect 15948 10918 17099 10920
rect 23152 10976 23244 10978
rect 23152 10920 23202 10976
rect 23152 10918 23244 10920
rect 15948 10916 15954 10918
rect 17033 10915 17099 10918
rect 23197 10916 23244 10918
rect 23308 10916 23314 10980
rect 24577 10978 24643 10981
rect 26233 10978 26299 10981
rect 24577 10976 26299 10978
rect 24577 10920 24582 10976
rect 24638 10920 26238 10976
rect 26294 10920 26299 10976
rect 24577 10918 26299 10920
rect 23197 10915 23263 10916
rect 24577 10915 24643 10918
rect 26233 10915 26299 10918
rect 26509 10976 26575 10981
rect 26509 10920 26514 10976
rect 26570 10920 26575 10976
rect 26509 10915 26575 10920
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 21725 10842 21791 10845
rect 26366 10842 26372 10844
rect 21725 10840 26372 10842
rect 21725 10784 21730 10840
rect 21786 10784 26372 10840
rect 21725 10782 26372 10784
rect 21725 10779 21791 10782
rect 26366 10780 26372 10782
rect 26436 10780 26442 10844
rect 25405 10706 25471 10709
rect 26969 10706 27035 10709
rect 25405 10704 27035 10706
rect 25405 10648 25410 10704
rect 25466 10648 26974 10704
rect 27030 10648 27035 10704
rect 25405 10646 27035 10648
rect 25405 10643 25471 10646
rect 26969 10643 27035 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 9489 10026 9555 10029
rect 11421 10026 11487 10029
rect 9489 10024 11487 10026
rect 9489 9968 9494 10024
rect 9550 9968 11426 10024
rect 11482 9968 11487 10024
rect 9489 9966 11487 9968
rect 9489 9963 9555 9966
rect 11421 9963 11487 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 20437 9618 20503 9621
rect 25589 9618 25655 9621
rect 20437 9616 25655 9618
rect 20437 9560 20442 9616
rect 20498 9560 25594 9616
rect 25650 9560 25655 9616
rect 20437 9558 25655 9560
rect 20437 9555 20503 9558
rect 25589 9555 25655 9558
rect 25865 9482 25931 9485
rect 26601 9482 26667 9485
rect 25865 9480 26667 9482
rect 25865 9424 25870 9480
rect 25926 9424 26606 9480
rect 26662 9424 26667 9480
rect 25865 9422 26667 9424
rect 25865 9419 25931 9422
rect 26601 9419 26667 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 15009 8530 15075 8533
rect 16021 8530 16087 8533
rect 17033 8530 17099 8533
rect 15009 8528 17099 8530
rect 15009 8472 15014 8528
rect 15070 8472 16026 8528
rect 16082 8472 17038 8528
rect 17094 8472 17099 8528
rect 15009 8470 17099 8472
rect 15009 8467 15075 8470
rect 16021 8467 16087 8470
rect 17033 8467 17099 8470
rect 41045 8258 41111 8261
rect 41720 8258 42520 8288
rect 41045 8256 42520 8258
rect 41045 8200 41050 8256
rect 41106 8200 42520 8256
rect 41045 8198 42520 8200
rect 41045 8195 41111 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 41720 8168 42520 8198
rect 34930 8127 35246 8128
rect 24761 7850 24827 7853
rect 25865 7850 25931 7853
rect 24761 7848 25931 7850
rect 24761 7792 24766 7848
rect 24822 7792 25870 7848
rect 25926 7792 25931 7848
rect 24761 7790 25931 7792
rect 24761 7787 24827 7790
rect 25865 7787 25931 7790
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 19885 7306 19951 7309
rect 22737 7306 22803 7309
rect 19885 7304 22803 7306
rect 19885 7248 19890 7304
rect 19946 7248 22742 7304
rect 22798 7248 22803 7304
rect 19885 7246 22803 7248
rect 19885 7243 19951 7246
rect 22737 7243 22803 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 9438 6700 9444 6764
rect 9508 6762 9514 6764
rect 9581 6762 9647 6765
rect 9508 6760 9647 6762
rect 9508 6704 9586 6760
rect 9642 6704 9647 6760
rect 9508 6702 9647 6704
rect 9508 6700 9514 6702
rect 9581 6699 9647 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 25957 5268 26023 5269
rect 25957 5266 26004 5268
rect 25912 5264 26004 5266
rect 25912 5208 25962 5264
rect 25912 5206 26004 5208
rect 25957 5204 26004 5206
rect 26068 5204 26074 5268
rect 25957 5203 26023 5204
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 17769 4858 17835 4861
rect 26550 4858 26556 4860
rect 17769 4856 26556 4858
rect 17769 4800 17774 4856
rect 17830 4800 26556 4856
rect 17769 4798 26556 4800
rect 17769 4795 17835 4798
rect 26550 4796 26556 4798
rect 26620 4796 26626 4860
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 41045 4178 41111 4181
rect 41720 4178 42520 4208
rect 41045 4176 42520 4178
rect 41045 4120 41050 4176
rect 41106 4120 42520 4176
rect 41045 4118 42520 4120
rect 41045 4115 41111 4118
rect 41720 4088 42520 4118
rect 15745 4042 15811 4045
rect 15878 4042 15884 4044
rect 15745 4040 15884 4042
rect 15745 3984 15750 4040
rect 15806 3984 15884 4040
rect 15745 3982 15884 3984
rect 15745 3979 15811 3982
rect 15878 3980 15884 3982
rect 15948 3980 15954 4044
rect 14590 3844 14596 3908
rect 14660 3906 14666 3908
rect 17861 3906 17927 3909
rect 14660 3904 17927 3906
rect 14660 3848 17866 3904
rect 17922 3848 17927 3904
rect 14660 3846 17927 3848
rect 14660 3844 14666 3846
rect 17861 3843 17927 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19517 2682 19583 2685
rect 20294 2682 20300 2684
rect 19517 2680 20300 2682
rect 19517 2624 19522 2680
rect 19578 2624 20300 2680
rect 19517 2622 20300 2624
rect 19517 2619 19583 2622
rect 20294 2620 20300 2622
rect 20364 2620 20370 2684
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 39941 98 40007 101
rect 41720 98 42520 128
rect 39941 96 42520 98
rect 39941 40 39946 96
rect 40002 40 42520 96
rect 39941 38 42520 40
rect 39941 35 40007 38
rect 41720 8 42520 38
<< via3 >>
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 14780 41788 14844 41852
rect 19380 41848 19444 41852
rect 19380 41792 19430 41848
rect 19430 41792 19444 41848
rect 19380 41788 19444 41792
rect 30604 41788 30668 41852
rect 20668 41712 20732 41716
rect 20668 41656 20718 41712
rect 20718 41656 20732 41712
rect 20668 41652 20732 41656
rect 10548 41380 10612 41444
rect 23612 41516 23676 41580
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 20116 41304 20180 41308
rect 20116 41248 20166 41304
rect 20166 41248 20180 41304
rect 20116 41244 20180 41248
rect 24900 40836 24964 40900
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19380 40352 19444 40356
rect 19380 40296 19394 40352
rect 19394 40296 19444 40352
rect 19380 40292 19444 40296
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 18460 40080 18524 40084
rect 18460 40024 18474 40080
rect 18474 40024 18524 40080
rect 18460 40020 18524 40024
rect 20116 40216 20180 40220
rect 20116 40160 20166 40216
rect 20166 40160 20180 40216
rect 20116 40156 20180 40160
rect 26188 40156 26252 40220
rect 27292 40216 27356 40220
rect 27292 40160 27306 40216
rect 27306 40160 27356 40216
rect 27292 40156 27356 40160
rect 28396 40080 28460 40084
rect 28396 40024 28410 40080
rect 28410 40024 28460 40080
rect 28396 40020 28460 40024
rect 29684 40020 29748 40084
rect 31156 40020 31220 40084
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 25268 39536 25332 39540
rect 25268 39480 25318 39536
rect 25318 39480 25332 39536
rect 25268 39476 25332 39480
rect 27108 39340 27172 39404
rect 24348 39204 24412 39268
rect 26004 39264 26068 39268
rect 26004 39208 26054 39264
rect 26054 39208 26068 39264
rect 26004 39204 26068 39208
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 23428 38796 23492 38860
rect 25268 38660 25332 38724
rect 28028 38720 28092 38724
rect 28028 38664 28042 38720
rect 28042 38664 28092 38720
rect 28028 38660 28092 38664
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 29500 37980 29564 38044
rect 24164 37904 24228 37908
rect 24164 37848 24178 37904
rect 24178 37848 24228 37904
rect 24164 37844 24228 37848
rect 23612 37708 23676 37772
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 10916 37300 10980 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 19196 36756 19260 36820
rect 15148 36620 15212 36684
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 17540 36076 17604 36140
rect 20116 36076 20180 36140
rect 18644 35940 18708 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 17724 35864 17788 35868
rect 17724 35808 17738 35864
rect 17738 35808 17788 35864
rect 17724 35804 17788 35808
rect 25268 35668 25332 35732
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 9260 34988 9324 35052
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 24900 34716 24964 34780
rect 27660 34716 27724 34780
rect 11100 34640 11164 34644
rect 11100 34584 11114 34640
rect 11114 34584 11164 34640
rect 11100 34580 11164 34584
rect 11468 34580 11532 34644
rect 16804 34580 16868 34644
rect 19196 34580 19260 34644
rect 21772 34580 21836 34644
rect 27476 34640 27540 34644
rect 27476 34584 27490 34640
rect 27490 34584 27540 34640
rect 27476 34580 27540 34584
rect 24716 34444 24780 34508
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 24348 34172 24412 34236
rect 26188 34172 26252 34236
rect 9628 33764 9692 33828
rect 26004 33764 26068 33828
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 25820 33280 25884 33284
rect 25820 33224 25834 33280
rect 25834 33224 25884 33280
rect 25820 33220 25884 33224
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 26924 33084 26988 33148
rect 23428 32948 23492 33012
rect 27108 32948 27172 33012
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 11284 32404 11348 32468
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 10364 31996 10428 32060
rect 16252 32132 16316 32196
rect 21404 32132 21468 32196
rect 29132 32268 29196 32332
rect 22140 32132 22204 32196
rect 23612 32132 23676 32196
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 24900 31724 24964 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 9628 31452 9692 31516
rect 27292 31588 27356 31652
rect 27108 31452 27172 31516
rect 28028 31044 28092 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 23612 30908 23676 30972
rect 24164 30772 24228 30836
rect 29316 30832 29380 30836
rect 29316 30776 29366 30832
rect 29366 30776 29380 30832
rect 29316 30772 29380 30776
rect 21036 30636 21100 30700
rect 21772 30636 21836 30700
rect 24532 30636 24596 30700
rect 20484 30500 20548 30564
rect 27292 30560 27356 30564
rect 27292 30504 27342 30560
rect 27342 30504 27356 30560
rect 27292 30500 27356 30504
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 16068 30364 16132 30428
rect 22692 30424 22756 30428
rect 22692 30368 22742 30424
rect 22742 30368 22756 30424
rect 22692 30364 22756 30368
rect 29500 30228 29564 30292
rect 11652 30092 11716 30156
rect 18644 30092 18708 30156
rect 12572 29956 12636 30020
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 14044 29684 14108 29748
rect 17908 29548 17972 29612
rect 22140 29548 22204 29612
rect 11652 29412 11716 29476
rect 29316 29684 29380 29748
rect 27660 29412 27724 29476
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 9996 29140 10060 29204
rect 19196 29200 19260 29204
rect 19196 29144 19210 29200
rect 19210 29144 19260 29200
rect 19196 29140 19260 29144
rect 16252 29004 16316 29068
rect 18460 29004 18524 29068
rect 20852 29004 20916 29068
rect 29684 28928 29748 28932
rect 29684 28872 29698 28928
rect 29698 28872 29748 28928
rect 29684 28868 29748 28872
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 31156 28732 31220 28796
rect 23428 28596 23492 28660
rect 24900 28324 24964 28388
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 14596 28188 14660 28252
rect 9260 28052 9324 28116
rect 15884 28112 15948 28116
rect 15884 28056 15898 28112
rect 15898 28056 15948 28112
rect 15884 28052 15948 28056
rect 16620 28052 16684 28116
rect 20300 28188 20364 28252
rect 22140 27916 22204 27980
rect 23428 27780 23492 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 16252 27644 16316 27708
rect 18092 27644 18156 27708
rect 12756 27508 12820 27572
rect 26924 27568 26988 27572
rect 26924 27512 26938 27568
rect 26938 27512 26988 27568
rect 26924 27508 26988 27512
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 26556 27100 26620 27164
rect 12572 26828 12636 26892
rect 28396 26888 28460 26892
rect 28396 26832 28410 26888
rect 28410 26832 28460 26888
rect 28396 26828 28460 26832
rect 15148 26692 15212 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 5028 26344 5092 26348
rect 5028 26288 5042 26344
rect 5042 26288 5092 26344
rect 5028 26284 5092 26288
rect 9996 26284 10060 26348
rect 10364 26148 10428 26212
rect 26556 26208 26620 26212
rect 26556 26152 26570 26208
rect 26570 26152 26620 26208
rect 26556 26148 26620 26152
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 18828 26072 18892 26076
rect 18828 26016 18842 26072
rect 18842 26016 18892 26072
rect 18828 26012 18892 26016
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 18092 25060 18156 25124
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 11652 24788 11716 24852
rect 25820 24788 25884 24852
rect 29316 24848 29380 24852
rect 29316 24792 29330 24848
rect 29330 24792 29380 24848
rect 29316 24788 29380 24792
rect 22692 24576 22756 24580
rect 22692 24520 22742 24576
rect 22742 24520 22756 24576
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 16068 24244 16132 24308
rect 22692 24516 22756 24520
rect 24900 24652 24964 24716
rect 25268 24652 25332 24716
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 30604 24304 30668 24308
rect 30604 24248 30618 24304
rect 30618 24248 30668 24304
rect 30604 24244 30668 24248
rect 20300 24168 20364 24172
rect 20300 24112 20350 24168
rect 20350 24112 20364 24168
rect 20300 24108 20364 24112
rect 16620 23972 16684 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 18092 23700 18156 23764
rect 12388 23428 12452 23492
rect 21404 23428 21468 23492
rect 29132 23428 29196 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 9444 23156 9508 23220
rect 21036 23080 21100 23084
rect 21036 23024 21086 23080
rect 21086 23024 21100 23080
rect 21036 23020 21100 23024
rect 17908 22884 17972 22948
rect 18828 22884 18892 22948
rect 19196 22944 19260 22948
rect 19196 22888 19246 22944
rect 19246 22888 19260 22944
rect 19196 22884 19260 22888
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 11468 21856 11532 21860
rect 11468 21800 11482 21856
rect 11482 21800 11532 21856
rect 11468 21796 11532 21800
rect 12388 21796 12452 21860
rect 22140 21796 22204 21860
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 20484 21524 20548 21588
rect 24532 21524 24596 21588
rect 14780 21312 14844 21316
rect 14780 21256 14794 21312
rect 14794 21256 14844 21312
rect 14780 21252 14844 21256
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 15884 21116 15948 21180
rect 18092 21176 18156 21180
rect 18092 21120 18142 21176
rect 18142 21120 18156 21176
rect 18092 21116 18156 21120
rect 20300 20844 20364 20908
rect 26372 20904 26436 20908
rect 26372 20848 26386 20904
rect 26386 20848 26436 20904
rect 26372 20844 26436 20848
rect 5212 20768 5276 20772
rect 5212 20712 5226 20768
rect 5226 20712 5276 20768
rect 5212 20708 5276 20712
rect 24716 20708 24780 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 12572 20572 12636 20636
rect 15148 20572 15212 20636
rect 28948 20572 29012 20636
rect 14044 20360 14108 20364
rect 14044 20304 14058 20360
rect 14058 20304 14108 20360
rect 14044 20300 14108 20304
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 23428 20028 23492 20092
rect 11284 19620 11348 19684
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 23428 19348 23492 19412
rect 16804 19272 16868 19276
rect 16804 19216 16818 19272
rect 16818 19216 16868 19272
rect 16804 19212 16868 19216
rect 20116 19212 20180 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 11100 18804 11164 18868
rect 20852 18668 20916 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 10548 18320 10612 18324
rect 10548 18264 10562 18320
rect 10562 18264 10612 18320
rect 10548 18260 10612 18264
rect 29132 18260 29196 18324
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 25452 17716 25516 17780
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 23244 17172 23308 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 17540 16764 17604 16828
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 25452 16084 25516 16148
rect 26004 16084 26068 16148
rect 5028 15812 5092 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 10916 15540 10980 15604
rect 18276 15540 18340 15604
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 14964 15192 15028 15196
rect 14964 15136 14978 15192
rect 14978 15136 15028 15192
rect 14964 15132 15028 15136
rect 17724 15132 17788 15196
rect 28948 15132 29012 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 18092 14588 18156 14652
rect 20668 14588 20732 14652
rect 23428 14588 23492 14652
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 5212 13696 5276 13700
rect 5212 13640 5262 13696
rect 5262 13640 5276 13696
rect 5212 13636 5276 13640
rect 18092 13636 18156 13700
rect 29132 13636 29196 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 26556 11460 26620 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 15884 10916 15948 10980
rect 23244 10976 23308 10980
rect 23244 10920 23258 10976
rect 23258 10920 23308 10976
rect 23244 10916 23308 10920
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 26372 10780 26436 10844
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 9444 6700 9508 6764
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 26004 5264 26068 5268
rect 26004 5208 26018 5264
rect 26018 5208 26068 5264
rect 26004 5204 26068 5208
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 26556 4796 26620 4860
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 15884 3980 15948 4044
rect 14596 3844 14660 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 20300 2620 20364 2684
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 41920 4528 42480
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 19568 42464 19888 42480
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 14779 41852 14845 41853
rect 14779 41788 14780 41852
rect 14844 41788 14845 41852
rect 14779 41787 14845 41788
rect 19379 41852 19445 41853
rect 19379 41788 19380 41852
rect 19444 41788 19445 41852
rect 19379 41787 19445 41788
rect 10547 41444 10613 41445
rect 10547 41380 10548 41444
rect 10612 41380 10613 41444
rect 10547 41379 10613 41380
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 9259 35052 9325 35053
rect 9259 34988 9260 35052
rect 9324 34988 9325 35052
rect 9259 34987 9325 34988
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 9262 28117 9322 34987
rect 9627 33828 9693 33829
rect 9627 33764 9628 33828
rect 9692 33764 9693 33828
rect 9627 33763 9693 33764
rect 9630 31517 9690 33763
rect 10363 32060 10429 32061
rect 10363 31996 10364 32060
rect 10428 31996 10429 32060
rect 10363 31995 10429 31996
rect 9627 31516 9693 31517
rect 9627 31452 9628 31516
rect 9692 31452 9693 31516
rect 9627 31451 9693 31452
rect 9995 29204 10061 29205
rect 9995 29140 9996 29204
rect 10060 29140 10061 29204
rect 9995 29139 10061 29140
rect 9259 28116 9325 28117
rect 9259 28052 9260 28116
rect 9324 28052 9325 28116
rect 9259 28051 9325 28052
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 9998 26349 10058 29139
rect 5027 26348 5093 26349
rect 5027 26284 5028 26348
rect 5092 26284 5093 26348
rect 5027 26283 5093 26284
rect 9995 26348 10061 26349
rect 9995 26284 9996 26348
rect 10060 26284 10061 26348
rect 9995 26283 10061 26284
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 5030 15877 5090 26283
rect 10366 26213 10426 31995
rect 10363 26212 10429 26213
rect 10363 26148 10364 26212
rect 10428 26148 10429 26212
rect 10363 26147 10429 26148
rect 9443 23220 9509 23221
rect 9443 23156 9444 23220
rect 9508 23156 9509 23220
rect 9443 23155 9509 23156
rect 5211 20772 5277 20773
rect 5211 20708 5212 20772
rect 5276 20708 5277 20772
rect 5211 20707 5277 20708
rect 5027 15876 5093 15877
rect 5027 15812 5028 15876
rect 5092 15812 5093 15876
rect 5027 15811 5093 15812
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 5214 13701 5274 20707
rect 5211 13700 5277 13701
rect 5211 13636 5212 13700
rect 5276 13636 5277 13700
rect 5211 13635 5277 13636
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 9446 6765 9506 23155
rect 10550 18325 10610 41379
rect 10915 37364 10981 37365
rect 10915 37300 10916 37364
rect 10980 37300 10981 37364
rect 10915 37299 10981 37300
rect 10547 18324 10613 18325
rect 10547 18260 10548 18324
rect 10612 18260 10613 18324
rect 10547 18259 10613 18260
rect 10918 15605 10978 37299
rect 11099 34644 11165 34645
rect 11099 34580 11100 34644
rect 11164 34580 11165 34644
rect 11099 34579 11165 34580
rect 11467 34644 11533 34645
rect 11467 34580 11468 34644
rect 11532 34580 11533 34644
rect 11467 34579 11533 34580
rect 11102 18869 11162 34579
rect 11283 32468 11349 32469
rect 11283 32404 11284 32468
rect 11348 32404 11349 32468
rect 11283 32403 11349 32404
rect 11286 19685 11346 32403
rect 11470 21861 11530 34579
rect 11651 30156 11717 30157
rect 11651 30092 11652 30156
rect 11716 30092 11717 30156
rect 11651 30091 11717 30092
rect 11654 29477 11714 30091
rect 12571 30020 12637 30021
rect 12571 29956 12572 30020
rect 12636 29956 12637 30020
rect 12571 29955 12637 29956
rect 11651 29476 11717 29477
rect 11651 29412 11652 29476
rect 11716 29412 11717 29476
rect 11651 29411 11717 29412
rect 11654 24853 11714 29411
rect 12574 26893 12634 29955
rect 14043 29748 14109 29749
rect 14043 29684 14044 29748
rect 14108 29684 14109 29748
rect 14043 29683 14109 29684
rect 12755 27572 12821 27573
rect 12755 27508 12756 27572
rect 12820 27508 12821 27572
rect 12755 27507 12821 27508
rect 12571 26892 12637 26893
rect 12571 26828 12572 26892
rect 12636 26828 12637 26892
rect 12571 26827 12637 26828
rect 11651 24852 11717 24853
rect 11651 24788 11652 24852
rect 11716 24788 11717 24852
rect 11651 24787 11717 24788
rect 12387 23492 12453 23493
rect 12387 23428 12388 23492
rect 12452 23490 12453 23492
rect 12452 23430 12634 23490
rect 12452 23428 12453 23430
rect 12387 23427 12453 23428
rect 12574 22810 12634 23430
rect 12390 22750 12634 22810
rect 12390 21861 12450 22750
rect 12758 22110 12818 27507
rect 12574 22050 12818 22110
rect 11467 21860 11533 21861
rect 11467 21796 11468 21860
rect 11532 21796 11533 21860
rect 11467 21795 11533 21796
rect 12387 21860 12453 21861
rect 12387 21796 12388 21860
rect 12452 21796 12453 21860
rect 12387 21795 12453 21796
rect 12574 20637 12634 22050
rect 12571 20636 12637 20637
rect 12571 20572 12572 20636
rect 12636 20572 12637 20636
rect 12571 20571 12637 20572
rect 14046 20365 14106 29683
rect 14595 28252 14661 28253
rect 14595 28188 14596 28252
rect 14660 28188 14661 28252
rect 14595 28187 14661 28188
rect 14043 20364 14109 20365
rect 14043 20300 14044 20364
rect 14108 20300 14109 20364
rect 14043 20299 14109 20300
rect 11283 19684 11349 19685
rect 11283 19620 11284 19684
rect 11348 19620 11349 19684
rect 11283 19619 11349 19620
rect 11099 18868 11165 18869
rect 11099 18804 11100 18868
rect 11164 18804 11165 18868
rect 11099 18803 11165 18804
rect 10915 15604 10981 15605
rect 10915 15540 10916 15604
rect 10980 15540 10981 15604
rect 10915 15539 10981 15540
rect 9443 6764 9509 6765
rect 9443 6700 9444 6764
rect 9508 6700 9509 6764
rect 9443 6699 9509 6700
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 14598 3909 14658 28187
rect 14782 21317 14842 41787
rect 19382 40357 19442 41787
rect 19568 41376 19888 42400
rect 34928 41920 35248 42480
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 30603 41852 30669 41853
rect 30603 41788 30604 41852
rect 30668 41788 30669 41852
rect 30603 41787 30669 41788
rect 20667 41716 20733 41717
rect 20667 41652 20668 41716
rect 20732 41652 20733 41716
rect 20667 41651 20733 41652
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19379 40356 19445 40357
rect 19379 40292 19380 40356
rect 19444 40292 19445 40356
rect 19379 40291 19445 40292
rect 19568 40288 19888 41312
rect 20115 41308 20181 41309
rect 20115 41244 20116 41308
rect 20180 41244 20181 41308
rect 20115 41243 20181 41244
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 18459 40084 18525 40085
rect 18459 40020 18460 40084
rect 18524 40020 18525 40084
rect 18459 40019 18525 40020
rect 15147 36684 15213 36685
rect 15147 36620 15148 36684
rect 15212 36620 15213 36684
rect 15147 36619 15213 36620
rect 15150 26890 15210 36619
rect 17539 36140 17605 36141
rect 17539 36076 17540 36140
rect 17604 36076 17605 36140
rect 17539 36075 17605 36076
rect 16803 34644 16869 34645
rect 16803 34580 16804 34644
rect 16868 34580 16869 34644
rect 16803 34579 16869 34580
rect 16251 32196 16317 32197
rect 16251 32132 16252 32196
rect 16316 32132 16317 32196
rect 16251 32131 16317 32132
rect 16067 30428 16133 30429
rect 16067 30364 16068 30428
rect 16132 30364 16133 30428
rect 16067 30363 16133 30364
rect 15883 28116 15949 28117
rect 15883 28052 15884 28116
rect 15948 28052 15949 28116
rect 15883 28051 15949 28052
rect 14966 26830 15210 26890
rect 14779 21316 14845 21317
rect 14779 21252 14780 21316
rect 14844 21252 14845 21316
rect 14779 21251 14845 21252
rect 14966 15197 15026 26830
rect 15147 26756 15213 26757
rect 15147 26692 15148 26756
rect 15212 26692 15213 26756
rect 15147 26691 15213 26692
rect 15150 20637 15210 26691
rect 15886 21181 15946 28051
rect 16070 24309 16130 30363
rect 16254 29069 16314 32131
rect 16251 29068 16317 29069
rect 16251 29004 16252 29068
rect 16316 29004 16317 29068
rect 16251 29003 16317 29004
rect 16254 27709 16314 29003
rect 16619 28116 16685 28117
rect 16619 28052 16620 28116
rect 16684 28052 16685 28116
rect 16619 28051 16685 28052
rect 16251 27708 16317 27709
rect 16251 27644 16252 27708
rect 16316 27644 16317 27708
rect 16251 27643 16317 27644
rect 16067 24308 16133 24309
rect 16067 24244 16068 24308
rect 16132 24244 16133 24308
rect 16067 24243 16133 24244
rect 16622 24037 16682 28051
rect 16619 24036 16685 24037
rect 16619 23972 16620 24036
rect 16684 23972 16685 24036
rect 16619 23971 16685 23972
rect 15883 21180 15949 21181
rect 15883 21116 15884 21180
rect 15948 21116 15949 21180
rect 15883 21115 15949 21116
rect 15147 20636 15213 20637
rect 15147 20572 15148 20636
rect 15212 20572 15213 20636
rect 15147 20571 15213 20572
rect 16806 19277 16866 34579
rect 16803 19276 16869 19277
rect 16803 19212 16804 19276
rect 16868 19212 16869 19276
rect 16803 19211 16869 19212
rect 17542 16829 17602 36075
rect 17723 35868 17789 35869
rect 17723 35804 17724 35868
rect 17788 35804 17789 35868
rect 17723 35803 17789 35804
rect 17539 16828 17605 16829
rect 17539 16764 17540 16828
rect 17604 16764 17605 16828
rect 17539 16763 17605 16764
rect 17726 15197 17786 35803
rect 17907 29612 17973 29613
rect 17907 29548 17908 29612
rect 17972 29548 17973 29612
rect 17907 29547 17973 29548
rect 17910 22949 17970 29547
rect 18462 29069 18522 40019
rect 19568 39200 19888 40224
rect 20118 40221 20178 41243
rect 20115 40220 20181 40221
rect 20115 40156 20116 40220
rect 20180 40156 20181 40220
rect 20115 40155 20181 40156
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19195 36820 19261 36821
rect 19195 36756 19196 36820
rect 19260 36756 19261 36820
rect 19195 36755 19261 36756
rect 18643 36004 18709 36005
rect 18643 35940 18644 36004
rect 18708 35940 18709 36004
rect 18643 35939 18709 35940
rect 18646 30157 18706 35939
rect 19198 34645 19258 36755
rect 19568 35936 19888 36960
rect 20115 36140 20181 36141
rect 20115 36076 20116 36140
rect 20180 36076 20181 36140
rect 20115 36075 20181 36076
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19195 34644 19261 34645
rect 19195 34580 19196 34644
rect 19260 34580 19261 34644
rect 19195 34579 19261 34580
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 18643 30156 18709 30157
rect 18643 30092 18644 30156
rect 18708 30092 18709 30156
rect 18643 30091 18709 30092
rect 18459 29068 18525 29069
rect 18459 29004 18460 29068
rect 18524 29004 18525 29068
rect 18459 29003 18525 29004
rect 18091 27708 18157 27709
rect 18091 27644 18092 27708
rect 18156 27644 18157 27708
rect 18091 27643 18157 27644
rect 18094 25125 18154 27643
rect 18091 25124 18157 25125
rect 18091 25060 18092 25124
rect 18156 25060 18157 25124
rect 18091 25059 18157 25060
rect 18091 23764 18157 23765
rect 18091 23700 18092 23764
rect 18156 23700 18157 23764
rect 18091 23699 18157 23700
rect 17907 22948 17973 22949
rect 17907 22884 17908 22948
rect 17972 22884 17973 22948
rect 17907 22883 17973 22884
rect 18094 21181 18154 23699
rect 18646 22110 18706 30091
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19195 29204 19261 29205
rect 19195 29140 19196 29204
rect 19260 29140 19261 29204
rect 19195 29139 19261 29140
rect 18827 26076 18893 26077
rect 18827 26012 18828 26076
rect 18892 26012 18893 26076
rect 18827 26011 18893 26012
rect 18830 22949 18890 26011
rect 19198 22949 19258 29139
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 18827 22948 18893 22949
rect 18827 22884 18828 22948
rect 18892 22884 18893 22948
rect 18827 22883 18893 22884
rect 19195 22948 19261 22949
rect 19195 22884 19196 22948
rect 19260 22884 19261 22948
rect 19195 22883 19261 22884
rect 18278 22050 18706 22110
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 18091 21180 18157 21181
rect 18091 21116 18092 21180
rect 18156 21116 18157 21180
rect 18091 21115 18157 21116
rect 18278 15605 18338 22050
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 20118 19277 20178 36075
rect 20483 30564 20549 30565
rect 20483 30500 20484 30564
rect 20548 30500 20549 30564
rect 20483 30499 20549 30500
rect 20299 28252 20365 28253
rect 20299 28188 20300 28252
rect 20364 28188 20365 28252
rect 20299 28187 20365 28188
rect 20302 24173 20362 28187
rect 20299 24172 20365 24173
rect 20299 24108 20300 24172
rect 20364 24108 20365 24172
rect 20299 24107 20365 24108
rect 20486 21589 20546 30499
rect 20483 21588 20549 21589
rect 20483 21524 20484 21588
rect 20548 21524 20549 21588
rect 20483 21523 20549 21524
rect 20299 20908 20365 20909
rect 20299 20844 20300 20908
rect 20364 20844 20365 20908
rect 20299 20843 20365 20844
rect 20115 19276 20181 19277
rect 20115 19212 20116 19276
rect 20180 19212 20181 19276
rect 20115 19211 20181 19212
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 18275 15604 18341 15605
rect 18275 15540 18276 15604
rect 18340 15540 18341 15604
rect 18275 15539 18341 15540
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 14963 15196 15029 15197
rect 14963 15132 14964 15196
rect 15028 15132 15029 15196
rect 14963 15131 15029 15132
rect 17723 15196 17789 15197
rect 17723 15132 17724 15196
rect 17788 15132 17789 15196
rect 17723 15131 17789 15132
rect 18091 14652 18157 14653
rect 18091 14588 18092 14652
rect 18156 14588 18157 14652
rect 18091 14587 18157 14588
rect 18094 13701 18154 14587
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 18091 13700 18157 13701
rect 18091 13636 18092 13700
rect 18156 13636 18157 13700
rect 18091 13635 18157 13636
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 15883 10980 15949 10981
rect 15883 10916 15884 10980
rect 15948 10916 15949 10980
rect 15883 10915 15949 10916
rect 15886 4045 15946 10915
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 15883 4044 15949 4045
rect 15883 3980 15884 4044
rect 15948 3980 15949 4044
rect 15883 3979 15949 3980
rect 14595 3908 14661 3909
rect 14595 3844 14596 3908
rect 14660 3844 14661 3908
rect 14595 3843 14661 3844
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 20302 2685 20362 20843
rect 20670 14653 20730 41651
rect 23611 41580 23677 41581
rect 23611 41516 23612 41580
rect 23676 41516 23677 41580
rect 23611 41515 23677 41516
rect 23427 38860 23493 38861
rect 23427 38796 23428 38860
rect 23492 38796 23493 38860
rect 23427 38795 23493 38796
rect 23430 35050 23490 38795
rect 23614 37773 23674 41515
rect 24899 40900 24965 40901
rect 24899 40836 24900 40900
rect 24964 40836 24965 40900
rect 24899 40835 24965 40836
rect 24347 39268 24413 39269
rect 24347 39204 24348 39268
rect 24412 39204 24413 39268
rect 24347 39203 24413 39204
rect 24163 37908 24229 37909
rect 24163 37844 24164 37908
rect 24228 37844 24229 37908
rect 24163 37843 24229 37844
rect 23611 37772 23677 37773
rect 23611 37708 23612 37772
rect 23676 37708 23677 37772
rect 23611 37707 23677 37708
rect 23430 34990 23674 35050
rect 21771 34644 21837 34645
rect 21771 34580 21772 34644
rect 21836 34580 21837 34644
rect 21771 34579 21837 34580
rect 21403 32196 21469 32197
rect 21403 32132 21404 32196
rect 21468 32132 21469 32196
rect 21403 32131 21469 32132
rect 21035 30700 21101 30701
rect 21035 30636 21036 30700
rect 21100 30636 21101 30700
rect 21035 30635 21101 30636
rect 20851 29068 20917 29069
rect 20851 29004 20852 29068
rect 20916 29004 20917 29068
rect 20851 29003 20917 29004
rect 20854 18733 20914 29003
rect 21038 23085 21098 30635
rect 21406 23493 21466 32131
rect 21774 30701 21834 34579
rect 23427 33012 23493 33013
rect 23427 32948 23428 33012
rect 23492 32948 23493 33012
rect 23427 32947 23493 32948
rect 22139 32196 22205 32197
rect 22139 32132 22140 32196
rect 22204 32132 22205 32196
rect 22139 32131 22205 32132
rect 21771 30700 21837 30701
rect 21771 30636 21772 30700
rect 21836 30636 21837 30700
rect 21771 30635 21837 30636
rect 22142 29613 22202 32131
rect 22691 30428 22757 30429
rect 22691 30364 22692 30428
rect 22756 30364 22757 30428
rect 22691 30363 22757 30364
rect 22139 29612 22205 29613
rect 22139 29548 22140 29612
rect 22204 29548 22205 29612
rect 22139 29547 22205 29548
rect 22139 27980 22205 27981
rect 22139 27916 22140 27980
rect 22204 27916 22205 27980
rect 22139 27915 22205 27916
rect 21403 23492 21469 23493
rect 21403 23428 21404 23492
rect 21468 23428 21469 23492
rect 21403 23427 21469 23428
rect 21035 23084 21101 23085
rect 21035 23020 21036 23084
rect 21100 23020 21101 23084
rect 21035 23019 21101 23020
rect 22142 21861 22202 27915
rect 22694 24581 22754 30363
rect 23430 28661 23490 32947
rect 23614 32197 23674 34990
rect 23611 32196 23677 32197
rect 23611 32132 23612 32196
rect 23676 32132 23677 32196
rect 23611 32131 23677 32132
rect 23614 30973 23674 32131
rect 23611 30972 23677 30973
rect 23611 30908 23612 30972
rect 23676 30908 23677 30972
rect 23611 30907 23677 30908
rect 24166 30837 24226 37843
rect 24350 34237 24410 39203
rect 24902 34781 24962 40835
rect 26187 40220 26253 40221
rect 26187 40156 26188 40220
rect 26252 40156 26253 40220
rect 26187 40155 26253 40156
rect 27291 40220 27357 40221
rect 27291 40156 27292 40220
rect 27356 40156 27357 40220
rect 27291 40155 27357 40156
rect 25267 39540 25333 39541
rect 25267 39476 25268 39540
rect 25332 39476 25333 39540
rect 25267 39475 25333 39476
rect 25270 38725 25330 39475
rect 26003 39268 26069 39269
rect 26003 39204 26004 39268
rect 26068 39204 26069 39268
rect 26003 39203 26069 39204
rect 25267 38724 25333 38725
rect 25267 38660 25268 38724
rect 25332 38660 25333 38724
rect 25267 38659 25333 38660
rect 25267 35732 25333 35733
rect 25267 35668 25268 35732
rect 25332 35668 25333 35732
rect 25267 35667 25333 35668
rect 24899 34780 24965 34781
rect 24899 34716 24900 34780
rect 24964 34716 24965 34780
rect 24899 34715 24965 34716
rect 24715 34508 24781 34509
rect 24715 34444 24716 34508
rect 24780 34444 24781 34508
rect 24715 34443 24781 34444
rect 24347 34236 24413 34237
rect 24347 34172 24348 34236
rect 24412 34172 24413 34236
rect 24347 34171 24413 34172
rect 24163 30836 24229 30837
rect 24163 30772 24164 30836
rect 24228 30772 24229 30836
rect 24163 30771 24229 30772
rect 24531 30700 24597 30701
rect 24531 30636 24532 30700
rect 24596 30636 24597 30700
rect 24531 30635 24597 30636
rect 23427 28660 23493 28661
rect 23427 28596 23428 28660
rect 23492 28596 23493 28660
rect 23427 28595 23493 28596
rect 23427 27844 23493 27845
rect 23427 27780 23428 27844
rect 23492 27780 23493 27844
rect 23427 27779 23493 27780
rect 22691 24580 22757 24581
rect 22691 24516 22692 24580
rect 22756 24516 22757 24580
rect 22691 24515 22757 24516
rect 22139 21860 22205 21861
rect 22139 21796 22140 21860
rect 22204 21796 22205 21860
rect 22139 21795 22205 21796
rect 23430 20093 23490 27779
rect 24534 21589 24594 30635
rect 24531 21588 24597 21589
rect 24531 21524 24532 21588
rect 24596 21524 24597 21588
rect 24531 21523 24597 21524
rect 24718 20773 24778 34443
rect 24902 31789 24962 34715
rect 24899 31788 24965 31789
rect 24899 31724 24900 31788
rect 24964 31724 24965 31788
rect 24899 31723 24965 31724
rect 24902 28389 24962 31723
rect 24899 28388 24965 28389
rect 24899 28324 24900 28388
rect 24964 28324 24965 28388
rect 24899 28323 24965 28324
rect 24902 24717 24962 28323
rect 25270 24717 25330 35667
rect 26006 33829 26066 39203
rect 26190 34237 26250 40155
rect 27107 39404 27173 39405
rect 27107 39340 27108 39404
rect 27172 39340 27173 39404
rect 27107 39339 27173 39340
rect 26187 34236 26253 34237
rect 26187 34172 26188 34236
rect 26252 34172 26253 34236
rect 26187 34171 26253 34172
rect 26003 33828 26069 33829
rect 26003 33764 26004 33828
rect 26068 33764 26069 33828
rect 26003 33763 26069 33764
rect 25819 33284 25885 33285
rect 25819 33220 25820 33284
rect 25884 33220 25885 33284
rect 25819 33219 25885 33220
rect 25822 24853 25882 33219
rect 26923 33148 26989 33149
rect 26923 33084 26924 33148
rect 26988 33084 26989 33148
rect 26923 33083 26989 33084
rect 26926 27573 26986 33083
rect 27110 33013 27170 39339
rect 27107 33012 27173 33013
rect 27107 32948 27108 33012
rect 27172 32948 27173 33012
rect 27107 32947 27173 32948
rect 27294 31653 27354 40155
rect 28395 40084 28461 40085
rect 28395 40020 28396 40084
rect 28460 40020 28461 40084
rect 28395 40019 28461 40020
rect 29683 40084 29749 40085
rect 29683 40020 29684 40084
rect 29748 40020 29749 40084
rect 29683 40019 29749 40020
rect 28027 38724 28093 38725
rect 28027 38660 28028 38724
rect 28092 38660 28093 38724
rect 28027 38659 28093 38660
rect 27659 34780 27725 34781
rect 27659 34716 27660 34780
rect 27724 34716 27725 34780
rect 27659 34715 27725 34716
rect 27475 34644 27541 34645
rect 27475 34580 27476 34644
rect 27540 34580 27541 34644
rect 27475 34579 27541 34580
rect 27291 31652 27357 31653
rect 27291 31588 27292 31652
rect 27356 31588 27357 31652
rect 27291 31587 27357 31588
rect 27107 31516 27173 31517
rect 27107 31452 27108 31516
rect 27172 31452 27173 31516
rect 27107 31451 27173 31452
rect 27110 30970 27170 31451
rect 27478 30970 27538 34579
rect 27110 30910 27538 30970
rect 27294 30565 27354 30910
rect 27291 30564 27357 30565
rect 27291 30500 27292 30564
rect 27356 30500 27357 30564
rect 27291 30499 27357 30500
rect 27662 29477 27722 34715
rect 28030 31109 28090 38659
rect 28027 31108 28093 31109
rect 28027 31044 28028 31108
rect 28092 31044 28093 31108
rect 28027 31043 28093 31044
rect 27659 29476 27725 29477
rect 27659 29412 27660 29476
rect 27724 29412 27725 29476
rect 27659 29411 27725 29412
rect 26923 27572 26989 27573
rect 26923 27508 26924 27572
rect 26988 27508 26989 27572
rect 26923 27507 26989 27508
rect 26555 27164 26621 27165
rect 26555 27100 26556 27164
rect 26620 27100 26621 27164
rect 26555 27099 26621 27100
rect 26558 26213 26618 27099
rect 28398 26893 28458 40019
rect 29499 38044 29565 38045
rect 29499 37980 29500 38044
rect 29564 37980 29565 38044
rect 29499 37979 29565 37980
rect 29131 32332 29197 32333
rect 29131 32268 29132 32332
rect 29196 32268 29197 32332
rect 29131 32267 29197 32268
rect 28395 26892 28461 26893
rect 28395 26828 28396 26892
rect 28460 26828 28461 26892
rect 28395 26827 28461 26828
rect 26555 26212 26621 26213
rect 26555 26148 26556 26212
rect 26620 26148 26621 26212
rect 26555 26147 26621 26148
rect 25819 24852 25885 24853
rect 25819 24788 25820 24852
rect 25884 24788 25885 24852
rect 25819 24787 25885 24788
rect 24899 24716 24965 24717
rect 24899 24652 24900 24716
rect 24964 24652 24965 24716
rect 24899 24651 24965 24652
rect 25267 24716 25333 24717
rect 25267 24652 25268 24716
rect 25332 24652 25333 24716
rect 25267 24651 25333 24652
rect 29134 23493 29194 32267
rect 29315 30836 29381 30837
rect 29315 30772 29316 30836
rect 29380 30772 29381 30836
rect 29315 30771 29381 30772
rect 29318 29749 29378 30771
rect 29502 30293 29562 37979
rect 29499 30292 29565 30293
rect 29499 30228 29500 30292
rect 29564 30228 29565 30292
rect 29499 30227 29565 30228
rect 29315 29748 29381 29749
rect 29315 29684 29316 29748
rect 29380 29684 29381 29748
rect 29315 29683 29381 29684
rect 29318 24853 29378 29683
rect 29686 28933 29746 40019
rect 29683 28932 29749 28933
rect 29683 28868 29684 28932
rect 29748 28868 29749 28932
rect 29683 28867 29749 28868
rect 29315 24852 29381 24853
rect 29315 24788 29316 24852
rect 29380 24788 29381 24852
rect 29315 24787 29381 24788
rect 30606 24309 30666 41787
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 31155 40084 31221 40085
rect 31155 40020 31156 40084
rect 31220 40020 31221 40084
rect 31155 40019 31221 40020
rect 31158 28797 31218 40019
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 31155 28796 31221 28797
rect 31155 28732 31156 28796
rect 31220 28732 31221 28796
rect 31155 28731 31221 28732
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 30603 24308 30669 24309
rect 30603 24244 30604 24308
rect 30668 24244 30669 24308
rect 30603 24243 30669 24244
rect 29131 23492 29197 23493
rect 29131 23428 29132 23492
rect 29196 23428 29197 23492
rect 29131 23427 29197 23428
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 26371 20908 26437 20909
rect 26371 20844 26372 20908
rect 26436 20844 26437 20908
rect 26371 20843 26437 20844
rect 24715 20772 24781 20773
rect 24715 20708 24716 20772
rect 24780 20708 24781 20772
rect 24715 20707 24781 20708
rect 23427 20092 23493 20093
rect 23427 20028 23428 20092
rect 23492 20028 23493 20092
rect 23427 20027 23493 20028
rect 23427 19412 23493 19413
rect 23427 19348 23428 19412
rect 23492 19348 23493 19412
rect 23427 19347 23493 19348
rect 20851 18732 20917 18733
rect 20851 18668 20852 18732
rect 20916 18668 20917 18732
rect 20851 18667 20917 18668
rect 23243 17236 23309 17237
rect 23243 17172 23244 17236
rect 23308 17172 23309 17236
rect 23243 17171 23309 17172
rect 20667 14652 20733 14653
rect 20667 14588 20668 14652
rect 20732 14588 20733 14652
rect 20667 14587 20733 14588
rect 23246 10981 23306 17171
rect 23430 14653 23490 19347
rect 25451 17780 25517 17781
rect 25451 17716 25452 17780
rect 25516 17716 25517 17780
rect 25451 17715 25517 17716
rect 25454 16149 25514 17715
rect 25451 16148 25517 16149
rect 25451 16084 25452 16148
rect 25516 16084 25517 16148
rect 25451 16083 25517 16084
rect 26003 16148 26069 16149
rect 26003 16084 26004 16148
rect 26068 16084 26069 16148
rect 26003 16083 26069 16084
rect 23427 14652 23493 14653
rect 23427 14588 23428 14652
rect 23492 14588 23493 14652
rect 23427 14587 23493 14588
rect 23243 10980 23309 10981
rect 23243 10916 23244 10980
rect 23308 10916 23309 10980
rect 23243 10915 23309 10916
rect 26006 5269 26066 16083
rect 26374 10845 26434 20843
rect 28947 20636 29013 20637
rect 28947 20572 28948 20636
rect 29012 20572 29013 20636
rect 28947 20571 29013 20572
rect 28950 15197 29010 20571
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 29131 18324 29197 18325
rect 29131 18260 29132 18324
rect 29196 18260 29197 18324
rect 29131 18259 29197 18260
rect 28947 15196 29013 15197
rect 28947 15132 28948 15196
rect 29012 15132 29013 15196
rect 28947 15131 29013 15132
rect 29134 13701 29194 18259
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 29131 13700 29197 13701
rect 29131 13636 29132 13700
rect 29196 13636 29197 13700
rect 29131 13635 29197 13636
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 26555 11524 26621 11525
rect 26555 11460 26556 11524
rect 26620 11460 26621 11524
rect 26555 11459 26621 11460
rect 26371 10844 26437 10845
rect 26371 10780 26372 10844
rect 26436 10780 26437 10844
rect 26371 10779 26437 10780
rect 26003 5268 26069 5269
rect 26003 5204 26004 5268
rect 26068 5204 26069 5268
rect 26003 5203 26069 5204
rect 26558 4861 26618 11459
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 26555 4860 26621 4861
rect 26555 4796 26556 4860
rect 26620 4796 26621 4860
rect 26555 4795 26621 4796
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 20299 2684 20365 2685
rect 20299 2620 20300 2684
rect 20364 2620 20365 2684
rect 20299 2619 20365 2620
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__clkbuf_2  _1503_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35052 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1504_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35420 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1505_
timestamp 1688980957
transform 1 0 35512 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1506_
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_1  _1507_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34868 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1508_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1509_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33488 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1510_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1511_
timestamp 1688980957
transform 1 0 33488 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1512_
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1513_
timestamp 1688980957
transform 1 0 32016 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1514_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27968 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _1515_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1516_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1517_
timestamp 1688980957
transform 1 0 33304 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1518_
timestamp 1688980957
transform 1 0 32660 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _1519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31004 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  _1520_
timestamp 1688980957
transform 1 0 28336 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1521_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_4  _1522_
timestamp 1688980957
transform 1 0 31004 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  _1523_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _1524_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27048 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1525_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1526_
timestamp 1688980957
transform 1 0 34040 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1527_
timestamp 1688980957
transform 1 0 33396 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1528_
timestamp 1688980957
transform 1 0 33488 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1529_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1530_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25392 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand4b_2  _1531_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1532_
timestamp 1688980957
transform 1 0 28336 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1533_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21344 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1534_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30544 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1535_
timestamp 1688980957
transform 1 0 30084 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1536_
timestamp 1688980957
transform 1 0 35144 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1537_
timestamp 1688980957
transform 1 0 34040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1538_
timestamp 1688980957
transform 1 0 29532 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1539_
timestamp 1688980957
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1540_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29716 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1541_
timestamp 1688980957
transform 1 0 28888 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1542_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21620 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1543_
timestamp 1688980957
transform 1 0 26312 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1544_
timestamp 1688980957
transform 1 0 34040 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1545_
timestamp 1688980957
transform 1 0 33856 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1546_
timestamp 1688980957
transform 1 0 25576 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1547_
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1548_
timestamp 1688980957
transform 1 0 34500 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1549_
timestamp 1688980957
transform 1 0 25852 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_4  _1550_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32752 0 -1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__or2b_1  _1551_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29624 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1552_
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1553_
timestamp 1688980957
transform 1 0 35236 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_4  _1554_
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__a41o_1  _1555_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1556_
timestamp 1688980957
transform 1 0 25576 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1557_
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  _1558_
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  _1559_
timestamp 1688980957
transform 1 0 27784 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1560_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23828 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1561_
timestamp 1688980957
transform 1 0 29992 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1562_
timestamp 1688980957
transform 1 0 31648 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1563_
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1564_
timestamp 1688980957
transform 1 0 27600 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1565_
timestamp 1688980957
transform 1 0 23828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1566_
timestamp 1688980957
transform 1 0 27048 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1567_
timestamp 1688980957
transform 1 0 20608 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1568_
timestamp 1688980957
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1569_
timestamp 1688980957
transform 1 0 12604 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1570_
timestamp 1688980957
transform 1 0 12512 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1571_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1572_
timestamp 1688980957
transform 1 0 7544 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1573_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30636 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1574_
timestamp 1688980957
transform 1 0 34408 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1575_
timestamp 1688980957
transform 1 0 33856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1576_
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1577_
timestamp 1688980957
transform 1 0 35144 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1578_
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1579_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29808 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1580_
timestamp 1688980957
transform 1 0 29900 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_2  _1581_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29900 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1582_
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1583_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29808 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1584_
timestamp 1688980957
transform 1 0 28612 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1585_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28244 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1586_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1587_
timestamp 1688980957
transform 1 0 28520 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_1  _1588_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1589_
timestamp 1688980957
transform 1 0 8280 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1590_
timestamp 1688980957
transform 1 0 8004 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1591_
timestamp 1688980957
transform 1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1592_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1593_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15088 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1594_
timestamp 1688980957
transform 1 0 31372 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1595_
timestamp 1688980957
transform 1 0 32292 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1596_
timestamp 1688980957
transform 1 0 33028 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1597_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31556 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1598_
timestamp 1688980957
transform 1 0 17848 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1599_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1600_
timestamp 1688980957
transform 1 0 28520 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1601_
timestamp 1688980957
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand4b_4  _1602_
timestamp 1688980957
transform 1 0 33396 0 -1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1603_
timestamp 1688980957
transform 1 0 29624 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1604_
timestamp 1688980957
transform 1 0 27784 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1605_
timestamp 1688980957
transform 1 0 28796 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1606_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23552 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _1607_
timestamp 1688980957
transform 1 0 19136 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1608_
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _1609_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21988 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1610_
timestamp 1688980957
transform 1 0 8924 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1611_
timestamp 1688980957
transform 1 0 24564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1612_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20884 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1613_
timestamp 1688980957
transform 1 0 26404 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1614_
timestamp 1688980957
transform 1 0 30912 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1615_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1616_
timestamp 1688980957
transform 1 0 27416 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1617_
timestamp 1688980957
transform 1 0 20240 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1618_
timestamp 1688980957
transform 1 0 19688 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_2  _1619_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25024 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_4  _1620_
timestamp 1688980957
transform 1 0 30820 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1621_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23276 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1622_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1623_
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _1624_
timestamp 1688980957
transform 1 0 17664 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1625_
timestamp 1688980957
transform 1 0 7728 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1626_
timestamp 1688980957
transform 1 0 22540 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1627_
timestamp 1688980957
transform 1 0 17480 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1628_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1629_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1630_
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1631_
timestamp 1688980957
transform 1 0 16928 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_2  _1632_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30360 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1633_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30544 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _1634_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22724 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_2  _1635_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1636_
timestamp 1688980957
transform 1 0 23000 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1637_
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1638_
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o41ai_2  _1639_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4_2  _1640_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_4  _1641_
timestamp 1688980957
transform 1 0 9936 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _1642_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _1643_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_2  _1644_
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1645_
timestamp 1688980957
transform 1 0 5704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1646_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1647_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20700 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1648_
timestamp 1688980957
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1649_
timestamp 1688980957
transform 1 0 15640 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1650_
timestamp 1688980957
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1651_
timestamp 1688980957
transform 1 0 18584 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1652_
timestamp 1688980957
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _1653_
timestamp 1688980957
transform 1 0 15364 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1654_
timestamp 1688980957
transform 1 0 17296 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1655_
timestamp 1688980957
transform 1 0 20056 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1656_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1657_
timestamp 1688980957
transform 1 0 12696 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1658_
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1659_
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1660_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1661_
timestamp 1688980957
transform 1 0 16744 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1662_
timestamp 1688980957
transform 1 0 17112 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1663_
timestamp 1688980957
transform 1 0 18584 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1664_
timestamp 1688980957
transform 1 0 10488 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1665_
timestamp 1688980957
transform 1 0 18492 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1666_
timestamp 1688980957
transform 1 0 19228 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1667_
timestamp 1688980957
transform 1 0 19688 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1668_
timestamp 1688980957
transform 1 0 19964 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1669_
timestamp 1688980957
transform 1 0 20700 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1670_
timestamp 1688980957
transform 1 0 19780 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1671_
timestamp 1688980957
transform 1 0 25116 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1672_
timestamp 1688980957
transform 1 0 30636 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1673_
timestamp 1688980957
transform 1 0 31556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1674_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1675_
timestamp 1688980957
transform 1 0 17020 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1676_
timestamp 1688980957
transform 1 0 17572 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1677_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13064 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _1678_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1679_
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1680_
timestamp 1688980957
transform 1 0 10488 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1681_
timestamp 1688980957
transform 1 0 8004 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1682_
timestamp 1688980957
transform 1 0 9844 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1683_
timestamp 1688980957
transform 1 0 9292 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1684_
timestamp 1688980957
transform 1 0 7728 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1685_
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1686_
timestamp 1688980957
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_1  _1687_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7636 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1688_
timestamp 1688980957
transform 1 0 9108 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1689_
timestamp 1688980957
transform 1 0 9844 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1690_
timestamp 1688980957
transform 1 0 7544 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1691_
timestamp 1688980957
transform 1 0 8648 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1692_
timestamp 1688980957
transform 1 0 9752 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1693_
timestamp 1688980957
transform 1 0 9200 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_2  _1694_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8004 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1695_
timestamp 1688980957
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1696_
timestamp 1688980957
transform 1 0 17020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1697_
timestamp 1688980957
transform 1 0 11684 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1698_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1699_
timestamp 1688980957
transform 1 0 6348 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1700_
timestamp 1688980957
transform 1 0 5428 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1701_
timestamp 1688980957
transform 1 0 13064 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1702_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1703_
timestamp 1688980957
transform 1 0 15272 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1704_
timestamp 1688980957
transform 1 0 14260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1705_
timestamp 1688980957
transform 1 0 11960 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1706_
timestamp 1688980957
transform 1 0 9016 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1707_
timestamp 1688980957
transform 1 0 11040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1708_
timestamp 1688980957
transform 1 0 11316 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1709_
timestamp 1688980957
transform 1 0 5612 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1710_
timestamp 1688980957
transform 1 0 5612 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1711_
timestamp 1688980957
transform 1 0 4968 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1712_
timestamp 1688980957
transform 1 0 6256 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1714_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1715_
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1716_
timestamp 1688980957
transform 1 0 15456 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1717_
timestamp 1688980957
transform 1 0 16652 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1718_
timestamp 1688980957
transform 1 0 18124 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1719_
timestamp 1688980957
transform 1 0 17940 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1720_
timestamp 1688980957
transform 1 0 10028 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1721_
timestamp 1688980957
transform 1 0 9752 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1722_
timestamp 1688980957
transform 1 0 15364 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1723_
timestamp 1688980957
transform 1 0 15272 0 1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__and4b_1  _1724_
timestamp 1688980957
transform 1 0 23920 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1725_
timestamp 1688980957
transform 1 0 25668 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1726_
timestamp 1688980957
transform 1 0 10580 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 1688980957
transform 1 0 9200 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1728_
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1729_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1730_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32476 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_2  _1731_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17572 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _1732_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1733_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1734_
timestamp 1688980957
transform 1 0 14904 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1735_
timestamp 1688980957
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 1688980957
transform 1 0 12328 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1737_
timestamp 1688980957
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1738_
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1739_
timestamp 1688980957
transform 1 0 14996 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1740_
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1741_
timestamp 1688980957
transform 1 0 15180 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1742_
timestamp 1688980957
transform 1 0 9936 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1743_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16192 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1744_
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1745_
timestamp 1688980957
transform 1 0 18124 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1746_
timestamp 1688980957
transform 1 0 17572 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1747_
timestamp 1688980957
transform 1 0 14076 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1748_
timestamp 1688980957
transform 1 0 16192 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1749_
timestamp 1688980957
transform 1 0 14996 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1750_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15548 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1751_
timestamp 1688980957
transform 1 0 8280 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1752_
timestamp 1688980957
transform 1 0 17572 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1753_
timestamp 1688980957
transform 1 0 18032 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1754_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1755_
timestamp 1688980957
transform 1 0 10948 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1756_
timestamp 1688980957
transform 1 0 17204 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1757_
timestamp 1688980957
transform 1 0 17204 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1758_
timestamp 1688980957
transform 1 0 16376 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 1688980957
transform 1 0 14260 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1760_
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1761_
timestamp 1688980957
transform 1 0 16100 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1762_
timestamp 1688980957
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1763_
timestamp 1688980957
transform 1 0 12880 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1764_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1765_
timestamp 1688980957
transform 1 0 25944 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1766_
timestamp 1688980957
transform 1 0 26128 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1767_
timestamp 1688980957
transform 1 0 23000 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1768_
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1769_
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1770_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1771_
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1772_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1773_
timestamp 1688980957
transform 1 0 27232 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1774_
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1775_
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1776_
timestamp 1688980957
transform 1 0 23092 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1777_
timestamp 1688980957
transform 1 0 23920 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1778_
timestamp 1688980957
transform 1 0 21528 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1779_
timestamp 1688980957
transform 1 0 22724 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1780_
timestamp 1688980957
transform 1 0 29992 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1781_
timestamp 1688980957
transform 1 0 31556 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1782_
timestamp 1688980957
transform 1 0 20792 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1783_
timestamp 1688980957
transform 1 0 27600 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1784_
timestamp 1688980957
transform 1 0 17848 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1785_
timestamp 1688980957
transform 1 0 17204 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1786_
timestamp 1688980957
transform 1 0 28152 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1787_
timestamp 1688980957
transform 1 0 23460 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1788_
timestamp 1688980957
transform 1 0 23000 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1789_
timestamp 1688980957
transform 1 0 29624 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1790_
timestamp 1688980957
transform 1 0 17848 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1791_
timestamp 1688980957
transform 1 0 21896 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1792_
timestamp 1688980957
transform 1 0 27876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1793_
timestamp 1688980957
transform 1 0 22080 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1794_
timestamp 1688980957
transform 1 0 22172 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1795_
timestamp 1688980957
transform 1 0 27784 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1796_
timestamp 1688980957
transform 1 0 23000 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_4  _1797_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22448 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__a31o_1  _1798_
timestamp 1688980957
transform 1 0 22540 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1799_
timestamp 1688980957
transform 1 0 22264 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_4  _1800_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30728 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _1801_
timestamp 1688980957
transform 1 0 24932 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1802_
timestamp 1688980957
transform 1 0 19964 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1803_
timestamp 1688980957
transform 1 0 20424 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1804_
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1805_
timestamp 1688980957
transform 1 0 24288 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1806_
timestamp 1688980957
transform 1 0 19320 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1807_
timestamp 1688980957
transform 1 0 26588 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1808_
timestamp 1688980957
transform 1 0 22264 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1809_
timestamp 1688980957
transform 1 0 23000 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1810_
timestamp 1688980957
transform 1 0 26772 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _1811_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _1812_
timestamp 1688980957
transform 1 0 27416 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1813_
timestamp 1688980957
transform 1 0 27600 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1814_
timestamp 1688980957
transform 1 0 27692 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1815_
timestamp 1688980957
transform 1 0 29164 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1816_
timestamp 1688980957
transform 1 0 31004 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1817_
timestamp 1688980957
transform 1 0 27784 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1818_
timestamp 1688980957
transform 1 0 13156 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1819_
timestamp 1688980957
transform 1 0 19872 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1820_
timestamp 1688980957
transform 1 0 19504 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1821_
timestamp 1688980957
transform 1 0 27416 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1822_
timestamp 1688980957
transform 1 0 27140 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1823_
timestamp 1688980957
transform 1 0 24564 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1824_
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1825_
timestamp 1688980957
transform 1 0 28060 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1826_
timestamp 1688980957
transform 1 0 28980 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1827_
timestamp 1688980957
transform 1 0 30268 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1828_
timestamp 1688980957
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _1829_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21988 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1830_
timestamp 1688980957
transform 1 0 19780 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _1831_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18952 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1832_
timestamp 1688980957
transform 1 0 21436 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1833_
timestamp 1688980957
transform 1 0 20424 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1834_
timestamp 1688980957
transform 1 0 20148 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1835_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1836_
timestamp 1688980957
transform 1 0 21896 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1837_
timestamp 1688980957
transform 1 0 25944 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1838_
timestamp 1688980957
transform 1 0 29716 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _1839_
timestamp 1688980957
transform 1 0 24840 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1840_
timestamp 1688980957
transform 1 0 25392 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1841_
timestamp 1688980957
transform 1 0 28612 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1842_
timestamp 1688980957
transform 1 0 28796 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1843_
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1844_
timestamp 1688980957
transform 1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1845_
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1846_
timestamp 1688980957
transform 1 0 31188 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1847_
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1848_
timestamp 1688980957
transform 1 0 25024 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1849_
timestamp 1688980957
transform 1 0 18584 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1850_
timestamp 1688980957
transform 1 0 19964 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1851_
timestamp 1688980957
transform 1 0 19412 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1852_
timestamp 1688980957
transform 1 0 19596 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1853_
timestamp 1688980957
transform 1 0 19504 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1854_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1855_
timestamp 1688980957
transform 1 0 20240 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1856_
timestamp 1688980957
transform 1 0 26128 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1857_
timestamp 1688980957
transform 1 0 28704 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1858_
timestamp 1688980957
transform 1 0 26956 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1859_
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1860_
timestamp 1688980957
transform 1 0 25852 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1861_
timestamp 1688980957
transform 1 0 25760 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1862_
timestamp 1688980957
transform 1 0 26772 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1863_
timestamp 1688980957
transform 1 0 28428 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1864_
timestamp 1688980957
transform 1 0 31556 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1865_
timestamp 1688980957
transform 1 0 32660 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1866_
timestamp 1688980957
transform 1 0 33304 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1867_
timestamp 1688980957
transform 1 0 25852 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1868_
timestamp 1688980957
transform 1 0 24288 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1869_
timestamp 1688980957
transform 1 0 24840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1870_
timestamp 1688980957
transform 1 0 23552 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1871_
timestamp 1688980957
transform 1 0 25944 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1872_
timestamp 1688980957
transform 1 0 25760 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1873_
timestamp 1688980957
transform 1 0 25208 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1874_
timestamp 1688980957
transform 1 0 25024 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1875_
timestamp 1688980957
transform 1 0 26220 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1876_
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1877_
timestamp 1688980957
transform 1 0 26956 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1878_
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1879_
timestamp 1688980957
transform 1 0 27968 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1880_
timestamp 1688980957
transform 1 0 23092 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1881_
timestamp 1688980957
transform 1 0 29532 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1882_
timestamp 1688980957
transform 1 0 29348 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1883_
timestamp 1688980957
transform 1 0 27508 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1884_
timestamp 1688980957
transform 1 0 28428 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1885_
timestamp 1688980957
transform 1 0 27968 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1886_
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1887_
timestamp 1688980957
transform 1 0 23736 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1888_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30452 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1889_
timestamp 1688980957
transform 1 0 30268 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1890_
timestamp 1688980957
transform 1 0 22908 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1891_
timestamp 1688980957
transform 1 0 24932 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1892_
timestamp 1688980957
transform 1 0 24564 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1893_
timestamp 1688980957
transform 1 0 23184 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1894_
timestamp 1688980957
transform 1 0 29440 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1895_
timestamp 1688980957
transform 1 0 31004 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1896_
timestamp 1688980957
transform 1 0 32200 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1897_
timestamp 1688980957
transform 1 0 32844 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1898_
timestamp 1688980957
transform 1 0 22172 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1899_
timestamp 1688980957
transform 1 0 18584 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1900_
timestamp 1688980957
transform 1 0 21712 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1901_
timestamp 1688980957
transform 1 0 20976 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1902_
timestamp 1688980957
transform 1 0 22172 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1903_
timestamp 1688980957
transform 1 0 31924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1904_
timestamp 1688980957
transform 1 0 31280 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1905_
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1906_
timestamp 1688980957
transform 1 0 30912 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1907_
timestamp 1688980957
transform 1 0 26496 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1908_
timestamp 1688980957
transform 1 0 24196 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1909_
timestamp 1688980957
transform 1 0 25208 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1910_
timestamp 1688980957
transform 1 0 30360 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1911_
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1912_
timestamp 1688980957
transform 1 0 25392 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1913_
timestamp 1688980957
transform 1 0 19688 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1914_
timestamp 1688980957
transform 1 0 28612 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1915_
timestamp 1688980957
transform 1 0 30912 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1916_
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1917_
timestamp 1688980957
transform 1 0 32016 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1918_
timestamp 1688980957
transform 1 0 33212 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1919_
timestamp 1688980957
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1920_
timestamp 1688980957
transform 1 0 26864 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1921_
timestamp 1688980957
transform 1 0 27140 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1922_
timestamp 1688980957
transform 1 0 27048 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1923_
timestamp 1688980957
transform 1 0 23552 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1924_
timestamp 1688980957
transform 1 0 23552 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1925_
timestamp 1688980957
transform 1 0 28612 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1926_
timestamp 1688980957
transform 1 0 31464 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1927_
timestamp 1688980957
transform 1 0 22264 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _1928_
timestamp 1688980957
transform 1 0 22356 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1929_
timestamp 1688980957
transform 1 0 30360 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1930_
timestamp 1688980957
transform 1 0 30820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1931_
timestamp 1688980957
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1932_
timestamp 1688980957
transform 1 0 32200 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1933_
timestamp 1688980957
transform 1 0 33396 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1934_
timestamp 1688980957
transform 1 0 28796 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1935_
timestamp 1688980957
transform 1 0 29256 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1936_
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1937_
timestamp 1688980957
transform 1 0 31004 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1938_
timestamp 1688980957
transform 1 0 29072 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1939_
timestamp 1688980957
transform 1 0 28612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1940_
timestamp 1688980957
transform 1 0 25208 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1941_
timestamp 1688980957
transform 1 0 25852 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1942_
timestamp 1688980957
transform 1 0 25852 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1943_
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1944_
timestamp 1688980957
transform 1 0 31188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1945_
timestamp 1688980957
transform 1 0 32292 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1946_
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1947_
timestamp 1688980957
transform 1 0 30176 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1948_
timestamp 1688980957
transform 1 0 26312 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1949_
timestamp 1688980957
transform 1 0 15364 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1950_
timestamp 1688980957
transform 1 0 20884 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1951_
timestamp 1688980957
transform 1 0 23644 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1952_
timestamp 1688980957
transform 1 0 26956 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1953_
timestamp 1688980957
transform 1 0 27876 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1954_
timestamp 1688980957
transform 1 0 28060 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1955_
timestamp 1688980957
transform 1 0 32108 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1956_
timestamp 1688980957
transform 1 0 33028 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1957_
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1958_
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1959_
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1960_
timestamp 1688980957
transform 1 0 40296 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1961_
timestamp 1688980957
transform 1 0 19780 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1962_
timestamp 1688980957
transform 1 0 2116 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1963_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1840 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _1964_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25852 0 1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__a311oi_2  _1965_
timestamp 1688980957
transform 1 0 24932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__a311oi_2  _1966_
timestamp 1688980957
transform 1 0 24932 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1967_
timestamp 1688980957
transform 1 0 11776 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1968_
timestamp 1688980957
transform 1 0 12604 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1969_
timestamp 1688980957
transform 1 0 20056 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1970_
timestamp 1688980957
transform 1 0 16652 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1971_
timestamp 1688980957
transform 1 0 17480 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1972_
timestamp 1688980957
transform 1 0 17204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1973_
timestamp 1688980957
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_1  _1974_
timestamp 1688980957
transform 1 0 18032 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1975_
timestamp 1688980957
transform 1 0 24288 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1976_
timestamp 1688980957
transform 1 0 20976 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1977_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1978_
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1979_
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1980_
timestamp 1688980957
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1981_
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1982_
timestamp 1688980957
transform 1 0 11316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1983_
timestamp 1688980957
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  _1984_
timestamp 1688980957
transform 1 0 20424 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__a22o_1  _1985_
timestamp 1688980957
transform 1 0 20976 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _1986_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23552 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1987_
timestamp 1688980957
transform 1 0 15732 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1988_
timestamp 1688980957
transform 1 0 21252 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1989_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _1990_
timestamp 1688980957
transform 1 0 11868 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1991_
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1992_
timestamp 1688980957
transform 1 0 22080 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1993_
timestamp 1688980957
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _1994_
timestamp 1688980957
transform 1 0 12696 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1995_
timestamp 1688980957
transform 1 0 21252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1996_
timestamp 1688980957
transform 1 0 22356 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1997_
timestamp 1688980957
transform 1 0 22356 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1998_
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__o31a_1  _1999_
timestamp 1688980957
transform 1 0 23460 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _2000_
timestamp 1688980957
transform 1 0 21988 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_4  _2001_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__and4b_1  _2002_
timestamp 1688980957
transform 1 0 31280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2003_
timestamp 1688980957
transform 1 0 22632 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2004_
timestamp 1688980957
transform 1 0 22448 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _2005_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21896 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2006_
timestamp 1688980957
transform 1 0 18676 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_4  _2007_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_2  _2008_
timestamp 1688980957
transform 1 0 19136 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2009_
timestamp 1688980957
transform 1 0 10304 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2010_
timestamp 1688980957
transform 1 0 10580 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2011_
timestamp 1688980957
transform 1 0 9200 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _2012_
timestamp 1688980957
transform 1 0 8648 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2013_
timestamp 1688980957
transform 1 0 9292 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2014_
timestamp 1688980957
transform 1 0 9476 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2015_
timestamp 1688980957
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _2016_
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _2017_
timestamp 1688980957
transform 1 0 15364 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _2018_
timestamp 1688980957
transform 1 0 20976 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2019_
timestamp 1688980957
transform 1 0 20148 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2020_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2021_
timestamp 1688980957
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2022_
timestamp 1688980957
transform 1 0 7912 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2023_
timestamp 1688980957
transform 1 0 10488 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2024_
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2025_
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2026_
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2027_
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _2028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19044 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _2029_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21528 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  _2030_
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _2031_
timestamp 1688980957
transform 1 0 20976 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2032_
timestamp 1688980957
transform 1 0 17020 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2033_
timestamp 1688980957
transform 1 0 17112 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2034_
timestamp 1688980957
transform 1 0 17756 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2035_
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2036_
timestamp 1688980957
transform 1 0 20240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2037_
timestamp 1688980957
transform 1 0 17296 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2038_
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _2039_
timestamp 1688980957
transform 1 0 23460 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2040_
timestamp 1688980957
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _2041_
timestamp 1688980957
transform 1 0 24196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_4  _2042_
timestamp 1688980957
transform 1 0 22264 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__and3_2  _2043_
timestamp 1688980957
transform 1 0 22448 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2044_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _2045_
timestamp 1688980957
transform 1 0 25116 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2046_
timestamp 1688980957
transform 1 0 23828 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2047_
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2048_
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2049_
timestamp 1688980957
transform 1 0 23368 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2050_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2051_
timestamp 1688980957
transform 1 0 17664 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _2052_
timestamp 1688980957
transform 1 0 17664 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _2053_
timestamp 1688980957
transform 1 0 19504 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__a31o_1  _2054_
timestamp 1688980957
transform 1 0 19412 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2055_
timestamp 1688980957
transform 1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2056_
timestamp 1688980957
transform 1 0 20148 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _2057_
timestamp 1688980957
transform 1 0 13248 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _2058_
timestamp 1688980957
transform 1 0 8924 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _2059_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2060_
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2061_
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_1  _2062_
timestamp 1688980957
transform 1 0 16192 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2063_
timestamp 1688980957
transform 1 0 23000 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2064_
timestamp 1688980957
transform 1 0 23736 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _2065_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _2066_
timestamp 1688980957
transform 1 0 24656 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _2067_
timestamp 1688980957
transform 1 0 23460 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _2068_
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _2069_
timestamp 1688980957
transform 1 0 17112 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2070_
timestamp 1688980957
transform 1 0 20976 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2071_
timestamp 1688980957
transform 1 0 12788 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2072_
timestamp 1688980957
transform 1 0 15088 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _2073_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2074_
timestamp 1688980957
transform 1 0 10396 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2075_
timestamp 1688980957
transform 1 0 11684 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _2076_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_4  _2077_
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_1  _2078_
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2079_
timestamp 1688980957
transform 1 0 15364 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2080_
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2081_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21988 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _2082_
timestamp 1688980957
transform 1 0 20884 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2083_
timestamp 1688980957
transform 1 0 18032 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2084_
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2085_
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _2086_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2087_
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2088_
timestamp 1688980957
transform 1 0 18492 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _2089_
timestamp 1688980957
transform 1 0 19320 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2090_
timestamp 1688980957
transform 1 0 19136 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2091_
timestamp 1688980957
transform 1 0 11040 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2092_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _2093_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2094_
timestamp 1688980957
transform 1 0 17940 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2095_
timestamp 1688980957
transform 1 0 17112 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2096_
timestamp 1688980957
transform 1 0 16376 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2097_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2098_
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _2099_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__and3b_2  _2100_
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _2101_
timestamp 1688980957
transform 1 0 18124 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _2102_
timestamp 1688980957
transform 1 0 19596 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2103_
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _2104_
timestamp 1688980957
transform 1 0 16468 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _2105_
timestamp 1688980957
transform 1 0 16928 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2106_
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2107_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2108_
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2109_
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2110_
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2111_
timestamp 1688980957
transform 1 0 12972 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2112_
timestamp 1688980957
transform 1 0 16652 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _2113_
timestamp 1688980957
transform 1 0 17020 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _2114_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _2115_
timestamp 1688980957
transform 1 0 19780 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2116_
timestamp 1688980957
transform 1 0 16652 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2117_
timestamp 1688980957
transform 1 0 22724 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2118_
timestamp 1688980957
transform 1 0 16468 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2119_
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2120_
timestamp 1688980957
transform 1 0 20792 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2121_
timestamp 1688980957
transform 1 0 20056 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2122_
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2123_
timestamp 1688980957
transform 1 0 18952 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2124_
timestamp 1688980957
transform 1 0 18032 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2125_
timestamp 1688980957
transform 1 0 18216 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2126_
timestamp 1688980957
transform 1 0 18308 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2127_
timestamp 1688980957
transform 1 0 12788 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2128_
timestamp 1688980957
transform 1 0 16100 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _2129_
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2130_
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2131_
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o41ai_2  _2132_
timestamp 1688980957
transform 1 0 20424 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _2133_
timestamp 1688980957
transform 1 0 16008 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2134_
timestamp 1688980957
transform 1 0 15640 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2135_
timestamp 1688980957
transform 1 0 17112 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2136_
timestamp 1688980957
transform 1 0 15548 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _2137_
timestamp 1688980957
transform 1 0 16008 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2138_
timestamp 1688980957
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2139_
timestamp 1688980957
transform 1 0 14076 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _2140_
timestamp 1688980957
transform 1 0 7728 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2141_
timestamp 1688980957
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2142_
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2143_
timestamp 1688980957
transform 1 0 11316 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2144_
timestamp 1688980957
transform 1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_2  _2145_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2146_
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _2147_
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2148_
timestamp 1688980957
transform 1 0 11960 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_4  _2149_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__a31o_1  _2150_
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2151_
timestamp 1688980957
transform 1 0 20424 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2152_
timestamp 1688980957
transform 1 0 18308 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2153_
timestamp 1688980957
transform 1 0 16836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _2154_
timestamp 1688980957
transform 1 0 15732 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2155_
timestamp 1688980957
transform 1 0 17112 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2156_
timestamp 1688980957
transform 1 0 18584 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2157_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2158_
timestamp 1688980957
transform 1 0 22172 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2159_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23920 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _2160_
timestamp 1688980957
transform 1 0 23092 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _2161_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2162_
timestamp 1688980957
transform 1 0 9476 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2163_
timestamp 1688980957
transform 1 0 9292 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2164_
timestamp 1688980957
transform 1 0 7820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _2165_
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2166_
timestamp 1688980957
transform 1 0 11684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2167_
timestamp 1688980957
transform 1 0 12788 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _2168_
timestamp 1688980957
transform 1 0 14076 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2169_
timestamp 1688980957
transform 1 0 13432 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2170_
timestamp 1688980957
transform 1 0 12328 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2171_
timestamp 1688980957
transform 1 0 16560 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2172_
timestamp 1688980957
transform 1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2173_
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2174_
timestamp 1688980957
transform 1 0 8832 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2175_
timestamp 1688980957
transform 1 0 9108 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2176_
timestamp 1688980957
transform 1 0 8740 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2177_
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2178_
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2179_
timestamp 1688980957
transform 1 0 20516 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2180_
timestamp 1688980957
transform 1 0 18676 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2181_
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2182_
timestamp 1688980957
transform 1 0 24196 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2183_
timestamp 1688980957
transform 1 0 18400 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2184_
timestamp 1688980957
transform 1 0 18216 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2185_
timestamp 1688980957
transform 1 0 18124 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _2186_
timestamp 1688980957
transform 1 0 10396 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2187_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2188_
timestamp 1688980957
transform 1 0 9200 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2189_
timestamp 1688980957
transform 1 0 13248 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2190_
timestamp 1688980957
transform 1 0 12696 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2191_
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2192_
timestamp 1688980957
transform 1 0 12328 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2193_
timestamp 1688980957
transform 1 0 12512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2194_
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2195_
timestamp 1688980957
transform 1 0 13616 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2196_
timestamp 1688980957
transform 1 0 15732 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2197_
timestamp 1688980957
transform 1 0 14904 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _2198_
timestamp 1688980957
transform 1 0 22724 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _2199_
timestamp 1688980957
transform 1 0 21988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2200_
timestamp 1688980957
transform 1 0 15916 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2201_
timestamp 1688980957
transform 1 0 23644 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2202_
timestamp 1688980957
transform 1 0 15272 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2203_
timestamp 1688980957
transform 1 0 17020 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2204_
timestamp 1688980957
transform 1 0 9752 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _2205_
timestamp 1688980957
transform 1 0 10488 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_2  _2206_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2207_
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2208_
timestamp 1688980957
transform 1 0 23184 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2209_
timestamp 1688980957
transform 1 0 23000 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2210_
timestamp 1688980957
transform 1 0 12512 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_2  _2211_
timestamp 1688980957
transform 1 0 12052 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a311o_1  _2212_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14996 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2213_
timestamp 1688980957
transform 1 0 14996 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2214_
timestamp 1688980957
transform 1 0 14904 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_2  _2215_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_2  _2216_
timestamp 1688980957
transform 1 0 14720 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2217_
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2218_
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2219_
timestamp 1688980957
transform 1 0 12236 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2220_
timestamp 1688980957
transform 1 0 12420 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2221_
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2222_
timestamp 1688980957
transform 1 0 10396 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2223_
timestamp 1688980957
transform 1 0 9660 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2224_
timestamp 1688980957
transform 1 0 9016 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o32ai_4  _2225_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__o211ai_1  _2226_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2227_
timestamp 1688980957
transform 1 0 12328 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2228_
timestamp 1688980957
transform 1 0 14076 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2229_
timestamp 1688980957
transform 1 0 14720 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2230_
timestamp 1688980957
transform 1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _2231_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_2  _2232_
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2233_
timestamp 1688980957
transform 1 0 14720 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_4  _2234_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__nand2b_2  _2235_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2236_
timestamp 1688980957
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _2237_
timestamp 1688980957
transform 1 0 15272 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2238_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _2239_
timestamp 1688980957
transform 1 0 14260 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _2240_
timestamp 1688980957
transform 1 0 18124 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _2241_
timestamp 1688980957
transform 1 0 17572 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _2242_
timestamp 1688980957
transform 1 0 17940 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2243_
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2244_
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2245_
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2246_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2247_
timestamp 1688980957
transform 1 0 9292 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2248_
timestamp 1688980957
transform 1 0 8096 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2249_
timestamp 1688980957
transform 1 0 25668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2250_
timestamp 1688980957
transform 1 0 15272 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2251_
timestamp 1688980957
transform 1 0 16376 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2252_
timestamp 1688980957
transform 1 0 25024 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2253_
timestamp 1688980957
transform 1 0 25024 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2254_
timestamp 1688980957
transform 1 0 25760 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2255_
timestamp 1688980957
transform 1 0 27324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2256_
timestamp 1688980957
transform 1 0 25944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2257_
timestamp 1688980957
transform 1 0 26680 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _2258_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26036 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2259_
timestamp 1688980957
transform 1 0 10672 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2260_
timestamp 1688980957
transform 1 0 21804 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2261_
timestamp 1688980957
transform 1 0 24840 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2262_
timestamp 1688980957
transform 1 0 12052 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2263_
timestamp 1688980957
transform 1 0 15180 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2264_
timestamp 1688980957
transform 1 0 18124 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _2265_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2266_
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2267_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2268_
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2269_
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2270_
timestamp 1688980957
transform 1 0 8096 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2271_
timestamp 1688980957
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2272_
timestamp 1688980957
transform 1 0 16652 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2273_
timestamp 1688980957
transform 1 0 17572 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2274_
timestamp 1688980957
transform 1 0 20884 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2275_
timestamp 1688980957
transform 1 0 20884 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2276_
timestamp 1688980957
transform 1 0 20424 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2277_
timestamp 1688980957
transform 1 0 28060 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2278_
timestamp 1688980957
transform 1 0 27140 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2279_
timestamp 1688980957
transform 1 0 27784 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2280_
timestamp 1688980957
transform 1 0 22724 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2281_
timestamp 1688980957
transform 1 0 22080 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _2282_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2283_
timestamp 1688980957
transform 1 0 10396 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _2284_
timestamp 1688980957
transform 1 0 20700 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2285_
timestamp 1688980957
transform 1 0 12880 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2286_
timestamp 1688980957
transform 1 0 16928 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2287_
timestamp 1688980957
transform 1 0 17480 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _2288_
timestamp 1688980957
transform 1 0 17020 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _2289_
timestamp 1688980957
transform 1 0 17940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2290_
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2291_
timestamp 1688980957
transform 1 0 9476 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2292_
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _2293_
timestamp 1688980957
transform 1 0 7268 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2294_
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2295_
timestamp 1688980957
transform 1 0 27876 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2296_
timestamp 1688980957
transform 1 0 26312 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2297_
timestamp 1688980957
transform 1 0 27048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2298_
timestamp 1688980957
transform 1 0 27416 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2299_
timestamp 1688980957
transform 1 0 20700 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2300_
timestamp 1688980957
transform 1 0 25760 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2301_
timestamp 1688980957
transform 1 0 15548 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2302_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _2303_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2304_
timestamp 1688980957
transform 1 0 24748 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _2305_
timestamp 1688980957
transform 1 0 23552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _2306_
timestamp 1688980957
transform 1 0 23184 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2307_
timestamp 1688980957
transform 1 0 10212 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _2308_
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2309_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2310_
timestamp 1688980957
transform 1 0 14628 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2311_
timestamp 1688980957
transform 1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _2312_
timestamp 1688980957
transform 1 0 14996 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2313_
timestamp 1688980957
transform 1 0 11960 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2314_
timestamp 1688980957
transform 1 0 9108 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2315_
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2316_
timestamp 1688980957
transform 1 0 7728 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2317_
timestamp 1688980957
transform 1 0 27600 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2318_
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2319_
timestamp 1688980957
transform 1 0 26956 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2320_
timestamp 1688980957
transform 1 0 26404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2321_
timestamp 1688980957
transform 1 0 24196 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2322_
timestamp 1688980957
transform 1 0 24932 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2323_
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2324_
timestamp 1688980957
transform 1 0 25024 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2325_
timestamp 1688980957
transform 1 0 25576 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2326_
timestamp 1688980957
transform 1 0 25668 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _2327_
timestamp 1688980957
transform 1 0 25208 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _2328_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _2329_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24932 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2330_
timestamp 1688980957
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _2331_
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2332_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _2333_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17572 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_2  _2334_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _2335_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _2336_
timestamp 1688980957
transform 1 0 19412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2337_
timestamp 1688980957
transform 1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2338_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2339_
timestamp 1688980957
transform 1 0 18768 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _2340_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2341_
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2342_
timestamp 1688980957
transform 1 0 16192 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2343_
timestamp 1688980957
transform 1 0 19320 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2344_
timestamp 1688980957
transform 1 0 22356 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2345_
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _2346_
timestamp 1688980957
transform 1 0 22264 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2347_
timestamp 1688980957
transform 1 0 19964 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _2348_
timestamp 1688980957
transform 1 0 20240 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2349_
timestamp 1688980957
transform 1 0 12512 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _2350_
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2351_
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2352_
timestamp 1688980957
transform 1 0 18216 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _2353_
timestamp 1688980957
transform 1 0 18216 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2354_
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2355_
timestamp 1688980957
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2356_
timestamp 1688980957
transform 1 0 19688 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _2357_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2358_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2359_
timestamp 1688980957
transform 1 0 23092 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _2360_
timestamp 1688980957
transform 1 0 20240 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o32ai_4  _2361_
timestamp 1688980957
transform 1 0 19688 0 -1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _2362_
timestamp 1688980957
transform 1 0 11960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2363_
timestamp 1688980957
transform 1 0 11868 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2364_
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2365_
timestamp 1688980957
transform 1 0 8464 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2366_
timestamp 1688980957
transform 1 0 11960 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2367_
timestamp 1688980957
transform 1 0 12972 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2368_
timestamp 1688980957
transform 1 0 25300 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2369_
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2370_
timestamp 1688980957
transform 1 0 11592 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2371_
timestamp 1688980957
transform 1 0 10028 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2372_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2373_
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _2374_
timestamp 1688980957
transform 1 0 9384 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2375_
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2376_
timestamp 1688980957
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _2377_
timestamp 1688980957
transform 1 0 23368 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2378_
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2379_
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2380_
timestamp 1688980957
transform 1 0 20976 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2381_
timestamp 1688980957
transform 1 0 15548 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o41ai_2  _2382_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _2383_
timestamp 1688980957
transform 1 0 23460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2384_
timestamp 1688980957
transform 1 0 23092 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2385_
timestamp 1688980957
transform 1 0 22632 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _2386_
timestamp 1688980957
transform 1 0 21896 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _2387_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2388_
timestamp 1688980957
transform 1 0 21896 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2389_
timestamp 1688980957
transform 1 0 12972 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2390_
timestamp 1688980957
transform 1 0 15180 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _2391_
timestamp 1688980957
transform 1 0 17480 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2392_
timestamp 1688980957
transform 1 0 16008 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _2393_
timestamp 1688980957
transform 1 0 15272 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _2394_
timestamp 1688980957
transform 1 0 11960 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _2395_
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _2396_
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _2397_
timestamp 1688980957
transform 1 0 10212 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2398_
timestamp 1688980957
transform 1 0 9200 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2399_
timestamp 1688980957
transform 1 0 7544 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2400_
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2401_
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2402_
timestamp 1688980957
transform 1 0 6256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2403_
timestamp 1688980957
transform 1 0 6532 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2404_
timestamp 1688980957
transform 1 0 6716 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2405_
timestamp 1688980957
transform 1 0 25668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2406_
timestamp 1688980957
transform 1 0 14904 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2407_
timestamp 1688980957
transform 1 0 24932 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2408_
timestamp 1688980957
transform 1 0 24840 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2409_
timestamp 1688980957
transform 1 0 26404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2410_
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2411_
timestamp 1688980957
transform 1 0 24748 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2412_
timestamp 1688980957
transform 1 0 25116 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2413_
timestamp 1688980957
transform 1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2414_
timestamp 1688980957
transform 1 0 27692 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2415_
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2416_
timestamp 1688980957
transform 1 0 26680 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _2417_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _2418_
timestamp 1688980957
transform 1 0 9292 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2419_
timestamp 1688980957
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2420_
timestamp 1688980957
transform 1 0 25944 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2421_
timestamp 1688980957
transform 1 0 12788 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2422_
timestamp 1688980957
transform 1 0 14536 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2423_
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _2424_
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2425_
timestamp 1688980957
transform 1 0 12512 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2426_
timestamp 1688980957
transform 1 0 11960 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _2427_
timestamp 1688980957
transform 1 0 9384 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2428_
timestamp 1688980957
transform 1 0 6532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2429_
timestamp 1688980957
transform 1 0 9844 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2430_
timestamp 1688980957
transform 1 0 7452 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _2431_
timestamp 1688980957
transform 1 0 20792 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2432_
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2433_
timestamp 1688980957
transform 1 0 6992 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2434_
timestamp 1688980957
transform 1 0 7176 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _2435_
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2436_
timestamp 1688980957
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2437_
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _2438_
timestamp 1688980957
transform 1 0 27232 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2439_
timestamp 1688980957
transform 1 0 27048 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2440_
timestamp 1688980957
transform 1 0 26864 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2441_
timestamp 1688980957
transform 1 0 27692 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2442_
timestamp 1688980957
transform 1 0 26036 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2443_
timestamp 1688980957
transform 1 0 6348 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _2444_
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2445_
timestamp 1688980957
transform 1 0 11684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2446_
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2447_
timestamp 1688980957
transform 1 0 28336 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2448_
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2449_
timestamp 1688980957
transform 1 0 27968 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2450_
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2451_
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2452_
timestamp 1688980957
transform 1 0 28888 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2453_
timestamp 1688980957
transform 1 0 28520 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2454_
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2455_
timestamp 1688980957
transform 1 0 30268 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2456_
timestamp 1688980957
transform 1 0 28336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2457_
timestamp 1688980957
transform 1 0 28428 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2458_
timestamp 1688980957
transform 1 0 29256 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2459_
timestamp 1688980957
transform 1 0 20700 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2460_
timestamp 1688980957
transform 1 0 24840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2461_
timestamp 1688980957
transform 1 0 25576 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2462_
timestamp 1688980957
transform 1 0 24932 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2463_
timestamp 1688980957
transform 1 0 24932 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _2464_
timestamp 1688980957
transform 1 0 25392 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2465_
timestamp 1688980957
transform 1 0 27048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2466_
timestamp 1688980957
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _2467_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2468_
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2469_
timestamp 1688980957
transform 1 0 20056 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2470_
timestamp 1688980957
transform 1 0 14076 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2471_
timestamp 1688980957
transform 1 0 17756 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2472_
timestamp 1688980957
transform 1 0 15272 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2473_
timestamp 1688980957
transform 1 0 16100 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2474_
timestamp 1688980957
transform 1 0 15548 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _2475_
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2476_
timestamp 1688980957
transform 1 0 12788 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _2477_
timestamp 1688980957
transform 1 0 12788 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _2478_
timestamp 1688980957
transform 1 0 6808 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2479_
timestamp 1688980957
transform 1 0 23000 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_4  _2480_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20976 0 1 29376
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_1  _2481_
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2482_
timestamp 1688980957
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_4  _2483_
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_4  _2484_
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__o22ai_2  _2485_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _2486_
timestamp 1688980957
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2487_
timestamp 1688980957
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _2488_
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2489_
timestamp 1688980957
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2490_
timestamp 1688980957
transform 1 0 5428 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _2491_
timestamp 1688980957
transform 1 0 5152 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _2492_
timestamp 1688980957
transform 1 0 4600 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2493_
timestamp 1688980957
transform 1 0 8464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2494_
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2495_
timestamp 1688980957
transform 1 0 5336 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _2496_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2497_
timestamp 1688980957
transform 1 0 5428 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2498_
timestamp 1688980957
transform 1 0 7452 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _2499_
timestamp 1688980957
transform 1 0 6256 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2500_
timestamp 1688980957
transform 1 0 6440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _2501_
timestamp 1688980957
transform 1 0 6716 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _2502_
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2503_
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 1688980957
transform 1 0 28060 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2505_
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2506_
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2507_
timestamp 1688980957
transform 1 0 27232 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2508_
timestamp 1688980957
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _2509_
timestamp 1688980957
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2510_
timestamp 1688980957
transform 1 0 15456 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2511_
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2512_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2513_
timestamp 1688980957
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2514_
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2515_
timestamp 1688980957
transform 1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2516_
timestamp 1688980957
transform 1 0 15456 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2517_
timestamp 1688980957
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2518_
timestamp 1688980957
transform 1 0 17296 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2519_
timestamp 1688980957
transform 1 0 17020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2520_
timestamp 1688980957
transform 1 0 15456 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2521_
timestamp 1688980957
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2522_
timestamp 1688980957
transform 1 0 17940 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2523_
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2524_
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2525_
timestamp 1688980957
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2526_
timestamp 1688980957
transform 1 0 20056 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2527_
timestamp 1688980957
transform 1 0 15456 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_2  _2528_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13156 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _2529_
timestamp 1688980957
transform 1 0 10396 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2530_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2531_
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2532_
timestamp 1688980957
transform 1 0 10488 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2533_
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2534_
timestamp 1688980957
transform 1 0 10948 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2535_
timestamp 1688980957
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2536_
timestamp 1688980957
transform 1 0 10488 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _2537_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2538_
timestamp 1688980957
transform 1 0 10948 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2539_
timestamp 1688980957
transform 1 0 10672 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2540_
timestamp 1688980957
transform 1 0 11224 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2541_
timestamp 1688980957
transform 1 0 11684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2542_
timestamp 1688980957
transform 1 0 10948 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2543_
timestamp 1688980957
transform 1 0 10488 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2544_
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2545_
timestamp 1688980957
transform 1 0 6532 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2546_
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2547_
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2548_
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2549_
timestamp 1688980957
transform 1 0 8740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2550_
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _2551_
timestamp 1688980957
transform 1 0 8004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2552_
timestamp 1688980957
transform 1 0 4876 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2553_
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2554_
timestamp 1688980957
transform 1 0 3864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2555_
timestamp 1688980957
transform 1 0 4600 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2556_
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2557_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2558_
timestamp 1688980957
transform 1 0 5704 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2559_
timestamp 1688980957
transform 1 0 5520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2560_
timestamp 1688980957
transform 1 0 4416 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2561_
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2562_
timestamp 1688980957
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2563_
timestamp 1688980957
transform 1 0 6072 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2564_
timestamp 1688980957
transform 1 0 6256 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2565_
timestamp 1688980957
transform 1 0 10304 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2566_
timestamp 1688980957
transform 1 0 9016 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2567_
timestamp 1688980957
transform 1 0 8188 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2568_
timestamp 1688980957
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2569_
timestamp 1688980957
transform 1 0 8004 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2570_
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2571_
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2572_
timestamp 1688980957
transform 1 0 6348 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2573_
timestamp 1688980957
transform 1 0 10212 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2574_
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2575_
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2576_
timestamp 1688980957
transform 1 0 7912 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2577_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _2578_
timestamp 1688980957
transform 1 0 5612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _2579_
timestamp 1688980957
transform 1 0 4508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a41oi_4  _2580_
timestamp 1688980957
transform 1 0 4140 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__a31o_1  _2581_
timestamp 1688980957
transform 1 0 4416 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2582_
timestamp 1688980957
transform 1 0 7268 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2583_
timestamp 1688980957
transform 1 0 7268 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2584_
timestamp 1688980957
transform 1 0 8648 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2585_
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2586_
timestamp 1688980957
transform 1 0 6532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _2587_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2588_
timestamp 1688980957
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2589_
timestamp 1688980957
transform 1 0 7544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2590_
timestamp 1688980957
transform 1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2591_
timestamp 1688980957
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2592_
timestamp 1688980957
transform 1 0 8648 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2593_
timestamp 1688980957
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _2594_
timestamp 1688980957
transform 1 0 7636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2595_
timestamp 1688980957
transform 1 0 6716 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _2596_
timestamp 1688980957
transform 1 0 4416 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2597_
timestamp 1688980957
transform 1 0 4968 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2598_
timestamp 1688980957
transform 1 0 5336 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _2599_
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _2600_
timestamp 1688980957
transform 1 0 5244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2601_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2602_
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2603_
timestamp 1688980957
transform 1 0 4232 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2604_
timestamp 1688980957
transform 1 0 4692 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2605_
timestamp 1688980957
transform 1 0 5060 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2606_
timestamp 1688980957
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2607_
timestamp 1688980957
transform 1 0 4692 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2608_
timestamp 1688980957
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2609_
timestamp 1688980957
transform 1 0 6900 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2610_
timestamp 1688980957
transform 1 0 9568 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2611_
timestamp 1688980957
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2612_
timestamp 1688980957
transform 1 0 7912 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2613_
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2614_
timestamp 1688980957
transform 1 0 3864 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _2615_
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2616_
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2617_
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2618_
timestamp 1688980957
transform 1 0 18216 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2619_
timestamp 1688980957
transform 1 0 15272 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2620_
timestamp 1688980957
transform 1 0 15824 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2621_
timestamp 1688980957
transform 1 0 15640 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2622_
timestamp 1688980957
transform 1 0 17480 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2623_
timestamp 1688980957
transform 1 0 14260 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2624_
timestamp 1688980957
transform 1 0 13432 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2625_
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2626_
timestamp 1688980957
transform 1 0 13984 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2627_
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2628_
timestamp 1688980957
transform 1 0 13248 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2629_
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _2630_
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2631_
timestamp 1688980957
transform 1 0 9384 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2632_
timestamp 1688980957
transform 1 0 9108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _2633_
timestamp 1688980957
transform 1 0 9384 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2634_
timestamp 1688980957
transform 1 0 9660 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _2635_
timestamp 1688980957
transform 1 0 10488 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2636_
timestamp 1688980957
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2637_
timestamp 1688980957
transform 1 0 2668 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2638_
timestamp 1688980957
transform 1 0 10948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2639_
timestamp 1688980957
transform 1 0 2392 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2640_
timestamp 1688980957
transform 1 0 29716 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2641_
timestamp 1688980957
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2642_
timestamp 1688980957
transform 1 0 35972 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2643_
timestamp 1688980957
transform 1 0 35512 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2644_
timestamp 1688980957
transform 1 0 5704 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2645_
timestamp 1688980957
transform 1 0 5060 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2646_
timestamp 1688980957
transform 1 0 8924 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2647_
timestamp 1688980957
transform 1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2648_
timestamp 1688980957
transform 1 0 36156 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2649_
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2650_
timestamp 1688980957
transform 1 0 26220 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2651_
timestamp 1688980957
transform 1 0 25944 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_4  _2652_
timestamp 1688980957
transform 1 0 25576 0 -1 26112
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2653_
timestamp 1688980957
transform 1 0 20516 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2654_
timestamp 1688980957
transform 1 0 21344 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2655_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2656_
timestamp 1688980957
transform 1 0 22172 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2657_
timestamp 1688980957
transform 1 0 24748 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2658_
timestamp 1688980957
transform 1 0 24748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2659_
timestamp 1688980957
transform 1 0 26220 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2660_
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2661_
timestamp 1688980957
transform 1 0 20884 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2662_
timestamp 1688980957
transform 1 0 20148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2663_
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2664_
timestamp 1688980957
transform 1 0 27784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2665_
timestamp 1688980957
transform 1 0 22264 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2666_
timestamp 1688980957
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2667_
timestamp 1688980957
transform 1 0 25576 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2668_
timestamp 1688980957
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2669_
timestamp 1688980957
transform 1 0 30084 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _2670_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31188 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_2  _2671_
timestamp 1688980957
transform 1 0 29992 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2672_
timestamp 1688980957
transform 1 0 14260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2673_
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2674_
timestamp 1688980957
transform 1 0 15456 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2675_
timestamp 1688980957
transform 1 0 13248 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2676_
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2677_
timestamp 1688980957
transform 1 0 14720 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2678_
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2679_
timestamp 1688980957
transform 1 0 12696 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2680_
timestamp 1688980957
transform 1 0 9292 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _2681_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8832 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _2682_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2683_
timestamp 1688980957
transform 1 0 30636 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2684_
timestamp 1688980957
transform 1 0 31464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2685_
timestamp 1688980957
transform 1 0 33764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2686_
timestamp 1688980957
transform 1 0 35880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2687_
timestamp 1688980957
transform 1 0 30360 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2688_
timestamp 1688980957
transform 1 0 12236 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2689_
timestamp 1688980957
transform 1 0 12420 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2690_
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_4  _2691_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16560 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _2692_
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2693_
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2694_
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2695_
timestamp 1688980957
transform 1 0 29348 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _2696_
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2697_
timestamp 1688980957
transform 1 0 31372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2698_
timestamp 1688980957
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2699_
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2700_
timestamp 1688980957
transform 1 0 30912 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2701_
timestamp 1688980957
transform 1 0 30728 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2702_
timestamp 1688980957
transform 1 0 31832 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2703_
timestamp 1688980957
transform 1 0 31188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _2704_
timestamp 1688980957
transform 1 0 33580 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2705_
timestamp 1688980957
transform 1 0 38272 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2706_
timestamp 1688980957
transform 1 0 37720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2707_
timestamp 1688980957
transform 1 0 36432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2708_
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2709_
timestamp 1688980957
transform 1 0 31004 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2710_
timestamp 1688980957
transform 1 0 31096 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2711_
timestamp 1688980957
transform 1 0 28336 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2712_
timestamp 1688980957
transform 1 0 28796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2713_
timestamp 1688980957
transform 1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2714_
timestamp 1688980957
transform 1 0 30452 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2715_
timestamp 1688980957
transform 1 0 31464 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2716_
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2717_
timestamp 1688980957
transform 1 0 29348 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2718_
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2719_
timestamp 1688980957
transform 1 0 30544 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _2720_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31004 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2721_
timestamp 1688980957
transform 1 0 32108 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2722_
timestamp 1688980957
transform 1 0 31648 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2723_
timestamp 1688980957
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2724_
timestamp 1688980957
transform 1 0 29532 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2725_
timestamp 1688980957
transform 1 0 29532 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2726_
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2727_
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2728_
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2729_
timestamp 1688980957
transform 1 0 31372 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2730_
timestamp 1688980957
transform 1 0 31832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2731_
timestamp 1688980957
transform 1 0 31832 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2732_
timestamp 1688980957
transform 1 0 31556 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2733_
timestamp 1688980957
transform 1 0 31188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _2734_
timestamp 1688980957
transform 1 0 31188 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2735_
timestamp 1688980957
transform 1 0 30544 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2736_
timestamp 1688980957
transform 1 0 29716 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2737_
timestamp 1688980957
transform 1 0 28520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2738_
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2739_
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2740_
timestamp 1688980957
transform 1 0 36156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2741_
timestamp 1688980957
transform 1 0 30820 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2742_
timestamp 1688980957
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2743_
timestamp 1688980957
transform 1 0 33396 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2744_
timestamp 1688980957
transform 1 0 33856 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2745_
timestamp 1688980957
transform 1 0 30544 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2746_
timestamp 1688980957
transform 1 0 33396 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2747_
timestamp 1688980957
transform 1 0 33948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _2748_
timestamp 1688980957
transform 1 0 29624 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _2749_
timestamp 1688980957
transform 1 0 32292 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2750_
timestamp 1688980957
transform 1 0 33304 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2751_
timestamp 1688980957
transform 1 0 33120 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2752_
timestamp 1688980957
transform 1 0 32752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2753_
timestamp 1688980957
transform 1 0 35144 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2754_
timestamp 1688980957
transform 1 0 34592 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2755_
timestamp 1688980957
transform 1 0 35328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2756_
timestamp 1688980957
transform 1 0 35604 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2757_
timestamp 1688980957
transform 1 0 34868 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2758_
timestamp 1688980957
transform 1 0 32292 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _2759_
timestamp 1688980957
transform 1 0 32568 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2760_
timestamp 1688980957
transform 1 0 34224 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2761_
timestamp 1688980957
transform 1 0 34408 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2762_
timestamp 1688980957
transform 1 0 35512 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2763_
timestamp 1688980957
transform 1 0 35512 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2764_
timestamp 1688980957
transform 1 0 33120 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2765_
timestamp 1688980957
transform 1 0 33580 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2766_
timestamp 1688980957
transform 1 0 33120 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2767_
timestamp 1688980957
transform 1 0 32936 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2768_
timestamp 1688980957
transform 1 0 35328 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2769_
timestamp 1688980957
transform 1 0 35420 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2770_
timestamp 1688980957
transform 1 0 35696 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2771_
timestamp 1688980957
transform 1 0 35604 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2772_
timestamp 1688980957
transform 1 0 34868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _2773_
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2774_
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2775_
timestamp 1688980957
transform 1 0 33488 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _2776_
timestamp 1688980957
transform 1 0 33212 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2777_
timestamp 1688980957
transform 1 0 33856 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2778_
timestamp 1688980957
transform 1 0 34776 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2779_
timestamp 1688980957
transform 1 0 35512 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2780_
timestamp 1688980957
transform 1 0 35788 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2781_
timestamp 1688980957
transform 1 0 35236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2782_
timestamp 1688980957
transform 1 0 35972 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2783_
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2784_
timestamp 1688980957
transform 1 0 35972 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2785_
timestamp 1688980957
transform 1 0 35604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2786_
timestamp 1688980957
transform 1 0 36432 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2787_
timestamp 1688980957
transform 1 0 37076 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2788_
timestamp 1688980957
transform 1 0 37904 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2789_
timestamp 1688980957
transform 1 0 21344 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _2790_
timestamp 1688980957
transform 1 0 21528 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2791_
timestamp 1688980957
transform 1 0 20700 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _2792_
timestamp 1688980957
transform 1 0 20516 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _2793_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2794_
timestamp 1688980957
transform 1 0 14536 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2795_
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2796_
timestamp 1688980957
transform 1 0 13064 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2797_
timestamp 1688980957
transform 1 0 13800 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2798_
timestamp 1688980957
transform 1 0 14536 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2799_
timestamp 1688980957
transform 1 0 14444 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2800_
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2801_
timestamp 1688980957
transform 1 0 10396 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _2802_
timestamp 1688980957
transform 1 0 10764 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _2803_
timestamp 1688980957
transform 1 0 36984 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2804_
timestamp 1688980957
transform 1 0 36708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2805_
timestamp 1688980957
transform 1 0 22724 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2806_
timestamp 1688980957
transform 1 0 23276 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _2807_
timestamp 1688980957
transform 1 0 23000 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2808_
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2809_
timestamp 1688980957
transform 1 0 34592 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2810_
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _2811_
timestamp 1688980957
transform 1 0 26036 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2812_
timestamp 1688980957
transform 1 0 17296 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2813_
timestamp 1688980957
transform 1 0 16744 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2814_
timestamp 1688980957
transform 1 0 24472 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2815_
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2816_
timestamp 1688980957
transform 1 0 26864 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2817_
timestamp 1688980957
transform 1 0 38088 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2818_
timestamp 1688980957
transform 1 0 38916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2819_
timestamp 1688980957
transform 1 0 21160 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2820_
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2821_
timestamp 1688980957
transform 1 0 4508 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2822_
timestamp 1688980957
transform 1 0 3956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2823_
timestamp 1688980957
transform 1 0 26404 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _2824_
timestamp 1688980957
transform 1 0 26864 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2825_
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2826_
timestamp 1688980957
transform 1 0 34224 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2827_
timestamp 1688980957
transform 1 0 23736 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _2828_
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2829_
timestamp 1688980957
transform 1 0 37168 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2830_
timestamp 1688980957
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2831_
timestamp 1688980957
transform 1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2832_
timestamp 1688980957
transform 1 0 25484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _2833_
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2834_
timestamp 1688980957
transform 1 0 37352 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2835_
timestamp 1688980957
transform 1 0 37076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2836_
timestamp 1688980957
transform 1 0 31556 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2837_
timestamp 1688980957
transform 1 0 32108 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2838_
timestamp 1688980957
transform 1 0 24472 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2839_
timestamp 1688980957
transform 1 0 24748 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2840_
timestamp 1688980957
transform 1 0 24656 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2841_
timestamp 1688980957
transform 1 0 25024 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2842_
timestamp 1688980957
transform 1 0 18952 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2843_
timestamp 1688980957
transform 1 0 18584 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2844_
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2845_
timestamp 1688980957
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2846_
timestamp 1688980957
transform 1 0 23000 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2847_
timestamp 1688980957
transform 1 0 22724 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2848_
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2849_
timestamp 1688980957
transform 1 0 28520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2850_
timestamp 1688980957
transform 1 0 20516 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2851_
timestamp 1688980957
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2852_
timestamp 1688980957
transform 1 0 26404 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2853_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2854_
timestamp 1688980957
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2855_
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2856_
timestamp 1688980957
transform 1 0 25668 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2857_
timestamp 1688980957
transform 1 0 25760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2858_
timestamp 1688980957
transform 1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2859_
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2860_
timestamp 1688980957
transform 1 0 20424 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_4  _2861_
timestamp 1688980957
transform 1 0 19044 0 -1 26112
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2862_
timestamp 1688980957
transform 1 0 14076 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2863_
timestamp 1688980957
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2864_
timestamp 1688980957
transform 1 0 14444 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2865_
timestamp 1688980957
transform 1 0 14168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2866_
timestamp 1688980957
transform 1 0 13064 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2867_
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2868_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2869_
timestamp 1688980957
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2870_
timestamp 1688980957
transform 1 0 15640 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2871_
timestamp 1688980957
transform 1 0 15272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2872_
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2873_
timestamp 1688980957
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2874_
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2875_
timestamp 1688980957
transform 1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2876_
timestamp 1688980957
transform 1 0 13156 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2877_
timestamp 1688980957
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2878_
timestamp 1688980957
transform 1 0 37720 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2879_
timestamp 1688980957
transform 1 0 36248 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2880_
timestamp 1688980957
transform 1 0 36156 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2881_
timestamp 1688980957
transform 1 0 38824 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2882_
timestamp 1688980957
transform 1 0 38916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2883_
timestamp 1688980957
transform 1 0 35604 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2884_
timestamp 1688980957
transform 1 0 34960 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2885_
timestamp 1688980957
transform 1 0 36432 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2886_
timestamp 1688980957
transform 1 0 36708 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2887_
timestamp 1688980957
transform 1 0 36616 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2888_
timestamp 1688980957
transform 1 0 38272 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2889_
timestamp 1688980957
transform 1 0 36248 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2890_
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2891_
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2892_
timestamp 1688980957
transform 1 0 38456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2893_
timestamp 1688980957
transform 1 0 38916 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2894_
timestamp 1688980957
transform 1 0 38548 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2895_
timestamp 1688980957
transform 1 0 39192 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2896_
timestamp 1688980957
transform 1 0 39192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2897_
timestamp 1688980957
transform 1 0 38732 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2898_
timestamp 1688980957
transform 1 0 39192 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2899_
timestamp 1688980957
transform 1 0 38364 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2900_
timestamp 1688980957
transform 1 0 38824 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2901_
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2902_
timestamp 1688980957
transform 1 0 38548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2903_
timestamp 1688980957
transform 1 0 38364 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2904_
timestamp 1688980957
transform 1 0 38640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _2905_
timestamp 1688980957
transform 1 0 39100 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2906_
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2907_
timestamp 1688980957
transform 1 0 36800 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2908_
timestamp 1688980957
transform 1 0 37720 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2909_
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2910_
timestamp 1688980957
transform 1 0 38640 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2911_
timestamp 1688980957
transform 1 0 38364 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2912_
timestamp 1688980957
transform 1 0 35880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2913_
timestamp 1688980957
transform 1 0 36156 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2914_
timestamp 1688980957
transform 1 0 36616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2915_
timestamp 1688980957
transform 1 0 37352 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2916_
timestamp 1688980957
transform 1 0 39468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2917_
timestamp 1688980957
transform 1 0 39008 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2918_
timestamp 1688980957
transform 1 0 39744 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _2919_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38916 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2920_
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2921_
timestamp 1688980957
transform 1 0 38640 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2922_
timestamp 1688980957
transform 1 0 38272 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2923_
timestamp 1688980957
transform 1 0 38456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2924_
timestamp 1688980957
transform 1 0 36800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2925_
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2926_
timestamp 1688980957
transform 1 0 38824 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_2  _2927_
timestamp 1688980957
transform 1 0 38916 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2928_
timestamp 1688980957
transform 1 0 37720 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2929_
timestamp 1688980957
transform 1 0 36064 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2930_
timestamp 1688980957
transform 1 0 35604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2931_
timestamp 1688980957
transform 1 0 35972 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2932_
timestamp 1688980957
transform 1 0 36432 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2933_
timestamp 1688980957
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2934_
timestamp 1688980957
transform 1 0 36064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2935_
timestamp 1688980957
transform 1 0 36616 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2936_
timestamp 1688980957
transform 1 0 33672 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2937_
timestamp 1688980957
transform 1 0 34132 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2938_
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _2939_
timestamp 1688980957
transform 1 0 38088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2940_
timestamp 1688980957
transform 1 0 34132 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2941_
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2942_
timestamp 1688980957
transform 1 0 35144 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2943_
timestamp 1688980957
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2944_
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2945_
timestamp 1688980957
transform 1 0 35144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2946_
timestamp 1688980957
transform 1 0 34776 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2947_
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2948_
timestamp 1688980957
transform 1 0 31096 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2949_
timestamp 1688980957
transform 1 0 30544 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2950_
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2951_
timestamp 1688980957
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2952_
timestamp 1688980957
transform 1 0 31004 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2953_
timestamp 1688980957
transform 1 0 32292 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2954_
timestamp 1688980957
transform 1 0 33120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2955_
timestamp 1688980957
transform 1 0 32476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2956_
timestamp 1688980957
transform 1 0 32200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2957_
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2958_
timestamp 1688980957
transform 1 0 33580 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2959_
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2960_
timestamp 1688980957
transform 1 0 33028 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2961_
timestamp 1688980957
transform 1 0 32752 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2962_
timestamp 1688980957
transform 1 0 31556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2963_
timestamp 1688980957
transform 1 0 30544 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2964_
timestamp 1688980957
transform 1 0 30544 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2965_
timestamp 1688980957
transform 1 0 30452 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2966_
timestamp 1688980957
transform 1 0 30912 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2967_
timestamp 1688980957
transform 1 0 29716 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2968_
timestamp 1688980957
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2969_
timestamp 1688980957
transform 1 0 12144 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2970_
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2971_
timestamp 1688980957
transform 1 0 12236 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2972_
timestamp 1688980957
transform 1 0 12696 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _2973_
timestamp 1688980957
transform 1 0 11776 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _2974_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2975_
timestamp 1688980957
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2976_
timestamp 1688980957
transform 1 0 30728 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2977_
timestamp 1688980957
transform 1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2978_
timestamp 1688980957
transform 1 0 29808 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2979_
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2980_
timestamp 1688980957
transform 1 0 40020 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2981_
timestamp 1688980957
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2982_
timestamp 1688980957
transform 1 0 4416 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2983_
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2984_
timestamp 1688980957
transform 1 0 10580 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2985_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2986_
timestamp 1688980957
transform 1 0 4232 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2987_
timestamp 1688980957
transform 1 0 3680 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2988_
timestamp 1688980957
transform 1 0 40020 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2989_
timestamp 1688980957
transform 1 0 39468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2990_
timestamp 1688980957
transform 1 0 30544 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2991_
timestamp 1688980957
transform 1 0 35420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2992_
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2993_
timestamp 1688980957
transform 1 0 33948 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2994_
timestamp 1688980957
transform 1 0 34868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2995_
timestamp 1688980957
transform 1 0 33212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2996_
timestamp 1688980957
transform 1 0 33304 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2997_
timestamp 1688980957
transform 1 0 5336 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2998_
timestamp 1688980957
transform 1 0 5060 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2999_
timestamp 1688980957
transform 1 0 32752 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _3000_
timestamp 1688980957
transform 1 0 33028 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _3001_
timestamp 1688980957
transform 1 0 31096 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _3002_
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _3003_
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _3004_
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3005_
timestamp 1688980957
transform 1 0 6900 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _3006_
timestamp 1688980957
transform 1 0 11960 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _3007_
timestamp 1688980957
transform 1 0 11316 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _3008_
timestamp 1688980957
transform 1 0 9844 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _3009_
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _3010_
timestamp 1688980957
transform 1 0 7360 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3011_
timestamp 1688980957
transform 1 0 6716 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _3012_
timestamp 1688980957
transform 1 0 10396 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _3013_
timestamp 1688980957
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _3014_
timestamp 1688980957
transform 1 0 20792 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _3015_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _3016_
timestamp 1688980957
transform 1 0 25484 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _3017_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3018_
timestamp 1688980957
transform 1 0 27232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _3019_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3020_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3021_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3022_
timestamp 1688980957
transform 1 0 9660 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3023_
timestamp 1688980957
transform 1 0 7268 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3024_
timestamp 1688980957
transform 1 0 9200 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3025_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3026_
timestamp 1688980957
transform 1 0 12236 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3027_
timestamp 1688980957
transform 1 0 11040 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3028_
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3029_
timestamp 1688980957
transform 1 0 9568 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3030_
timestamp 1688980957
transform 1 0 7636 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3031_
timestamp 1688980957
transform 1 0 8004 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3032_
timestamp 1688980957
transform 1 0 14720 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3033_
timestamp 1688980957
transform 1 0 18308 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3034_
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3035_
timestamp 1688980957
transform 1 0 14628 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3036_
timestamp 1688980957
transform 1 0 16560 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3037_
timestamp 1688980957
transform 1 0 13616 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3038_
timestamp 1688980957
transform 1 0 16744 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3039_
timestamp 1688980957
transform 1 0 23460 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3040_
timestamp 1688980957
transform 1 0 2668 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3041_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3042_
timestamp 1688980957
transform 1 0 12144 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3043_
timestamp 1688980957
transform 1 0 9568 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3044_
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3045_
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3046_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3047_
timestamp 1688980957
transform 1 0 2668 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3048_
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3049_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3050_
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3051_
timestamp 1688980957
transform 1 0 10212 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3052_
timestamp 1688980957
transform 1 0 1656 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3053_
timestamp 1688980957
transform 1 0 29256 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3054_
timestamp 1688980957
transform 1 0 35788 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3055_
timestamp 1688980957
transform 1 0 4324 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3056_
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3057_
timestamp 1688980957
transform 1 0 36248 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3058_
timestamp 1688980957
transform 1 0 20516 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3059_
timestamp 1688980957
transform 1 0 22264 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3060_
timestamp 1688980957
transform 1 0 25024 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3061_
timestamp 1688980957
transform 1 0 27048 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3062_
timestamp 1688980957
transform 1 0 20424 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3063_
timestamp 1688980957
transform 1 0 27232 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3064_
timestamp 1688980957
transform 1 0 22356 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3065_
timestamp 1688980957
transform 1 0 26404 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3066_
timestamp 1688980957
transform 1 0 29900 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3067_
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3068_
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3069_
timestamp 1688980957
transform 1 0 28244 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3070_
timestamp 1688980957
transform 1 0 33028 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3071_
timestamp 1688980957
transform 1 0 36248 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3072_
timestamp 1688980957
transform 1 0 33304 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3073_
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3074_
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3075_
timestamp 1688980957
transform 1 0 34224 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3076_
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3077_
timestamp 1688980957
transform 1 0 38824 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3078_
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3079_
timestamp 1688980957
transform 1 0 34500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3080_
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3081_
timestamp 1688980957
transform 1 0 37352 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3082_
timestamp 1688980957
transform 1 0 32476 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3083_
timestamp 1688980957
transform 1 0 17940 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3084_
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3085_
timestamp 1688980957
transform 1 0 22264 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3086_
timestamp 1688980957
transform 1 0 27324 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3087_
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3088_
timestamp 1688980957
transform 1 0 27324 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3089_
timestamp 1688980957
transform 1 0 18584 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3090_
timestamp 1688980957
transform 1 0 25208 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3091_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3092_
timestamp 1688980957
transform 1 0 13800 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3093_
timestamp 1688980957
transform 1 0 12144 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3094_
timestamp 1688980957
transform 1 0 12144 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3095_
timestamp 1688980957
transform 1 0 14720 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3096_
timestamp 1688980957
transform 1 0 13248 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3097_
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3098_
timestamp 1688980957
transform 1 0 12696 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3099_
timestamp 1688980957
transform 1 0 38364 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3100_
timestamp 1688980957
transform 1 0 39192 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3101_
timestamp 1688980957
transform 1 0 39008 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3102_
timestamp 1688980957
transform 1 0 38088 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3103_
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3104_
timestamp 1688980957
transform 1 0 34684 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3105_
timestamp 1688980957
transform 1 0 31648 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3106_
timestamp 1688980957
transform 1 0 28612 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3107_
timestamp 1688980957
transform 1 0 5060 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3108_
timestamp 1688980957
transform 1 0 31556 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3109_
timestamp 1688980957
transform 1 0 29992 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3110_
timestamp 1688980957
transform 1 0 39284 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3111_
timestamp 1688980957
transform 1 0 3220 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3112_
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3113_
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3114_
timestamp 1688980957
transform 1 0 39284 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3115_
timestamp 1688980957
transform 1 0 32568 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3116_
timestamp 1688980957
transform 1 0 30636 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3117_
timestamp 1688980957
transform 1 0 37904 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3118_
timestamp 1688980957
transform 1 0 37628 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3119_
timestamp 1688980957
transform 1 0 34776 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3120_
timestamp 1688980957
transform 1 0 34776 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3121_
timestamp 1688980957
transform 1 0 33580 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3122_
timestamp 1688980957
transform 1 0 4416 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3123_
timestamp 1688980957
transform 1 0 33672 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _3124_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3125_
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _3126_
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3127_
timestamp 1688980957
transform 1 0 4140 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3128_
timestamp 1688980957
transform 1 0 5612 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3129_
timestamp 1688980957
transform 1 0 4324 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3130_
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3131_
timestamp 1688980957
transform 1 0 4048 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3132_
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3133_
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3134_
timestamp 1688980957
transform 1 0 25760 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3135_
timestamp 1688980957
transform 1 0 32660 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3136_
timestamp 1688980957
transform 1 0 28244 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3137_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3138_
timestamp 1688980957
transform 1 0 33488 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3139_
timestamp 1688980957
transform 1 0 32752 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3140_
timestamp 1688980957
transform 1 0 33580 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3141_
timestamp 1688980957
transform 1 0 33764 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3142_
timestamp 1688980957
transform 1 0 32384 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3143_
timestamp 1688980957
transform 1 0 33304 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3144_
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _3145_
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3146_
timestamp 1688980957
transform 1 0 8464 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3147_
timestamp 1688980957
transform 1 0 27508 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _3148_
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 31188 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform 1 0 15732 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 17020 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform 1 0 4600 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform 1 0 4232 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 6624 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform 1 0 10672 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform 1 0 25668 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 28796 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform 1 0 36616 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 37628 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform 1 0 37720 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform 1 0 37352 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 33488 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 1688980957
transform 1 0 11592 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 1688980957
transform 1 0 13616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 1688980957
transform 1 0 14904 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout60
timestamp 1688980957
transform 1 0 9660 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout61
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout64
timestamp 1688980957
transform 1 0 21712 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout65
timestamp 1688980957
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout66
timestamp 1688980957
transform 1 0 27416 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1688980957
transform 1 0 10396 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout68
timestamp 1688980957
transform 1 0 13616 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 1688980957
transform 1 0 37628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout71
timestamp 1688980957
transform 1 0 32108 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 1688980957
transform 1 0 14536 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_79
timestamp 1688980957
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_163
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_210
timestamp 1688980957
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp 1688980957
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_247
timestamp 1688980957
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_289
timestamp 1688980957
transform 1 0 27692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_301
timestamp 1688980957
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_331
timestamp 1688980957
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_373
timestamp 1688980957
transform 1 0 35420 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_385
timestamp 1688980957
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1688980957
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_415
timestamp 1688980957
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_419
timestamp 1688980957
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_146
timestamp 1688980957
transform 1 0 14536 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_189
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_197
timestamp 1688980957
transform 1 0 19228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_220
timestamp 1688980957
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_232
timestamp 1688980957
transform 1 0 22448 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_240
timestamp 1688980957
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_263
timestamp 1688980957
transform 1 0 25300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_276
timestamp 1688980957
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_9
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_21
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_127
timestamp 1688980957
transform 1 0 12788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_157
timestamp 1688980957
transform 1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_170
timestamp 1688980957
transform 1 0 16744 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_174
timestamp 1688980957
transform 1 0 17112 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_206
timestamp 1688980957
transform 1 0 20056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_282
timestamp 1688980957
transform 1 0 27048 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_294
timestamp 1688980957
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_306
timestamp 1688980957
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_185
timestamp 1688980957
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_234
timestamp 1688980957
transform 1 0 22632 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_246
timestamp 1688980957
transform 1 0 23736 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_251
timestamp 1688980957
transform 1 0 24196 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_259
timestamp 1688980957
transform 1 0 24932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_271
timestamp 1688980957
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_278
timestamp 1688980957
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_413
timestamp 1688980957
transform 1 0 39100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_425
timestamp 1688980957
transform 1 0 40204 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_433
timestamp 1688980957
transform 1 0 40940 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_117
timestamp 1688980957
transform 1 0 11868 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_128
timestamp 1688980957
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_226
timestamp 1688980957
transform 1 0 21896 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_238
timestamp 1688980957
transform 1 0 23000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_295
timestamp 1688980957
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_385
timestamp 1688980957
transform 1 0 36524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_399
timestamp 1688980957
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_403
timestamp 1688980957
transform 1 0 38180 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_412
timestamp 1688980957
transform 1 0 39008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_43
timestamp 1688980957
transform 1 0 5060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1688980957
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_74
timestamp 1688980957
transform 1 0 7912 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_86
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_94
timestamp 1688980957
transform 1 0 9752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_116
timestamp 1688980957
transform 1 0 11776 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_140
timestamp 1688980957
transform 1 0 13984 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_152
timestamp 1688980957
transform 1 0 15088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_164
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_220
timestamp 1688980957
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_357
timestamp 1688980957
transform 1 0 33948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_383
timestamp 1688980957
transform 1 0 36340 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_63
timestamp 1688980957
transform 1 0 6900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_78
timestamp 1688980957
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_119
timestamp 1688980957
transform 1 0 12052 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_127
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_167
timestamp 1688980957
transform 1 0 16468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_182
timestamp 1688980957
transform 1 0 17848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_231
timestamp 1688980957
transform 1 0 22356 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_250
timestamp 1688980957
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_262
timestamp 1688980957
transform 1 0 25208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_266
timestamp 1688980957
transform 1 0 25576 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_278
timestamp 1688980957
transform 1 0 26680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_290
timestamp 1688980957
transform 1 0 27784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_302
timestamp 1688980957
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_351
timestamp 1688980957
transform 1 0 33396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_374
timestamp 1688980957
transform 1 0 35512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_384
timestamp 1688980957
transform 1 0 36432 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_94
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_123
timestamp 1688980957
transform 1 0 12420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_127
timestamp 1688980957
transform 1 0 12788 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_131
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_135
timestamp 1688980957
transform 1 0 13524 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_142
timestamp 1688980957
transform 1 0 14168 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_150
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_155
timestamp 1688980957
transform 1 0 15364 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_210
timestamp 1688980957
transform 1 0 20424 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1688980957
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_229
timestamp 1688980957
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_266
timestamp 1688980957
transform 1 0 25576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 1688980957
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_284
timestamp 1688980957
transform 1 0 27232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_326
timestamp 1688980957
transform 1 0 31096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_334
timestamp 1688980957
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_421
timestamp 1688980957
transform 1 0 39836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_433
timestamp 1688980957
transform 1 0 40940 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_98
timestamp 1688980957
transform 1 0 10120 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_106
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_113
timestamp 1688980957
transform 1 0 11500 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_119
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_150
timestamp 1688980957
transform 1 0 14904 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_162
timestamp 1688980957
transform 1 0 16008 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_172
timestamp 1688980957
transform 1 0 16928 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_180
timestamp 1688980957
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_192
timestamp 1688980957
transform 1 0 18768 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_228
timestamp 1688980957
transform 1 0 22080 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_240
timestamp 1688980957
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_264
timestamp 1688980957
transform 1 0 25392 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_272
timestamp 1688980957
transform 1 0 26128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_302
timestamp 1688980957
transform 1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_320
timestamp 1688980957
transform 1 0 30544 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_329
timestamp 1688980957
transform 1 0 31372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_341
timestamp 1688980957
transform 1 0 32476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_353
timestamp 1688980957
transform 1 0 33580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_361
timestamp 1688980957
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_385
timestamp 1688980957
transform 1 0 36524 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_397
timestamp 1688980957
transform 1 0 37628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_409
timestamp 1688980957
transform 1 0 38732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_417
timestamp 1688980957
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_164
timestamp 1688980957
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_175
timestamp 1688980957
transform 1 0 17204 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_185
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_197
timestamp 1688980957
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_209
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_215
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_238
timestamp 1688980957
transform 1 0 23000 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_250
timestamp 1688980957
transform 1 0 24104 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_266
timestamp 1688980957
transform 1 0 25576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_276
timestamp 1688980957
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_301
timestamp 1688980957
transform 1 0 28796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_313
timestamp 1688980957
transform 1 0 29900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_325
timestamp 1688980957
transform 1 0 31004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_333
timestamp 1688980957
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_386
timestamp 1688980957
transform 1 0 36616 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_409
timestamp 1688980957
transform 1 0 38732 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_430
timestamp 1688980957
transform 1 0 40664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_434
timestamp 1688980957
transform 1 0 41032 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 1688980957
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_49
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_59
timestamp 1688980957
transform 1 0 6532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_71
timestamp 1688980957
transform 1 0 7636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_93
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_104
timestamp 1688980957
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_120
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_127
timestamp 1688980957
transform 1 0 12788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1688980957
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_154
timestamp 1688980957
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_164
timestamp 1688980957
transform 1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_168
timestamp 1688980957
transform 1 0 16560 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_183
timestamp 1688980957
transform 1 0 17940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_204
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_212
timestamp 1688980957
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_229
timestamp 1688980957
transform 1 0 22172 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_239
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_275
timestamp 1688980957
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_287
timestamp 1688980957
transform 1 0 27508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_299
timestamp 1688980957
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_317
timestamp 1688980957
transform 1 0 30268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_355
timestamp 1688980957
transform 1 0 33764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_359
timestamp 1688980957
transform 1 0 34132 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_370
timestamp 1688980957
transform 1 0 35144 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_382
timestamp 1688980957
transform 1 0 36248 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_394
timestamp 1688980957
transform 1 0 37352 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_414
timestamp 1688980957
transform 1 0 39192 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_429
timestamp 1688980957
transform 1 0 40572 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_37
timestamp 1688980957
transform 1 0 4508 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_66
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_78
timestamp 1688980957
transform 1 0 8280 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_99
timestamp 1688980957
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_139
timestamp 1688980957
transform 1 0 13892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_153
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_165
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_211
timestamp 1688980957
transform 1 0 20516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_251
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_257
timestamp 1688980957
transform 1 0 24748 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_263
timestamp 1688980957
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_275
timestamp 1688980957
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_284
timestamp 1688980957
transform 1 0 27232 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 1688980957
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_353
timestamp 1688980957
transform 1 0 33580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_382
timestamp 1688980957
transform 1 0 36248 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_416
timestamp 1688980957
transform 1 0 39376 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_428
timestamp 1688980957
transform 1 0 40480 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_42
timestamp 1688980957
transform 1 0 4968 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_54
timestamp 1688980957
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_64
timestamp 1688980957
transform 1 0 6992 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_76
timestamp 1688980957
transform 1 0 8096 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1688980957
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_101
timestamp 1688980957
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_146
timestamp 1688980957
transform 1 0 14536 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_158
timestamp 1688980957
transform 1 0 15640 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_164
timestamp 1688980957
transform 1 0 16192 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_179
timestamp 1688980957
transform 1 0 17572 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_187
timestamp 1688980957
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 1688980957
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_202
timestamp 1688980957
transform 1 0 19688 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_210
timestamp 1688980957
transform 1 0 20424 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_231
timestamp 1688980957
transform 1 0 22356 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_243
timestamp 1688980957
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_273
timestamp 1688980957
transform 1 0 26220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_304
timestamp 1688980957
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_351
timestamp 1688980957
transform 1 0 33396 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_362
timestamp 1688980957
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_368
timestamp 1688980957
transform 1 0 34960 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_415
timestamp 1688980957
transform 1 0 39284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_52
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_88
timestamp 1688980957
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_135
timestamp 1688980957
transform 1 0 13524 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1688980957
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_176
timestamp 1688980957
transform 1 0 17296 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_188
timestamp 1688980957
transform 1 0 18400 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_203
timestamp 1688980957
transform 1 0 19780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_231
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_243
timestamp 1688980957
transform 1 0 23460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_255
timestamp 1688980957
transform 1 0 24564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_259
timestamp 1688980957
transform 1 0 24932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_266
timestamp 1688980957
transform 1 0 25576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_275
timestamp 1688980957
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_298
timestamp 1688980957
transform 1 0 28520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_327
timestamp 1688980957
transform 1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_342
timestamp 1688980957
transform 1 0 32568 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_354
timestamp 1688980957
transform 1 0 33672 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_366
timestamp 1688980957
transform 1 0 34776 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_378
timestamp 1688980957
transform 1 0 35880 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_390
timestamp 1688980957
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_401
timestamp 1688980957
transform 1 0 37996 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_409
timestamp 1688980957
transform 1 0 38732 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_423
timestamp 1688980957
transform 1 0 40020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_63
timestamp 1688980957
transform 1 0 6900 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_69
timestamp 1688980957
transform 1 0 7452 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_126
timestamp 1688980957
transform 1 0 12696 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1688980957
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_172
timestamp 1688980957
transform 1 0 16928 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_184
timestamp 1688980957
transform 1 0 18032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_188
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_239
timestamp 1688980957
transform 1 0 23092 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_243
timestamp 1688980957
transform 1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_275
timestamp 1688980957
transform 1 0 26404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_287
timestamp 1688980957
transform 1 0 27508 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_293
timestamp 1688980957
transform 1 0 28060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_317
timestamp 1688980957
transform 1 0 30268 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_326
timestamp 1688980957
transform 1 0 31096 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_338
timestamp 1688980957
transform 1 0 32200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_351
timestamp 1688980957
transform 1 0 33396 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_359
timestamp 1688980957
transform 1 0 34132 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_374
timestamp 1688980957
transform 1 0 35512 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_386
timestamp 1688980957
transform 1 0 36616 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_398
timestamp 1688980957
transform 1 0 37720 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_410
timestamp 1688980957
transform 1 0 38824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_428
timestamp 1688980957
transform 1 0 40480 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_434
timestamp 1688980957
transform 1 0 41032 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_89
timestamp 1688980957
transform 1 0 9292 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_97
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1688980957
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_119
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_131
timestamp 1688980957
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_152
timestamp 1688980957
transform 1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_173
timestamp 1688980957
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_180
timestamp 1688980957
transform 1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_184
timestamp 1688980957
transform 1 0 18032 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_206
timestamp 1688980957
transform 1 0 20056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_218
timestamp 1688980957
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_247
timestamp 1688980957
transform 1 0 23828 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_255
timestamp 1688980957
transform 1 0 24564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_274
timestamp 1688980957
transform 1 0 26312 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_320
timestamp 1688980957
transform 1 0 30544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_333
timestamp 1688980957
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_346
timestamp 1688980957
transform 1 0 32936 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_358
timestamp 1688980957
transform 1 0 34040 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_373
timestamp 1688980957
transform 1 0 35420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_384
timestamp 1688980957
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_405
timestamp 1688980957
transform 1 0 38364 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 1688980957
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_429
timestamp 1688980957
transform 1 0 40572 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_9
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_21
timestamp 1688980957
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_49
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_55
timestamp 1688980957
transform 1 0 6164 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_67
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 1688980957
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_127
timestamp 1688980957
transform 1 0 12788 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_135
timestamp 1688980957
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_156
timestamp 1688980957
transform 1 0 15456 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_164
timestamp 1688980957
transform 1 0 16192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_191
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_227
timestamp 1688980957
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_341
timestamp 1688980957
transform 1 0 32476 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_351
timestamp 1688980957
transform 1 0 33396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_372
timestamp 1688980957
transform 1 0 35328 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_378
timestamp 1688980957
transform 1 0 35880 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_393
timestamp 1688980957
transform 1 0 37260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_401
timestamp 1688980957
transform 1 0 37996 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_413
timestamp 1688980957
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 1688980957
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_433
timestamp 1688980957
transform 1 0 40940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_26
timestamp 1688980957
transform 1 0 3496 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_34
timestamp 1688980957
transform 1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_48
timestamp 1688980957
transform 1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_63
timestamp 1688980957
transform 1 0 6900 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_84
timestamp 1688980957
transform 1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_95
timestamp 1688980957
transform 1 0 9844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_122
timestamp 1688980957
transform 1 0 12328 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_128
timestamp 1688980957
transform 1 0 12880 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_138
timestamp 1688980957
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_150
timestamp 1688980957
transform 1 0 14904 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_160
timestamp 1688980957
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_173
timestamp 1688980957
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_180
timestamp 1688980957
transform 1 0 17664 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_198
timestamp 1688980957
transform 1 0 19320 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_234
timestamp 1688980957
transform 1 0 22632 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_245
timestamp 1688980957
transform 1 0 23644 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_267
timestamp 1688980957
transform 1 0 25668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_286
timestamp 1688980957
transform 1 0 27416 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_294
timestamp 1688980957
transform 1 0 28152 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_318
timestamp 1688980957
transform 1 0 30360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_330
timestamp 1688980957
transform 1 0 31464 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_373
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_390
timestamp 1688980957
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_401
timestamp 1688980957
transform 1 0 37996 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_423
timestamp 1688980957
transform 1 0 40020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_11
timestamp 1688980957
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_61
timestamp 1688980957
transform 1 0 6716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_73
timestamp 1688980957
transform 1 0 7820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_94
timestamp 1688980957
transform 1 0 9752 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_100
timestamp 1688980957
transform 1 0 10304 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_106
timestamp 1688980957
transform 1 0 10856 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_136
timestamp 1688980957
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_150
timestamp 1688980957
transform 1 0 14904 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_154
timestamp 1688980957
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_168
timestamp 1688980957
transform 1 0 16560 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_180
timestamp 1688980957
transform 1 0 17664 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_192
timestamp 1688980957
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_204
timestamp 1688980957
transform 1 0 19872 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_216
timestamp 1688980957
transform 1 0 20976 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_228
timestamp 1688980957
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1688980957
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_266
timestamp 1688980957
transform 1 0 25576 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_274
timestamp 1688980957
transform 1 0 26312 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_278
timestamp 1688980957
transform 1 0 26680 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_297
timestamp 1688980957
transform 1 0 28428 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_337
timestamp 1688980957
transform 1 0 32108 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_349
timestamp 1688980957
transform 1 0 33212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_361
timestamp 1688980957
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_401
timestamp 1688980957
transform 1 0 37996 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_405
timestamp 1688980957
transform 1 0 38364 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_409
timestamp 1688980957
transform 1 0 38732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_432
timestamp 1688980957
transform 1 0 40848 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_64
timestamp 1688980957
transform 1 0 6992 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_89
timestamp 1688980957
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_101
timestamp 1688980957
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_119
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_131
timestamp 1688980957
transform 1 0 13156 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_143
timestamp 1688980957
transform 1 0 14260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_147
timestamp 1688980957
transform 1 0 14628 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_187
timestamp 1688980957
transform 1 0 18308 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_210
timestamp 1688980957
transform 1 0 20424 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_219
timestamp 1688980957
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_243
timestamp 1688980957
transform 1 0 23460 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_252
timestamp 1688980957
transform 1 0 24288 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_264
timestamp 1688980957
transform 1 0 25392 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_276
timestamp 1688980957
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_312
timestamp 1688980957
transform 1 0 29808 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_324
timestamp 1688980957
transform 1 0 30912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_334
timestamp 1688980957
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_345
timestamp 1688980957
transform 1 0 32844 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_368
timestamp 1688980957
transform 1 0 34960 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_380
timestamp 1688980957
transform 1 0 36064 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_400
timestamp 1688980957
transform 1 0 37904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_412
timestamp 1688980957
transform 1 0 39008 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_49
timestamp 1688980957
transform 1 0 5612 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_59
timestamp 1688980957
transform 1 0 6532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_71
timestamp 1688980957
transform 1 0 7636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_117
timestamp 1688980957
transform 1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1688980957
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_161
timestamp 1688980957
transform 1 0 15916 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_181
timestamp 1688980957
transform 1 0 17756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1688980957
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_205
timestamp 1688980957
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_215
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_227
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_239
timestamp 1688980957
transform 1 0 23092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_269
timestamp 1688980957
transform 1 0 25852 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_291
timestamp 1688980957
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_303
timestamp 1688980957
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_339
timestamp 1688980957
transform 1 0 32292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_354
timestamp 1688980957
transform 1 0 33672 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_360
timestamp 1688980957
transform 1 0 34224 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_380
timestamp 1688980957
transform 1 0 36064 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_384
timestamp 1688980957
transform 1 0 36432 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_396
timestamp 1688980957
transform 1 0 37536 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_37
timestamp 1688980957
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_49
timestamp 1688980957
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_122
timestamp 1688980957
transform 1 0 12328 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_134
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_146
timestamp 1688980957
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_150
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1688980957
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_176
timestamp 1688980957
transform 1 0 17296 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_201
timestamp 1688980957
transform 1 0 19596 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_210
timestamp 1688980957
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_214
timestamp 1688980957
transform 1 0 20792 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_246
timestamp 1688980957
transform 1 0 23736 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_275
timestamp 1688980957
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_298
timestamp 1688980957
transform 1 0 28520 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_310
timestamp 1688980957
transform 1 0 29624 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_322
timestamp 1688980957
transform 1 0 30728 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_342
timestamp 1688980957
transform 1 0 32568 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_363
timestamp 1688980957
transform 1 0 34500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_381
timestamp 1688980957
transform 1 0 36156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_23
timestamp 1688980957
transform 1 0 3220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_45
timestamp 1688980957
transform 1 0 5244 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_79
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_90
timestamp 1688980957
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_118
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_126
timestamp 1688980957
transform 1 0 12696 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_135
timestamp 1688980957
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_169
timestamp 1688980957
transform 1 0 16652 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_205
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_219
timestamp 1688980957
transform 1 0 21252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_225
timestamp 1688980957
transform 1 0 21804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_239
timestamp 1688980957
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_273
timestamp 1688980957
transform 1 0 26220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_297
timestamp 1688980957
transform 1 0 28428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_305
timestamp 1688980957
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_340
timestamp 1688980957
transform 1 0 32384 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_352
timestamp 1688980957
transform 1 0 33488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_429
timestamp 1688980957
transform 1 0 40572 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_43
timestamp 1688980957
transform 1 0 5060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_50
timestamp 1688980957
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_64
timestamp 1688980957
transform 1 0 6992 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_70
timestamp 1688980957
transform 1 0 7544 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_117
timestamp 1688980957
transform 1 0 11868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_140
timestamp 1688980957
transform 1 0 13984 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_153
timestamp 1688980957
transform 1 0 15180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_165
timestamp 1688980957
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_176
timestamp 1688980957
transform 1 0 17296 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_182
timestamp 1688980957
transform 1 0 17848 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_189
timestamp 1688980957
transform 1 0 18492 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_197
timestamp 1688980957
transform 1 0 19228 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_233
timestamp 1688980957
transform 1 0 22540 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_238
timestamp 1688980957
transform 1 0 23000 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_246
timestamp 1688980957
transform 1 0 23736 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_254
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_266
timestamp 1688980957
transform 1 0 25576 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1688980957
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_295
timestamp 1688980957
transform 1 0 28244 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_307
timestamp 1688980957
transform 1 0 29348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_315
timestamp 1688980957
transform 1 0 30084 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_319
timestamp 1688980957
transform 1 0 30452 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_369
timestamp 1688980957
transform 1 0 35052 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_375
timestamp 1688980957
transform 1 0 35604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_387
timestamp 1688980957
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1688980957
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_405
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_412
timestamp 1688980957
transform 1 0 39008 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_424
timestamp 1688980957
transform 1 0 40112 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_432
timestamp 1688980957
transform 1 0 40848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_46
timestamp 1688980957
transform 1 0 5336 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_58
timestamp 1688980957
transform 1 0 6440 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_70
timestamp 1688980957
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_112
timestamp 1688980957
transform 1 0 11408 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_124
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_136
timestamp 1688980957
transform 1 0 13616 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_161
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_173
timestamp 1688980957
transform 1 0 17020 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_192
timestamp 1688980957
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_230
timestamp 1688980957
transform 1 0 22264 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_236
timestamp 1688980957
transform 1 0 22816 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_261
timestamp 1688980957
transform 1 0 25116 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_273
timestamp 1688980957
transform 1 0 26220 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_285
timestamp 1688980957
transform 1 0 27324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_297
timestamp 1688980957
transform 1 0 28428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_305
timestamp 1688980957
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_316
timestamp 1688980957
transform 1 0 30176 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_328
timestamp 1688980957
transform 1 0 31280 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_340
timestamp 1688980957
transform 1 0 32384 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_348
timestamp 1688980957
transform 1 0 33120 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_373
timestamp 1688980957
transform 1 0 35420 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1688980957
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1688980957
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 1688980957
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 1688980957
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1688980957
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_433
timestamp 1688980957
transform 1 0 40940 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_6
timestamp 1688980957
transform 1 0 1656 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_18
timestamp 1688980957
transform 1 0 2760 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_26
timestamp 1688980957
transform 1 0 3496 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_41
timestamp 1688980957
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_74
timestamp 1688980957
transform 1 0 7912 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_86
timestamp 1688980957
transform 1 0 9016 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_91
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_103
timestamp 1688980957
transform 1 0 10580 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_124
timestamp 1688980957
transform 1 0 12512 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_136
timestamp 1688980957
transform 1 0 13616 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_148
timestamp 1688980957
transform 1 0 14720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_152
timestamp 1688980957
transform 1 0 15088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_160
timestamp 1688980957
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_176
timestamp 1688980957
transform 1 0 17296 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_182
timestamp 1688980957
transform 1 0 17848 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_189
timestamp 1688980957
transform 1 0 18492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_201
timestamp 1688980957
transform 1 0 19596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_207
timestamp 1688980957
transform 1 0 20148 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_221
timestamp 1688980957
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_233
timestamp 1688980957
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_246
timestamp 1688980957
transform 1 0 23736 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_259
timestamp 1688980957
transform 1 0 24932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_268
timestamp 1688980957
transform 1 0 25760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_272
timestamp 1688980957
transform 1 0 26128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_290
timestamp 1688980957
transform 1 0 27784 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_298
timestamp 1688980957
transform 1 0 28520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_304
timestamp 1688980957
transform 1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_314
timestamp 1688980957
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_326
timestamp 1688980957
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_334
timestamp 1688980957
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_346
timestamp 1688980957
transform 1 0 32936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_360
timestamp 1688980957
transform 1 0 34224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_369
timestamp 1688980957
transform 1 0 35052 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_381
timestamp 1688980957
transform 1 0 36156 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1688980957
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_403
timestamp 1688980957
transform 1 0 38180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_412
timestamp 1688980957
transform 1 0 39008 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_37
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_49
timestamp 1688980957
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_61
timestamp 1688980957
transform 1 0 6716 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_69
timestamp 1688980957
transform 1 0 7452 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1688980957
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_92
timestamp 1688980957
transform 1 0 9568 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_104
timestamp 1688980957
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_108
timestamp 1688980957
transform 1 0 11040 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_170
timestamp 1688980957
transform 1 0 16744 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_184
timestamp 1688980957
transform 1 0 18032 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_234
timestamp 1688980957
transform 1 0 22632 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_238
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_246
timestamp 1688980957
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_295
timestamp 1688980957
transform 1 0 28244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_334
timestamp 1688980957
transform 1 0 31832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_338
timestamp 1688980957
transform 1 0 32200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1688980957
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_377
timestamp 1688980957
transform 1 0 35788 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_381
timestamp 1688980957
transform 1 0 36156 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_393
timestamp 1688980957
transform 1 0 37260 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_397
timestamp 1688980957
transform 1 0 37628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_402
timestamp 1688980957
transform 1 0 38088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_406
timestamp 1688980957
transform 1 0 38456 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_421
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_432
timestamp 1688980957
transform 1 0 40848 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_35
timestamp 1688980957
transform 1 0 4324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_48
timestamp 1688980957
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_67
timestamp 1688980957
transform 1 0 7268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_95
timestamp 1688980957
transform 1 0 9844 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_107
timestamp 1688980957
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_118
timestamp 1688980957
transform 1 0 11960 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_145
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_164
timestamp 1688980957
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_195
timestamp 1688980957
transform 1 0 19044 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_203
timestamp 1688980957
transform 1 0 19780 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_211
timestamp 1688980957
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_219
timestamp 1688980957
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_244
timestamp 1688980957
transform 1 0 23552 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_248
timestamp 1688980957
transform 1 0 23920 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_253
timestamp 1688980957
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_266
timestamp 1688980957
transform 1 0 25576 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_274
timestamp 1688980957
transform 1 0 26312 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 1688980957
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_316
timestamp 1688980957
transform 1 0 30176 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_326
timestamp 1688980957
transform 1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_334
timestamp 1688980957
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_345
timestamp 1688980957
transform 1 0 32844 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_355
timestamp 1688980957
transform 1 0 33764 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_367
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_379
timestamp 1688980957
transform 1 0 35972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_405
timestamp 1688980957
transform 1 0 38364 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_418
timestamp 1688980957
transform 1 0 39560 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_426
timestamp 1688980957
transform 1 0 40296 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_23
timestamp 1688980957
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_55
timestamp 1688980957
transform 1 0 6164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_67
timestamp 1688980957
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_79
timestamp 1688980957
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_92
timestamp 1688980957
transform 1 0 9568 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_96
timestamp 1688980957
transform 1 0 9936 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_100
timestamp 1688980957
transform 1 0 10304 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_108
timestamp 1688980957
transform 1 0 11040 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_118
timestamp 1688980957
transform 1 0 11960 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_126
timestamp 1688980957
transform 1 0 12696 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_144
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_162
timestamp 1688980957
transform 1 0 16008 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_174
timestamp 1688980957
transform 1 0 17112 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_212
timestamp 1688980957
transform 1 0 20608 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_224
timestamp 1688980957
transform 1 0 21712 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_230
timestamp 1688980957
transform 1 0 22264 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_239
timestamp 1688980957
transform 1 0 23092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_277
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_285
timestamp 1688980957
transform 1 0 27324 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_297
timestamp 1688980957
transform 1 0 28428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_305
timestamp 1688980957
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_317
timestamp 1688980957
transform 1 0 30268 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_332
timestamp 1688980957
transform 1 0 31648 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_344
timestamp 1688980957
transform 1 0 32752 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_356
timestamp 1688980957
transform 1 0 33856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_392
timestamp 1688980957
transform 1 0 37168 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_404
timestamp 1688980957
transform 1 0 38272 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_412
timestamp 1688980957
transform 1 0 39008 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 1688980957
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_23
timestamp 1688980957
transform 1 0 3220 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_35
timestamp 1688980957
transform 1 0 4324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_52
timestamp 1688980957
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_68
timestamp 1688980957
transform 1 0 7360 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_80
timestamp 1688980957
transform 1 0 8464 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_92
timestamp 1688980957
transform 1 0 9568 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_100
timestamp 1688980957
transform 1 0 10304 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_117
timestamp 1688980957
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_127
timestamp 1688980957
transform 1 0 12788 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_139
timestamp 1688980957
transform 1 0 13892 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_147
timestamp 1688980957
transform 1 0 14628 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_163
timestamp 1688980957
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_200
timestamp 1688980957
transform 1 0 19504 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_204
timestamp 1688980957
transform 1 0 19872 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_209
timestamp 1688980957
transform 1 0 20332 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_215
timestamp 1688980957
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_229
timestamp 1688980957
transform 1 0 22172 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_239
timestamp 1688980957
transform 1 0 23092 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_257
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_269
timestamp 1688980957
transform 1 0 25852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_277
timestamp 1688980957
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_296
timestamp 1688980957
transform 1 0 28336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_304
timestamp 1688980957
transform 1 0 29072 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_314
timestamp 1688980957
transform 1 0 29992 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_326
timestamp 1688980957
transform 1 0 31096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_333
timestamp 1688980957
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_343
timestamp 1688980957
transform 1 0 32660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_347
timestamp 1688980957
transform 1 0 33028 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_360
timestamp 1688980957
transform 1 0 34224 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_371
timestamp 1688980957
transform 1 0 35236 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_383
timestamp 1688980957
transform 1 0 36340 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_400
timestamp 1688980957
transform 1 0 37904 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_404
timestamp 1688980957
transform 1 0 38272 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_52
timestamp 1688980957
transform 1 0 5888 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_75
timestamp 1688980957
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_79
timestamp 1688980957
transform 1 0 8372 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_100
timestamp 1688980957
transform 1 0 10304 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_112
timestamp 1688980957
transform 1 0 11408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_120
timestamp 1688980957
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_127
timestamp 1688980957
transform 1 0 12788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_158
timestamp 1688980957
transform 1 0 15640 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_162
timestamp 1688980957
transform 1 0 16008 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_182
timestamp 1688980957
transform 1 0 17848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_186
timestamp 1688980957
transform 1 0 18216 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_193
timestamp 1688980957
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_206
timestamp 1688980957
transform 1 0 20056 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_218
timestamp 1688980957
transform 1 0 21160 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_226
timestamp 1688980957
transform 1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_232
timestamp 1688980957
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_243
timestamp 1688980957
transform 1 0 23460 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_267
timestamp 1688980957
transform 1 0 25668 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_279
timestamp 1688980957
transform 1 0 26772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_283
timestamp 1688980957
transform 1 0 27140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_318
timestamp 1688980957
transform 1 0 30360 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_326
timestamp 1688980957
transform 1 0 31096 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_342
timestamp 1688980957
transform 1 0 32568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_359
timestamp 1688980957
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_374
timestamp 1688980957
transform 1 0 35512 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_394
timestamp 1688980957
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_406
timestamp 1688980957
transform 1 0 38456 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 1688980957
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_424
timestamp 1688980957
transform 1 0 40112 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_432
timestamp 1688980957
transform 1 0 40848 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_49
timestamp 1688980957
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_70
timestamp 1688980957
transform 1 0 7544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_95
timestamp 1688980957
transform 1 0 9844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_119
timestamp 1688980957
transform 1 0 12052 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_130
timestamp 1688980957
transform 1 0 13064 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_138
timestamp 1688980957
transform 1 0 13800 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_153
timestamp 1688980957
transform 1 0 15180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_182
timestamp 1688980957
transform 1 0 17848 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_194
timestamp 1688980957
transform 1 0 18952 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_245
timestamp 1688980957
transform 1 0 23644 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_257
timestamp 1688980957
transform 1 0 24748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_263
timestamp 1688980957
transform 1 0 25300 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_272
timestamp 1688980957
transform 1 0 26128 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_290
timestamp 1688980957
transform 1 0 27784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_302
timestamp 1688980957
transform 1 0 28888 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_310
timestamp 1688980957
transform 1 0 29624 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_334
timestamp 1688980957
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_340
timestamp 1688980957
transform 1 0 32384 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_352
timestamp 1688980957
transform 1 0 33488 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 1688980957
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 1688980957
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 1688980957
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 1688980957
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_429
timestamp 1688980957
transform 1 0 40572 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 1688980957
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_35
timestamp 1688980957
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_42
timestamp 1688980957
transform 1 0 4968 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_54
timestamp 1688980957
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_58
timestamp 1688980957
transform 1 0 6440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_74
timestamp 1688980957
transform 1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_82
timestamp 1688980957
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_103
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_128
timestamp 1688980957
transform 1 0 12880 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_151
timestamp 1688980957
transform 1 0 14996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_163
timestamp 1688980957
transform 1 0 16100 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_172
timestamp 1688980957
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_186
timestamp 1688980957
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1688980957
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_215
timestamp 1688980957
transform 1 0 20884 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_238
timestamp 1688980957
transform 1 0 23000 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_242
timestamp 1688980957
transform 1 0 23368 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_248
timestamp 1688980957
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_261
timestamp 1688980957
transform 1 0 25116 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_332
timestamp 1688980957
transform 1 0 31648 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_344
timestamp 1688980957
transform 1 0 32752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_360
timestamp 1688980957
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_371
timestamp 1688980957
transform 1 0 35236 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_387
timestamp 1688980957
transform 1 0 36708 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_399
timestamp 1688980957
transform 1 0 37812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_403
timestamp 1688980957
transform 1 0 38180 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_414
timestamp 1688980957
transform 1 0 39192 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_433
timestamp 1688980957
transform 1 0 40940 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_49
timestamp 1688980957
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_135
timestamp 1688980957
transform 1 0 13524 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_156
timestamp 1688980957
transform 1 0 15456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_160
timestamp 1688980957
transform 1 0 15824 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_179
timestamp 1688980957
transform 1 0 17572 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_186
timestamp 1688980957
transform 1 0 18216 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_194
timestamp 1688980957
transform 1 0 18952 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_212
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_242
timestamp 1688980957
transform 1 0 23368 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_254
timestamp 1688980957
transform 1 0 24472 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_266
timestamp 1688980957
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_318
timestamp 1688980957
transform 1 0 30360 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_330
timestamp 1688980957
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_345
timestamp 1688980957
transform 1 0 32844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_389
timestamp 1688980957
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_397
timestamp 1688980957
transform 1 0 37628 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_428
timestamp 1688980957
transform 1 0 40480 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_434
timestamp 1688980957
transform 1 0 41032 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_40
timestamp 1688980957
transform 1 0 4784 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_48
timestamp 1688980957
transform 1 0 5520 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_74
timestamp 1688980957
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1688980957
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_99
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_106
timestamp 1688980957
transform 1 0 10856 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_118
timestamp 1688980957
transform 1 0 11960 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_135
timestamp 1688980957
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_159
timestamp 1688980957
transform 1 0 15732 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_176
timestamp 1688980957
transform 1 0 17296 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_188
timestamp 1688980957
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_206
timestamp 1688980957
transform 1 0 20056 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_218
timestamp 1688980957
transform 1 0 21160 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_230
timestamp 1688980957
transform 1 0 22264 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_242
timestamp 1688980957
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_250
timestamp 1688980957
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_261
timestamp 1688980957
transform 1 0 25116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_273
timestamp 1688980957
transform 1 0 26220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_281
timestamp 1688980957
transform 1 0 26956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_285
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_296
timestamp 1688980957
transform 1 0 28336 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_304
timestamp 1688980957
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_314
timestamp 1688980957
transform 1 0 29992 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_341
timestamp 1688980957
transform 1 0 32476 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_353
timestamp 1688980957
transform 1 0 33580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_361
timestamp 1688980957
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_371
timestamp 1688980957
transform 1 0 35236 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_382
timestamp 1688980957
transform 1 0 36248 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_394
timestamp 1688980957
transform 1 0 37352 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_402
timestamp 1688980957
transform 1 0 38088 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_415
timestamp 1688980957
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 1688980957
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_37
timestamp 1688980957
transform 1 0 4508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 1688980957
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1688980957
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_117
timestamp 1688980957
transform 1 0 11868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_129
timestamp 1688980957
transform 1 0 12972 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_141
timestamp 1688980957
transform 1 0 14076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_153
timestamp 1688980957
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1688980957
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_197
timestamp 1688980957
transform 1 0 19228 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_209
timestamp 1688980957
transform 1 0 20332 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1688980957
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_238
timestamp 1688980957
transform 1 0 23000 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_242
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_248
timestamp 1688980957
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_260
timestamp 1688980957
transform 1 0 25024 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_311
timestamp 1688980957
transform 1 0 29716 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_319
timestamp 1688980957
transform 1 0 30452 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_360
timestamp 1688980957
transform 1 0 34224 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_372
timestamp 1688980957
transform 1 0 35328 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1688980957
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1688980957
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 1688980957
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_429
timestamp 1688980957
transform 1 0 40572 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_17
timestamp 1688980957
transform 1 0 2668 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_25
timestamp 1688980957
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_49
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_61
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_76
timestamp 1688980957
transform 1 0 8096 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_82
timestamp 1688980957
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_93
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_102
timestamp 1688980957
transform 1 0 10488 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_147
timestamp 1688980957
transform 1 0 14628 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_160
timestamp 1688980957
transform 1 0 15824 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_172
timestamp 1688980957
transform 1 0 16928 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_176
timestamp 1688980957
transform 1 0 17296 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_200
timestamp 1688980957
transform 1 0 19504 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_206
timestamp 1688980957
transform 1 0 20056 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_262
timestamp 1688980957
transform 1 0 25208 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_274
timestamp 1688980957
transform 1 0 26312 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_292
timestamp 1688980957
transform 1 0 27968 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_302
timestamp 1688980957
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_320
timestamp 1688980957
transform 1 0 30544 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_332
timestamp 1688980957
transform 1 0 31648 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_344
timestamp 1688980957
transform 1 0 32752 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_356
timestamp 1688980957
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_373
timestamp 1688980957
transform 1 0 35420 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_381
timestamp 1688980957
transform 1 0 36156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_389
timestamp 1688980957
transform 1 0 36892 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_403
timestamp 1688980957
transform 1 0 38180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_415
timestamp 1688980957
transform 1 0 39284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1688980957
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_433
timestamp 1688980957
transform 1 0 40940 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_35
timestamp 1688980957
transform 1 0 4324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_90
timestamp 1688980957
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_108
timestamp 1688980957
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_124
timestamp 1688980957
transform 1 0 12512 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_162
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_173
timestamp 1688980957
transform 1 0 17020 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_185
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_196
timestamp 1688980957
transform 1 0 19136 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_204
timestamp 1688980957
transform 1 0 19872 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_216
timestamp 1688980957
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_256
timestamp 1688980957
transform 1 0 24656 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_268
timestamp 1688980957
transform 1 0 25760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_313
timestamp 1688980957
transform 1 0 29900 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_325
timestamp 1688980957
transform 1 0 31004 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_333
timestamp 1688980957
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_367
timestamp 1688980957
transform 1 0 34868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_379
timestamp 1688980957
transform 1 0 35972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_416
timestamp 1688980957
transform 1 0 39376 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_428
timestamp 1688980957
transform 1 0 40480 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_434
timestamp 1688980957
transform 1 0 41032 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_7
timestamp 1688980957
transform 1 0 1748 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_11
timestamp 1688980957
transform 1 0 2116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_23
timestamp 1688980957
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_46
timestamp 1688980957
transform 1 0 5336 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_59
timestamp 1688980957
transform 1 0 6532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_74
timestamp 1688980957
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 1688980957
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_90
timestamp 1688980957
transform 1 0 9384 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_98
timestamp 1688980957
transform 1 0 10120 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_114
timestamp 1688980957
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_126
timestamp 1688980957
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1688980957
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_166
timestamp 1688980957
transform 1 0 16376 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_178
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_186
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_205
timestamp 1688980957
transform 1 0 19964 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_220
timestamp 1688980957
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_232
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1688980957
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_273
timestamp 1688980957
transform 1 0 26220 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_295
timestamp 1688980957
transform 1 0 28244 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_305
timestamp 1688980957
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_324
timestamp 1688980957
transform 1 0 30912 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_374
timestamp 1688980957
transform 1 0 35512 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_386
timestamp 1688980957
transform 1 0 36616 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_398
timestamp 1688980957
transform 1 0 37720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_410
timestamp 1688980957
transform 1 0 38824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_418
timestamp 1688980957
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_421
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_433
timestamp 1688980957
transform 1 0 40940 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_85
timestamp 1688980957
transform 1 0 8924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_108
timestamp 1688980957
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_121
timestamp 1688980957
transform 1 0 12236 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_131
timestamp 1688980957
transform 1 0 13156 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_143
timestamp 1688980957
transform 1 0 14260 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_157
timestamp 1688980957
transform 1 0 15548 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_166
timestamp 1688980957
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_179
timestamp 1688980957
transform 1 0 17572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_187
timestamp 1688980957
transform 1 0 18308 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_195
timestamp 1688980957
transform 1 0 19044 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_207
timestamp 1688980957
transform 1 0 20148 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_212
timestamp 1688980957
transform 1 0 20608 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_221
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_256
timestamp 1688980957
transform 1 0 24656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_272
timestamp 1688980957
transform 1 0 26128 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_294
timestamp 1688980957
transform 1 0 28152 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_306
timestamp 1688980957
transform 1 0 29256 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_334
timestamp 1688980957
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_358
timestamp 1688980957
transform 1 0 34040 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_390
timestamp 1688980957
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_396
timestamp 1688980957
transform 1 0 37536 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_409
timestamp 1688980957
transform 1 0 38732 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_421
timestamp 1688980957
transform 1 0 39836 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_433
timestamp 1688980957
transform 1 0 40940 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_9
timestamp 1688980957
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_21
timestamp 1688980957
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_66
timestamp 1688980957
transform 1 0 7176 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_78
timestamp 1688980957
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_106
timestamp 1688980957
transform 1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_116
timestamp 1688980957
transform 1 0 11776 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_120
timestamp 1688980957
transform 1 0 12144 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_136
timestamp 1688980957
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_147
timestamp 1688980957
transform 1 0 14628 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_155
timestamp 1688980957
transform 1 0 15364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_166
timestamp 1688980957
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_187
timestamp 1688980957
transform 1 0 18308 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_194
timestamp 1688980957
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_206
timestamp 1688980957
transform 1 0 20056 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_222
timestamp 1688980957
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_226
timestamp 1688980957
transform 1 0 21896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 1688980957
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_261
timestamp 1688980957
transform 1 0 25116 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_269
timestamp 1688980957
transform 1 0 25852 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_292
timestamp 1688980957
transform 1 0 27968 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_304
timestamp 1688980957
transform 1 0 29072 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_313
timestamp 1688980957
transform 1 0 29900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_326
timestamp 1688980957
transform 1 0 31096 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_332
timestamp 1688980957
transform 1 0 31648 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_336
timestamp 1688980957
transform 1 0 32016 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_348
timestamp 1688980957
transform 1 0 33120 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_360
timestamp 1688980957
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_377
timestamp 1688980957
transform 1 0 35788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_381
timestamp 1688980957
transform 1 0 36156 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_402
timestamp 1688980957
transform 1 0 38088 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_414
timestamp 1688980957
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_433
timestamp 1688980957
transform 1 0 40940 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_31
timestamp 1688980957
transform 1 0 3956 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_43
timestamp 1688980957
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_88
timestamp 1688980957
transform 1 0 9200 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_100
timestamp 1688980957
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_117
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_148
timestamp 1688980957
transform 1 0 14720 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_162
timestamp 1688980957
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_173
timestamp 1688980957
transform 1 0 17020 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_180
timestamp 1688980957
transform 1 0 17664 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_192
timestamp 1688980957
transform 1 0 18768 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_238
timestamp 1688980957
transform 1 0 23000 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_253
timestamp 1688980957
transform 1 0 24380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_265
timestamp 1688980957
transform 1 0 25484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 1688980957
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_288
timestamp 1688980957
transform 1 0 27600 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_300
timestamp 1688980957
transform 1 0 28704 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_312
timestamp 1688980957
transform 1 0 29808 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_324
timestamp 1688980957
transform 1 0 30912 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_331
timestamp 1688980957
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1688980957
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 1688980957
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1688980957
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 1688980957
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 1688980957
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_429
timestamp 1688980957
transform 1 0 40572 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_49
timestamp 1688980957
transform 1 0 5612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_64
timestamp 1688980957
transform 1 0 6992 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_72
timestamp 1688980957
transform 1 0 7728 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_96
timestamp 1688980957
transform 1 0 9936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_108
timestamp 1688980957
transform 1 0 11040 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_112
timestamp 1688980957
transform 1 0 11408 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_124
timestamp 1688980957
transform 1 0 12512 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_136
timestamp 1688980957
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_145
timestamp 1688980957
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_176
timestamp 1688980957
transform 1 0 17296 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_182
timestamp 1688980957
transform 1 0 17848 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_191
timestamp 1688980957
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_215
timestamp 1688980957
transform 1 0 20884 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_223
timestamp 1688980957
transform 1 0 21620 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_231
timestamp 1688980957
transform 1 0 22356 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_239
timestamp 1688980957
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_266
timestamp 1688980957
transform 1 0 25576 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_278
timestamp 1688980957
transform 1 0 26680 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_290
timestamp 1688980957
transform 1 0 27784 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_297
timestamp 1688980957
transform 1 0 28428 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_312
timestamp 1688980957
transform 1 0 29808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_316
timestamp 1688980957
transform 1 0 30176 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_320
timestamp 1688980957
transform 1 0 30544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_324
timestamp 1688980957
transform 1 0 30912 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_329
timestamp 1688980957
transform 1 0 31372 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 1688980957
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 1688980957
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1688980957
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_433
timestamp 1688980957
transform 1 0 40940 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_35
timestamp 1688980957
transform 1 0 4324 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_87
timestamp 1688980957
transform 1 0 9108 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_102
timestamp 1688980957
transform 1 0 10488 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_131
timestamp 1688980957
transform 1 0 13156 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_191
timestamp 1688980957
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_209
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_221
timestamp 1688980957
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_257
timestamp 1688980957
transform 1 0 24748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_301
timestamp 1688980957
transform 1 0 28796 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_313
timestamp 1688980957
transform 1 0 29900 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_319
timestamp 1688980957
transform 1 0 30452 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_325
timestamp 1688980957
transform 1 0 31004 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_389
timestamp 1688980957
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1688980957
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_429
timestamp 1688980957
transform 1 0 40572 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_55
timestamp 1688980957
transform 1 0 6164 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_67
timestamp 1688980957
transform 1 0 7268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_76
timestamp 1688980957
transform 1 0 8096 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_93
timestamp 1688980957
transform 1 0 9660 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_101
timestamp 1688980957
transform 1 0 10396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_106
timestamp 1688980957
transform 1 0 10856 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_110
timestamp 1688980957
transform 1 0 11224 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_114
timestamp 1688980957
transform 1 0 11592 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_126
timestamp 1688980957
transform 1 0 12696 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_138
timestamp 1688980957
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_149
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_164
timestamp 1688980957
transform 1 0 16192 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_176
timestamp 1688980957
transform 1 0 17296 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_207
timestamp 1688980957
transform 1 0 20148 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_217
timestamp 1688980957
transform 1 0 21068 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_225
timestamp 1688980957
transform 1 0 21804 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_231
timestamp 1688980957
transform 1 0 22356 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_235
timestamp 1688980957
transform 1 0 22724 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_240
timestamp 1688980957
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_280
timestamp 1688980957
transform 1 0 26864 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_292
timestamp 1688980957
transform 1 0 27968 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_304
timestamp 1688980957
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_353
timestamp 1688980957
transform 1 0 33580 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_361
timestamp 1688980957
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_381
timestamp 1688980957
transform 1 0 36156 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_393
timestamp 1688980957
transform 1 0 37260 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_405
timestamp 1688980957
transform 1 0 38364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_417
timestamp 1688980957
transform 1 0 39468 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_433
timestamp 1688980957
transform 1 0 40940 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_34
timestamp 1688980957
transform 1 0 4232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_46
timestamp 1688980957
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 1688980957
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_80
timestamp 1688980957
transform 1 0 8464 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_98
timestamp 1688980957
transform 1 0 10120 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_110
timestamp 1688980957
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_131
timestamp 1688980957
transform 1 0 13156 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_139
timestamp 1688980957
transform 1 0 13892 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_147
timestamp 1688980957
transform 1 0 14628 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_172
timestamp 1688980957
transform 1 0 16928 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_179
timestamp 1688980957
transform 1 0 17572 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_187
timestamp 1688980957
transform 1 0 18308 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_194
timestamp 1688980957
transform 1 0 18952 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_201
timestamp 1688980957
transform 1 0 19596 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_254
timestamp 1688980957
transform 1 0 24472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_271
timestamp 1688980957
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_306
timestamp 1688980957
transform 1 0 29256 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_312
timestamp 1688980957
transform 1 0 29808 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_323
timestamp 1688980957
transform 1 0 30820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_345
timestamp 1688980957
transform 1 0 32844 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_374
timestamp 1688980957
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_386
timestamp 1688980957
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1688980957
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_429
timestamp 1688980957
transform 1 0 40572 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_64
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_76
timestamp 1688980957
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_92
timestamp 1688980957
transform 1 0 9568 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_104
timestamp 1688980957
transform 1 0 10672 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_116
timestamp 1688980957
transform 1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_120
timestamp 1688980957
transform 1 0 12144 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_138
timestamp 1688980957
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_148
timestamp 1688980957
transform 1 0 14720 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_159
timestamp 1688980957
transform 1 0 15732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_166
timestamp 1688980957
transform 1 0 16376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_170
timestamp 1688980957
transform 1 0 16744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_178
timestamp 1688980957
transform 1 0 17480 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_186
timestamp 1688980957
transform 1 0 18216 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_222
timestamp 1688980957
transform 1 0 21528 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_226
timestamp 1688980957
transform 1 0 21896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_242
timestamp 1688980957
transform 1 0 23368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_271
timestamp 1688980957
transform 1 0 26036 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_275
timestamp 1688980957
transform 1 0 26404 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_294
timestamp 1688980957
transform 1 0 28152 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_335
timestamp 1688980957
transform 1 0 31924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_347
timestamp 1688980957
transform 1 0 33028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_359
timestamp 1688980957
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1688980957
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_401
timestamp 1688980957
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_413
timestamp 1688980957
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 1688980957
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_433
timestamp 1688980957
transform 1 0 40940 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_6
timestamp 1688980957
transform 1 0 1656 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_18
timestamp 1688980957
transform 1 0 2760 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_30
timestamp 1688980957
transform 1 0 3864 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_45
timestamp 1688980957
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_53
timestamp 1688980957
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_101
timestamp 1688980957
transform 1 0 10396 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_109
timestamp 1688980957
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_129
timestamp 1688980957
transform 1 0 12972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_141
timestamp 1688980957
transform 1 0 14076 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_145
timestamp 1688980957
transform 1 0 14444 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_154
timestamp 1688980957
transform 1 0 15272 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_158
timestamp 1688980957
transform 1 0 15640 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_166
timestamp 1688980957
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_177
timestamp 1688980957
transform 1 0 17388 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_201
timestamp 1688980957
transform 1 0 19596 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_213
timestamp 1688980957
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_221
timestamp 1688980957
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_291
timestamp 1688980957
transform 1 0 27876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_303
timestamp 1688980957
transform 1 0 28980 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_311
timestamp 1688980957
transform 1 0 29716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_326
timestamp 1688980957
transform 1 0 31096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_330
timestamp 1688980957
transform 1 0 31464 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_355
timestamp 1688980957
transform 1 0 33764 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_364
timestamp 1688980957
transform 1 0 34592 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_375
timestamp 1688980957
transform 1 0 35604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_387
timestamp 1688980957
transform 1 0 36708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1688980957
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_403
timestamp 1688980957
transform 1 0 38180 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_414
timestamp 1688980957
transform 1 0 39192 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_426
timestamp 1688980957
transform 1 0 40296 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_434
timestamp 1688980957
transform 1 0 41032 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_69
timestamp 1688980957
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 1688980957
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_90
timestamp 1688980957
transform 1 0 9384 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_98
timestamp 1688980957
transform 1 0 10120 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_116
timestamp 1688980957
transform 1 0 11776 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_123
timestamp 1688980957
transform 1 0 12420 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_131
timestamp 1688980957
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_148
timestamp 1688980957
transform 1 0 14720 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_160
timestamp 1688980957
transform 1 0 15824 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_172
timestamp 1688980957
transform 1 0 16928 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_184
timestamp 1688980957
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_203
timestamp 1688980957
transform 1 0 19780 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_214
timestamp 1688980957
transform 1 0 20792 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_218
timestamp 1688980957
transform 1 0 21160 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_226
timestamp 1688980957
transform 1 0 21896 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_239
timestamp 1688980957
transform 1 0 23092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_260
timestamp 1688980957
transform 1 0 25024 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_268
timestamp 1688980957
transform 1 0 25760 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_297
timestamp 1688980957
transform 1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_312
timestamp 1688980957
transform 1 0 29808 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_318
timestamp 1688980957
transform 1 0 30360 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_330
timestamp 1688980957
transform 1 0 31464 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_342
timestamp 1688980957
transform 1 0 32568 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_354
timestamp 1688980957
transform 1 0 33672 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_362
timestamp 1688980957
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 1688980957
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_389
timestamp 1688980957
transform 1 0 36892 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_414
timestamp 1688980957
transform 1 0 39192 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 1688980957
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_433
timestamp 1688980957
transform 1 0 40940 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_31
timestamp 1688980957
transform 1 0 3956 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_91
timestamp 1688980957
transform 1 0 9476 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_106
timestamp 1688980957
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_129
timestamp 1688980957
transform 1 0 12972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_141
timestamp 1688980957
transform 1 0 14076 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_156
timestamp 1688980957
transform 1 0 15456 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_164
timestamp 1688980957
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_176
timestamp 1688980957
transform 1 0 17296 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_184
timestamp 1688980957
transform 1 0 18032 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_203
timestamp 1688980957
transform 1 0 19780 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_213
timestamp 1688980957
transform 1 0 20700 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1688980957
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_259
timestamp 1688980957
transform 1 0 24932 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_268
timestamp 1688980957
transform 1 0 25760 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_301
timestamp 1688980957
transform 1 0 28796 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_307
timestamp 1688980957
transform 1 0 29348 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_326
timestamp 1688980957
transform 1 0 31096 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_343
timestamp 1688980957
transform 1 0 32660 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_363
timestamp 1688980957
transform 1 0 34500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_375
timestamp 1688980957
transform 1 0 35604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_388
timestamp 1688980957
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_405
timestamp 1688980957
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_417
timestamp 1688980957
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_429
timestamp 1688980957
transform 1 0 40572 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_54
timestamp 1688980957
transform 1 0 6072 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_66
timestamp 1688980957
transform 1 0 7176 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_70
timestamp 1688980957
transform 1 0 7544 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_78
timestamp 1688980957
transform 1 0 8280 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_91
timestamp 1688980957
transform 1 0 9476 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_101
timestamp 1688980957
transform 1 0 10396 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_114
timestamp 1688980957
transform 1 0 11592 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_122
timestamp 1688980957
transform 1 0 12328 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_131
timestamp 1688980957
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_156
timestamp 1688980957
transform 1 0 15456 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_210
timestamp 1688980957
transform 1 0 20424 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_230
timestamp 1688980957
transform 1 0 22264 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_237
timestamp 1688980957
transform 1 0 22908 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_242
timestamp 1688980957
transform 1 0 23368 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_250
timestamp 1688980957
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_257
timestamp 1688980957
transform 1 0 24748 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_261
timestamp 1688980957
transform 1 0 25116 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_273
timestamp 1688980957
transform 1 0 26220 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_285
timestamp 1688980957
transform 1 0 27324 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_294
timestamp 1688980957
transform 1 0 28152 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_306
timestamp 1688980957
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_403
timestamp 1688980957
transform 1 0 38180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_415
timestamp 1688980957
transform 1 0 39284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_419
timestamp 1688980957
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 1688980957
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_433
timestamp 1688980957
transform 1 0 40940 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_77
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_83
timestamp 1688980957
transform 1 0 8740 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_88
timestamp 1688980957
transform 1 0 9200 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_100
timestamp 1688980957
transform 1 0 10304 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_119
timestamp 1688980957
transform 1 0 12052 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_131
timestamp 1688980957
transform 1 0 13156 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_165
timestamp 1688980957
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_174
timestamp 1688980957
transform 1 0 17112 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_210
timestamp 1688980957
transform 1 0 20424 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_218
timestamp 1688980957
transform 1 0 21160 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_222
timestamp 1688980957
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_233
timestamp 1688980957
transform 1 0 22540 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_247
timestamp 1688980957
transform 1 0 23828 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_259
timestamp 1688980957
transform 1 0 24932 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_275
timestamp 1688980957
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_309
timestamp 1688980957
transform 1 0 29532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_333
timestamp 1688980957
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_379
timestamp 1688980957
transform 1 0 35972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1688980957
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 1688980957
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_429
timestamp 1688980957
transform 1 0 40572 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_63
timestamp 1688980957
transform 1 0 6900 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_71
timestamp 1688980957
transform 1 0 7636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_89
timestamp 1688980957
transform 1 0 9292 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_100
timestamp 1688980957
transform 1 0 10304 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_108
timestamp 1688980957
transform 1 0 11040 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_156
timestamp 1688980957
transform 1 0 15456 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_170
timestamp 1688980957
transform 1 0 16744 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_178
timestamp 1688980957
transform 1 0 17480 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_186
timestamp 1688980957
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_194
timestamp 1688980957
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_204
timestamp 1688980957
transform 1 0 19872 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_216
timestamp 1688980957
transform 1 0 20976 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_220
timestamp 1688980957
transform 1 0 21344 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_224
timestamp 1688980957
transform 1 0 21712 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_232
timestamp 1688980957
transform 1 0 22448 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_241
timestamp 1688980957
transform 1 0 23276 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_280
timestamp 1688980957
transform 1 0 26864 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_294
timestamp 1688980957
transform 1 0 28152 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_313
timestamp 1688980957
transform 1 0 29900 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_325
timestamp 1688980957
transform 1 0 31004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_337
timestamp 1688980957
transform 1 0 32108 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1688980957
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1688980957
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_401
timestamp 1688980957
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_413
timestamp 1688980957
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 1688980957
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 1688980957
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_433
timestamp 1688980957
transform 1 0 40940 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_47
timestamp 1688980957
transform 1 0 5428 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_88
timestamp 1688980957
transform 1 0 9200 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_96
timestamp 1688980957
transform 1 0 9936 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_108
timestamp 1688980957
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_133
timestamp 1688980957
transform 1 0 13340 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_209
timestamp 1688980957
transform 1 0 20332 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_232
timestamp 1688980957
transform 1 0 22448 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_264
timestamp 1688980957
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_278
timestamp 1688980957
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_319
timestamp 1688980957
transform 1 0 30452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_323
timestamp 1688980957
transform 1 0 30820 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_359
timestamp 1688980957
transform 1 0 34132 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_371
timestamp 1688980957
transform 1 0 35236 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_383
timestamp 1688980957
transform 1 0 36340 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1688980957
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 1688980957
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 1688980957
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_429
timestamp 1688980957
transform 1 0 40572 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_56
timestamp 1688980957
transform 1 0 6256 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_68
timestamp 1688980957
transform 1 0 7360 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_82
timestamp 1688980957
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_106
timestamp 1688980957
transform 1 0 10856 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_118
timestamp 1688980957
transform 1 0 11960 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_122
timestamp 1688980957
transform 1 0 12328 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_131
timestamp 1688980957
transform 1 0 13156 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_157
timestamp 1688980957
transform 1 0 15548 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_164
timestamp 1688980957
transform 1 0 16192 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_168
timestamp 1688980957
transform 1 0 16560 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_175
timestamp 1688980957
transform 1 0 17204 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_192
timestamp 1688980957
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_213
timestamp 1688980957
transform 1 0 20700 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_262
timestamp 1688980957
transform 1 0 25208 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_296
timestamp 1688980957
transform 1 0 28336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_313
timestamp 1688980957
transform 1 0 29900 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_338
timestamp 1688980957
transform 1 0 32200 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_358
timestamp 1688980957
transform 1 0 34040 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_371
timestamp 1688980957
transform 1 0 35236 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_383
timestamp 1688980957
transform 1 0 36340 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_395
timestamp 1688980957
transform 1 0 37444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_407
timestamp 1688980957
transform 1 0 38548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 1688980957
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1688980957
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_433
timestamp 1688980957
transform 1 0 40940 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_9
timestamp 1688980957
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_21
timestamp 1688980957
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_33
timestamp 1688980957
transform 1 0 4140 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_60
timestamp 1688980957
transform 1 0 6624 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_94
timestamp 1688980957
transform 1 0 9752 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_109
timestamp 1688980957
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_119
timestamp 1688980957
transform 1 0 12052 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_129
timestamp 1688980957
transform 1 0 12972 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_145
timestamp 1688980957
transform 1 0 14444 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_190
timestamp 1688980957
transform 1 0 18584 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_213
timestamp 1688980957
transform 1 0 20700 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_221
timestamp 1688980957
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_231
timestamp 1688980957
transform 1 0 22356 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_243
timestamp 1688980957
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_254
timestamp 1688980957
transform 1 0 24472 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_266
timestamp 1688980957
transform 1 0 25576 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_278
timestamp 1688980957
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_290
timestamp 1688980957
transform 1 0 27784 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_298
timestamp 1688980957
transform 1 0 28520 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_304
timestamp 1688980957
transform 1 0 29072 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_312
timestamp 1688980957
transform 1 0 29808 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_376
timestamp 1688980957
transform 1 0 35696 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_388
timestamp 1688980957
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1688980957
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1688980957
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_429
timestamp 1688980957
transform 1 0 40572 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_47
timestamp 1688980957
transform 1 0 5428 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_63
timestamp 1688980957
transform 1 0 6900 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_71
timestamp 1688980957
transform 1 0 7636 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_117
timestamp 1688980957
transform 1 0 11868 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_125
timestamp 1688980957
transform 1 0 12604 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_138
timestamp 1688980957
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_149
timestamp 1688980957
transform 1 0 14812 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_157
timestamp 1688980957
transform 1 0 15548 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_167
timestamp 1688980957
transform 1 0 16468 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_179
timestamp 1688980957
transform 1 0 17572 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_183
timestamp 1688980957
transform 1 0 17940 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_191
timestamp 1688980957
transform 1 0 18676 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_217
timestamp 1688980957
transform 1 0 21068 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_226
timestamp 1688980957
transform 1 0 21896 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_238
timestamp 1688980957
transform 1 0 23000 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_250
timestamp 1688980957
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_258
timestamp 1688980957
transform 1 0 24840 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_283
timestamp 1688980957
transform 1 0 27140 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_302
timestamp 1688980957
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_342
timestamp 1688980957
transform 1 0 32568 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_362
timestamp 1688980957
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_378
timestamp 1688980957
transform 1 0 35880 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_390
timestamp 1688980957
transform 1 0 36984 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_402
timestamp 1688980957
transform 1 0 38088 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_414
timestamp 1688980957
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_421
timestamp 1688980957
transform 1 0 39836 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_429
timestamp 1688980957
transform 1 0 40572 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_78
timestamp 1688980957
transform 1 0 8280 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_99
timestamp 1688980957
transform 1 0 10212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_117
timestamp 1688980957
transform 1 0 11868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_136
timestamp 1688980957
transform 1 0 13616 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_145
timestamp 1688980957
transform 1 0 14444 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_153
timestamp 1688980957
transform 1 0 15180 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_185
timestamp 1688980957
transform 1 0 18124 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_195
timestamp 1688980957
transform 1 0 19044 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_207
timestamp 1688980957
transform 1 0 20148 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_211
timestamp 1688980957
transform 1 0 20516 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_218
timestamp 1688980957
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_250
timestamp 1688980957
transform 1 0 24104 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_262
timestamp 1688980957
transform 1 0 25208 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_274
timestamp 1688980957
transform 1 0 26312 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_289
timestamp 1688980957
transform 1 0 27692 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_296
timestamp 1688980957
transform 1 0 28336 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_312
timestamp 1688980957
transform 1 0 29808 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_324
timestamp 1688980957
transform 1 0 30912 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_328
timestamp 1688980957
transform 1 0 31280 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_377
timestamp 1688980957
transform 1 0 35788 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_389
timestamp 1688980957
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1688980957
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1688980957
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_429
timestamp 1688980957
transform 1 0 40572 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_69
timestamp 1688980957
transform 1 0 7452 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_76
timestamp 1688980957
transform 1 0 8096 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_89
timestamp 1688980957
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_98
timestamp 1688980957
transform 1 0 10120 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_106
timestamp 1688980957
transform 1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_123
timestamp 1688980957
transform 1 0 12420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_137
timestamp 1688980957
transform 1 0 13708 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_146
timestamp 1688980957
transform 1 0 14536 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_160
timestamp 1688980957
transform 1 0 15824 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_168
timestamp 1688980957
transform 1 0 16560 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_174
timestamp 1688980957
transform 1 0 17112 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_184
timestamp 1688980957
transform 1 0 18032 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_193
timestamp 1688980957
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_204
timestamp 1688980957
transform 1 0 19872 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_220
timestamp 1688980957
transform 1 0 21344 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_227
timestamp 1688980957
transform 1 0 21988 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_235
timestamp 1688980957
transform 1 0 22724 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_240
timestamp 1688980957
transform 1 0 23184 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_267
timestamp 1688980957
transform 1 0 25668 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_279
timestamp 1688980957
transform 1 0 26772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_291
timestamp 1688980957
transform 1 0 27876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_303
timestamp 1688980957
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_336
timestamp 1688980957
transform 1 0 32016 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_348
timestamp 1688980957
transform 1 0 33120 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_373
timestamp 1688980957
transform 1 0 35420 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_385
timestamp 1688980957
transform 1 0 36524 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_397
timestamp 1688980957
transform 1 0 37628 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_409
timestamp 1688980957
transform 1 0 38732 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_417
timestamp 1688980957
transform 1 0 39468 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1688980957
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_433
timestamp 1688980957
transform 1 0 40940 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_71
timestamp 1688980957
transform 1 0 7636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_83
timestamp 1688980957
transform 1 0 8740 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_100
timestamp 1688980957
transform 1 0 10304 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_121
timestamp 1688980957
transform 1 0 12236 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_151
timestamp 1688980957
transform 1 0 14996 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_163
timestamp 1688980957
transform 1 0 16100 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_186
timestamp 1688980957
transform 1 0 18216 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_200
timestamp 1688980957
transform 1 0 19504 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_212
timestamp 1688980957
transform 1 0 20608 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_222
timestamp 1688980957
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_233
timestamp 1688980957
transform 1 0 22540 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_245
timestamp 1688980957
transform 1 0 23644 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_257
timestamp 1688980957
transform 1 0 24748 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_269
timestamp 1688980957
transform 1 0 25852 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_285
timestamp 1688980957
transform 1 0 27324 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_313
timestamp 1688980957
transform 1 0 29900 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_325
timestamp 1688980957
transform 1 0 31004 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_340
timestamp 1688980957
transform 1 0 32384 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_352
timestamp 1688980957
transform 1 0 33488 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_378
timestamp 1688980957
transform 1 0 35880 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_390
timestamp 1688980957
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1688980957
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_429
timestamp 1688980957
transform 1 0 40572 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_64
timestamp 1688980957
transform 1 0 6992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_122
timestamp 1688980957
transform 1 0 12328 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_131
timestamp 1688980957
transform 1 0 13156 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_144
timestamp 1688980957
transform 1 0 14352 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_171
timestamp 1688980957
transform 1 0 16836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_183
timestamp 1688980957
transform 1 0 17940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_229
timestamp 1688980957
transform 1 0 22172 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_234
timestamp 1688980957
transform 1 0 22632 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_246
timestamp 1688980957
transform 1 0 23736 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_269
timestamp 1688980957
transform 1 0 25852 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_281
timestamp 1688980957
transform 1 0 26956 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_285
timestamp 1688980957
transform 1 0 27324 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_293
timestamp 1688980957
transform 1 0 28060 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_316
timestamp 1688980957
transform 1 0 30176 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_326
timestamp 1688980957
transform 1 0 31096 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_338
timestamp 1688980957
transform 1 0 32200 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_360
timestamp 1688980957
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_369
timestamp 1688980957
transform 1 0 35052 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_381
timestamp 1688980957
transform 1 0 36156 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_393
timestamp 1688980957
transform 1 0 37260 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_405
timestamp 1688980957
transform 1 0 38364 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_417
timestamp 1688980957
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1688980957
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_433
timestamp 1688980957
transform 1 0 40940 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_78
timestamp 1688980957
transform 1 0 8280 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_84
timestamp 1688980957
transform 1 0 8832 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_90
timestamp 1688980957
transform 1 0 9384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_108
timestamp 1688980957
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_121
timestamp 1688980957
transform 1 0 12236 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_131
timestamp 1688980957
transform 1 0 13156 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_143
timestamp 1688980957
transform 1 0 14260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_155
timestamp 1688980957
transform 1 0 15364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_199
timestamp 1688980957
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_206
timestamp 1688980957
transform 1 0 20056 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_218
timestamp 1688980957
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_248
timestamp 1688980957
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_260
timestamp 1688980957
transform 1 0 25024 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_268
timestamp 1688980957
transform 1 0 25760 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_276
timestamp 1688980957
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_297
timestamp 1688980957
transform 1 0 28428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_316
timestamp 1688980957
transform 1 0 30176 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_326
timestamp 1688980957
transform 1 0 31096 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_334
timestamp 1688980957
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_342
timestamp 1688980957
transform 1 0 32568 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_370
timestamp 1688980957
transform 1 0 35144 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_382
timestamp 1688980957
transform 1 0 36248 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_390
timestamp 1688980957
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1688980957
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_429
timestamp 1688980957
transform 1 0 40572 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_9
timestamp 1688980957
transform 1 0 1932 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_21
timestamp 1688980957
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_57
timestamp 1688980957
transform 1 0 6348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_79
timestamp 1688980957
transform 1 0 8372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_91
timestamp 1688980957
transform 1 0 9476 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_103
timestamp 1688980957
transform 1 0 10580 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_161
timestamp 1688980957
transform 1 0 15916 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_168
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_176
timestamp 1688980957
transform 1 0 17296 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_185
timestamp 1688980957
transform 1 0 18124 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_218
timestamp 1688980957
transform 1 0 21160 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_236
timestamp 1688980957
transform 1 0 22816 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_257
timestamp 1688980957
transform 1 0 24748 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_266
timestamp 1688980957
transform 1 0 25576 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_278
timestamp 1688980957
transform 1 0 26680 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_282
timestamp 1688980957
transform 1 0 27048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_290
timestamp 1688980957
transform 1 0 27784 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_304
timestamp 1688980957
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_351
timestamp 1688980957
transform 1 0 33396 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1688980957
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1688980957
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1688980957
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1688980957
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_433
timestamp 1688980957
transform 1 0 40940 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_99
timestamp 1688980957
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_110
timestamp 1688980957
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_120
timestamp 1688980957
transform 1 0 12144 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_144
timestamp 1688980957
transform 1 0 14352 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_152
timestamp 1688980957
transform 1 0 15088 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_160
timestamp 1688980957
transform 1 0 15824 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_172
timestamp 1688980957
transform 1 0 16928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_201
timestamp 1688980957
transform 1 0 19596 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_211
timestamp 1688980957
transform 1 0 20516 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_220
timestamp 1688980957
transform 1 0 21344 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_240
timestamp 1688980957
transform 1 0 23184 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_257
timestamp 1688980957
transform 1 0 24748 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_263
timestamp 1688980957
transform 1 0 25300 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_272
timestamp 1688980957
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_289
timestamp 1688980957
transform 1 0 27692 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_297
timestamp 1688980957
transform 1 0 28428 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_306
timestamp 1688980957
transform 1 0 29256 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_318
timestamp 1688980957
transform 1 0 30360 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_324
timestamp 1688980957
transform 1 0 30912 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_342
timestamp 1688980957
transform 1 0 32568 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_346
timestamp 1688980957
transform 1 0 32936 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_350
timestamp 1688980957
transform 1 0 33304 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_354
timestamp 1688980957
transform 1 0 33672 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_375
timestamp 1688980957
transform 1 0 35604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_387
timestamp 1688980957
transform 1 0 36708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1688980957
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1688980957
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_429
timestamp 1688980957
transform 1 0 40572 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_93
timestamp 1688980957
transform 1 0 9660 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_114
timestamp 1688980957
transform 1 0 11592 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_122
timestamp 1688980957
transform 1 0 12328 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1688980957
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_149
timestamp 1688980957
transform 1 0 14812 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_167
timestamp 1688980957
transform 1 0 16468 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_175
timestamp 1688980957
transform 1 0 17204 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_182
timestamp 1688980957
transform 1 0 17848 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_192
timestamp 1688980957
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_213
timestamp 1688980957
transform 1 0 20700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_225
timestamp 1688980957
transform 1 0 21804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_237
timestamp 1688980957
transform 1 0 22908 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_244
timestamp 1688980957
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_261
timestamp 1688980957
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_271
timestamp 1688980957
transform 1 0 26036 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_288
timestamp 1688980957
transform 1 0 27600 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_300
timestamp 1688980957
transform 1 0 28704 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_322
timestamp 1688980957
transform 1 0 30728 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_343
timestamp 1688980957
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_354
timestamp 1688980957
transform 1 0 33672 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_362
timestamp 1688980957
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1688980957
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 1688980957
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 1688980957
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_421
timestamp 1688980957
transform 1 0 39836 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_429
timestamp 1688980957
transform 1 0 40572 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_65
timestamp 1688980957
transform 1 0 7084 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_87
timestamp 1688980957
transform 1 0 9108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_91
timestamp 1688980957
transform 1 0 9476 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_136
timestamp 1688980957
transform 1 0 13616 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_148
timestamp 1688980957
transform 1 0 14720 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_175
timestamp 1688980957
transform 1 0 17204 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_187
timestamp 1688980957
transform 1 0 18308 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_195
timestamp 1688980957
transform 1 0 19044 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_210
timestamp 1688980957
transform 1 0 20424 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_222
timestamp 1688980957
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_237
timestamp 1688980957
transform 1 0 22908 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_246
timestamp 1688980957
transform 1 0 23736 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_258
timestamp 1688980957
transform 1 0 24840 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_270
timestamp 1688980957
transform 1 0 25944 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_278
timestamp 1688980957
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_289
timestamp 1688980957
transform 1 0 27692 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_300
timestamp 1688980957
transform 1 0 28704 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_311
timestamp 1688980957
transform 1 0 29716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_323
timestamp 1688980957
transform 1 0 30820 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_329
timestamp 1688980957
transform 1 0 31372 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_343
timestamp 1688980957
transform 1 0 32660 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_351
timestamp 1688980957
transform 1 0 33396 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_372
timestamp 1688980957
transform 1 0 35328 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_384
timestamp 1688980957
transform 1 0 36432 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1688980957
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 1688980957
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_429
timestamp 1688980957
transform 1 0 40572 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_136
timestamp 1688980957
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_163
timestamp 1688980957
transform 1 0 16100 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_171
timestamp 1688980957
transform 1 0 16836 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_180
timestamp 1688980957
transform 1 0 17664 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_188
timestamp 1688980957
transform 1 0 18400 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_209
timestamp 1688980957
transform 1 0 20332 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_224
timestamp 1688980957
transform 1 0 21712 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_236
timestamp 1688980957
transform 1 0 22816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_244
timestamp 1688980957
transform 1 0 23552 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_259
timestamp 1688980957
transform 1 0 24932 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_267
timestamp 1688980957
transform 1 0 25668 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_275
timestamp 1688980957
transform 1 0 26404 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_287
timestamp 1688980957
transform 1 0 27508 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_304
timestamp 1688980957
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_317
timestamp 1688980957
transform 1 0 30268 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_329
timestamp 1688980957
transform 1 0 31372 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_341
timestamp 1688980957
transform 1 0 32476 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_353
timestamp 1688980957
transform 1 0 33580 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_361
timestamp 1688980957
transform 1 0 34316 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1688980957
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1688980957
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1688980957
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 1688980957
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 1688980957
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 1688980957
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_433
timestamp 1688980957
transform 1 0 40940 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_91
timestamp 1688980957
transform 1 0 9476 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_101
timestamp 1688980957
transform 1 0 10396 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_109
timestamp 1688980957
transform 1 0 11132 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_146
timestamp 1688980957
transform 1 0 14536 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_158
timestamp 1688980957
transform 1 0 15640 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_166
timestamp 1688980957
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_194
timestamp 1688980957
transform 1 0 18952 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_207
timestamp 1688980957
transform 1 0 20148 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_238
timestamp 1688980957
transform 1 0 23000 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_247
timestamp 1688980957
transform 1 0 23828 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_270
timestamp 1688980957
transform 1 0 25944 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_281
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_296
timestamp 1688980957
transform 1 0 28336 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_315
timestamp 1688980957
transform 1 0 30084 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_322
timestamp 1688980957
transform 1 0 30728 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_348
timestamp 1688980957
transform 1 0 33120 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_352
timestamp 1688980957
transform 1 0 33488 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 1688980957
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 1688980957
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1688980957
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1688980957
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_429
timestamp 1688980957
transform 1 0 40572 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_91
timestamp 1688980957
transform 1 0 9476 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1688980957
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_164
timestamp 1688980957
transform 1 0 16192 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_176
timestamp 1688980957
transform 1 0 17296 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_187
timestamp 1688980957
transform 1 0 18308 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_207
timestamp 1688980957
transform 1 0 20148 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_219
timestamp 1688980957
transform 1 0 21252 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_231
timestamp 1688980957
transform 1 0 22356 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_243
timestamp 1688980957
transform 1 0 23460 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 1688980957
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_261
timestamp 1688980957
transform 1 0 25116 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_268
timestamp 1688980957
transform 1 0 25760 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_280
timestamp 1688980957
transform 1 0 26864 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_292
timestamp 1688980957
transform 1 0 27968 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 1688980957
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 1688980957
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_314
timestamp 1688980957
transform 1 0 29992 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_322
timestamp 1688980957
transform 1 0 30728 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_330
timestamp 1688980957
transform 1 0 31464 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_342
timestamp 1688980957
transform 1 0 32568 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_353
timestamp 1688980957
transform 1 0 33580 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_361
timestamp 1688980957
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1688980957
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1688980957
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_389
timestamp 1688980957
transform 1 0 36892 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_397
timestamp 1688980957
transform 1 0 37628 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 1688980957
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_433
timestamp 1688980957
transform 1 0 40940 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_77
timestamp 1688980957
transform 1 0 8188 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_87
timestamp 1688980957
transform 1 0 9108 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_102
timestamp 1688980957
transform 1 0 10488 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_110
timestamp 1688980957
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_134
timestamp 1688980957
transform 1 0 13432 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_140
timestamp 1688980957
transform 1 0 13984 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_148
timestamp 1688980957
transform 1 0 14720 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_164
timestamp 1688980957
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_208
timestamp 1688980957
transform 1 0 20240 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_220
timestamp 1688980957
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_232
timestamp 1688980957
transform 1 0 22448 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_244
timestamp 1688980957
transform 1 0 23552 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_253
timestamp 1688980957
transform 1 0 24380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_265
timestamp 1688980957
transform 1 0 25484 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_275
timestamp 1688980957
transform 1 0 26404 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1688980957
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_286
timestamp 1688980957
transform 1 0 27416 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_298
timestamp 1688980957
transform 1 0 28520 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_310
timestamp 1688980957
transform 1 0 29624 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_322
timestamp 1688980957
transform 1 0 30728 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_331
timestamp 1688980957
transform 1 0 31556 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 1688980957
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_337
timestamp 1688980957
transform 1 0 32108 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_348
timestamp 1688980957
transform 1 0 33120 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_360
timestamp 1688980957
transform 1 0 34224 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_372
timestamp 1688980957
transform 1 0 35328 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_384
timestamp 1688980957
transform 1 0 36432 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1688980957
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1688980957
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 1688980957
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_429
timestamp 1688980957
transform 1 0 40572 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_13
timestamp 1688980957
transform 1 0 2300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_25
timestamp 1688980957
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_93
timestamp 1688980957
transform 1 0 9660 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_102
timestamp 1688980957
transform 1 0 10488 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_128
timestamp 1688980957
transform 1 0 12880 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_138
timestamp 1688980957
transform 1 0 13800 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_151
timestamp 1688980957
transform 1 0 14996 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_174
timestamp 1688980957
transform 1 0 17112 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_178
timestamp 1688980957
transform 1 0 17480 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_187
timestamp 1688980957
transform 1 0 18308 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_204
timestamp 1688980957
transform 1 0 19872 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_212
timestamp 1688980957
transform 1 0 20608 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_220
timestamp 1688980957
transform 1 0 21344 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_242
timestamp 1688980957
transform 1 0 23368 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_260
timestamp 1688980957
transform 1 0 25024 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_265
timestamp 1688980957
transform 1 0 25484 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_275
timestamp 1688980957
transform 1 0 26404 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_287
timestamp 1688980957
transform 1 0 27508 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_295
timestamp 1688980957
transform 1 0 28244 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_304
timestamp 1688980957
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_316
timestamp 1688980957
transform 1 0 30176 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_322
timestamp 1688980957
transform 1 0 30728 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_334
timestamp 1688980957
transform 1 0 31832 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_343
timestamp 1688980957
transform 1 0 32660 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1688980957
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1688980957
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_389
timestamp 1688980957
transform 1 0 36892 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_417
timestamp 1688980957
transform 1 0 39468 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_429
timestamp 1688980957
transform 1 0 40572 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_87
timestamp 1688980957
transform 1 0 9108 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_108
timestamp 1688980957
transform 1 0 11040 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_121
timestamp 1688980957
transform 1 0 12236 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_131
timestamp 1688980957
transform 1 0 13156 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_152
timestamp 1688980957
transform 1 0 15088 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_207
timestamp 1688980957
transform 1 0 20148 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_222
timestamp 1688980957
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_231
timestamp 1688980957
transform 1 0 22356 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_247
timestamp 1688980957
transform 1 0 23828 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_256
timestamp 1688980957
transform 1 0 24656 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_273
timestamp 1688980957
transform 1 0 26220 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_313
timestamp 1688980957
transform 1 0 29900 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_327
timestamp 1688980957
transform 1 0 31188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 1688980957
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_343
timestamp 1688980957
transform 1 0 32660 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_355
timestamp 1688980957
transform 1 0 33764 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_367
timestamp 1688980957
transform 1 0 34868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_379
timestamp 1688980957
transform 1 0 35972 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 1688980957
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1688980957
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1688980957
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_417
timestamp 1688980957
transform 1 0 39468 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_425
timestamp 1688980957
transform 1 0 40204 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_107
timestamp 1688980957
transform 1 0 10948 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_129
timestamp 1688980957
transform 1 0 12972 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_175
timestamp 1688980957
transform 1 0 17204 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_183
timestamp 1688980957
transform 1 0 17940 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_208
timestamp 1688980957
transform 1 0 20240 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_215
timestamp 1688980957
transform 1 0 20884 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_239
timestamp 1688980957
transform 1 0 23092 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_245
timestamp 1688980957
transform 1 0 23644 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_262
timestamp 1688980957
transform 1 0 25208 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_270
timestamp 1688980957
transform 1 0 25944 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_283
timestamp 1688980957
transform 1 0 27140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_295
timestamp 1688980957
transform 1 0 28244 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_303
timestamp 1688980957
transform 1 0 28980 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 1688980957
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1688980957
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_341
timestamp 1688980957
transform 1 0 32476 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_362
timestamp 1688980957
transform 1 0 34408 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1688980957
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 1688980957
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 1688980957
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 1688980957
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 1688980957
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 1688980957
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 1688980957
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_433
timestamp 1688980957
transform 1 0 40940 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_9
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_21
timestamp 1688980957
transform 1 0 3036 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_29
timestamp 1688980957
transform 1 0 3772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_41
timestamp 1688980957
transform 1 0 4876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_53
timestamp 1688980957
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_65
timestamp 1688980957
transform 1 0 7084 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_70
timestamp 1688980957
transform 1 0 7544 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_82
timestamp 1688980957
transform 1 0 8648 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_85
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_97
timestamp 1688980957
transform 1 0 10028 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_116
timestamp 1688980957
transform 1 0 11776 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_128
timestamp 1688980957
transform 1 0 12880 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_141
timestamp 1688980957
transform 1 0 14076 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_145
timestamp 1688980957
transform 1 0 14444 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_156
timestamp 1688980957
transform 1 0 15456 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_193
timestamp 1688980957
transform 1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_203
timestamp 1688980957
transform 1 0 19780 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_215
timestamp 1688980957
transform 1 0 20884 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1688980957
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_225
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_233
timestamp 1688980957
transform 1 0 22540 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_238
timestamp 1688980957
transform 1 0 23000 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_250
timestamp 1688980957
transform 1 0 24104 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_253
timestamp 1688980957
transform 1 0 24380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_265
timestamp 1688980957
transform 1 0 25484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_277
timestamp 1688980957
transform 1 0 26588 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 1688980957
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 1688980957
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_305
timestamp 1688980957
transform 1 0 29164 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_309
timestamp 1688980957
transform 1 0 29532 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_317
timestamp 1688980957
transform 1 0 30268 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_324
timestamp 1688980957
transform 1 0 30912 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_337
timestamp 1688980957
transform 1 0 32108 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_351
timestamp 1688980957
transform 1 0 33396 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_363
timestamp 1688980957
transform 1 0 34500 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_371
timestamp 1688980957
transform 1 0 35236 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_383
timestamp 1688980957
transform 1 0 36340 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 1688980957
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_393
timestamp 1688980957
transform 1 0 37260 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_401
timestamp 1688980957
transform 1 0 37996 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_408
timestamp 1688980957
transform 1 0 38640 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_421
timestamp 1688980957
transform 1 0 39836 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_429
timestamp 1688980957
transform 1 0 40572 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32660 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 39836 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 13064 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 33396 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 14444 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 11684 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 12788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 6164 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 11500 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 10212 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 40388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 40388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 6440 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 24840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 9752 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 10580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 1932 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 4508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 15640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 20240 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 38272 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 27784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 20148 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 24104 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 16192 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 21620 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 18492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 6164 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 15916 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 35696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 9844 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 8188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 32844 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 38456 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 9108 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 39100 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 35512 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 7176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 5612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 21160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 3956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 25024 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 37352 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 36340 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 40848 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1688980957
transform 1 0 34684 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1688980957
transform 1 0 40572 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1688980957
transform 1 0 7176 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1688980957
transform 1 0 22632 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1688980957
transform 1 0 40756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1688980957
transform 1 0 3312 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 40848 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 11040 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1688980957
transform 1 0 15088 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  max_cap1
timestamp 1688980957
transform 1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap44
timestamp 1688980957
transform 1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  max_cap46
timestamp 1688980957
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap47
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap48
timestamp 1688980957
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  max_cap49
timestamp 1688980957
transform 1 0 17572 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap50
timestamp 1688980957
transform 1 0 17940 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap52
timestamp 1688980957
transform 1 0 16100 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap54
timestamp 1688980957
transform 1 0 8464 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap56
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output15
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1688980957
transform 1 0 38732 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 19228 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 15548 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform 1 0 40572 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform 1 0 40572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform 1 0 40572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1688980957
transform 1 0 40756 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform 1 0 31004 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1688980957
transform 1 0 40756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 38088 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 34868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform 1 0 30360 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 3956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform 1 0 11684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 40572 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 19412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output41
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 27140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform 1 0 40572 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 41400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 41400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 41400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 41400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 41400 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 41400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 41400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 41400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 41400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 41400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 41400 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 41400 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 41400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 41400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 41400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 41400 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 41400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 41400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 41400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 41400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 41400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 41400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 41400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 41400 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 41400 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 41400 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 41400 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 41400 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 41400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 41400 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 41400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 41400 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 41400 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 41400 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 41400 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 41400 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 41400 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 41400 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 41400 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 41400 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 41400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 41400 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 41400 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 41400 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 41400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 41400 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 41400 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 41400 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 41400 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 41400 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 41400 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 41400 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 41400 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 41400 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 41400 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 41400 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 41400 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 41400 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 41400 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 41400 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 41400 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 41400 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 41400 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 41400 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 41400 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 41400 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 41400 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 41400 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 41400 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 41400 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 41400 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 41400 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1688980957
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1688980957
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1688980957
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1688980957
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1688980957
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1688980957
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1688980957
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1688980957
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1688980957
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1688980957
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1688980957
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1688980957
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1688980957
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1688980957
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1688980957
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1688980957
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1688980957
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1688980957
transform 1 0 8832 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1688980957
transform 1 0 13984 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1688980957
transform 1 0 19136 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1688980957
transform 1 0 24288 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1688980957
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1688980957
transform 1 0 29440 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1688980957
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1688980957
transform 1 0 34592 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1688980957
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1688980957
transform 1 0 39744 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire2
timestamp 1688980957
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  wire45
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  wire51
timestamp 1688980957
transform 1 0 19504 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  wire53
timestamp 1688980957
transform 1 0 27232 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  wire55
timestamp 1688980957
transform 1 0 29440 0 -1 29376
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 M10ClkOut
port 0 nsew signal tristate
flabel metal4 s 19568 2128 19888 42480 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 42480 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 34928 2128 35248 42480 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 addressBusHigh[0]
port 3 nsew signal tristate
flabel metal2 s 18694 43864 18750 44664 0 FreeSans 224 90 0 0 addressBusHigh[1]
port 4 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 addressBusHigh[2]
port 5 nsew signal tristate
flabel metal3 s 41720 8168 42520 8288 0 FreeSans 480 0 0 0 addressBusHigh[3]
port 6 nsew signal tristate
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 addressBusHigh[4]
port 7 nsew signal tristate
flabel metal3 s 41720 4088 42520 4208 0 FreeSans 480 0 0 0 addressBusHigh[5]
port 8 nsew signal tristate
flabel metal3 s 41720 8 42520 128 0 FreeSans 480 0 0 0 addressBusHigh[6]
port 9 nsew signal tristate
flabel metal3 s 41720 32648 42520 32768 0 FreeSans 480 0 0 0 addressBusHigh[7]
port 10 nsew signal tristate
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 addressBusLow[0]
port 11 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 addressBusLow[1]
port 12 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 addressBusLow[2]
port 13 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 addressBusLow[3]
port 14 nsew signal tristate
flabel metal3 s 41720 36728 42520 36848 0 FreeSans 480 0 0 0 addressBusLow[4]
port 15 nsew signal tristate
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 addressBusLow[5]
port 16 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 addressBusLow[6]
port 17 nsew signal tristate
flabel metal2 s 38014 43864 38070 44664 0 FreeSans 224 90 0 0 addressBusLow[7]
port 18 nsew signal tristate
flabel metal2 s 26422 43864 26478 44664 0 FreeSans 224 90 0 0 clk
port 19 nsew signal input
flabel metal3 s 41720 24488 42520 24608 0 FreeSans 480 0 0 0 dataBusEnable
port 20 nsew signal input
flabel metal2 s 34150 43864 34206 44664 0 FreeSans 224 90 0 0 dataBusInput[0]
port 21 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 dataBusInput[1]
port 22 nsew signal input
flabel metal3 s 41720 40808 42520 40928 0 FreeSans 480 0 0 0 dataBusInput[2]
port 23 nsew signal input
flabel metal2 s 7102 43864 7158 44664 0 FreeSans 224 90 0 0 dataBusInput[3]
port 24 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 dataBusInput[4]
port 25 nsew signal input
flabel metal2 s 22558 43864 22614 44664 0 FreeSans 224 90 0 0 dataBusInput[5]
port 26 nsew signal input
flabel metal3 s 41720 28568 42520 28688 0 FreeSans 480 0 0 0 dataBusInput[6]
port 27 nsew signal input
flabel metal2 s 3238 43864 3294 44664 0 FreeSans 224 90 0 0 dataBusInput[7]
port 28 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 dataBusOutput[0]
port 29 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 dataBusOutput[1]
port 30 nsew signal tristate
flabel metal2 s 30286 43864 30342 44664 0 FreeSans 224 90 0 0 dataBusOutput[2]
port 31 nsew signal tristate
flabel metal3 s 41720 12248 42520 12368 0 FreeSans 480 0 0 0 dataBusOutput[3]
port 32 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 dataBusOutput[4]
port 33 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 dataBusOutput[5]
port 34 nsew signal tristate
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 dataBusOutput[6]
port 35 nsew signal tristate
flabel metal3 s 41720 16328 42520 16448 0 FreeSans 480 0 0 0 dataBusOutput[7]
port 36 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 dataBusSelect
port 37 nsew signal tristate
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 functionalClockOut
port 38 nsew signal tristate
flabel metal2 s 41878 43864 41934 44664 0 FreeSans 224 90 0 0 interruptRequest
port 39 nsew signal input
flabel metal2 s 10966 43864 11022 44664 0 FreeSans 224 90 0 0 nonMaskableInterrupt
port 40 nsew signal input
flabel metal2 s 14830 43864 14886 44664 0 FreeSans 224 90 0 0 nrst
port 41 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 readNotWrite
port 42 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 ready
port 43 nsew signal input
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 setOverflow
port 44 nsew signal input
flabel metal3 s 41720 20408 42520 20528 0 FreeSans 480 0 0 0 sync
port 45 nsew signal tristate
rlabel metal1 21252 42432 21252 42432 0 VGND
rlabel metal1 21252 41888 21252 41888 0 VPWR
rlabel metal3 820 15708 820 15708 0 M10ClkOut
rlabel metal1 11316 41242 11316 41242 0 _0000_
rlabel metal2 11546 37604 11546 37604 0 _0001_
rlabel metal1 8142 38998 8142 38998 0 _0002_
rlabel metal1 9154 36686 9154 36686 0 _0003_
rlabel metal1 9423 36346 9423 36346 0 _0004_
rlabel metal1 13018 39032 13018 39032 0 _0005_
rlabel metal1 10166 39066 10166 39066 0 _0006_
rlabel metal1 7958 37434 7958 37434 0 _0007_
rlabel metal1 9752 40698 9752 40698 0 _0008_
rlabel metal2 11822 38114 11822 38114 0 _0009_
rlabel metal2 12558 37094 12558 37094 0 _0010_
rlabel metal1 12788 40154 12788 40154 0 _0011_
rlabel metal1 13892 41514 13892 41514 0 _0012_
rlabel metal1 6164 33082 6164 33082 0 _0013_
rlabel metal1 5658 30566 5658 30566 0 _0014_
rlabel metal1 5740 28730 5740 28730 0 _0015_
rlabel metal2 6210 32164 6210 32164 0 _0016_
rlabel metal1 6440 31382 6440 31382 0 _0017_
rlabel metal1 5191 28934 5191 28934 0 _0018_
rlabel metal1 6670 27064 6670 27064 0 _0019_
rlabel metal1 33764 37910 33764 37910 0 _0020_
rlabel metal1 32982 40154 32982 40154 0 _0021_
rlabel metal1 33580 38862 33580 38862 0 _0022_
rlabel metal1 34086 36856 34086 36856 0 _0023_
rlabel metal1 32512 35258 32512 35258 0 _0024_
rlabel metal1 33442 35598 33442 35598 0 _0025_
rlabel via1 15035 12614 15035 12614 0 _0026_
rlabel metal1 18814 3706 18814 3706 0 _0027_
rlabel metal1 23230 5304 23230 5304 0 _0028_
rlabel metal1 14996 5746 14996 5746 0 _0029_
rlabel metal1 16974 4250 16974 4250 0 _0030_
rlabel metal1 14122 9146 14122 9146 0 _0031_
rlabel metal1 17342 5882 17342 5882 0 _0032_
rlabel metal1 23828 3094 23828 3094 0 _0033_
rlabel metal2 12466 14756 12466 14756 0 _0034_
rlabel metal1 9890 7480 9890 7480 0 _0035_
rlabel via1 5559 6970 5559 6970 0 _0036_
rlabel metal2 8050 7582 8050 7582 0 _0037_
rlabel metal1 4508 11866 4508 11866 0 _0038_
rlabel metal1 2990 14008 2990 14008 0 _0039_
rlabel metal1 4646 15606 4646 15606 0 _0040_
rlabel metal1 4370 7922 4370 7922 0 _0041_
rlabel metal1 2208 17850 2208 17850 0 _0042_
rlabel metal1 10757 5882 10757 5882 0 _0043_
rlabel metal1 2116 11798 2116 11798 0 _0044_
rlabel metal1 29578 6392 29578 6392 0 _0045_
rlabel metal1 35834 29546 35834 29546 0 _0046_
rlabel metal1 4876 23290 4876 23290 0 _0047_
rlabel metal1 7728 5882 7728 5882 0 _0048_
rlabel metal1 36938 23834 36938 23834 0 _0049_
rlabel metal1 21160 9010 21160 9010 0 _0050_
rlabel metal1 22402 3162 22402 3162 0 _0051_
rlabel metal1 25070 5270 25070 5270 0 _0052_
rlabel metal2 27002 6562 27002 6562 0 _0053_
rlabel metal1 20470 2618 20470 2618 0 _0054_
rlabel metal1 27692 8874 27692 8874 0 _0055_
rlabel metal1 22402 8534 22402 8534 0 _0056_
rlabel metal1 26588 4250 26588 4250 0 _0057_
rlabel metal1 30084 18394 30084 18394 0 _0058_
rlabel metal1 32660 20570 32660 20570 0 _0059_
rlabel metal1 29762 14450 29762 14450 0 _0060_
rlabel metal2 28566 11934 28566 11934 0 _0061_
rlabel metal1 33304 12886 33304 12886 0 _0062_
rlabel metal1 36386 14450 36386 14450 0 _0063_
rlabel metal1 33902 20026 33902 20026 0 _0064_
rlabel metal1 37766 22202 37766 22202 0 _0065_
rlabel metal1 37536 4182 37536 4182 0 _0066_
rlabel metal1 34592 22746 34592 22746 0 _0067_
rlabel metal1 16974 3128 16974 3128 0 _0068_
rlabel metal2 39146 7514 39146 7514 0 _0069_
rlabel metal1 4048 27098 4048 27098 0 _0070_
rlabel metal1 34546 5134 34546 5134 0 _0071_
rlabel metal1 37582 6392 37582 6392 0 _0072_
rlabel metal1 37398 28458 37398 28458 0 _0073_
rlabel metal1 32752 25194 32752 25194 0 _0074_
rlabel metal1 18262 8568 18262 8568 0 _0075_
rlabel metal1 20010 2958 20010 2958 0 _0076_
rlabel metal1 22678 5882 22678 5882 0 _0077_
rlabel metal1 27646 6392 27646 6392 0 _0078_
rlabel metal1 20240 5338 20240 5338 0 _0079_
rlabel metal1 27324 8398 27324 8398 0 _0080_
rlabel metal2 18906 6426 18906 6426 0 _0081_
rlabel metal1 25576 3570 25576 3570 0 _0082_
rlabel metal1 14122 15402 14122 15402 0 _0083_
rlabel metal1 14168 3706 14168 3706 0 _0084_
rlabel metal1 12558 4794 12558 4794 0 _0085_
rlabel metal1 12696 6426 12696 6426 0 _0086_
rlabel metal1 15180 3094 15180 3094 0 _0087_
rlabel metal1 13570 10744 13570 10744 0 _0088_
rlabel metal1 12512 8058 12512 8058 0 _0089_
rlabel metal1 12972 3094 12972 3094 0 _0090_
rlabel metal1 38502 20026 38502 20026 0 _0091_
rlabel metal1 39514 18360 39514 18360 0 _0092_
rlabel metal2 39330 14110 39330 14110 0 _0093_
rlabel metal1 38456 11662 38456 11662 0 _0094_
rlabel metal1 37582 8568 37582 8568 0 _0095_
rlabel metal1 35236 7310 35236 7310 0 _0096_
rlabel metal1 32108 7786 32108 7786 0 _0097_
rlabel metal1 29072 9622 29072 9622 0 _0098_
rlabel metal2 5658 5474 5658 5474 0 _0099_
rlabel metal2 31878 5474 31878 5474 0 _0100_
rlabel metal2 30682 23426 30682 23426 0 _0101_
rlabel metal1 39560 12410 39560 12410 0 _0102_
rlabel metal1 3542 5304 3542 5304 0 _0103_
rlabel metal1 10941 4794 10941 4794 0 _0104_
rlabel metal1 3910 24922 3910 24922 0 _0105_
rlabel metal1 39606 16184 39606 16184 0 _0106_
rlabel metal1 35604 25330 35604 25330 0 _0107_
rlabel metal1 35321 27642 35321 27642 0 _0108_
rlabel metal1 33672 25942 33672 25942 0 _0109_
rlabel metal1 4738 25976 4738 25976 0 _0110_
rlabel metal1 33810 26894 33810 26894 0 _0111_
rlabel metal1 32154 23630 32154 23630 0 _0112_
rlabel metal1 6854 23630 6854 23630 0 _0113_
rlabel metal1 9798 21862 9798 21862 0 _0114_
rlabel metal2 6762 35428 6762 35428 0 _0115_
rlabel metal1 9614 21454 9614 21454 0 _0116_
rlabel metal1 27554 18666 27554 18666 0 _0117_
rlabel metal1 13478 19822 13478 19822 0 _0118_
rlabel metal1 15778 18292 15778 18292 0 _0119_
rlabel metal1 14996 19414 14996 19414 0 _0120_
rlabel metal2 15594 17986 15594 17986 0 _0121_
rlabel metal1 17250 16660 17250 16660 0 _0122_
rlabel metal1 15824 14382 15824 14382 0 _0123_
rlabel metal1 13800 19958 13800 19958 0 _0124_
rlabel metal1 15686 16082 15686 16082 0 _0125_
rlabel metal1 17434 9418 17434 9418 0 _0126_
rlabel metal1 15134 17204 15134 17204 0 _0127_
rlabel metal1 17618 15504 17618 15504 0 _0128_
rlabel metal2 20746 16337 20746 16337 0 _0129_
rlabel metal1 10350 6358 10350 6358 0 _0130_
rlabel metal1 11362 17612 11362 17612 0 _0131_
rlabel metal1 9430 17272 9430 17272 0 _0132_
rlabel metal1 8970 16524 8970 16524 0 _0133_
rlabel metal1 5198 19482 5198 19482 0 _0134_
rlabel metal1 8786 17102 8786 17102 0 _0135_
rlabel metal1 8556 16558 8556 16558 0 _0136_
rlabel metal2 26358 9146 26358 9146 0 _0137_
rlabel metal1 16238 10030 16238 10030 0 _0138_
rlabel metal2 21482 9792 21482 9792 0 _0139_
rlabel metal1 26588 10030 26588 10030 0 _0140_
rlabel metal1 25668 13158 25668 13158 0 _0141_
rlabel metal1 26404 10234 26404 10234 0 _0142_
rlabel metal1 27186 13328 27186 13328 0 _0143_
rlabel metal1 27278 13260 27278 13260 0 _0144_
rlabel metal1 26680 11050 26680 11050 0 _0145_
rlabel metal2 10902 11526 10902 11526 0 _0146_
rlabel metal1 10028 11526 10028 11526 0 _0147_
rlabel metal1 21896 12070 21896 12070 0 _0148_
rlabel metal1 18538 12920 18538 12920 0 _0149_
rlabel metal1 12006 13498 12006 13498 0 _0150_
rlabel via1 16261 14382 16261 14382 0 _0151_
rlabel metal1 17894 14280 17894 14280 0 _0152_
rlabel metal2 15594 15419 15594 15419 0 _0153_
rlabel metal1 11500 16082 11500 16082 0 _0154_
rlabel metal1 8970 14280 8970 14280 0 _0155_
rlabel metal1 8188 14926 8188 14926 0 _0156_
rlabel metal1 8832 14926 8832 14926 0 _0157_
rlabel metal2 8050 14586 8050 14586 0 _0158_
rlabel metal1 21528 7514 21528 7514 0 _0159_
rlabel metal1 17526 7378 17526 7378 0 _0160_
rlabel metal1 19458 7514 19458 7514 0 _0161_
rlabel metal1 21022 11050 21022 11050 0 _0162_
rlabel metal1 21390 12206 21390 12206 0 _0163_
rlabel metal1 22310 11628 22310 11628 0 _0164_
rlabel metal1 27738 25466 27738 25466 0 _0165_
rlabel metal1 27646 14314 27646 14314 0 _0166_
rlabel metal2 22770 13991 22770 13991 0 _0167_
rlabel metal1 23046 13294 23046 13294 0 _0168_
rlabel metal1 22264 11866 22264 11866 0 _0169_
rlabel via1 21937 11866 21937 11866 0 _0170_
rlabel metal1 10488 12818 10488 12818 0 _0171_
rlabel metal2 4922 7514 4922 7514 0 _0172_
rlabel metal1 12834 12954 12834 12954 0 _0173_
rlabel metal1 17388 14586 17388 14586 0 _0174_
rlabel metal2 17066 14501 17066 14501 0 _0175_
rlabel metal1 18170 15028 18170 15028 0 _0176_
rlabel metal1 17434 14858 17434 14858 0 _0177_
rlabel metal1 11178 12886 11178 12886 0 _0178_
rlabel metal1 8510 12784 8510 12784 0 _0179_
rlabel metal1 9982 12648 9982 12648 0 _0180_
rlabel metal1 7866 12750 7866 12750 0 _0181_
rlabel metal1 6670 13158 6670 13158 0 _0182_
rlabel metal1 28014 13702 28014 13702 0 _0183_
rlabel metal1 27186 13906 27186 13906 0 _0184_
rlabel metal1 27186 13702 27186 13702 0 _0185_
rlabel metal1 24426 12206 24426 12206 0 _0186_
rlabel metal2 23690 14076 23690 14076 0 _0187_
rlabel metal1 26036 7514 26036 7514 0 _0188_
rlabel metal1 16514 7378 16514 7378 0 _0189_
rlabel metal1 17894 7174 17894 7174 0 _0190_
rlabel metal1 24840 8058 24840 8058 0 _0191_
rlabel metal1 24794 12886 24794 12886 0 _0192_
rlabel metal2 23966 12444 23966 12444 0 _0193_
rlabel metal1 11822 11696 11822 11696 0 _0194_
rlabel metal2 9154 10880 9154 10880 0 _0195_
rlabel metal1 20056 12342 20056 12342 0 _0196_
rlabel metal1 12650 12138 12650 12138 0 _0197_
rlabel metal2 15594 13163 15594 13163 0 _0198_
rlabel metal1 15732 13770 15732 13770 0 _0199_
rlabel metal1 29670 16694 29670 16694 0 _0200_
rlabel metal1 9614 11764 9614 11764 0 _0201_
rlabel metal1 6578 11764 6578 11764 0 _0202_
rlabel metal1 8832 11594 8832 11594 0 _0203_
rlabel metal1 6440 11866 6440 11866 0 _0204_
rlabel metal1 27600 14518 27600 14518 0 _0205_
rlabel metal1 27462 14586 27462 14586 0 _0206_
rlabel metal2 27002 12988 27002 12988 0 _0207_
rlabel metal1 25208 11730 25208 11730 0 _0208_
rlabel metal1 24886 7480 24886 7480 0 _0209_
rlabel metal2 25346 7344 25346 7344 0 _0210_
rlabel metal1 21666 7990 21666 7990 0 _0211_
rlabel metal2 26082 9350 26082 9350 0 _0212_
rlabel metal1 26450 11696 26450 11696 0 _0213_
rlabel metal1 26404 10778 26404 10778 0 _0214_
rlabel metal1 13478 5610 13478 5610 0 _0215_
rlabel metal2 11362 10234 11362 10234 0 _0216_
rlabel metal1 28934 19346 28934 19346 0 _0217_
rlabel metal1 11914 11832 11914 11832 0 _0218_
rlabel metal2 17296 15878 17296 15878 0 _0219_
rlabel metal1 17342 8364 17342 8364 0 _0220_
rlabel metal1 2622 12308 2622 12308 0 _0221_
rlabel metal2 9614 10132 9614 10132 0 _0222_
rlabel metal1 8280 9894 8280 9894 0 _0223_
rlabel metal1 19734 9622 19734 9622 0 _0224_
rlabel metal1 19688 11118 19688 11118 0 _0225_
rlabel metal1 20838 9554 20838 9554 0 _0226_
rlabel metal2 19642 11356 19642 11356 0 _0227_
rlabel metal1 19734 12274 19734 12274 0 _0228_
rlabel metal1 16238 13328 16238 13328 0 _0229_
rlabel metal1 20102 12852 20102 12852 0 _0230_
rlabel metal1 21298 13430 21298 13430 0 _0231_
rlabel metal1 22586 17850 22586 17850 0 _0232_
rlabel metal1 23138 18122 23138 18122 0 _0233_
rlabel metal1 21648 15470 21648 15470 0 _0234_
rlabel metal2 20194 14178 20194 14178 0 _0235_
rlabel metal1 20746 13328 20746 13328 0 _0236_
rlabel metal1 12489 16422 12489 16422 0 _0237_
rlabel metal1 18768 17646 18768 17646 0 _0238_
rlabel metal1 17618 15130 17618 15130 0 _0239_
rlabel metal1 18262 17680 18262 17680 0 _0240_
rlabel metal1 4646 17748 4646 17748 0 _0241_
rlabel metal1 12144 16218 12144 16218 0 _0242_
rlabel metal1 12190 16014 12190 16014 0 _0243_
rlabel metal1 20240 12954 20240 12954 0 _0244_
rlabel via2 20930 16099 20930 16099 0 _0245_
rlabel metal1 20700 16422 20700 16422 0 _0246_
rlabel metal1 21068 16490 21068 16490 0 _0247_
rlabel metal1 20378 14994 20378 14994 0 _0248_
rlabel metal1 19642 14858 19642 14858 0 _0249_
rlabel metal1 12466 16592 12466 16592 0 _0250_
rlabel metal2 10810 16116 10810 16116 0 _0251_
rlabel via1 8676 24786 8676 24786 0 _0252_
rlabel metal2 9154 24038 9154 24038 0 _0253_
rlabel metal2 13294 24378 13294 24378 0 _0254_
rlabel metal2 12006 23868 12006 23868 0 _0255_
rlabel via3 25829 33252 25829 33252 0 _0256_
rlabel metal1 24380 24174 24380 24174 0 _0257_
rlabel metal1 12190 23800 12190 23800 0 _0258_
rlabel metal1 9798 19380 9798 19380 0 _0259_
rlabel metal1 11684 16558 11684 16558 0 _0260_
rlabel metal1 11270 15028 11270 15028 0 _0261_
rlabel metal1 10304 10778 10304 10778 0 _0262_
rlabel metal1 24104 18122 24104 18122 0 _0263_
rlabel metal1 23690 18258 23690 18258 0 _0264_
rlabel metal1 22586 15436 22586 15436 0 _0265_
rlabel metal1 22218 14382 22218 14382 0 _0266_
rlabel metal2 22586 7174 22586 7174 0 _0267_
rlabel metal2 21390 6528 21390 6528 0 _0268_
rlabel metal1 16974 7378 16974 7378 0 _0269_
rlabel metal1 22862 13192 22862 13192 0 _0270_
rlabel metal1 23138 13838 23138 13838 0 _0271_
rlabel metal1 22816 16082 22816 16082 0 _0272_
rlabel metal2 22586 14824 22586 14824 0 _0273_
rlabel metal2 16054 13566 16054 13566 0 _0274_
rlabel metal1 12098 10030 12098 10030 0 _0275_
rlabel metal2 13662 11713 13662 11713 0 _0276_
rlabel metal1 12466 11220 12466 11220 0 _0277_
rlabel metal1 15824 16218 15824 16218 0 _0278_
rlabel metal1 16238 16490 16238 16490 0 _0279_
rlabel metal1 16008 16558 16008 16558 0 _0280_
rlabel metal1 11178 6800 11178 6800 0 _0281_
rlabel metal2 12098 10744 12098 10744 0 _0282_
rlabel via1 11160 10030 11160 10030 0 _0283_
rlabel metal1 10534 10608 10534 10608 0 _0284_
rlabel metal1 8050 10098 8050 10098 0 _0285_
rlabel viali 8234 10030 8234 10030 0 _0286_
rlabel metal1 6348 11730 6348 11730 0 _0287_
rlabel metal1 5842 11084 5842 11084 0 _0288_
rlabel metal1 7314 14280 7314 14280 0 _0289_
rlabel metal1 6808 14314 6808 14314 0 _0290_
rlabel metal2 7498 15606 7498 15606 0 _0291_
rlabel metal1 7268 18258 7268 18258 0 _0292_
rlabel metal1 25438 7412 25438 7412 0 _0293_
rlabel metal1 19274 7208 19274 7208 0 _0294_
rlabel metal2 24978 7990 24978 7990 0 _0295_
rlabel metal1 25392 8534 25392 8534 0 _0296_
rlabel metal1 25346 17204 25346 17204 0 _0297_
rlabel metal1 24794 17136 24794 17136 0 _0298_
rlabel metal1 25622 16660 25622 16660 0 _0299_
rlabel metal1 25898 16116 25898 16116 0 _0300_
rlabel metal1 26312 15946 26312 15946 0 _0301_
rlabel metal1 27002 18224 27002 18224 0 _0302_
rlabel metal1 27186 17680 27186 17680 0 _0303_
rlabel metal1 26680 16082 26680 16082 0 _0304_
rlabel metal1 19642 2890 19642 2890 0 _0305_
rlabel metal1 9568 18666 9568 18666 0 _0306_
rlabel metal1 26542 16218 26542 16218 0 _0307_
rlabel metal1 13478 17748 13478 17748 0 _0308_
rlabel metal1 12650 17850 12650 17850 0 _0309_
rlabel metal1 14904 16966 14904 16966 0 _0310_
rlabel metal1 15824 17034 15824 17034 0 _0311_
rlabel metal1 22080 17816 22080 17816 0 _0312_
rlabel metal1 12190 18326 12190 18326 0 _0313_
rlabel metal1 11040 18734 11040 18734 0 _0314_
rlabel metal1 9246 18802 9246 18802 0 _0315_
rlabel metal1 6624 20910 6624 20910 0 _0316_
rlabel metal1 7866 19822 7866 19822 0 _0317_
rlabel metal1 7038 19890 7038 19890 0 _0318_
rlabel metal3 18147 22100 18147 22100 0 _0319_
rlabel metal1 7820 20910 7820 20910 0 _0320_
rlabel metal1 4554 11696 4554 11696 0 _0321_
rlabel metal1 7038 25330 7038 25330 0 _0322_
rlabel metal2 21574 29682 21574 29682 0 _0323_
rlabel metal1 28474 24242 28474 24242 0 _0324_
rlabel metal1 5382 20400 5382 20400 0 _0325_
rlabel metal1 26772 24038 26772 24038 0 _0326_
rlabel metal1 27002 24174 27002 24174 0 _0327_
rlabel metal1 26956 23834 26956 23834 0 _0328_
rlabel metal1 27462 23494 27462 23494 0 _0329_
rlabel metal2 6854 25313 6854 25313 0 _0330_
rlabel metal2 6486 21529 6486 21529 0 _0331_
rlabel metal2 23874 22321 23874 22321 0 _0332_
rlabel via1 26151 21522 26151 21522 0 _0333_
rlabel via1 28750 25262 28750 25262 0 _0334_
rlabel metal1 28980 21590 28980 21590 0 _0335_
rlabel metal1 28934 20842 28934 20842 0 _0336_
rlabel metal1 29670 21114 29670 21114 0 _0337_
rlabel metal1 29670 30566 29670 30566 0 _0338_
rlabel metal1 28842 20910 28842 20910 0 _0339_
rlabel metal1 30314 25296 30314 25296 0 _0340_
rlabel metal1 30084 25126 30084 25126 0 _0341_
rlabel metal2 28842 23834 28842 23834 0 _0342_
rlabel metal1 29854 22644 29854 22644 0 _0343_
rlabel metal1 21206 12716 21206 12716 0 _0344_
rlabel metal1 26082 25738 26082 25738 0 _0345_
rlabel metal1 25576 25262 25576 25262 0 _0346_
rlabel metal1 25714 23562 25714 23562 0 _0347_
rlabel metal1 25208 19414 25208 19414 0 _0348_
rlabel metal1 25806 19482 25806 19482 0 _0349_
rlabel metal1 26542 20468 26542 20468 0 _0350_
rlabel metal1 25714 19890 25714 19890 0 _0351_
rlabel metal2 25898 21284 25898 21284 0 _0352_
rlabel metal2 15134 22525 15134 22525 0 _0353_
rlabel metal1 14996 22610 14996 22610 0 _0354_
rlabel metal1 17618 24310 17618 24310 0 _0355_
rlabel metal2 15962 24480 15962 24480 0 _0356_
rlabel metal1 16054 23834 16054 23834 0 _0357_
rlabel metal2 14858 23358 14858 23358 0 _0358_
rlabel metal1 14168 21862 14168 21862 0 _0359_
rlabel metal2 13202 22304 13202 22304 0 _0360_
rlabel metal1 6486 12206 6486 12206 0 _0361_
rlabel metal1 6915 19346 6915 19346 0 _0362_
rlabel metal1 21758 29580 21758 29580 0 _0363_
rlabel metal3 16836 27336 16836 27336 0 _0364_
rlabel metal1 8602 19482 8602 19482 0 _0365_
rlabel metal1 5198 11526 5198 11526 0 _0366_
rlabel metal2 4646 8738 4646 8738 0 _0367_
rlabel metal1 5658 10132 5658 10132 0 _0368_
rlabel metal1 5252 11798 5252 11798 0 _0369_
rlabel metal2 4922 12172 4922 12172 0 _0370_
rlabel metal1 5566 14926 5566 14926 0 _0371_
rlabel metal1 5290 19142 5290 19142 0 _0372_
rlabel metal2 5290 16354 5290 16354 0 _0373_
rlabel metal2 5842 14790 5842 14790 0 _0374_
rlabel viali 5565 16536 5565 16536 0 _0375_
rlabel metal1 4416 16558 4416 16558 0 _0376_
rlabel metal1 8786 18734 8786 18734 0 _0377_
rlabel metal1 5014 19380 5014 19380 0 _0378_
rlabel metal1 5520 18054 5520 18054 0 _0379_
rlabel metal1 5620 18326 5620 18326 0 _0380_
rlabel metal1 5934 18394 5934 18394 0 _0381_
rlabel metal1 6256 12206 6256 12206 0 _0382_
rlabel metal1 6164 19346 6164 19346 0 _0383_
rlabel metal1 6992 19210 6992 19210 0 _0384_
rlabel metal1 7590 21454 7590 21454 0 _0385_
rlabel metal2 28290 21488 28290 21488 0 _0386_
rlabel metal1 28842 22134 28842 22134 0 _0387_
rlabel metal1 27922 21862 27922 21862 0 _0388_
rlabel metal1 16146 12138 16146 12138 0 _0389_
rlabel metal3 28221 32300 28221 32300 0 _0390_
rlabel metal1 27278 23120 27278 23120 0 _0391_
rlabel metal2 16146 10880 16146 10880 0 _0392_
rlabel metal1 15272 12206 15272 12206 0 _0393_
rlabel metal1 19182 3502 19182 3502 0 _0394_
rlabel metal1 24242 5678 24242 5678 0 _0395_
rlabel metal1 15410 6290 15410 6290 0 _0396_
rlabel metal1 17296 4114 17296 4114 0 _0397_
rlabel metal1 14996 8942 14996 8942 0 _0398_
rlabel metal1 17802 5712 17802 5712 0 _0399_
rlabel metal1 24288 3706 24288 3706 0 _0400_
rlabel metal1 18400 29002 18400 29002 0 _0401_
rlabel metal1 14858 21522 14858 21522 0 _0402_
rlabel metal1 14122 15606 14122 15606 0 _0403_
rlabel metal1 10580 15334 10580 15334 0 _0404_
rlabel metal1 11546 14280 11546 14280 0 _0405_
rlabel metal1 9062 8432 9062 8432 0 _0406_
rlabel metal2 8602 18938 8602 18938 0 _0407_
rlabel metal1 8970 10710 8970 10710 0 _0408_
rlabel metal1 11178 18258 11178 18258 0 _0409_
rlabel metal2 8464 9962 8464 9962 0 _0410_
rlabel metal1 11040 14586 11040 14586 0 _0411_
rlabel metal2 8418 11815 8418 11815 0 _0412_
rlabel metal1 11086 14994 11086 14994 0 _0413_
rlabel metal1 11270 14450 11270 14450 0 _0414_
rlabel metal1 10994 10064 10994 10064 0 _0415_
rlabel metal1 10994 8976 10994 8976 0 _0416_
rlabel metal2 10258 8330 10258 8330 0 _0417_
rlabel metal1 6348 8942 6348 8942 0 _0418_
rlabel metal1 7130 8432 7130 8432 0 _0419_
rlabel metal2 10074 8092 10074 8092 0 _0420_
rlabel metal2 8602 9894 8602 9894 0 _0421_
rlabel metal1 8556 10506 8556 10506 0 _0422_
rlabel metal1 8602 10234 8602 10234 0 _0423_
rlabel metal2 8050 10030 8050 10030 0 _0424_
rlabel metal1 5152 9622 5152 9622 0 _0425_
rlabel metal1 4876 9146 4876 9146 0 _0426_
rlabel metal1 4508 9554 4508 9554 0 _0427_
rlabel metal1 5244 9486 5244 9486 0 _0428_
rlabel metal1 5842 9486 5842 9486 0 _0429_
rlabel metal1 6256 7854 6256 7854 0 _0430_
rlabel metal1 5750 7446 5750 7446 0 _0431_
rlabel metal1 4186 9520 4186 9520 0 _0432_
rlabel metal1 6670 8976 6670 8976 0 _0433_
rlabel metal2 6762 9554 6762 9554 0 _0434_
rlabel metal1 6670 9996 6670 9996 0 _0435_
rlabel metal2 7682 8296 7682 8296 0 _0436_
rlabel metal1 9430 12410 9430 12410 0 _0437_
rlabel metal1 8924 11730 8924 11730 0 _0438_
rlabel metal1 8418 11866 8418 11866 0 _0439_
rlabel metal1 8648 7854 8648 7854 0 _0440_
rlabel metal1 5152 11594 5152 11594 0 _0441_
rlabel metal1 6716 12886 6716 12886 0 _0442_
rlabel metal1 6532 12410 6532 12410 0 _0443_
rlabel metal2 8418 14892 8418 14892 0 _0444_
rlabel metal1 8096 12818 8096 12818 0 _0445_
rlabel metal1 8234 12852 8234 12852 0 _0446_
rlabel metal1 6394 12920 6394 12920 0 _0447_
rlabel metal2 6348 12274 6348 12274 0 _0448_
rlabel metal1 5014 11798 5014 11798 0 _0449_
rlabel metal2 4140 16082 4140 16082 0 _0450_
rlabel metal2 3450 15776 3450 15776 0 _0451_
rlabel metal1 6762 14450 6762 14450 0 _0452_
rlabel via1 7051 14314 7051 14314 0 _0453_
rlabel metal1 8326 14416 8326 14416 0 _0454_
rlabel metal1 7498 14382 7498 14382 0 _0455_
rlabel metal1 4186 14450 4186 14450 0 _0456_
rlabel metal1 3818 14450 3818 14450 0 _0457_
rlabel metal1 7222 16048 7222 16048 0 _0458_
rlabel metal1 6946 15912 6946 15912 0 _0459_
rlabel metal1 8188 16694 8188 16694 0 _0460_
rlabel metal1 8372 16626 8372 16626 0 _0461_
rlabel metal2 8142 16762 8142 16762 0 _0462_
rlabel metal1 6762 16116 6762 16116 0 _0463_
rlabel metal1 4922 15504 4922 15504 0 _0464_
rlabel metal1 4830 19346 4830 19346 0 _0465_
rlabel metal1 4876 19278 4876 19278 0 _0466_
rlabel metal1 4738 19482 4738 19482 0 _0467_
rlabel metal1 4186 16524 4186 16524 0 _0468_
rlabel metal1 4278 16592 4278 16592 0 _0469_
rlabel metal2 4554 16218 4554 16218 0 _0470_
rlabel metal1 4278 16116 4278 16116 0 _0471_
rlabel metal1 4784 15470 4784 15470 0 _0472_
rlabel metal1 5198 17306 5198 17306 0 _0473_
rlabel metal1 5109 18802 5109 18802 0 _0474_
rlabel metal1 4508 18666 4508 18666 0 _0475_
rlabel metal1 7590 18394 7590 18394 0 _0476_
rlabel metal1 6992 18666 6992 18666 0 _0477_
rlabel metal1 8786 19380 8786 19380 0 _0478_
rlabel metal1 8970 19210 8970 19210 0 _0479_
rlabel metal1 7728 18734 7728 18734 0 _0480_
rlabel via2 4370 18717 4370 18717 0 _0481_
rlabel metal1 3864 8602 3864 8602 0 _0482_
rlabel metal2 14858 28515 14858 28515 0 _0483_
rlabel metal2 15962 32096 15962 32096 0 _0484_
rlabel metal1 16238 31858 16238 31858 0 _0485_
rlabel metal1 15916 32538 15916 32538 0 _0486_
rlabel metal2 15686 32266 15686 32266 0 _0487_
rlabel via1 15318 29750 15318 29750 0 _0488_
rlabel metal1 15364 34578 15364 34578 0 _0489_
rlabel metal2 14812 32028 14812 32028 0 _0490_
rlabel metal1 14168 33898 14168 33898 0 _0491_
rlabel via1 14584 32878 14584 32878 0 _0492_
rlabel metal2 14398 33082 14398 33082 0 _0493_
rlabel metal1 14076 33830 14076 33830 0 _0494_
rlabel metal1 14122 32912 14122 32912 0 _0495_
rlabel metal1 14582 32742 14582 32742 0 _0496_
rlabel metal1 11362 29512 11362 29512 0 _0497_
rlabel metal1 9844 30770 9844 30770 0 _0498_
rlabel metal1 9062 29750 9062 29750 0 _0499_
rlabel metal1 9706 29648 9706 29648 0 _0500_
rlabel metal1 10810 29648 10810 29648 0 _0501_
rlabel metal1 9522 6256 9522 6256 0 _0502_
rlabel metal1 5934 11016 5934 11016 0 _0503_
rlabel metal1 29440 6766 29440 6766 0 _0504_
rlabel metal1 35880 29274 35880 29274 0 _0505_
rlabel metal1 5520 23086 5520 23086 0 _0506_
rlabel metal1 8602 5678 8602 5678 0 _0507_
rlabel metal1 37490 23630 37490 23630 0 _0508_
rlabel metal2 26450 26044 26450 26044 0 _0509_
rlabel metal3 26082 31756 26082 31756 0 _0510_
rlabel metal1 21574 4080 21574 4080 0 _0511_
rlabel metal1 21390 9486 21390 9486 0 _0512_
rlabel metal2 21850 3536 21850 3536 0 _0513_
rlabel metal1 24886 4794 24886 4794 0 _0514_
rlabel metal1 26726 6290 26726 6290 0 _0515_
rlabel metal1 20608 2414 20608 2414 0 _0516_
rlabel metal1 27508 9418 27508 9418 0 _0517_
rlabel metal1 22264 8058 22264 8058 0 _0518_
rlabel metal1 26450 4114 26450 4114 0 _0519_
rlabel metal2 30314 26316 30314 26316 0 _0520_
rlabel metal2 31602 23664 31602 23664 0 _0521_
rlabel metal1 30268 17170 30268 17170 0 _0522_
rlabel metal1 14398 26010 14398 26010 0 _0523_
rlabel metal1 14536 27642 14536 27642 0 _0524_
rlabel metal1 15042 32232 15042 32232 0 _0525_
rlabel metal1 13846 32470 13846 32470 0 _0526_
rlabel metal1 14766 32504 14766 32504 0 _0527_
rlabel metal1 15134 27982 15134 27982 0 _0528_
rlabel metal1 8510 26758 8510 26758 0 _0529_
rlabel metal1 10120 28050 10120 28050 0 _0530_
rlabel metal1 8878 28084 8878 28084 0 _0531_
rlabel metal1 13754 28016 13754 28016 0 _0532_
rlabel via2 14674 27931 14674 27931 0 _0533_
rlabel metal1 31510 16524 31510 16524 0 _0534_
rlabel metal1 33902 19448 33902 19448 0 _0535_
rlabel metal2 38870 16660 38870 16660 0 _0536_
rlabel viali 34965 11118 34965 11118 0 _0537_
rlabel metal1 33994 18802 33994 18802 0 _0538_
rlabel metal2 12926 29444 12926 29444 0 _0539_
rlabel metal1 17894 29580 17894 29580 0 _0540_
rlabel metal2 17066 29818 17066 29818 0 _0541_
rlabel metal2 17894 28781 17894 28781 0 _0542_
rlabel metal2 32246 18938 32246 18938 0 _0543_
rlabel metal2 34270 14025 34270 14025 0 _0544_
rlabel metal1 29486 18292 29486 18292 0 _0545_
rlabel metal1 38318 19822 38318 19822 0 _0546_
rlabel metal2 31510 20468 31510 20468 0 _0547_
rlabel metal1 31648 21590 31648 21590 0 _0548_
rlabel metal1 31050 20944 31050 20944 0 _0549_
rlabel metal1 31326 20910 31326 20910 0 _0550_
rlabel metal1 32154 20876 32154 20876 0 _0551_
rlabel viali 32616 20434 32616 20434 0 _0552_
rlabel metal1 39008 13294 39008 13294 0 _0553_
rlabel metal1 36386 12614 36386 12614 0 _0554_
rlabel via1 37124 8942 37124 8942 0 _0555_
rlabel metal1 39514 13362 39514 13362 0 _0556_
rlabel metal2 36662 16592 36662 16592 0 _0557_
rlabel metal1 32108 8806 32108 8806 0 _0558_
rlabel metal1 31372 16626 31372 16626 0 _0559_
rlabel metal1 30912 17646 30912 17646 0 _0560_
rlabel metal1 30820 16541 30820 16541 0 _0561_
rlabel metal1 29992 16422 29992 16422 0 _0562_
rlabel metal1 30866 17306 30866 17306 0 _0563_
rlabel metal1 31234 17850 31234 17850 0 _0564_
rlabel metal1 31878 18394 31878 18394 0 _0565_
rlabel metal1 29440 15538 29440 15538 0 _0566_
rlabel metal1 30084 14994 30084 14994 0 _0567_
rlabel metal1 32108 14314 32108 14314 0 _0568_
rlabel metal2 31510 16065 31510 16065 0 _0569_
rlabel metal1 31510 14960 31510 14960 0 _0570_
rlabel metal1 31740 14586 31740 14586 0 _0571_
rlabel metal1 29762 14926 29762 14926 0 _0572_
rlabel viali 29302 16576 29302 16576 0 _0573_
rlabel metal1 28842 12274 28842 12274 0 _0574_
rlabel metal1 30924 12206 30924 12206 0 _0575_
rlabel metal1 31970 13804 31970 13804 0 _0576_
rlabel metal2 31326 12988 31326 12988 0 _0577_
rlabel metal1 31832 12410 31832 12410 0 _0578_
rlabel metal2 32246 13022 32246 13022 0 _0579_
rlabel metal1 31602 12750 31602 12750 0 _0580_
rlabel metal2 30774 12512 30774 12512 0 _0581_
rlabel metal1 30636 12206 30636 12206 0 _0582_
rlabel metal1 30360 12138 30360 12138 0 _0583_
rlabel metal1 28750 12172 28750 12172 0 _0584_
rlabel metal2 35558 13719 35558 13719 0 _0585_
rlabel metal1 36064 13294 36064 13294 0 _0586_
rlabel metal2 34178 13600 34178 13600 0 _0587_
rlabel metal1 31372 13906 31372 13906 0 _0588_
rlabel metal1 33212 13294 33212 13294 0 _0589_
rlabel metal1 33304 13498 33304 13498 0 _0590_
rlabel metal1 33120 13702 33120 13702 0 _0591_
rlabel metal1 33258 17102 33258 17102 0 _0592_
rlabel metal1 33902 16048 33902 16048 0 _0593_
rlabel metal1 33902 15878 33902 15878 0 _0594_
rlabel metal1 32338 16490 32338 16490 0 _0595_
rlabel metal1 33212 16082 33212 16082 0 _0596_
rlabel metal1 33718 13906 33718 13906 0 _0597_
rlabel metal1 33120 13838 33120 13838 0 _0598_
rlabel metal1 35604 13498 35604 13498 0 _0599_
rlabel metal2 34730 14518 34730 14518 0 _0600_
rlabel metal1 35282 14382 35282 14382 0 _0601_
rlabel metal1 35512 13974 35512 13974 0 _0602_
rlabel metal1 35558 14314 35558 14314 0 _0603_
rlabel metal1 32798 16524 32798 16524 0 _0604_
rlabel metal1 34178 16558 34178 16558 0 _0605_
rlabel metal1 34500 16014 34500 16014 0 _0606_
rlabel metal1 35466 15470 35466 15470 0 _0607_
rlabel metal2 35558 14858 35558 14858 0 _0608_
rlabel metal1 33258 17306 33258 17306 0 _0609_
rlabel metal1 33550 18326 33550 18326 0 _0610_
rlabel metal1 33396 18394 33396 18394 0 _0611_
rlabel metal1 33672 18938 33672 18938 0 _0612_
rlabel viali 35923 20910 35923 20910 0 _0613_
rlabel viali 35745 20910 35745 20910 0 _0614_
rlabel metal1 36570 20400 36570 20400 0 _0615_
rlabel metal1 35972 13498 35972 13498 0 _0616_
rlabel metal1 34868 13770 34868 13770 0 _0617_
rlabel metal1 34868 19822 34868 19822 0 _0618_
rlabel metal1 33534 19856 33534 19856 0 _0619_
rlabel metal1 34868 17510 34868 17510 0 _0620_
rlabel metal1 34600 18394 34600 18394 0 _0621_
rlabel metal1 35328 18394 35328 18394 0 _0622_
rlabel metal1 36478 22066 36478 22066 0 _0623_
rlabel metal1 36294 20434 36294 20434 0 _0624_
rlabel metal1 35604 18938 35604 18938 0 _0625_
rlabel metal1 36156 21522 36156 21522 0 _0626_
rlabel metal1 36018 21624 36018 21624 0 _0627_
rlabel metal1 36524 21590 36524 21590 0 _0628_
rlabel metal1 36064 21386 36064 21386 0 _0629_
rlabel metal1 37260 21658 37260 21658 0 _0630_
rlabel metal1 37122 21896 37122 21896 0 _0631_
rlabel metal1 21712 16626 21712 16626 0 _0632_
rlabel metal2 26404 11730 26404 11730 0 _0633_
rlabel metal2 21758 16218 21758 16218 0 _0634_
rlabel metal2 21482 16048 21482 16048 0 _0635_
rlabel metal2 36570 17068 36570 17068 0 _0636_
rlabel metal2 14582 34646 14582 34646 0 _0637_
rlabel metal2 13754 34782 13754 34782 0 _0638_
rlabel metal1 13846 34646 13846 34646 0 _0639_
rlabel metal1 14536 34578 14536 34578 0 _0640_
rlabel metal1 14582 29206 14582 29206 0 _0641_
rlabel metal1 10626 28968 10626 28968 0 _0642_
rlabel metal1 10496 29274 10496 29274 0 _0643_
rlabel metal2 10810 28730 10810 28730 0 _0644_
rlabel metal3 16261 3876 16261 3876 0 _0645_
rlabel metal1 36984 4590 36984 4590 0 _0646_
rlabel metal1 23138 15130 23138 15130 0 _0647_
rlabel metal1 23000 15470 23000 15470 0 _0648_
rlabel metal2 37444 20604 37444 20604 0 _0649_
rlabel metal1 34776 22610 34776 22610 0 _0650_
rlabel metal1 26082 11764 26082 11764 0 _0651_
rlabel metal2 17802 4199 17802 4199 0 _0652_
rlabel metal1 17158 3706 17158 3706 0 _0653_
rlabel metal1 24610 15878 24610 15878 0 _0654_
rlabel metal1 25346 11526 25346 11526 0 _0655_
rlabel metal1 37812 11118 37812 11118 0 _0656_
rlabel metal1 39146 7922 39146 7922 0 _0657_
rlabel metal1 21436 11730 21436 11730 0 _0658_
rlabel metal2 21206 11679 21206 11679 0 _0659_
rlabel metal1 4370 26962 4370 26962 0 _0660_
rlabel metal1 26864 10778 26864 10778 0 _0661_
rlabel metal1 34868 9962 34868 9962 0 _0662_
rlabel metal1 34454 5270 34454 5270 0 _0663_
rlabel metal1 24288 11118 24288 11118 0 _0664_
rlabel metal1 32798 10030 32798 10030 0 _0665_
rlabel metal1 37168 5882 37168 5882 0 _0666_
rlabel metal1 26910 16150 26910 16150 0 _0667_
rlabel metal1 27002 16048 27002 16048 0 _0668_
rlabel metal2 32246 16099 32246 16099 0 _0669_
rlabel metal1 37352 28186 37352 28186 0 _0670_
rlabel metal1 32154 26282 32154 26282 0 _0671_
rlabel metal1 24840 31382 24840 31382 0 _0672_
rlabel metal3 24725 21556 24725 21556 0 _0673_
rlabel metal1 25116 20502 25116 20502 0 _0674_
rlabel metal1 20102 6868 20102 6868 0 _0675_
rlabel metal1 18814 8942 18814 8942 0 _0676_
rlabel metal2 20378 3978 20378 3978 0 _0677_
rlabel metal1 23000 5678 23000 5678 0 _0678_
rlabel metal1 28750 7310 28750 7310 0 _0679_
rlabel metal1 20516 5202 20516 5202 0 _0680_
rlabel metal1 26818 8466 26818 8466 0 _0681_
rlabel metal1 19274 6766 19274 6766 0 _0682_
rlabel metal2 25714 3638 25714 3638 0 _0683_
rlabel metal1 14766 15062 14766 15062 0 _0684_
rlabel metal1 20930 26418 20930 26418 0 _0685_
rlabel metal1 19826 25908 19826 25908 0 _0686_
rlabel metal1 14674 14892 14674 14892 0 _0687_
rlabel metal1 14030 15130 14030 15130 0 _0688_
rlabel metal1 14444 3502 14444 3502 0 _0689_
rlabel metal1 12972 4590 12972 4590 0 _0690_
rlabel metal1 13110 6324 13110 6324 0 _0691_
rlabel metal1 15594 3502 15594 3502 0 _0692_
rlabel metal1 13938 11152 13938 11152 0 _0693_
rlabel metal1 12834 7854 12834 7854 0 _0694_
rlabel metal1 13156 3502 13156 3502 0 _0695_
rlabel metal1 39100 19822 39100 19822 0 _0696_
rlabel metal1 36708 20026 36708 20026 0 _0697_
rlabel metal2 38870 20706 38870 20706 0 _0698_
rlabel metal1 38916 19890 38916 19890 0 _0699_
rlabel metal1 38778 19958 38778 19958 0 _0700_
rlabel metal1 35788 17578 35788 17578 0 _0701_
rlabel metal1 36202 18258 36202 18258 0 _0702_
rlabel metal1 36708 18394 36708 18394 0 _0703_
rlabel metal1 36984 18394 36984 18394 0 _0704_
rlabel metal1 37168 18938 37168 18938 0 _0705_
rlabel metal1 36892 17646 36892 17646 0 _0706_
rlabel metal1 37490 17510 37490 17510 0 _0707_
rlabel metal1 38318 18394 38318 18394 0 _0708_
rlabel metal1 38778 17272 38778 17272 0 _0709_
rlabel via2 39422 16541 39422 16541 0 _0710_
rlabel metal1 39146 15878 39146 15878 0 _0711_
rlabel via1 39236 17238 39236 17238 0 _0712_
rlabel metal1 39330 16966 39330 16966 0 _0713_
rlabel metal1 39238 17034 39238 17034 0 _0714_
rlabel metal1 39238 17850 39238 17850 0 _0715_
rlabel metal1 38594 18122 38594 18122 0 _0716_
rlabel metal1 39468 18734 39468 18734 0 _0717_
rlabel metal1 38732 14790 38732 14790 0 _0718_
rlabel metal2 39422 14212 39422 14212 0 _0719_
rlabel metal2 38686 14501 38686 14501 0 _0720_
rlabel metal1 38558 14416 38558 14416 0 _0721_
rlabel metal1 37720 15878 37720 15878 0 _0722_
rlabel metal1 37766 16116 37766 16116 0 _0723_
rlabel metal2 37398 14348 37398 14348 0 _0724_
rlabel metal1 37858 12852 37858 12852 0 _0725_
rlabel metal1 38824 13430 38824 13430 0 _0726_
rlabel metal1 36478 11866 36478 11866 0 _0727_
rlabel metal1 36938 11764 36938 11764 0 _0728_
rlabel metal1 36386 11050 36386 11050 0 _0729_
rlabel metal1 38916 10778 38916 10778 0 _0730_
rlabel metal2 39606 9724 39606 9724 0 _0731_
rlabel metal1 39790 9588 39790 9588 0 _0732_
rlabel metal2 39882 9860 39882 9860 0 _0733_
rlabel metal1 39652 13158 39652 13158 0 _0734_
rlabel metal1 39744 10234 39744 10234 0 _0735_
rlabel metal2 38686 10880 38686 10880 0 _0736_
rlabel metal1 38502 11322 38502 11322 0 _0737_
rlabel metal1 37812 8806 37812 8806 0 _0738_
rlabel metal1 39054 8976 39054 8976 0 _0739_
rlabel metal1 38134 8942 38134 8942 0 _0740_
rlabel metal1 37766 9520 37766 9520 0 _0741_
rlabel metal1 36938 8942 36938 8942 0 _0742_
rlabel viali 36754 8942 36754 8942 0 _0743_
rlabel metal1 36202 11322 36202 11322 0 _0744_
rlabel metal1 36624 11050 36624 11050 0 _0745_
rlabel metal1 36386 10676 36386 10676 0 _0746_
rlabel metal1 36064 10710 36064 10710 0 _0747_
rlabel metal1 36662 8908 36662 8908 0 _0748_
rlabel metal2 34086 8738 34086 8738 0 _0749_
rlabel metal1 34730 8976 34730 8976 0 _0750_
rlabel metal1 34362 8500 34362 8500 0 _0751_
rlabel metal1 34362 8398 34362 8398 0 _0752_
rlabel metal1 34914 8330 34914 8330 0 _0753_
rlabel metal1 35236 10642 35236 10642 0 _0754_
rlabel metal1 34776 10030 34776 10030 0 _0755_
rlabel metal1 35374 10064 35374 10064 0 _0756_
rlabel metal1 35466 9996 35466 9996 0 _0757_
rlabel metal1 34776 8466 34776 8466 0 _0758_
rlabel metal1 30774 8432 30774 8432 0 _0759_
rlabel metal1 30774 7820 30774 7820 0 _0760_
rlabel metal1 31096 7854 31096 7854 0 _0761_
rlabel metal1 34546 7786 34546 7786 0 _0762_
rlabel metal2 31142 8092 31142 8092 0 _0763_
rlabel metal2 32062 8058 32062 8058 0 _0764_
rlabel metal1 32936 10438 32936 10438 0 _0765_
rlabel metal1 32890 10166 32890 10166 0 _0766_
rlabel metal1 32522 9622 32522 9622 0 _0767_
rlabel metal1 32154 8500 32154 8500 0 _0768_
rlabel metal1 33258 10540 33258 10540 0 _0769_
rlabel metal1 32982 10234 32982 10234 0 _0770_
rlabel metal2 33534 10812 33534 10812 0 _0771_
rlabel metal2 32154 10982 32154 10982 0 _0772_
rlabel metal1 31142 8398 31142 8398 0 _0773_
rlabel metal1 30636 8602 30636 8602 0 _0774_
rlabel metal1 30958 10098 30958 10098 0 _0775_
rlabel metal1 31188 10234 31188 10234 0 _0776_
rlabel metal1 30544 10778 30544 10778 0 _0777_
rlabel metal1 29578 10030 29578 10030 0 _0778_
rlabel metal1 12788 26758 12788 26758 0 _0779_
rlabel metal1 12604 27574 12604 27574 0 _0780_
rlabel via1 12934 27098 12934 27098 0 _0781_
rlabel metal2 13110 26350 13110 26350 0 _0782_
rlabel metal2 6486 5814 6486 5814 0 _0783_
rlabel metal1 6118 5202 6118 5202 0 _0784_
rlabel metal2 31786 5406 31786 5406 0 _0785_
rlabel metal1 30360 23086 30360 23086 0 _0786_
rlabel metal1 39882 12206 39882 12206 0 _0787_
rlabel metal1 4278 6290 4278 6290 0 _0788_
rlabel metal1 11730 5134 11730 5134 0 _0789_
rlabel metal1 4094 24786 4094 24786 0 _0790_
rlabel metal1 39882 16558 39882 16558 0 _0791_
rlabel metal1 35742 25806 35742 25806 0 _0792_
rlabel metal1 35788 26010 35788 26010 0 _0793_
rlabel metal1 34730 28186 34730 28186 0 _0794_
rlabel metal1 33304 25874 33304 25874 0 _0795_
rlabel metal1 5336 26350 5336 26350 0 _0796_
rlabel metal2 33166 26758 33166 26758 0 _0797_
rlabel metal2 31510 24378 31510 24378 0 _0798_
rlabel metal1 7820 23154 7820 23154 0 _0799_
rlabel metal2 7130 23732 7130 23732 0 _0800_
rlabel metal1 11224 21522 11224 21522 0 _0801_
rlabel metal1 10074 22032 10074 22032 0 _0802_
rlabel metal1 8050 34918 8050 34918 0 _0803_
rlabel metal1 7176 35054 7176 35054 0 _0804_
rlabel metal1 10764 21114 10764 21114 0 _0805_
rlabel metal1 25668 23698 25668 23698 0 _0806_
rlabel metal1 26772 23562 26772 23562 0 _0807_
rlabel metal1 27140 19210 27140 19210 0 _0808_
rlabel metal1 27232 18734 27232 18734 0 _0809_
rlabel metal2 34822 33116 34822 33116 0 _0810_
rlabel metal1 35466 33082 35466 33082 0 _0811_
rlabel metal2 35006 32572 35006 32572 0 _0812_
rlabel metal1 34546 34442 34546 34442 0 _0813_
rlabel metal1 35190 31790 35190 31790 0 _0814_
rlabel metal1 34776 31858 34776 31858 0 _0815_
rlabel metal1 27370 32436 27370 32436 0 _0816_
rlabel metal1 33534 33898 33534 33898 0 _0817_
rlabel metal2 30222 33456 30222 33456 0 _0818_
rlabel metal2 30682 33218 30682 33218 0 _0819_
rlabel metal1 32039 32810 32039 32810 0 _0820_
rlabel metal2 25852 28764 25852 28764 0 _0821_
rlabel metal1 19182 30260 19182 30260 0 _0822_
rlabel metal1 21758 30702 21758 30702 0 _0823_
rlabel metal1 33350 31926 33350 31926 0 _0824_
rlabel metal2 32890 27608 32890 27608 0 _0825_
rlabel metal1 30038 32946 30038 32946 0 _0826_
rlabel metal1 27830 32912 27830 32912 0 _0827_
rlabel metal1 21528 31994 21528 31994 0 _0828_
rlabel metal2 30314 31994 30314 31994 0 _0829_
rlabel metal1 27462 31382 27462 31382 0 _0830_
rlabel metal1 23828 39270 23828 39270 0 _0831_
rlabel metal1 33212 30226 33212 30226 0 _0832_
rlabel metal1 21298 28458 21298 28458 0 _0833_
rlabel metal2 32706 30498 32706 30498 0 _0834_
rlabel metal1 34040 29478 34040 29478 0 _0835_
rlabel metal1 30268 30158 30268 30158 0 _0836_
rlabel metal2 24610 33626 24610 33626 0 _0837_
rlabel metal1 28658 30668 28658 30668 0 _0838_
rlabel via1 17618 34578 17618 34578 0 _0839_
rlabel metal2 21666 26163 21666 26163 0 _0840_
rlabel metal1 31786 31824 31786 31824 0 _0841_
rlabel metal1 30268 32538 30268 32538 0 _0842_
rlabel metal1 34270 33898 34270 33898 0 _0843_
rlabel metal1 27232 26962 27232 26962 0 _0844_
rlabel metal1 29256 41242 29256 41242 0 _0845_
rlabel metal2 26174 34595 26174 34595 0 _0846_
rlabel metal2 19458 33983 19458 33983 0 _0847_
rlabel metal2 21390 32912 21390 32912 0 _0848_
rlabel metal1 21574 31858 21574 31858 0 _0849_
rlabel metal1 26082 30736 26082 30736 0 _0850_
rlabel metal1 34592 32538 34592 32538 0 _0851_
rlabel metal1 34086 32980 34086 32980 0 _0852_
rlabel metal1 25622 33422 25622 33422 0 _0853_
rlabel metal1 35052 33014 35052 33014 0 _0854_
rlabel metal2 31878 33728 31878 33728 0 _0855_
rlabel metal1 25576 28934 25576 28934 0 _0856_
rlabel metal1 32706 28050 32706 28050 0 _0857_
rlabel metal2 30130 29818 30130 29818 0 _0858_
rlabel metal2 35466 30260 35466 30260 0 _0859_
rlabel metal1 34822 30770 34822 30770 0 _0860_
rlabel metal1 27600 28050 27600 28050 0 _0861_
rlabel metal1 26542 29682 26542 29682 0 _0862_
rlabel metal1 22034 31246 22034 31246 0 _0863_
rlabel metal1 33442 32538 33442 32538 0 _0864_
rlabel metal1 33304 32810 33304 32810 0 _0865_
rlabel metal2 27738 26367 27738 26367 0 _0866_
rlabel metal1 24748 32470 24748 32470 0 _0867_
rlabel metal2 20930 34204 20930 34204 0 _0868_
rlabel metal1 31602 31994 31602 31994 0 _0869_
rlabel metal2 26542 27200 26542 27200 0 _0870_
rlabel metal2 24702 26656 24702 26656 0 _0871_
rlabel metal1 23920 38862 23920 38862 0 _0872_
rlabel metal1 22034 39542 22034 39542 0 _0873_
rlabel metal1 21160 31994 21160 31994 0 _0874_
rlabel metal1 8740 32946 8740 32946 0 _0875_
rlabel metal1 22126 31348 22126 31348 0 _0876_
rlabel metal1 12650 28526 12650 28526 0 _0877_
rlabel metal3 21137 23460 21137 23460 0 _0878_
rlabel metal3 14398 33932 14398 33932 0 _0879_
rlabel metal3 30935 40052 30935 40052 0 _0880_
rlabel metal1 33902 34612 33902 34612 0 _0881_
rlabel metal1 32246 34476 32246 34476 0 _0882_
rlabel metal1 30912 26894 30912 26894 0 _0883_
rlabel metal2 35926 30464 35926 30464 0 _0884_
rlabel metal1 33626 28050 33626 28050 0 _0885_
rlabel metal1 30268 27098 30268 27098 0 _0886_
rlabel metal1 30406 26962 30406 26962 0 _0887_
rlabel metal2 30038 26605 30038 26605 0 _0888_
rlabel metal3 29785 40052 29785 40052 0 _0889_
rlabel metal3 24380 28900 24380 28900 0 _0890_
rlabel metal1 27332 27302 27332 27302 0 _0891_
rlabel metal1 28888 27574 28888 27574 0 _0892_
rlabel metal1 28980 27098 28980 27098 0 _0893_
rlabel metal1 28704 27098 28704 27098 0 _0894_
rlabel metal1 28014 27506 28014 27506 0 _0895_
rlabel metal1 19366 28492 19366 28492 0 _0896_
rlabel metal1 20884 24718 20884 24718 0 _0897_
rlabel metal1 14766 25228 14766 25228 0 _0898_
rlabel metal1 15180 25330 15180 25330 0 _0899_
rlabel metal1 15318 25466 15318 25466 0 _0900_
rlabel metal1 32476 28050 32476 28050 0 _0901_
rlabel metal1 32108 28050 32108 28050 0 _0902_
rlabel metal1 31694 28084 31694 28084 0 _0903_
rlabel via2 31970 27965 31970 27965 0 _0904_
rlabel metal1 14260 27914 14260 27914 0 _0905_
rlabel metal2 21022 23137 21022 23137 0 _0906_
rlabel metal1 28014 31858 28014 31858 0 _0907_
rlabel metal1 29118 30906 29118 30906 0 _0908_
rlabel metal1 32338 30056 32338 30056 0 _0909_
rlabel metal1 28382 39406 28382 39406 0 _0910_
rlabel metal1 21022 31824 21022 31824 0 _0911_
rlabel metal1 17802 24786 17802 24786 0 _0912_
rlabel metal1 19642 32198 19642 32198 0 _0913_
rlabel metal1 20010 32436 20010 32436 0 _0914_
rlabel metal1 24196 27302 24196 27302 0 _0915_
rlabel metal1 21390 27472 21390 27472 0 _0916_
rlabel metal1 17112 29138 17112 29138 0 _0917_
rlabel metal2 24610 26350 24610 26350 0 _0918_
rlabel metal1 20930 27608 20930 27608 0 _0919_
rlabel metal1 18492 32402 18492 32402 0 _0920_
rlabel metal2 31142 37162 31142 37162 0 _0921_
rlabel metal1 18262 32538 18262 32538 0 _0922_
rlabel metal1 29026 37196 29026 37196 0 _0923_
rlabel metal1 19596 26894 19596 26894 0 _0924_
rlabel metal1 18860 31994 18860 31994 0 _0925_
rlabel metal1 20562 29614 20562 29614 0 _0926_
rlabel metal1 21666 21420 21666 21420 0 _0927_
rlabel metal1 18262 30294 18262 30294 0 _0928_
rlabel metal1 18630 30022 18630 30022 0 _0929_
rlabel metal1 12926 25874 12926 25874 0 _0930_
rlabel metal1 18032 30906 18032 30906 0 _0931_
rlabel metal1 7958 32436 7958 32436 0 _0932_
rlabel metal1 21298 33320 21298 33320 0 _0933_
rlabel metal1 16928 32402 16928 32402 0 _0934_
rlabel via2 21114 23069 21114 23069 0 _0935_
rlabel metal1 14260 28730 14260 28730 0 _0936_
rlabel metal1 16238 30668 16238 30668 0 _0937_
rlabel metal1 17342 29002 17342 29002 0 _0938_
rlabel metal1 29624 32198 29624 32198 0 _0939_
rlabel metal1 30176 28526 30176 28526 0 _0940_
rlabel metal1 17986 23120 17986 23120 0 _0941_
rlabel metal1 18538 29274 18538 29274 0 _0942_
rlabel metal1 20608 28526 20608 28526 0 _0943_
rlabel metal2 19918 29801 19918 29801 0 _0944_
rlabel metal1 12098 27098 12098 27098 0 _0945_
rlabel metal2 19366 30022 19366 30022 0 _0946_
rlabel metal1 9522 34952 9522 34952 0 _0947_
rlabel metal1 20608 20434 20608 20434 0 _0948_
rlabel metal2 20010 30464 20010 30464 0 _0949_
rlabel metal1 19826 20876 19826 20876 0 _0950_
rlabel metal1 16284 20026 16284 20026 0 _0951_
rlabel metal1 21436 20502 21436 20502 0 _0952_
rlabel metal2 28014 23494 28014 23494 0 _0953_
rlabel metal2 15318 37281 15318 37281 0 _0954_
rlabel metal1 30866 25466 30866 25466 0 _0955_
rlabel metal2 16790 40868 16790 40868 0 _0956_
rlabel via1 14950 14382 14950 14382 0 _0957_
rlabel metal1 16560 40154 16560 40154 0 _0958_
rlabel metal1 17296 20502 17296 20502 0 _0959_
rlabel metal1 17986 20230 17986 20230 0 _0960_
rlabel metal2 13018 21165 13018 21165 0 _0961_
rlabel metal1 16652 36754 16652 36754 0 _0962_
rlabel metal2 16698 36312 16698 36312 0 _0963_
rlabel metal2 19274 40953 19274 40953 0 _0964_
rlabel metal1 17572 38318 17572 38318 0 _0965_
rlabel metal1 13202 37808 13202 37808 0 _0966_
rlabel metal1 19596 38930 19596 38930 0 _0967_
rlabel metal2 18906 37502 18906 37502 0 _0968_
rlabel metal1 18768 36550 18768 36550 0 _0969_
rlabel metal1 19918 37876 19918 37876 0 _0970_
rlabel metal1 19918 38318 19918 38318 0 _0971_
rlabel metal2 13110 37910 13110 37910 0 _0972_
rlabel metal1 20102 36142 20102 36142 0 _0973_
rlabel metal1 25300 40494 25300 40494 0 _0974_
rlabel metal1 25392 40358 25392 40358 0 _0975_
rlabel via1 27556 35666 27556 35666 0 _0976_
rlabel metal1 14306 40052 14306 40052 0 _0977_
rlabel metal1 18400 36074 18400 36074 0 _0978_
rlabel metal1 18078 36210 18078 36210 0 _0979_
rlabel metal1 12558 37196 12558 37196 0 _0980_
rlabel metal1 5980 29614 5980 29614 0 _0981_
rlabel metal2 18262 29546 18262 29546 0 _0982_
rlabel metal2 8602 32606 8602 32606 0 _0983_
rlabel metal2 9430 34850 9430 34850 0 _0984_
rlabel metal1 8418 32402 8418 32402 0 _0985_
rlabel metal1 8142 32300 8142 32300 0 _0986_
rlabel metal1 9338 32368 9338 32368 0 _0987_
rlabel metal1 9154 26860 9154 26860 0 _0988_
rlabel metal1 8510 30260 8510 30260 0 _0989_
rlabel metal1 8970 32402 8970 32402 0 _0990_
rlabel metal2 9614 34272 9614 34272 0 _0991_
rlabel metal1 8418 33558 8418 33558 0 _0992_
rlabel metal1 10810 26384 10810 26384 0 _0993_
rlabel via1 9545 33490 9545 33490 0 _0994_
rlabel metal1 9154 33286 9154 33286 0 _0995_
rlabel metal1 8878 32538 8878 32538 0 _0996_
rlabel metal1 17342 18734 17342 18734 0 _0997_
rlabel metal2 17710 18598 17710 18598 0 _0998_
rlabel metal1 15870 38352 15870 38352 0 _0999_
rlabel metal2 6394 32071 6394 32071 0 _1000_
rlabel metal1 14076 23834 14076 23834 0 _1001_
rlabel metal1 14536 24038 14536 24038 0 _1002_
rlabel metal1 16744 22746 16744 22746 0 _1003_
rlabel metal2 12098 27710 12098 27710 0 _1004_
rlabel metal1 19458 22032 19458 22032 0 _1005_
rlabel metal2 16054 23273 16054 23273 0 _1006_
rlabel metal2 13386 35020 13386 35020 0 _1007_
rlabel metal1 20746 26316 20746 26316 0 _1008_
rlabel metal2 6486 32674 6486 32674 0 _1009_
rlabel metal2 21850 41202 21850 41202 0 _1010_
rlabel metal2 15962 38964 15962 38964 0 _1011_
rlabel metal1 25852 18394 25852 18394 0 _1012_
rlabel via2 18630 39389 18630 39389 0 _1013_
rlabel metal1 15594 41140 15594 41140 0 _1014_
rlabel metal1 9844 38930 9844 38930 0 _1015_
rlabel metal2 15778 37026 15778 37026 0 _1016_
rlabel metal1 17802 39440 17802 39440 0 _1017_
rlabel metal1 25254 41208 25254 41208 0 _1018_
rlabel metal1 25622 41242 25622 41242 0 _1019_
rlabel metal2 9246 39678 9246 39678 0 _1020_
rlabel metal1 8970 39610 8970 39610 0 _1021_
rlabel metal1 18354 36788 18354 36788 0 _1022_
rlabel metal1 18170 38352 18170 38352 0 _1023_
rlabel metal1 17250 40528 17250 40528 0 _1024_
rlabel metal1 16514 41072 16514 41072 0 _1025_
rlabel metal1 15456 37774 15456 37774 0 _1026_
rlabel via2 12834 41021 12834 41021 0 _1027_
rlabel metal1 11868 41106 11868 41106 0 _1028_
rlabel metal1 15456 37842 15456 37842 0 _1029_
rlabel metal1 15088 37162 15088 37162 0 _1030_
rlabel metal1 13662 40392 13662 40392 0 _1031_
rlabel metal2 16790 39185 16790 39185 0 _1032_
rlabel metal1 19826 39440 19826 39440 0 _1033_
rlabel metal1 19872 38522 19872 38522 0 _1034_
rlabel metal1 17112 39610 17112 39610 0 _1035_
rlabel metal1 15226 37876 15226 37876 0 _1036_
rlabel metal1 15364 37706 15364 37706 0 _1037_
rlabel metal2 15778 37536 15778 37536 0 _1038_
rlabel metal1 18446 36720 18446 36720 0 _1039_
rlabel metal1 18216 38930 18216 38930 0 _1040_
rlabel metal1 16928 36210 16928 36210 0 _1041_
rlabel via1 16606 40477 16606 40477 0 _1042_
rlabel metal1 17204 40154 17204 40154 0 _1043_
rlabel metal1 15594 40698 15594 40698 0 _1044_
rlabel metal1 14076 41242 14076 41242 0 _1045_
rlabel metal2 16514 36550 16514 36550 0 _1046_
rlabel metal1 15732 36890 15732 36890 0 _1047_
rlabel metal2 26542 39270 26542 39270 0 _1048_
rlabel metal1 25921 38930 25921 38930 0 _1049_
rlabel metal1 27462 39032 27462 39032 0 _1050_
rlabel metal3 24725 39236 24725 39236 0 _1051_
rlabel metal1 23322 38998 23322 38998 0 _1052_
rlabel metal1 18906 36890 18906 36890 0 _1053_
rlabel metal1 25990 39984 25990 39984 0 _1054_
rlabel metal2 31326 35105 31326 35105 0 _1055_
rlabel metal1 26588 38998 26588 38998 0 _1056_
rlabel metal1 30636 38318 30636 38318 0 _1057_
rlabel metal1 24242 38862 24242 38862 0 _1058_
rlabel metal1 25668 39882 25668 39882 0 _1059_
rlabel metal1 23736 38522 23736 38522 0 _1060_
rlabel metal1 25530 39474 25530 39474 0 _1061_
rlabel metal2 22356 41548 22356 41548 0 _1062_
rlabel metal1 21528 38318 21528 38318 0 _1063_
rlabel metal1 31786 36788 31786 36788 0 _1064_
rlabel metal1 31234 39338 31234 39338 0 _1065_
rlabel metal1 20884 40358 20884 40358 0 _1066_
rlabel metal1 28106 38896 28106 38896 0 _1067_
rlabel metal2 17986 38760 17986 38760 0 _1068_
rlabel metal2 20654 38879 20654 38879 0 _1069_
rlabel metal1 28612 38726 28612 38726 0 _1070_
rlabel metal1 24472 30634 24472 30634 0 _1071_
rlabel metal2 29670 39100 29670 39100 0 _1072_
rlabel metal1 30866 38522 30866 38522 0 _1073_
rlabel metal1 18906 37128 18906 37128 0 _1074_
rlabel metal1 22218 37230 22218 37230 0 _1075_
rlabel metal1 27784 28662 27784 28662 0 _1076_
rlabel metal2 21574 37077 21574 37077 0 _1077_
rlabel metal1 23368 37230 23368 37230 0 _1078_
rlabel metal1 28298 26010 28298 26010 0 _1079_
rlabel metal1 22586 40392 22586 40392 0 _1080_
rlabel metal1 30544 40970 30544 40970 0 _1081_
rlabel metal1 22540 36142 22540 36142 0 _1082_
rlabel metal1 22494 35666 22494 35666 0 _1083_
rlabel via2 30958 29563 30958 29563 0 _1084_
rlabel metal2 25162 35122 25162 35122 0 _1085_
rlabel metal1 20608 41582 20608 41582 0 _1086_
rlabel metal2 24610 40630 24610 40630 0 _1087_
rlabel metal1 24932 38318 24932 38318 0 _1088_
rlabel metal1 23598 36176 23598 36176 0 _1089_
rlabel metal2 22494 40409 22494 40409 0 _1090_
rlabel metal1 29946 40562 29946 40562 0 _1091_
rlabel metal1 22494 38862 22494 38862 0 _1092_
rlabel metal2 23506 37536 23506 37536 0 _1093_
rlabel metal2 16054 32997 16054 32997 0 _1094_
rlabel metal1 20562 41208 20562 41208 0 _1095_
rlabel metal1 28244 36550 28244 36550 0 _1096_
rlabel via3 28037 38692 28037 38692 0 _1097_
rlabel metal1 28520 38862 28520 38862 0 _1098_
rlabel metal1 30544 38998 30544 38998 0 _1099_
rlabel metal2 32798 39678 32798 39678 0 _1100_
rlabel metal1 27646 36176 27646 36176 0 _1101_
rlabel metal1 20332 35598 20332 35598 0 _1102_
rlabel metal1 19826 35666 19826 35666 0 _1103_
rlabel metal1 28152 35122 28152 35122 0 _1104_
rlabel metal1 27600 35258 27600 35258 0 _1105_
rlabel metal1 30498 38352 30498 38352 0 _1106_
rlabel metal1 26266 38794 26266 38794 0 _1107_
rlabel metal2 28198 35768 28198 35768 0 _1108_
rlabel metal1 28842 37842 28842 37842 0 _1109_
rlabel metal1 29900 37978 29900 37978 0 _1110_
rlabel metal1 32522 39406 32522 39406 0 _1111_
rlabel metal2 22218 36516 22218 36516 0 _1112_
rlabel metal3 22724 38420 22724 38420 0 _1113_
rlabel metal2 19918 19091 19918 19091 0 _1114_
rlabel metal1 19366 36278 19366 36278 0 _1115_
rlabel metal2 20562 38080 20562 38080 0 _1116_
rlabel metal1 20378 36074 20378 36074 0 _1117_
rlabel metal2 20654 36516 20654 36516 0 _1118_
rlabel metal1 22402 36652 22402 36652 0 _1119_
rlabel metal2 21942 36533 21942 36533 0 _1120_
rlabel metal1 25714 33490 25714 33490 0 _1121_
rlabel metal2 25254 29291 25254 29291 0 _1122_
rlabel metal3 25369 38692 25369 38692 0 _1123_
rlabel metal1 27922 36720 27922 36720 0 _1124_
rlabel metal1 28750 35258 28750 35258 0 _1125_
rlabel metal2 31510 36669 31510 36669 0 _1126_
rlabel metal1 31694 34170 31694 34170 0 _1127_
rlabel metal2 26358 33150 26358 33150 0 _1128_
rlabel metal1 31234 35088 31234 35088 0 _1129_
rlabel metal1 32016 38726 32016 38726 0 _1130_
rlabel metal1 19826 28594 19826 28594 0 _1131_
rlabel metal1 26312 40902 26312 40902 0 _1132_
rlabel metal1 19964 39338 19964 39338 0 _1133_
rlabel metal1 20148 39882 20148 39882 0 _1134_
rlabel metal1 19412 41038 19412 41038 0 _1135_
rlabel metal1 19550 39338 19550 39338 0 _1136_
rlabel metal1 20286 38930 20286 38930 0 _1137_
rlabel metal1 21022 38862 21022 38862 0 _1138_
rlabel metal2 20286 39236 20286 39236 0 _1139_
rlabel metal1 29486 41174 29486 41174 0 _1140_
rlabel metal2 29302 40358 29302 40358 0 _1141_
rlabel metal1 28014 41072 28014 41072 0 _1142_
rlabel metal1 27140 33626 27140 33626 0 _1143_
rlabel via3 26059 39236 26059 39236 0 _1144_
rlabel metal1 26680 40494 26680 40494 0 _1145_
rlabel metal1 27508 40358 27508 40358 0 _1146_
rlabel metal1 30268 41446 30268 41446 0 _1147_
rlabel metal1 32706 38896 32706 38896 0 _1148_
rlabel metal1 33304 39066 33304 39066 0 _1149_
rlabel metal1 20746 32776 20746 32776 0 _1150_
rlabel metal1 23874 36754 23874 36754 0 _1151_
rlabel metal1 24380 24718 24380 24718 0 _1152_
rlabel metal2 25990 36346 25990 36346 0 _1153_
rlabel metal2 27278 37162 27278 37162 0 _1154_
rlabel metal1 26680 40358 26680 40358 0 _1155_
rlabel metal2 25392 32878 25392 32878 0 _1156_
rlabel metal1 25438 39542 25438 39542 0 _1157_
rlabel metal1 26910 37264 26910 37264 0 _1158_
rlabel metal2 27646 38148 27646 38148 0 _1159_
rlabel metal1 32062 39916 32062 39916 0 _1160_
rlabel via3 28405 40052 28405 40052 0 _1161_
rlabel metal1 29394 40936 29394 40936 0 _1162_
rlabel metal1 26266 41106 26266 41106 0 _1163_
rlabel metal1 30314 40358 30314 40358 0 _1164_
rlabel metal1 30728 39814 30728 39814 0 _1165_
rlabel metal1 20424 28526 20424 28526 0 _1166_
rlabel metal1 29486 40358 29486 40358 0 _1167_
rlabel metal3 21804 32164 21804 32164 0 _1168_
rlabel metal1 23966 40528 23966 40528 0 _1169_
rlabel metal2 23782 40681 23782 40681 0 _1170_
rlabel metal1 30314 40528 30314 40528 0 _1171_
rlabel metal1 31464 39950 31464 39950 0 _1172_
rlabel metal1 23184 34170 23184 34170 0 _1173_
rlabel metal2 24978 34102 24978 34102 0 _1174_
rlabel metal1 23230 35632 23230 35632 0 _1175_
rlabel metal1 29486 35632 29486 35632 0 _1176_
rlabel metal1 30912 40086 30912 40086 0 _1177_
rlabel metal2 32246 40290 32246 40290 0 _1178_
rlabel metal1 33074 40052 33074 40052 0 _1179_
rlabel metal1 22310 34714 22310 34714 0 _1180_
rlabel metal1 21206 38828 21206 38828 0 _1181_
rlabel metal1 21482 34578 21482 34578 0 _1182_
rlabel metal1 22448 38726 22448 38726 0 _1183_
rlabel metal1 22172 38726 22172 38726 0 _1184_
rlabel metal1 31924 34578 31924 34578 0 _1185_
rlabel metal1 32154 34544 32154 34544 0 _1186_
rlabel metal2 30866 36346 30866 36346 0 _1187_
rlabel metal1 32154 39508 32154 39508 0 _1188_
rlabel metal1 30636 34918 30636 34918 0 _1189_
rlabel metal2 24334 33864 24334 33864 0 _1190_
rlabel metal1 30544 35598 30544 35598 0 _1191_
rlabel metal2 32154 38012 32154 38012 0 _1192_
rlabel metal2 30314 37808 30314 37808 0 _1193_
rlabel metal1 28796 38250 28796 38250 0 _1194_
rlabel metal1 23736 37706 23736 37706 0 _1195_
rlabel metal1 29072 38522 29072 38522 0 _1196_
rlabel metal2 32154 38726 32154 38726 0 _1197_
rlabel metal2 32614 39202 32614 39202 0 _1198_
rlabel metal1 33442 38964 33442 38964 0 _1199_
rlabel metal1 26680 33626 26680 33626 0 _1200_
rlabel metal1 31418 37774 31418 37774 0 _1201_
rlabel metal2 21114 31127 21114 31127 0 _1202_
rlabel metal1 28244 35802 28244 35802 0 _1203_
rlabel metal1 20930 27506 20930 27506 0 _1204_
rlabel metal1 28520 36210 28520 36210 0 _1205_
rlabel metal1 31418 36142 31418 36142 0 _1206_
rlabel metal1 32338 37876 32338 37876 0 _1207_
rlabel metal1 22632 35258 22632 35258 0 _1208_
rlabel metal2 22402 35717 22402 35717 0 _1209_
rlabel metal1 32246 37672 32246 37672 0 _1210_
rlabel metal1 31510 36822 31510 36822 0 _1211_
rlabel metal1 32108 36890 32108 36890 0 _1212_
rlabel metal1 33396 37230 33396 37230 0 _1213_
rlabel via2 11914 32419 11914 32419 0 _1214_
rlabel metal1 30268 35462 30268 35462 0 _1215_
rlabel metal1 30774 35802 30774 35802 0 _1216_
rlabel metal1 31786 36618 31786 36618 0 _1217_
rlabel metal2 29670 39644 29670 39644 0 _1218_
rlabel metal1 29348 39066 29348 39066 0 _1219_
rlabel metal1 25852 38386 25852 38386 0 _1220_
rlabel metal2 25898 37026 25898 37026 0 _1221_
rlabel metal2 29026 38896 29026 38896 0 _1222_
rlabel metal1 30590 36074 30590 36074 0 _1223_
rlabel metal2 32522 35836 32522 35836 0 _1224_
rlabel metal1 32476 36890 32476 36890 0 _1225_
rlabel metal1 32154 37332 32154 37332 0 _1226_
rlabel metal1 26910 39814 26910 39814 0 _1227_
rlabel metal1 20654 38318 20654 38318 0 _1228_
rlabel metal2 20930 39236 20930 39236 0 _1229_
rlabel metal1 27002 40052 27002 40052 0 _1230_
rlabel metal2 32338 38573 32338 38573 0 _1231_
rlabel metal1 28060 36142 28060 36142 0 _1232_
rlabel metal1 32154 36210 32154 36210 0 _1233_
rlabel metal1 32936 36754 32936 36754 0 _1234_
rlabel metal1 5198 20910 5198 20910 0 _1235_
rlabel metal1 2208 22202 2208 22202 0 _1236_
rlabel metal1 25116 25942 25116 25942 0 _1237_
rlabel metal1 25162 27302 25162 27302 0 _1238_
rlabel metal1 25346 26826 25346 26826 0 _1239_
rlabel metal1 12972 35054 12972 35054 0 _1240_
rlabel metal1 13110 20808 13110 20808 0 _1241_
rlabel metal1 19366 26792 19366 26792 0 _1242_
rlabel metal2 17066 34612 17066 34612 0 _1243_
rlabel metal3 13754 28900 13754 28900 0 _1244_
rlabel metal1 17802 27302 17802 27302 0 _1245_
rlabel metal1 18262 28084 18262 28084 0 _1246_
rlabel viali 19368 28050 19368 28050 0 _1247_
rlabel metal1 20654 23562 20654 23562 0 _1248_
rlabel metal1 21114 29138 21114 29138 0 _1249_
rlabel metal2 19182 28220 19182 28220 0 _1250_
rlabel metal1 19044 27642 19044 27642 0 _1251_
rlabel metal1 19435 27846 19435 27846 0 _1252_
rlabel metal1 11086 25942 11086 25942 0 _1253_
rlabel metal1 12190 26996 12190 26996 0 _1254_
rlabel metal1 18906 26418 18906 26418 0 _1255_
rlabel metal1 19596 14994 19596 14994 0 _1256_
rlabel metal2 26818 15963 26818 15963 0 _1257_
rlabel metal1 21482 21522 21482 21522 0 _1258_
rlabel metal1 20838 32878 20838 32878 0 _1259_
rlabel metal2 16146 28679 16146 28679 0 _1260_
rlabel metal1 22080 21522 22080 21522 0 _1261_
rlabel metal1 22034 20400 22034 20400 0 _1262_
rlabel metal1 15870 27438 15870 27438 0 _1263_
rlabel metal1 21022 22644 21022 22644 0 _1264_
rlabel metal1 20240 18122 20240 18122 0 _1265_
rlabel metal1 20102 26418 20102 26418 0 _1266_
rlabel metal2 18446 24735 18446 24735 0 _1267_
rlabel metal1 22678 30192 22678 30192 0 _1268_
rlabel metal1 22632 24786 22632 24786 0 _1269_
rlabel metal1 22586 24650 22586 24650 0 _1270_
rlabel metal1 24518 22066 24518 22066 0 _1271_
rlabel metal1 22816 24038 22816 24038 0 _1272_
rlabel metal2 22310 30073 22310 30073 0 _1273_
rlabel metal2 20654 24837 20654 24837 0 _1274_
rlabel metal1 15686 28696 15686 28696 0 _1275_
rlabel metal2 23046 26826 23046 26826 0 _1276_
rlabel metal2 22218 24956 22218 24956 0 _1277_
rlabel metal1 20950 24174 20950 24174 0 _1278_
rlabel metal1 20056 24786 20056 24786 0 _1279_
rlabel metal1 20562 24038 20562 24038 0 _1280_
rlabel metal2 11086 24429 11086 24429 0 _1281_
rlabel metal2 10902 28152 10902 28152 0 _1282_
rlabel metal1 11132 27982 11132 27982 0 _1283_
rlabel metal1 9890 25296 9890 25296 0 _1284_
rlabel metal1 9522 31246 9522 31246 0 _1285_
rlabel metal1 9936 26962 9936 26962 0 _1286_
rlabel metal1 9798 25908 9798 25908 0 _1287_
rlabel metal1 9752 25466 9752 25466 0 _1288_
rlabel metal1 22034 20502 22034 20502 0 _1289_
rlabel metal1 17342 29614 17342 29614 0 _1290_
rlabel metal2 20654 22100 20654 22100 0 _1291_
rlabel metal2 21942 19958 21942 19958 0 _1292_
rlabel metal1 22724 20434 22724 20434 0 _1293_
rlabel metal1 24853 19822 24853 19822 0 _1294_
rlabel viali 17342 25896 17342 25896 0 _1295_
rlabel metal1 12006 32436 12006 32436 0 _1296_
rlabel via2 19550 20451 19550 20451 0 _1297_
rlabel metal1 23276 24378 23276 24378 0 _1298_
rlabel metal1 21666 21318 21666 21318 0 _1299_
rlabel metal1 19964 20570 19964 20570 0 _1300_
rlabel metal1 21022 19924 21022 19924 0 _1301_
rlabel metal1 22637 19686 22637 19686 0 _1302_
rlabel metal2 21390 19142 21390 19142 0 _1303_
rlabel metal2 22310 19686 22310 19686 0 _1304_
rlabel metal1 17250 21896 17250 21896 0 _1305_
rlabel metal1 17388 23086 17388 23086 0 _1306_
rlabel metal1 18216 21998 18216 21998 0 _1307_
rlabel metal2 18170 21896 18170 21896 0 _1308_
rlabel metal1 18814 21556 18814 21556 0 _1309_
rlabel metal1 17572 19686 17572 19686 0 _1310_
rlabel metal2 18630 21216 18630 21216 0 _1311_
rlabel metal1 23414 18734 23414 18734 0 _1312_
rlabel metal2 22678 18122 22678 18122 0 _1313_
rlabel metal1 25944 18122 25944 18122 0 _1314_
rlabel metal1 22678 18258 22678 18258 0 _1315_
rlabel metal1 23782 19346 23782 19346 0 _1316_
rlabel metal2 24702 19448 24702 19448 0 _1317_
rlabel metal1 27922 18360 27922 18360 0 _1318_
rlabel metal2 24426 15300 24426 15300 0 _1319_
rlabel metal2 24978 14314 24978 14314 0 _1320_
rlabel metal2 24472 12818 24472 12818 0 _1321_
rlabel metal2 23230 11322 23230 11322 0 _1322_
rlabel metal2 19826 20026 19826 20026 0 _1323_
rlabel metal1 18952 21998 18952 21998 0 _1324_
rlabel metal1 19872 19278 19872 19278 0 _1325_
rlabel metal1 19918 16524 19918 16524 0 _1326_
rlabel metal1 19412 14994 19412 14994 0 _1327_
rlabel metal1 20056 14382 20056 14382 0 _1328_
rlabel metal1 23276 16082 23276 16082 0 _1329_
rlabel metal1 19550 12784 19550 12784 0 _1330_
rlabel metal1 9430 35632 9430 35632 0 _1331_
rlabel metal2 16606 19737 16606 19737 0 _1332_
rlabel metal4 17940 26248 17940 26248 0 _1333_
rlabel metal1 16606 20026 16606 20026 0 _1334_
rlabel metal1 16192 18734 16192 18734 0 _1335_
rlabel metal2 23736 21522 23736 21522 0 _1336_
rlabel metal1 23644 22066 23644 22066 0 _1337_
rlabel metal1 23690 21522 23690 21522 0 _1338_
rlabel metal2 23552 21828 23552 21828 0 _1339_
rlabel metal1 19550 20944 19550 20944 0 _1340_
rlabel metal2 16974 14705 16974 14705 0 _1341_
rlabel metal1 17986 11866 17986 11866 0 _1342_
rlabel metal2 21482 34850 21482 34850 0 _1343_
rlabel metal1 15134 35088 15134 35088 0 _1344_
rlabel metal1 15410 34986 15410 34986 0 _1345_
rlabel metal2 16744 18802 16744 18802 0 _1346_
rlabel metal1 11362 35088 11362 35088 0 _1347_
rlabel metal1 11270 35020 11270 35020 0 _1348_
rlabel via2 16606 18819 16606 18819 0 _1349_
rlabel metal1 19642 11050 19642 11050 0 _1350_
rlabel viali 18538 21517 18538 21517 0 _1351_
rlabel metal1 16882 25364 16882 25364 0 _1352_
rlabel metal2 25806 26469 25806 26469 0 _1353_
rlabel metal1 21712 26758 21712 26758 0 _1354_
rlabel metal1 19136 25874 19136 25874 0 _1355_
rlabel metal1 18124 25262 18124 25262 0 _1356_
rlabel metal1 19366 24242 19366 24242 0 _1357_
rlabel metal3 20539 28220 20539 28220 0 _1358_
rlabel metal2 19274 23936 19274 23936 0 _1359_
rlabel metal2 23322 26996 23322 26996 0 _1360_
rlabel metal1 18860 26758 18860 26758 0 _1361_
rlabel metal1 19688 26214 19688 26214 0 _1362_
rlabel metal1 18906 25330 18906 25330 0 _1363_
rlabel metal1 9246 24752 9246 24752 0 _1364_
rlabel metal2 18446 21879 18446 21879 0 _1365_
rlabel metal1 18308 21318 18308 21318 0 _1366_
rlabel metal1 19412 11118 19412 11118 0 _1367_
rlabel metal1 18354 11322 18354 11322 0 _1368_
rlabel metal1 18492 11730 18492 11730 0 _1369_
rlabel metal2 18630 10506 18630 10506 0 _1370_
rlabel via1 19274 7395 19274 7395 0 _1371_
rlabel metal1 18722 12614 18722 12614 0 _1372_
rlabel metal1 19918 10438 19918 10438 0 _1373_
rlabel metal1 19688 10778 19688 10778 0 _1374_
rlabel metal1 19826 8500 19826 8500 0 _1375_
rlabel metal2 19734 8058 19734 8058 0 _1376_
rlabel metal1 16284 10642 16284 10642 0 _1377_
rlabel metal1 16192 13226 16192 13226 0 _1378_
rlabel metal1 19918 7854 19918 7854 0 _1379_
rlabel metal1 23000 10030 23000 10030 0 _1380_
rlabel metal1 19182 29002 19182 29002 0 _1381_
rlabel metal2 17342 18105 17342 18105 0 _1382_
rlabel metal1 21160 17170 21160 17170 0 _1383_
rlabel metal1 13156 28730 13156 28730 0 _1384_
rlabel metal1 17250 25908 17250 25908 0 _1385_
rlabel metal1 18354 16592 18354 16592 0 _1386_
rlabel metal1 20424 13906 20424 13906 0 _1387_
rlabel metal1 20332 12818 20332 12818 0 _1388_
rlabel metal2 16698 32096 16698 32096 0 _1389_
rlabel via1 16514 30685 16514 30685 0 _1390_
rlabel metal1 16744 32334 16744 32334 0 _1391_
rlabel metal1 15870 32470 15870 32470 0 _1392_
rlabel metal1 20102 34000 20102 34000 0 _1393_
rlabel metal1 16238 33320 16238 33320 0 _1394_
rlabel metal1 18722 33898 18722 33898 0 _1395_
rlabel metal1 18906 33966 18906 33966 0 _1396_
rlabel metal1 18584 33082 18584 33082 0 _1397_
rlabel metal1 17204 33422 17204 33422 0 _1398_
rlabel metal1 17526 34612 17526 34612 0 _1399_
rlabel metal1 14904 35054 14904 35054 0 _1400_
rlabel metal1 16882 34578 16882 34578 0 _1401_
rlabel metal1 15962 33592 15962 33592 0 _1402_
rlabel metal1 15962 30226 15962 30226 0 _1403_
rlabel metal1 20838 31280 20838 31280 0 _1404_
rlabel metal1 16008 30022 16008 30022 0 _1405_
rlabel metal1 16238 30362 16238 30362 0 _1406_
rlabel metal1 16790 20978 16790 20978 0 _1407_
rlabel metal1 17066 20910 17066 20910 0 _1408_
rlabel metal1 15778 25126 15778 25126 0 _1409_
rlabel metal1 16652 20910 16652 20910 0 _1410_
rlabel metal1 13662 31858 13662 31858 0 _1411_
rlabel metal1 16698 30260 16698 30260 0 _1412_
rlabel metal1 8372 29274 8372 29274 0 _1413_
rlabel metal1 11500 30022 11500 30022 0 _1414_
rlabel metal1 11454 29614 11454 29614 0 _1415_
rlabel metal1 11408 29818 11408 29818 0 _1416_
rlabel metal2 16330 29937 16330 29937 0 _1417_
rlabel metal2 16054 21063 16054 21063 0 _1418_
rlabel metal2 12282 20706 12282 20706 0 _1419_
rlabel metal2 12190 20706 12190 20706 0 _1420_
rlabel metal1 15042 20842 15042 20842 0 _1421_
rlabel metal2 16422 20060 16422 20060 0 _1422_
rlabel metal1 20148 18258 20148 18258 0 _1423_
rlabel metal1 23184 16558 23184 16558 0 _1424_
rlabel metal2 18078 17884 18078 17884 0 _1425_
rlabel metal1 17342 26792 17342 26792 0 _1426_
rlabel metal1 16100 27846 16100 27846 0 _1427_
rlabel metal2 17572 22080 17572 22080 0 _1428_
rlabel metal1 22218 16558 22218 16558 0 _1429_
rlabel metal1 21068 16082 21068 16082 0 _1430_
rlabel metal1 23966 13872 23966 13872 0 _1431_
rlabel metal1 24748 11118 24748 11118 0 _1432_
rlabel metal1 23000 10642 23000 10642 0 _1433_
rlabel metal1 9246 11322 9246 11322 0 _1434_
rlabel metal1 9292 34646 9292 34646 0 _1435_
rlabel metal1 8418 24310 8418 24310 0 _1436_
rlabel metal1 8050 24752 8050 24752 0 _1437_
rlabel metal1 10350 23086 10350 23086 0 _1438_
rlabel metal1 11730 23698 11730 23698 0 _1439_
rlabel metal2 13018 24922 13018 24922 0 _1440_
rlabel metal1 14444 27098 14444 27098 0 _1441_
rlabel metal1 12926 24208 12926 24208 0 _1442_
rlabel metal1 12236 24174 12236 24174 0 _1443_
rlabel metal1 16330 24242 16330 24242 0 _1444_
rlabel metal1 11638 24242 11638 24242 0 _1445_
rlabel metal1 9430 26962 9430 26962 0 _1446_
rlabel metal2 8878 26316 8878 26316 0 _1447_
rlabel metal1 8970 25466 8970 25466 0 _1448_
rlabel metal1 8970 25704 8970 25704 0 _1449_
rlabel metal2 10718 23562 10718 23562 0 _1450_
rlabel metal1 18630 21964 18630 21964 0 _1451_
rlabel metal1 20102 22508 20102 22508 0 _1452_
rlabel metal1 18492 20910 18492 20910 0 _1453_
rlabel metal1 20286 22406 20286 22406 0 _1454_
rlabel metal2 17710 23392 17710 23392 0 _1455_
rlabel metal1 18400 22610 18400 22610 0 _1456_
rlabel metal2 18584 22406 18584 22406 0 _1457_
rlabel metal1 16376 21046 16376 21046 0 _1458_
rlabel metal1 11316 18326 11316 18326 0 _1459_
rlabel metal1 10902 11662 10902 11662 0 _1460_
rlabel metal1 9522 16592 9522 16592 0 _1461_
rlabel metal2 13018 23188 13018 23188 0 _1462_
rlabel metal1 13248 23698 13248 23698 0 _1463_
rlabel metal2 12466 20407 12466 20407 0 _1464_
rlabel metal1 12742 18292 12742 18292 0 _1465_
rlabel metal2 12742 19958 12742 19958 0 _1466_
rlabel metal1 13340 17646 13340 17646 0 _1467_
rlabel metal1 13478 17578 13478 17578 0 _1468_
rlabel metal1 15318 25806 15318 25806 0 _1469_
rlabel metal1 15272 23086 15272 23086 0 _1470_
rlabel metal1 22402 24276 22402 24276 0 _1471_
rlabel metal2 15042 23205 15042 23205 0 _1472_
rlabel metal1 15778 23120 15778 23120 0 _1473_
rlabel metal1 22126 22542 22126 22542 0 _1474_
rlabel metal1 15410 22950 15410 22950 0 _1475_
rlabel metal1 16008 23290 16008 23290 0 _1476_
rlabel metal1 10580 23698 10580 23698 0 _1477_
rlabel metal1 13478 21998 13478 21998 0 _1478_
rlabel metal2 14582 22508 14582 22508 0 _1479_
rlabel metal1 13754 17510 13754 17510 0 _1480_
rlabel metal2 23874 10676 23874 10676 0 _1481_
rlabel metal2 13202 17153 13202 17153 0 _1482_
rlabel metal2 11638 17476 11638 17476 0 _1483_
rlabel metal2 13846 20400 13846 20400 0 _1484_
rlabel metal1 15226 27574 15226 27574 0 _1485_
rlabel metal1 15042 29614 15042 29614 0 _1486_
rlabel metal1 14352 29682 14352 29682 0 _1487_
rlabel metal1 13984 19822 13984 19822 0 _1488_
rlabel metal1 15962 26894 15962 26894 0 _1489_
rlabel metal2 14306 20060 14306 20060 0 _1490_
rlabel metal1 12558 31314 12558 31314 0 _1491_
rlabel metal1 12374 31790 12374 31790 0 _1492_
rlabel metal1 12880 31654 12880 31654 0 _1493_
rlabel metal1 12374 30804 12374 30804 0 _1494_
rlabel metal1 9798 30872 9798 30872 0 _1495_
rlabel metal1 9665 31768 9665 31768 0 _1496_
rlabel metal1 11822 30770 11822 30770 0 _1497_
rlabel metal1 13110 20434 13110 20434 0 _1498_
rlabel metal1 12834 21896 12834 21896 0 _1499_
rlabel metal1 14352 19414 14352 19414 0 _1500_
rlabel metal1 14858 18360 14858 18360 0 _1501_
rlabel metal1 18630 18224 18630 18224 0 _1502_
rlabel metal2 38686 1520 38686 1520 0 addressBusHigh[0]
rlabel metal1 19090 42330 19090 42330 0 addressBusHigh[1]
rlabel metal2 15502 1520 15502 1520 0 addressBusHigh[2]
rlabel metal1 41032 8330 41032 8330 0 addressBusHigh[3]
rlabel metal3 820 32028 820 32028 0 addressBusHigh[4]
rlabel metal1 41032 4454 41032 4454 0 addressBusHigh[5]
rlabel metal1 40388 2278 40388 2278 0 addressBusHigh[6]
rlabel via2 40986 32725 40986 32725 0 addressBusHigh[7]
rlabel metal3 1740 44268 1740 44268 0 addressBusLow[0]
rlabel metal2 23230 1571 23230 1571 0 addressBusLow[1]
rlabel metal3 820 11628 820 11628 0 addressBusLow[2]
rlabel metal2 30958 1520 30958 1520 0 addressBusLow[3]
rlabel metal2 40986 36941 40986 36941 0 addressBusLow[4]
rlabel metal3 820 23868 820 23868 0 addressBusLow[5]
rlabel metal2 7774 1520 7774 1520 0 addressBusLow[6]
rlabel metal2 38318 43163 38318 43163 0 addressBusLow[7]
rlabel metal1 14352 21998 14352 21998 0 branch_ff.branchBackward
rlabel metal3 19412 21896 19412 21896 0 branch_ff.branchForward
rlabel metal2 21850 30617 21850 30617 0 clk
rlabel metal1 35880 12886 35880 12886 0 clknet_0_clk
rlabel metal1 10442 5746 10442 5746 0 clknet_4_0_0_clk
rlabel metal1 34684 7378 34684 7378 0 clknet_4_10_0_clk
rlabel metal1 36248 14382 36248 14382 0 clknet_4_11_0_clk
rlabel metal1 33074 20434 33074 20434 0 clknet_4_12_0_clk
rlabel metal1 38824 18326 38824 18326 0 clknet_4_13_0_clk
rlabel metal1 37812 39474 37812 39474 0 clknet_4_14_0_clk
rlabel metal1 32706 40562 32706 40562 0 clknet_4_15_0_clk
rlabel metal1 12190 14892 12190 14892 0 clknet_4_1_0_clk
rlabel metal1 20286 3570 20286 3570 0 clknet_4_2_0_clk
rlabel metal1 16790 6358 16790 6358 0 clknet_4_3_0_clk
rlabel metal1 2070 21454 2070 21454 0 clknet_4_4_0_clk
rlabel metal1 4140 25806 4140 25806 0 clknet_4_5_0_clk
rlabel metal1 4370 32266 4370 32266 0 clknet_4_6_0_clk
rlabel metal1 9108 37774 9108 37774 0 clknet_4_7_0_clk
rlabel metal2 29302 6052 29302 6052 0 clknet_4_8_0_clk
rlabel metal1 29624 19346 29624 19346 0 clknet_4_9_0_clk
rlabel metal1 41124 24786 41124 24786 0 dataBusEnable
rlabel metal1 34684 42262 34684 42262 0 dataBusInput[0]
rlabel metal3 820 7548 820 7548 0 dataBusInput[1]
rlabel metal1 40940 41106 40940 41106 0 dataBusInput[2]
rlabel metal1 7222 42262 7222 42262 0 dataBusInput[3]
rlabel metal2 46 1554 46 1554 0 dataBusInput[4]
rlabel metal1 22632 42194 22632 42194 0 dataBusInput[5]
rlabel metal1 41078 29138 41078 29138 0 dataBusInput[6]
rlabel metal1 3312 42194 3312 42194 0 dataBusInput[7]
rlabel metal3 820 3468 820 3468 0 dataBusOutput[0]
rlabel metal2 34822 1520 34822 1520 0 dataBusOutput[1]
rlabel metal1 30498 42330 30498 42330 0 dataBusOutput[2]
rlabel metal1 39974 13158 39974 13158 0 dataBusOutput[3]
rlabel metal2 3910 1571 3910 1571 0 dataBusOutput[4]
rlabel metal2 11638 1520 11638 1520 0 dataBusOutput[5]
rlabel metal3 820 36108 820 36108 0 dataBusOutput[6]
rlabel metal1 41262 17510 41262 17510 0 dataBusOutput[7]
rlabel metal2 19366 1520 19366 1520 0 dataBusSelect
rlabel metal1 29210 26826 29210 26826 0 demux.PSR_C
rlabel metal1 29440 18938 29440 18938 0 demux.PSR_N
rlabel metal3 20148 21624 20148 21624 0 demux.PSR_V
rlabel metal1 27278 20944 27278 20944 0 demux.PSR_Z
rlabel metal1 8050 35190 8050 35190 0 demux.isAddressing
rlabel metal2 17802 17442 17802 17442 0 demux.nmi
rlabel metal2 16836 19346 16836 19346 0 demux.reset
rlabel metal1 34684 26350 34684 26350 0 demux.setInterruptFlag
rlabel metal1 13110 41106 13110 41106 0 demux.state_machine.currentAddress\[0\]
rlabel metal2 10350 37468 10350 37468 0 demux.state_machine.currentAddress\[10\]
rlabel metal1 9522 39066 9522 39066 0 demux.state_machine.currentAddress\[11\]
rlabel metal2 9798 34272 9798 34272 0 demux.state_machine.currentAddress\[12\]
rlabel metal1 8234 36040 8234 36040 0 demux.state_machine.currentAddress\[1\]
rlabel metal2 14582 39984 14582 39984 0 demux.state_machine.currentAddress\[2\]
rlabel metal1 11500 39474 11500 39474 0 demux.state_machine.currentAddress\[3\]
rlabel metal2 9062 37434 9062 37434 0 demux.state_machine.currentAddress\[4\]
rlabel metal1 11362 40902 11362 40902 0 demux.state_machine.currentAddress\[5\]
rlabel metal2 9614 25534 9614 25534 0 demux.state_machine.currentAddress\[6\]
rlabel metal1 11178 26894 11178 26894 0 demux.state_machine.currentAddress\[7\]
rlabel metal1 13662 40494 13662 40494 0 demux.state_machine.currentAddress\[8\]
rlabel metal1 14996 40494 14996 40494 0 demux.state_machine.currentAddress\[9\]
rlabel metal2 34822 36346 34822 36346 0 demux.state_machine.currentInstruction\[0\]
rlabel metal2 34914 34850 34914 34850 0 demux.state_machine.currentInstruction\[1\]
rlabel metal2 35374 36550 35374 36550 0 demux.state_machine.currentInstruction\[2\]
rlabel metal2 35558 35564 35558 35564 0 demux.state_machine.currentInstruction\[3\]
rlabel metal1 32246 32878 32246 32878 0 demux.state_machine.currentInstruction\[4\]
rlabel metal1 33442 35496 33442 35496 0 demux.state_machine.currentInstruction\[5\]
rlabel metal2 8234 33575 8234 33575 0 demux.state_machine.timeState\[0\]
rlabel metal1 13202 32742 13202 32742 0 demux.state_machine.timeState\[1\]
rlabel metal1 7636 29138 7636 29138 0 demux.state_machine.timeState\[2\]
rlabel metal1 7268 32878 7268 32878 0 demux.state_machine.timeState\[3\]
rlabel metal1 16744 33898 16744 33898 0 demux.state_machine.timeState\[4\]
rlabel metal1 19412 32402 19412 32402 0 demux.state_machine.timeState\[5\]
rlabel metal1 8418 27064 8418 27064 0 demux.state_machine.timeState\[6\]
rlabel metal1 8556 23698 8556 23698 0 free_carry_ff.freeCarry
rlabel metal3 820 27948 820 27948 0 functionalClockOut
rlabel metal1 38456 40562 38456 40562 0 instructionLoader.interruptInjector.interruptRequest
rlabel metal1 31050 25228 31050 25228 0 instructionLoader.interruptInjector.irqGenerated
rlabel metal1 37582 26418 37582 26418 0 instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
rlabel metal1 39652 40562 39652 40562 0 instructionLoader.interruptInjector.irqSync.nextQ2
rlabel metal2 34362 27370 34362 27370 0 instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
rlabel metal1 34132 41446 34132 41446 0 instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
rlabel metal1 11638 42296 11638 42296 0 instructionLoader.interruptInjector.nmiSync.in
rlabel metal1 32568 41786 32568 41786 0 instructionLoader.interruptInjector.nmiSync.nextQ2
rlabel metal1 27692 14994 27692 14994 0 instructionLoader.interruptInjector.processStatusRegIFlag
rlabel metal2 32430 23290 32430 23290 0 instructionLoader.interruptInjector.resetDetected
rlabel metal1 22402 9146 22402 9146 0 internalDataflow.accRegToDB\[0\]
rlabel metal1 21482 6698 21482 6698 0 internalDataflow.accRegToDB\[1\]
rlabel metal2 27922 13707 27922 13707 0 internalDataflow.accRegToDB\[2\]
rlabel metal1 28336 13838 28336 13838 0 internalDataflow.accRegToDB\[3\]
rlabel via1 21114 7378 21114 7378 0 internalDataflow.accRegToDB\[4\]
rlabel metal2 26358 12823 26358 12823 0 internalDataflow.accRegToDB\[5\]
rlabel metal1 20010 8398 20010 8398 0 internalDataflow.accRegToDB\[6\]
rlabel metal2 28014 15339 28014 15339 0 internalDataflow.accRegToDB\[7\]
rlabel metal1 37352 18802 37352 18802 0 internalDataflow.addressHighBusModule.busInputs\[16\]
rlabel metal1 23690 16524 23690 16524 0 internalDataflow.addressHighBusModule.busInputs\[17\]
rlabel metal1 28566 15062 28566 15062 0 internalDataflow.addressHighBusModule.busInputs\[18\]
rlabel metal2 32614 12517 32614 12517 0 internalDataflow.addressHighBusModule.busInputs\[19\]
rlabel metal1 35328 9554 35328 9554 0 internalDataflow.addressHighBusModule.busInputs\[20\]
rlabel metal2 32246 12551 32246 12551 0 internalDataflow.addressHighBusModule.busInputs\[21\]
rlabel metal1 24702 13396 24702 13396 0 internalDataflow.addressHighBusModule.busInputs\[22\]
rlabel metal1 26956 17170 26956 17170 0 internalDataflow.addressHighBusModule.busInputs\[23\]
rlabel metal1 18538 18326 18538 18326 0 internalDataflow.addressLowBusModule.busInputs\[16\]
rlabel metal2 21942 17374 21942 17374 0 internalDataflow.addressLowBusModule.busInputs\[17\]
rlabel metal1 27370 14246 27370 14246 0 internalDataflow.addressLowBusModule.busInputs\[18\]
rlabel metal1 31970 13362 31970 13362 0 internalDataflow.addressLowBusModule.busInputs\[19\]
rlabel metal2 17802 14127 17802 14127 0 internalDataflow.addressLowBusModule.busInputs\[20\]
rlabel metal1 27738 13260 27738 13260 0 internalDataflow.addressLowBusModule.busInputs\[21\]
rlabel metal2 18446 15521 18446 15521 0 internalDataflow.addressLowBusModule.busInputs\[22\]
rlabel metal2 15226 17340 15226 17340 0 internalDataflow.addressLowBusModule.busInputs\[23\]
rlabel metal1 16744 14994 16744 14994 0 internalDataflow.addressLowBusModule.busInputs\[24\]
rlabel metal1 11178 7854 11178 7854 0 internalDataflow.addressLowBusModule.busInputs\[25\]
rlabel metal2 7958 7990 7958 7990 0 internalDataflow.addressLowBusModule.busInputs\[26\]
rlabel metal1 10396 7174 10396 7174 0 internalDataflow.addressLowBusModule.busInputs\[27\]
rlabel metal1 5978 12206 5978 12206 0 internalDataflow.addressLowBusModule.busInputs\[28\]
rlabel metal1 15226 11696 15226 11696 0 internalDataflow.addressLowBusModule.busInputs\[29\]
rlabel metal2 7958 10064 7958 10064 0 internalDataflow.addressLowBusModule.busInputs\[30\]
rlabel metal2 5566 8194 5566 8194 0 internalDataflow.addressLowBusModule.busInputs\[31\]
rlabel metal1 16652 15062 16652 15062 0 internalDataflow.addressLowBusModule.busInputs\[32\]
rlabel metal1 15594 7922 15594 7922 0 internalDataflow.addressLowBusModule.busInputs\[33\]
rlabel metal2 17342 8194 17342 8194 0 internalDataflow.addressLowBusModule.busInputs\[34\]
rlabel metal1 14444 6630 14444 6630 0 internalDataflow.addressLowBusModule.busInputs\[35\]
rlabel metal1 16744 7854 16744 7854 0 internalDataflow.addressLowBusModule.busInputs\[36\]
rlabel metal1 15318 10676 15318 10676 0 internalDataflow.addressLowBusModule.busInputs\[37\]
rlabel metal1 16330 8976 16330 8976 0 internalDataflow.addressLowBusModule.busInputs\[38\]
rlabel metal1 14904 7378 14904 7378 0 internalDataflow.addressLowBusModule.busInputs\[39\]
rlabel metal1 7544 20978 7544 20978 0 internalDataflow.dataBusModule.busInputs\[43\]
rlabel metal1 27186 21454 27186 21454 0 internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
rlabel metal1 25852 19754 25852 19754 0 internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
rlabel metal1 29900 22746 29900 22746 0 internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
rlabel metal2 28566 20638 28566 20638 0 internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
rlabel metal1 6486 21114 6486 21114 0 internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
rlabel metal1 16560 12954 16560 12954 0 internalDataflow.stackBusModule.busInputs\[32\]
rlabel metal1 20378 4114 20378 4114 0 internalDataflow.stackBusModule.busInputs\[33\]
rlabel metal2 24886 5678 24886 5678 0 internalDataflow.stackBusModule.busInputs\[34\]
rlabel metal1 16698 6834 16698 6834 0 internalDataflow.stackBusModule.busInputs\[35\]
rlabel metal2 18354 6120 18354 6120 0 internalDataflow.stackBusModule.busInputs\[36\]
rlabel metal1 15686 9962 15686 9962 0 internalDataflow.stackBusModule.busInputs\[37\]
rlabel metal2 18630 7582 18630 7582 0 internalDataflow.stackBusModule.busInputs\[38\]
rlabel metal1 25208 4114 25208 4114 0 internalDataflow.stackBusModule.busInputs\[39\]
rlabel metal1 19596 8398 19596 8398 0 internalDataflow.stackBusModule.busInputs\[40\]
rlabel metal1 21528 4658 21528 4658 0 internalDataflow.stackBusModule.busInputs\[41\]
rlabel metal1 24426 6290 24426 6290 0 internalDataflow.stackBusModule.busInputs\[42\]
rlabel metal1 28244 7310 28244 7310 0 internalDataflow.stackBusModule.busInputs\[43\]
rlabel metal1 21528 5882 21528 5882 0 internalDataflow.stackBusModule.busInputs\[44\]
rlabel metal2 27922 9044 27922 9044 0 internalDataflow.stackBusModule.busInputs\[45\]
rlabel metal1 20240 6834 20240 6834 0 internalDataflow.stackBusModule.busInputs\[46\]
rlabel metal2 26082 5474 26082 5474 0 internalDataflow.stackBusModule.busInputs\[47\]
rlabel metal1 41492 42194 41492 42194 0 interruptRequest
rlabel metal1 6348 25806 6348 25806 0 negEdgeDetector.q1
rlabel metal1 20148 20910 20148 20910 0 net1
rlabel metal1 40618 41174 40618 41174 0 net10
rlabel metal1 20378 6698 20378 6698 0 net100
rlabel metal1 10304 40494 10304 40494 0 net101
rlabel metal1 38180 4522 38180 4522 0 net102
rlabel metal2 26818 9146 26818 9146 0 net103
rlabel metal1 19642 3604 19642 3604 0 net104
rlabel metal1 23598 5542 23598 5542 0 net105
rlabel metal2 15870 6528 15870 6528 0 net106
rlabel metal2 22310 5440 22310 5440 0 net107
rlabel metal1 18262 3434 18262 3434 0 net108
rlabel metal1 18768 6698 18768 6698 0 net109
rlabel metal1 11546 42160 11546 42160 0 net11
rlabel metal1 27922 7378 27922 7378 0 net110
rlabel metal1 6486 23086 6486 23086 0 net111
rlabel metal1 4738 14314 4738 14314 0 net112
rlabel metal1 14858 41242 14858 41242 0 net113
rlabel metal1 18078 4250 18078 4250 0 net114
rlabel metal1 35742 5610 35742 5610 0 net115
rlabel metal1 5382 6290 5382 6290 0 net116
rlabel metal1 10764 5202 10764 5202 0 net117
rlabel metal1 8234 23086 8234 23086 0 net118
rlabel metal1 33028 8534 33028 8534 0 net119
rlabel metal3 17963 21284 17963 21284 0 net12
rlabel metal1 34270 19754 34270 19754 0 net120
rlabel metal1 38456 28186 38456 28186 0 net121
rlabel metal1 30728 6698 30728 6698 0 net122
rlabel metal1 9568 6426 9568 6426 0 net123
rlabel metal1 38686 5678 38686 5678 0 net124
rlabel metal1 35696 8534 35696 8534 0 net125
rlabel metal1 7314 5202 7314 5202 0 net126
rlabel metal1 5612 27098 5612 27098 0 net127
rlabel metal1 21298 4522 21298 4522 0 net128
rlabel metal1 5014 15368 5014 15368 0 net129
rlabel via2 1702 19771 1702 19771 0 net13
rlabel via1 38778 14365 38778 14365 0 net130
rlabel metal1 24794 3604 24794 3604 0 net131
rlabel metal1 37536 8874 37536 8874 0 net132
rlabel metal1 36478 14042 36478 14042 0 net133
rlabel metal1 22586 13328 22586 13328 0 net134
rlabel metal1 17618 18700 17618 18700 0 net135
rlabel metal1 1702 26316 1702 26316 0 net14
rlabel metal1 1518 15674 1518 15674 0 net15
rlabel metal1 38962 2414 38962 2414 0 net16
rlabel metal1 32982 42296 32982 42296 0 net17
rlabel metal1 16698 2414 16698 2414 0 net18
rlabel metal1 40664 7514 40664 7514 0 net19
rlabel metal1 34914 42024 34914 42024 0 net2
rlabel metal1 1518 32504 1518 32504 0 net20
rlabel metal2 36294 4896 36294 4896 0 net21
rlabel metal1 39974 6222 39974 6222 0 net22
rlabel metal1 39974 32878 39974 32878 0 net23
rlabel metal1 1748 17714 1748 17714 0 net24
rlabel metal1 23414 2448 23414 2448 0 net25
rlabel metal1 2484 11526 2484 11526 0 net26
rlabel metal1 31096 6086 31096 6086 0 net27
rlabel metal1 39192 37230 39192 37230 0 net28
rlabel metal2 6118 24004 6118 24004 0 net29
rlabel metal1 5382 7752 5382 7752 0 net3
rlabel metal2 8878 4250 8878 4250 0 net30
rlabel metal2 38226 41797 38226 41797 0 net31
rlabel metal2 5566 4250 5566 4250 0 net32
rlabel metal1 34822 2414 34822 2414 0 net33
rlabel metal1 31832 23562 31832 23562 0 net34
rlabel metal1 40986 13294 40986 13294 0 net35
rlabel metal2 5014 3672 5014 3672 0 net36
rlabel metal1 11592 4726 11592 4726 0 net37
rlabel metal1 3174 36074 3174 36074 0 net38
rlabel metal2 40526 16660 40526 16660 0 net39
rlabel metal1 18078 40494 18078 40494 0 net4
rlabel metal3 19941 2652 19941 2652 0 net40
rlabel metal1 1748 23290 1748 23290 0 net41
rlabel metal1 23966 2346 23966 2346 0 net42
rlabel metal1 40710 20978 40710 20978 0 net43
rlabel metal2 22954 13804 22954 13804 0 net44
rlabel metal1 5796 12070 5796 12070 0 net45
rlabel metal1 17066 15062 17066 15062 0 net46
rlabel metal1 23046 15980 23046 15980 0 net47
rlabel metal1 23506 18190 23506 18190 0 net48
rlabel metal2 17802 18428 17802 18428 0 net49
rlabel metal1 7498 42024 7498 42024 0 net5
rlabel metal2 16974 13022 16974 13022 0 net50
rlabel metal1 18170 19856 18170 19856 0 net51
rlabel metal2 16330 27132 16330 27132 0 net52
rlabel metal1 16238 26350 16238 26350 0 net53
rlabel metal1 9614 32436 9614 32436 0 net54
rlabel metal2 18722 40698 18722 40698 0 net55
rlabel metal1 10258 35700 10258 35700 0 net56
rlabel metal1 11737 5678 11737 5678 0 net57
rlabel metal2 13846 6562 13846 6562 0 net58
rlabel metal1 14865 10642 14865 10642 0 net59
rlabel metal1 4301 2414 4301 2414 0 net6
rlabel metal1 14175 14994 14175 14994 0 net60
rlabel metal1 5842 11288 5842 11288 0 net61
rlabel metal1 22018 3434 22018 3434 0 net62
rlabel metal1 21942 9051 21942 9051 0 net63
rlabel metal1 21988 9554 21988 9554 0 net64
rlabel metal2 31786 19822 31786 19822 0 net65
rlabel metal2 39146 20808 39146 20808 0 net66
rlabel metal2 7130 33014 7130 33014 0 net67
rlabel metal2 13570 40120 13570 40120 0 net68
rlabel metal2 7314 31144 7314 31144 0 net69
rlabel metal3 19849 41684 19849 41684 0 net7
rlabel metal1 37359 29546 37359 29546 0 net70
rlabel metal2 38686 38989 38686 38989 0 net71
rlabel metal2 34638 40052 34638 40052 0 net72
rlabel metal1 33120 41650 33120 41650 0 net73
rlabel metal1 38778 39474 38778 39474 0 net74
rlabel metal1 3220 12070 3220 12070 0 net75
rlabel metal1 13524 40154 13524 40154 0 net76
rlabel metal1 33074 27030 33074 27030 0 net77
rlabel metal1 14766 39610 14766 39610 0 net78
rlabel metal1 11868 6426 11868 6426 0 net79
rlabel metal2 18170 15521 18170 15521 0 net8
rlabel metal1 12558 14314 12558 14314 0 net80
rlabel metal1 9200 37298 9200 37298 0 net81
rlabel metal1 8326 7888 8326 7888 0 net82
rlabel metal1 4876 8466 4876 8466 0 net83
rlabel metal1 5888 32878 5888 32878 0 net84
rlabel metal1 11132 38998 11132 38998 0 net85
rlabel metal1 11270 37128 11270 37128 0 net86
rlabel metal1 40756 16558 40756 16558 0 net87
rlabel metal1 40756 12206 40756 12206 0 net88
rlabel metal1 6854 25806 6854 25806 0 net89
rlabel metal1 5221 41990 5221 41990 0 net9
rlabel metal1 36340 25874 36340 25874 0 net90
rlabel metal1 39514 7786 39514 7786 0 net91
rlabel metal1 34316 26282 34316 26282 0 net92
rlabel metal1 25162 5678 25162 5678 0 net93
rlabel metal1 10304 22406 10304 22406 0 net94
rlabel metal1 11132 21590 11132 21590 0 net95
rlabel metal1 10948 7786 10948 7786 0 net96
rlabel metal1 2852 17578 2852 17578 0 net97
rlabel metal1 5382 22474 5382 22474 0 net98
rlabel metal1 16100 9690 16100 9690 0 net99
rlabel metal1 11178 42194 11178 42194 0 nonMaskableInterrupt
rlabel metal1 15042 42194 15042 42194 0 nrst
rlabel metal1 5658 21488 5658 21488 0 pulse_slower.currentEnableState\[0\]
rlabel metal1 5704 21862 5704 21862 0 pulse_slower.currentEnableState\[1\]
rlabel metal2 15962 20740 15962 20740 0 pulse_slower.nextEnableState\[0\]
rlabel metal1 4600 21114 4600 21114 0 pulse_slower.nextEnableState\[1\]
rlabel metal2 27094 1520 27094 1520 0 readNotWrite
rlabel metal3 820 19788 820 19788 0 ready
rlabel metal3 820 40188 820 40188 0 setOverflow
rlabel metal1 41262 20774 41262 20774 0 sync
<< properties >>
string FIXED_BBOX 0 0 42520 44664
<< end >>
