VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sass_synth
  CLASS BLOCK ;
  FOREIGN sass_synth ;
  ORIGIN 0.000 0.000 ;
  SIZE 367.785 BY 378.505 ;
  PIN beat_led[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END beat_led[0]
  PIN beat_led[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END beat_led[1]
  PIN beat_led[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END beat_led[2]
  PIN beat_led[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 374.505 22.910 378.505 ;
    END
  END beat_led[3]
  PIN beat_led[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 363.785 190.440 367.785 191.040 ;
    END
  END beat_led[4]
  PIN beat_led[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END beat_led[5]
  PIN beat_led[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END beat_led[6]
  PIN beat_led[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END beat_led[7]
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END cs
  PIN hwclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 363.785 44.240 367.785 44.840 ;
    END
  END hwclk
  PIN mode_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 374.505 245.090 378.505 ;
    END
  END mode_out[0]
  PIN mode_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 363.785 13.640 367.785 14.240 ;
    END
  END mode_out[1]
  PIN multi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 374.505 299.830 378.505 ;
    END
  END multi[0]
  PIN multi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 363.785 74.840 367.785 75.440 ;
    END
  END multi[1]
  PIN multi[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 374.505 51.890 378.505 ;
    END
  END multi[2]
  PIN multi[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 363.785 102.040 367.785 102.640 ;
    END
  END multi[3]
  PIN n_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END n_rst
  PIN note1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 363.785 336.640 367.785 337.240 ;
    END
  END note1[0]
  PIN note1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END note1[1]
  PIN note1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END note1[2]
  PIN note1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END note1[3]
  PIN note2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END note2[0]
  PIN note2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END note2[1]
  PIN note2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 363.785 278.840 367.785 279.440 ;
    END
  END note2[2]
  PIN note2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END note2[3]
  PIN note3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 215.830 374.505 216.110 378.505 ;
    END
  END note3[0]
  PIN note3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END note3[1]
  PIN note3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 363.785 363.840 367.785 364.440 ;
    END
  END note3[2]
  PIN note3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 161.090 374.505 161.370 378.505 ;
    END
  END note3[3]
  PIN note4[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 363.785 217.640 367.785 218.240 ;
    END
  END note4[0]
  PIN note4[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 273.790 374.505 274.070 378.505 ;
    END
  END note4[1]
  PIN note4[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END note4[2]
  PIN note4[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END note4[3]
  PIN piano_keys[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 374.505 106.630 378.505 ;
    END
  END piano_keys[0]
  PIN piano_keys[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 363.785 306.040 367.785 306.640 ;
    END
  END piano_keys[10]
  PIN piano_keys[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END piano_keys[11]
  PIN piano_keys[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 363.785 248.240 367.785 248.840 ;
    END
  END piano_keys[12]
  PIN piano_keys[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END piano_keys[13]
  PIN piano_keys[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 374.505 190.350 378.505 ;
    END
  END piano_keys[14]
  PIN piano_keys[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 363.785 132.640 367.785 133.240 ;
    END
  END piano_keys[1]
  PIN piano_keys[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END piano_keys[2]
  PIN piano_keys[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END piano_keys[3]
  PIN piano_keys[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END piano_keys[4]
  PIN piano_keys[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END piano_keys[5]
  PIN piano_keys[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END piano_keys[6]
  PIN piano_keys[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 354.290 374.505 354.570 378.505 ;
    END
  END piano_keys[7]
  PIN piano_keys[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 328.530 374.505 328.810 378.505 ;
    END
  END piano_keys[8]
  PIN piano_keys[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 374.505 80.870 378.505 ;
    END
  END piano_keys[9]
  PIN pwm_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.330 374.505 135.610 378.505 ;
    END
  END pwm_o
  PIN seq_led_on
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END seq_led_on
  PIN seq_play
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END seq_play
  PIN seq_power
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END seq_power
  PIN tempo_select
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 363.785 159.840 367.785 160.440 ;
    END
  END tempo_select
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 367.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 367.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 367.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 367.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 367.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 362.020 367.285 ;
      LAYER met1 ;
        RECT 0.070 9.900 362.870 367.440 ;
      LAYER met2 ;
        RECT 0.100 374.225 22.350 377.245 ;
        RECT 23.190 374.225 51.330 377.245 ;
        RECT 52.170 374.225 80.310 377.245 ;
        RECT 81.150 374.225 106.070 377.245 ;
        RECT 106.910 374.225 135.050 377.245 ;
        RECT 135.890 374.225 160.810 377.245 ;
        RECT 161.650 374.225 189.790 377.245 ;
        RECT 190.630 374.225 215.550 377.245 ;
        RECT 216.390 374.225 244.530 377.245 ;
        RECT 245.370 374.225 273.510 377.245 ;
        RECT 274.350 374.225 299.270 377.245 ;
        RECT 300.110 374.225 328.250 377.245 ;
        RECT 329.090 374.225 354.010 377.245 ;
        RECT 354.850 374.225 362.850 377.245 ;
        RECT 0.100 4.280 362.850 374.225 ;
        RECT 0.650 3.670 25.570 4.280 ;
        RECT 26.410 3.670 54.550 4.280 ;
        RECT 55.390 3.670 80.310 4.280 ;
        RECT 81.150 3.670 109.290 4.280 ;
        RECT 110.130 3.670 135.050 4.280 ;
        RECT 135.890 3.670 164.030 4.280 ;
        RECT 164.870 3.670 189.790 4.280 ;
        RECT 190.630 3.670 218.770 4.280 ;
        RECT 219.610 3.670 247.750 4.280 ;
        RECT 248.590 3.670 273.510 4.280 ;
        RECT 274.350 3.670 302.490 4.280 ;
        RECT 303.330 3.670 328.250 4.280 ;
        RECT 329.090 3.670 357.230 4.280 ;
        RECT 358.070 3.670 362.850 4.280 ;
      LAYER met3 ;
        RECT 4.400 377.040 363.785 377.890 ;
        RECT 3.990 364.840 363.785 377.040 ;
        RECT 3.990 363.440 363.385 364.840 ;
        RECT 3.990 347.840 363.785 363.440 ;
        RECT 4.400 346.440 363.785 347.840 ;
        RECT 3.990 337.640 363.785 346.440 ;
        RECT 3.990 336.240 363.385 337.640 ;
        RECT 3.990 320.640 363.785 336.240 ;
        RECT 4.400 319.240 363.785 320.640 ;
        RECT 3.990 307.040 363.785 319.240 ;
        RECT 3.990 305.640 363.385 307.040 ;
        RECT 3.990 290.040 363.785 305.640 ;
        RECT 4.400 288.640 363.785 290.040 ;
        RECT 3.990 279.840 363.785 288.640 ;
        RECT 3.990 278.440 363.385 279.840 ;
        RECT 3.990 262.840 363.785 278.440 ;
        RECT 4.400 261.440 363.785 262.840 ;
        RECT 3.990 249.240 363.785 261.440 ;
        RECT 3.990 247.840 363.385 249.240 ;
        RECT 3.990 232.240 363.785 247.840 ;
        RECT 4.400 230.840 363.785 232.240 ;
        RECT 3.990 218.640 363.785 230.840 ;
        RECT 3.990 217.240 363.385 218.640 ;
        RECT 3.990 201.640 363.785 217.240 ;
        RECT 4.400 200.240 363.785 201.640 ;
        RECT 3.990 191.440 363.785 200.240 ;
        RECT 3.990 190.040 363.385 191.440 ;
        RECT 3.990 174.440 363.785 190.040 ;
        RECT 4.400 173.040 363.785 174.440 ;
        RECT 3.990 160.840 363.785 173.040 ;
        RECT 3.990 159.440 363.385 160.840 ;
        RECT 3.990 143.840 363.785 159.440 ;
        RECT 4.400 142.440 363.785 143.840 ;
        RECT 3.990 133.640 363.785 142.440 ;
        RECT 3.990 132.240 363.385 133.640 ;
        RECT 3.990 116.640 363.785 132.240 ;
        RECT 4.400 115.240 363.785 116.640 ;
        RECT 3.990 103.040 363.785 115.240 ;
        RECT 3.990 101.640 363.385 103.040 ;
        RECT 3.990 86.040 363.785 101.640 ;
        RECT 4.400 84.640 363.785 86.040 ;
        RECT 3.990 75.840 363.785 84.640 ;
        RECT 3.990 74.440 363.385 75.840 ;
        RECT 3.990 58.840 363.785 74.440 ;
        RECT 4.400 57.440 363.785 58.840 ;
        RECT 3.990 45.240 363.785 57.440 ;
        RECT 3.990 43.840 363.385 45.240 ;
        RECT 3.990 28.240 363.785 43.840 ;
        RECT 4.400 26.840 363.785 28.240 ;
        RECT 3.990 14.640 363.785 26.840 ;
        RECT 3.990 13.240 363.385 14.640 ;
        RECT 3.990 10.715 363.785 13.240 ;
      LAYER met4 ;
        RECT 75.735 27.375 97.440 313.985 ;
        RECT 99.840 27.375 174.240 313.985 ;
        RECT 176.640 27.375 244.425 313.985 ;
  END
END sass_synth
END LIBRARY

