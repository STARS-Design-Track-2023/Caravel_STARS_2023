VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO calculator
  CLASS BLOCK ;
  FOREIGN calculator ;
  ORIGIN 0.000 0.000 ;
  SIZE 137.325 BY 148.045 ;
  PIN blue
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END blue
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 144.045 135.610 148.045 ;
    END
  END clk
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END nrst
  PIN pb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END pb[0]
  PIN pb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 144.045 35.790 148.045 ;
    END
  END pb[1]
  PIN pb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 144.045 58.330 148.045 ;
    END
  END pb[2]
  PIN pb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 133.325 40.840 137.325 41.440 ;
    END
  END pb[3]
  PIN pb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 144.045 116.290 148.045 ;
    END
  END pb[4]
  PIN pb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END pb[5]
  PIN pb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 133.325 85.040 137.325 85.640 ;
    END
  END pb[6]
  PIN pb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 144.045 96.970 148.045 ;
    END
  END pb[7]
  PIN pb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 133.325 0.040 137.325 0.640 ;
    END
  END pb[8]
  PIN pb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END pb[9]
  PIN red
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 144.045 16.470 148.045 ;
    END
  END red
  PIN ss[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END ss[0]
  PIN ss[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END ss[10]
  PIN ss[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END ss[11]
  PIN ss[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END ss[12]
  PIN ss[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 133.325 20.440 137.325 21.040 ;
    END
  END ss[13]
  PIN ss[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END ss[1]
  PIN ss[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 133.325 105.440 137.325 106.040 ;
    END
  END ss[2]
  PIN ss[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 133.325 125.840 137.325 126.440 ;
    END
  END ss[3]
  PIN ss[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END ss[4]
  PIN ss[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 144.045 77.650 148.045 ;
    END
  END ss[5]
  PIN ss[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END ss[6]
  PIN ss[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END ss[7]
  PIN ss[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END ss[8]
  PIN ss[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 133.325 64.640 137.325 65.240 ;
    END
  END ss[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.475 10.640 22.075 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.985 10.640 53.585 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.495 10.640 85.095 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.005 10.640 116.605 136.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 36.230 10.640 37.830 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.740 10.640 69.340 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.250 10.640 100.850 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 130.760 10.640 132.360 136.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 131.560 136.085 ;
      LAYER met1 ;
        RECT 0.070 10.640 135.630 136.240 ;
      LAYER met2 ;
        RECT 0.100 143.765 15.910 146.725 ;
        RECT 16.750 143.765 35.230 146.725 ;
        RECT 36.070 143.765 57.770 146.725 ;
        RECT 58.610 143.765 77.090 146.725 ;
        RECT 77.930 143.765 96.410 146.725 ;
        RECT 97.250 143.765 115.730 146.725 ;
        RECT 116.570 143.765 135.050 146.725 ;
        RECT 0.100 4.280 135.600 143.765 ;
        RECT 0.650 0.155 19.130 4.280 ;
        RECT 19.970 0.155 38.450 4.280 ;
        RECT 39.290 0.155 57.770 4.280 ;
        RECT 58.610 0.155 77.090 4.280 ;
        RECT 77.930 0.155 99.630 4.280 ;
        RECT 100.470 0.155 118.950 4.280 ;
        RECT 119.790 0.155 135.600 4.280 ;
      LAYER met3 ;
        RECT 4.400 145.840 134.010 146.705 ;
        RECT 3.990 126.840 134.010 145.840 ;
        RECT 4.400 125.440 132.925 126.840 ;
        RECT 3.990 106.440 134.010 125.440 ;
        RECT 4.400 105.040 132.925 106.440 ;
        RECT 3.990 86.040 134.010 105.040 ;
        RECT 3.990 84.640 132.925 86.040 ;
        RECT 3.990 82.640 134.010 84.640 ;
        RECT 4.400 81.240 134.010 82.640 ;
        RECT 3.990 65.640 134.010 81.240 ;
        RECT 3.990 64.240 132.925 65.640 ;
        RECT 3.990 62.240 134.010 64.240 ;
        RECT 4.400 60.840 134.010 62.240 ;
        RECT 3.990 41.840 134.010 60.840 ;
        RECT 4.400 40.440 132.925 41.840 ;
        RECT 3.990 21.440 134.010 40.440 ;
        RECT 4.400 20.040 132.925 21.440 ;
        RECT 3.990 1.040 134.010 20.040 ;
        RECT 3.990 0.175 132.925 1.040 ;
      LAYER met4 ;
        RECT 32.495 74.295 32.825 123.585 ;
  END
END calculator
END LIBRARY

