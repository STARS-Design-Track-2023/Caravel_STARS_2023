magic
tech sky130A
magscale 1 2
timestamp 1691553077
<< obsli1 >>
rect 1104 2159 147016 147985
<< obsm1 >>
rect 14 2128 147076 148016
<< metal2 >>
rect 2594 149514 2650 150314
rect 20626 149514 20682 150314
rect 38658 149514 38714 150314
rect 57334 149514 57390 150314
rect 75366 149514 75422 150314
rect 93398 149514 93454 150314
rect 111430 149514 111486 150314
rect 129462 149514 129518 150314
rect 147494 149514 147550 150314
rect 18 0 74 800
rect 18050 0 18106 800
rect 36082 0 36138 800
rect 54114 0 54170 800
rect 72146 0 72202 800
rect 90178 0 90234 800
rect 108854 0 108910 800
rect 126886 0 126942 800
rect 144918 0 144974 800
<< obsm2 >>
rect 20 149458 2538 149514
rect 2706 149458 20570 149514
rect 20738 149458 38602 149514
rect 38770 149458 57278 149514
rect 57446 149458 75310 149514
rect 75478 149458 93342 149514
rect 93510 149458 111374 149514
rect 111542 149458 129406 149514
rect 129574 149458 147438 149514
rect 20 856 147550 149458
rect 130 734 17994 856
rect 18162 734 36026 856
rect 36194 734 54058 856
rect 54226 734 72090 856
rect 72258 734 90122 856
rect 90290 734 108798 856
rect 108966 734 126830 856
rect 126998 734 144862 856
rect 145030 734 147550 856
<< metal3 >>
rect 0 133968 800 134088
rect 147370 130568 148170 130688
rect 0 114928 800 115048
rect 147370 111528 148170 111648
rect 0 95208 800 95328
rect 147370 92488 148170 92608
rect 0 76168 800 76288
rect 147370 73448 148170 73568
rect 0 57128 800 57248
rect 147370 54408 148170 54528
rect 0 38088 800 38208
rect 147370 34688 148170 34808
rect 0 19048 800 19168
rect 147370 15648 148170 15768
<< obsm3 >>
rect 800 134168 147555 148001
rect 880 133888 147555 134168
rect 800 130768 147555 133888
rect 800 130488 147290 130768
rect 800 115128 147555 130488
rect 880 114848 147555 115128
rect 800 111728 147555 114848
rect 800 111448 147290 111728
rect 800 95408 147555 111448
rect 880 95128 147555 95408
rect 800 92688 147555 95128
rect 800 92408 147290 92688
rect 800 76368 147555 92408
rect 880 76088 147555 76368
rect 800 73648 147555 76088
rect 800 73368 147290 73648
rect 800 57328 147555 73368
rect 880 57048 147555 57328
rect 800 54608 147555 57048
rect 800 54328 147290 54608
rect 800 38288 147555 54328
rect 880 38008 147555 38288
rect 800 34888 147555 38008
rect 800 34608 147290 34888
rect 800 19248 147555 34608
rect 880 18968 147555 19248
rect 800 15848 147555 18968
rect 800 15568 147290 15848
rect 800 2143 147555 15568
<< metal4 >>
rect 4208 2128 4528 148016
rect 4868 2128 5188 148016
rect 34928 2128 35248 148016
rect 35588 2128 35908 148016
rect 65648 2128 65968 148016
rect 66308 2128 66628 148016
rect 96368 2128 96688 148016
rect 97028 2128 97348 148016
rect 127088 2128 127408 148016
rect 127748 2128 128068 148016
<< obsm4 >>
rect 4659 3979 4788 147797
rect 5268 3979 34848 147797
rect 35328 3979 35508 147797
rect 35988 3979 65568 147797
rect 66048 3979 66228 147797
rect 66708 3979 96288 147797
rect 96768 3979 96948 147797
rect 97428 3979 127008 147797
rect 127488 3979 127668 147797
rect 128148 3979 143093 147797
<< metal5 >>
rect 1056 128550 147064 128870
rect 1056 127890 147064 128210
rect 1056 97914 147064 98234
rect 1056 97254 147064 97574
rect 1056 67278 147064 67598
rect 1056 66618 147064 66938
rect 1056 36642 147064 36962
rect 1056 35982 147064 36302
rect 1056 6006 147064 6326
rect 1056 5346 147064 5666
<< obsm5 >>
rect 26796 129190 137332 141260
rect 26796 98554 137332 127570
rect 26796 67918 137332 96934
rect 26796 37282 137332 66298
rect 26796 21940 137332 35662
<< labels >>
rlabel metal4 s 4868 2128 5188 148016 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 148016 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 148016 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97028 2128 97348 148016 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127748 2128 128068 148016 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 147064 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 147064 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 147064 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 97914 147064 98234 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 128550 147064 128870 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 148016 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 148016 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 148016 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 148016 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 148016 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 147064 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 147064 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 147064 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 147064 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 127890 147064 128210 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 147494 149514 147550 150314 6 clk
port 3 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 color[0]
port 4 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 color[10]
port 5 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 color[11]
port 6 nsew signal output
rlabel metal2 s 38658 149514 38714 150314 6 color[12]
port 7 nsew signal output
rlabel metal2 s 93398 149514 93454 150314 6 color[13]
port 8 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 color[14]
port 9 nsew signal output
rlabel metal3 s 147370 73448 148170 73568 6 color[15]
port 10 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 color[16]
port 11 nsew signal output
rlabel metal3 s 147370 92488 148170 92608 6 color[17]
port 12 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 color[18]
port 13 nsew signal output
rlabel metal2 s 18 0 74 800 6 color[19]
port 14 nsew signal output
rlabel metal2 s 111430 149514 111486 150314 6 color[1]
port 15 nsew signal output
rlabel metal2 s 129462 149514 129518 150314 6 color[20]
port 16 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 color[21]
port 17 nsew signal output
rlabel metal3 s 147370 15648 148170 15768 6 color[22]
port 18 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 color[23]
port 19 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 color[2]
port 20 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 color[3]
port 21 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 color[4]
port 22 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 color[5]
port 23 nsew signal output
rlabel metal2 s 20626 149514 20682 150314 6 color[6]
port 24 nsew signal output
rlabel metal3 s 147370 34688 148170 34808 6 color[7]
port 25 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 color[8]
port 26 nsew signal output
rlabel metal3 s 147370 111528 148170 111648 6 color[9]
port 27 nsew signal output
rlabel metal3 s 147370 130568 148170 130688 6 cs
port 28 nsew signal input
rlabel metal2 s 57334 149514 57390 150314 6 is_mandelbrot
port 29 nsew signal output
rlabel metal2 s 75366 149514 75422 150314 6 nrst
port 30 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 spi_clk
port 31 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 spi_data
port 32 nsew signal input
rlabel metal2 s 2594 149514 2650 150314 6 spi_en
port 33 nsew signal input
rlabel metal3 s 147370 54408 148170 54528 6 valid_out
port 34 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 148170 150314
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 67395098
string GDS_FILE /home/designer-25/CUP/openlane/DigiDoggs/runs/23_08_08_20_14/results/signoff/pushing_pixels.magic.gds
string GDS_START 1510688
<< end >>

