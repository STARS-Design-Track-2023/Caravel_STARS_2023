* NGSPICE file created from sass_synth.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt sass_synth beat_led[0] beat_led[1] beat_led[2] beat_led[3] beat_led[4] beat_led[5]
+ beat_led[6] beat_led[7] cs hwclk mode_out[0] mode_out[1] multi[0] multi[1] multi[2]
+ multi[3] n_rst note1[0] note1[1] note1[2] note1[3] note2[0] note2[1] note2[2] note2[3]
+ note3[0] note3[1] note3[2] note3[3] note4[0] note4[1] note4[2] note4[3] piano_keys[0]
+ piano_keys[10] piano_keys[11] piano_keys[12] piano_keys[13] piano_keys[14] piano_keys[1]
+ piano_keys[2] piano_keys[3] piano_keys[4] piano_keys[5] piano_keys[6] piano_keys[7]
+ piano_keys[8] piano_keys[9] pwm_o seq_led_on seq_play seq_power tempo_select vccd1
+ vssd1
X_7963_ clknet_leaf_21_hwclk net430 net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_6914_ _3184_ _3186_ vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__nor2_1
X_7894_ clknet_leaf_1_hwclk net594 net70 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6845_ net772 _1469_ _2864_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__mux2_1
X_3988_ pm.count\[1\] pm.count\[0\] net547 vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__and3_1
X_6776_ sound1.sdiv.Q\[3\] _2895_ sound1.sdiv.next_dived net392 vssd1 vssd1 vccd1
+ vccd1 _0144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5727_ net239 _2182_ _2185_ net401 _2194_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5658_ sound4.sdiv.A\[12\] _2062_ _2069_ _2140_ _2067_ vssd1 vssd1 vccd1 vccd1 _2141_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4609_ _0983_ _0978_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5589_ sound4.divisor_m\[11\] _2071_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7328_ _3486_ _3490_ _3497_ vssd1 vssd1 vccd1 vccd1 _3498_ sky130_fd_sc_hd__nand3_1
Xhold340 net895 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold351 sound4.count_m\[9\] vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold362 net912 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__dlymetal6s2s_1
X_7259_ _2843_ _1618_ _3436_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__o21ai_1
Xhold384 sound1.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 sound1.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 sound2.count_m\[17\] vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4960_ _1470_ _1506_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__nand2_1
X_4891_ sound2.count\[4\] _1441_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__xor2_1
X_3911_ _0575_ net63 vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__nor2_8
XFILLER_0_117_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6630_ sound1.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3842_ _0478_ _0485_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6561_ _2927_ _2929_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5512_ _0550_ net168 vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[2\] sky130_fd_sc_hd__nor2_1
X_3773_ inputcont.INTERNAL_SYNCED_I\[5\] vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
X_8300_ clknet_leaf_66_hwclk _0400_ net80 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6492_ net782 _2875_ _2864_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8231_ clknet_leaf_33_hwclk sound3.osc.next_count\[12\] net88 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[12\] sky130_fd_sc_hd__dfrtp_2
X_5443_ _1779_ _1936_ _1948_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8162_ clknet_leaf_42_hwclk net213 net98 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_5374_ sound4.count\[6\] _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__xor2_1
X_7113_ net520 _3168_ sound2.sdiv.next_dived _3364_ vssd1 vssd1 vccd1 vccd1 _0231_
+ sky130_fd_sc_hd__a22o_1
X_4325_ _0894_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nand2_1
X_8093_ clknet_leaf_77_hwclk net551 net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_7044_ _3302_ _3303_ vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__or2_1
X_4256_ _0838_ _0813_ _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__and3b_1
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4187_ seq.tempo_select.state\[1\] seq.clk_div.count\[12\] _0779_ seq.clk_div.count\[6\]
+ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7946_ clknet_leaf_32_hwclk _0109_ net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7877_ clknet_leaf_96_hwclk net110 net68 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_sync\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6828_ net482 _2857_ _3128_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6759_ net590 net888 net596 vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold170 sound3.sdiv.Q\[23\] vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _0320_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 sound1.sdiv.Q\[14\] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5090_ _1584_ _1595_ _1602_ _1620_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__or4_1
X_4110_ seq.player_6.state\[0\] _0729_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4041_ _0675_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__buf_12
X_5992_ _2402_ _2427_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__and2_1
X_7800_ clknet_leaf_7_hwclk oct.next_state\[1\] net71 vssd1 vssd1 vccd1 vccd1 oct.state\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_87_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7731_ clknet_leaf_84_hwclk net240 net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_4943_ _1004_ _1321_ _1338_ _1158_ _1493_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__o221a_1
X_7662_ _3722_ _2156_ vssd1 vssd1 vccd1 vccd1 _3723_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6613_ _2903_ _2977_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__and2_1
X_4874_ _0683_ _1323_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3825_ _0485_ _0501_ _0492_ _0502_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__a211o_1
X_7593_ _3675_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_1
X_6544_ _2909_ _2915_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6475_ net709 _2005_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8214_ clknet_leaf_46_hwclk _0335_ net98 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5426_ net414 _1779_ _1936_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[0\] sky130_fd_sc_hd__nand3_1
XFILLER_0_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5357_ sound4.count\[4\] _1866_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8145_ clknet_leaf_82_hwclk _0266_ net74 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8076_ clknet_leaf_79_hwclk _0218_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_4308_ seq.beat\[1\] seq.beat\[0\] seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__nor3b_1
X_5288_ _1773_ _1775_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__or2_1
X_4239_ seq.clk_div.count\[8\] _0824_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__nand2_1
X_7027_ _3277_ _3280_ _3288_ vssd1 vssd1 vccd1 vccd1 _3289_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7929_ clknet_leaf_10_hwclk _0092_ net83 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4590_ _0680_ _0958_ _1154_ _0950_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6260_ sound1.sdiv.Q\[5\] _0579_ _2690_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5211_ net702 _1732_ _1721_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__o21ai_1
X_6191_ sound2.sdiv.Q\[0\] sound2.sdiv.Q\[1\] sound2.sdiv.Q\[2\] _0578_ _2499_ vssd1
+ vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__o311a_1
X_5142_ _0948_ _1578_ _1617_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__o211a_2
X_5073_ _1018_ _1556_ _1603_ _0971_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__a22o_1
X_4024_ _0581_ _0583_ _0671_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__o21a_1
X_5975_ _2409_ sound1.divisor_m\[4\] _2410_ sound1.divisor_m\[3\] vssd1 vssd1 vccd1
+ vccd1 _2411_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7714_ _3756_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4926_ _0993_ _1383_ _1471_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4857_ _0685_ _1323_ _1338_ _1165_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__o221a_1
X_7645_ _2069_ _2140_ vssd1 vssd1 vccd1 vccd1 _3711_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7576_ _3665_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__clkbuf_1
X_3808_ _0473_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6527_ _2897_ sound1.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4788_ net38 _1316_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__nand2_4
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6458_ net464 _2836_ _2854_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__a21o_1
X_6389_ net711 _2812_ _2808_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5409_ net59 _1784_ _1781_ _1038_ _1769_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__o221a_1
X_8128_ clknet_leaf_83_hwclk _0249_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8059_ clknet_leaf_92_hwclk _0201_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5760_ _2207_ _2212_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ net985 _1272_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2_1
X_5691_ _2169_ _2170_ _2171_ _2172_ _2173_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7430_ _3586_ _3588_ vssd1 vssd1 vccd1 vccd1 _3589_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4642_ _0695_ _0977_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__or2_4
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7361_ _3448_ _3526_ vssd1 vssd1 vccd1 vccd1 _3527_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4573_ _1136_ _1137_ _1143_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold703 seq.player_8.state\[2\] vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7292_ sound3.divisor_m\[3\] sound3.divisor_m\[2\] sound3.divisor_m\[1\] sound3.divisor_m\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3465_ sky130_fd_sc_hd__or4_1
X_6312_ _2740_ _2742_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__xor2_1
Xhold725 seq.player_1.state\[1\] vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold714 rate_clk.count\[0\] vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 sound2.count\[17\] vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6243_ _2672_ _2675_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__xnor2_1
Xhold758 sound3.count\[0\] vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold769 sound4.count\[12\] vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 sound4.count\[8\] vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__dlygate4sd3_1
X_6174_ _2374_ _2574_ _2608_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__a21o_1
X_5125_ _1642_ _1649_ _1655_ sound3.count\[2\] vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5056_ _0677_ _1574_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__or2_1
X_4007_ net805 net118 _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5958_ _2377_ _2380_ _2388_ _2393_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4909_ sound2.count\[16\] _1459_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5889_ sound4.count_m\[13\] _2142_ sound4.divisor_m\[13\] _2324_ vssd1 vssd1 vccd1
+ vccd1 _2325_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7628_ _2132_ _3697_ vssd1 vssd1 vccd1 vccd1 _3699_ sky130_fd_sc_hd__or2b_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7559_ _3655_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold30 sound3.sdiv.Q\[15\] vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 sound2.sdiv.Q\[22\] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 _0369_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 rate_clk.count\[2\] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold52 _0267_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 sound3.count_m\[3\] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 _0153_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_5 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6930_ _1311_ _3201_ vssd1 vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6861_ net759 _3147_ _3142_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5812_ _2256_ _2257_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6792_ net376 _2893_ _0867_ net371 _2849_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5743_ sound4.count\[15\] _2201_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5674_ _2154_ _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__nor2_1
X_7413_ _3570_ _3572_ vssd1 vssd1 vccd1 vccd1 _3574_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4625_ _0959_ _1082_ _1192_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7344_ _3510_ _3511_ _3503_ _3507_ vssd1 vssd1 vccd1 vccd1 _3512_ sky130_fd_sc_hd__o211ai_1
Xhold500 _0345_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold511 _0041_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _1025_ _1038_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__nor2_4
Xhold522 sound1.sdiv.Q\[5\] vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 seq.player_1.state\[0\] vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold533 seq.player_4.state\[0\] vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 sound1.sdiv.A\[23\] vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 pm.count\[4\] vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__dlygate4sd3_1
X_7275_ sound3.divisor_m\[2\] _3449_ vssd1 vssd1 vccd1 vccd1 _3450_ sky130_fd_sc_hd__xnor2_1
Xhold577 sound3.count\[12\] vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 sound2.sdiv.Q\[5\] vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4487_ _0685_ _0977_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__nand2_4
Xhold599 pm.current_waveform\[5\] vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ sound1.sdiv.Q\[5\] _2293_ _2658_ _2292_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__o2bb2a_1
X_6157_ sound2.sdiv.Q\[2\] _0578_ _2591_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__and3_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _1189_ _1565_ _1637_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__o211a_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ sound3.count_m\[11\] vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__inv_2
X_5039_ _1569_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_1_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 multi[0] sky130_fd_sc_hd__clkbuf_4
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 note3[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4410_ _0980_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5390_ _0973_ _1777_ _1800_ _1016_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4341_ seq.player_5.state\[0\] _0890_ _0892_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4272_ _0850_ _0813_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__and3b_1
X_7060_ sound2.divisor_m\[17\] _3308_ _3177_ vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__o21a_1
X_6011_ sound2.count_m\[15\] _2446_ sound2.count_m\[14\] _2440_ vssd1 vssd1 vccd1
+ vccd1 _2447_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7962_ clknet_leaf_23_hwclk _0125_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6913_ sound2.divisor_m\[3\] _3185_ vssd1 vssd1 vccd1 vccd1 _3186_ sky130_fd_sc_hd__xnor2_1
X_7893_ clknet_leaf_7_hwclk net657 net72 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6844_ _3137_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
X_3987_ net535 net197 vssd1 vssd1 vccd1 vccd1 pm.next_count\[1\] sky130_fd_sc_hd__xor2_1
X_6775_ _2435_ _0866_ _2588_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5726_ net409 _2186_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5657_ _2073_ _2138_ _2139_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__a21o_1
X_4608_ _0943_ _1028_ _1175_ _0976_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5588_ sound4.divisor_m\[10\] _2030_ _2036_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7327_ _3495_ _3496_ vssd1 vssd1 vccd1 vccd1 _3497_ sky130_fd_sc_hd__nand2_1
Xhold330 _0356_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 sound4.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _0944_ _1012_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__nor2_2
Xhold341 sound2.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7258_ _2543_ _2005_ vssd1 vssd1 vccd1 vccd1 _3436_ sky130_fd_sc_hd__or2_1
Xhold363 sound1.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _0108_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold385 sound2.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _0186_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6209_ _2640_ _2642_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__xor2_1
X_7189_ net412 _3132_ _3395_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3910_ _0577_ vssd1 vssd1 vccd1 vccd1 sound3.sdiv.next_start sky130_fd_sc_hd__inv_2
X_4890_ _1139_ _1327_ _1435_ _1440_ _1317_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_86_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ _0500_ _0491_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6560_ _2927_ _2929_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3772_ inputcont.INTERNAL_SYNCED_I\[9\] inputcont.INTERNAL_SYNCED_I\[10\] _0454_
+ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5511_ rate_clk.count\[1\] net154 net167 vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__a21oi_1
X_6491_ _1157_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8230_ clknet_leaf_33_hwclk sound3.osc.next_count\[11\] net88 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[11\] sky130_fd_sc_hd__dfrtp_1
X_5442_ sound4.count\[4\] _1944_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8161_ clknet_leaf_30_hwclk net196 net91 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_5373_ _1880_ _1883_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7112_ _3360_ _3363_ vssd1 vssd1 vccd1 vccd1 _3364_ sky130_fd_sc_hd__xor2_1
X_8092_ clknet_leaf_84_hwclk _0234_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4324_ seq.player_6.state\[0\] seq.player_6.state\[1\] seq.player_6.state\[2\] seq.player_6.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__or4_1
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7043_ _3299_ _3301_ vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__and2_1
X_4255_ seq.clk_div.count\[12\] _0835_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__or2_1
X_4186_ seq.clk_div.count\[10\] vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7945_ clknet_leaf_12_hwclk net500 net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7876_ clknet_leaf_96_hwclk net217 net64 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_6827_ sound2.count\[13\] _2855_ vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_81_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_6758_ _2890_ _3103_ _3104_ _2894_ net590 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6689_ sound1.divisor_m\[17\] _3036_ _2903_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__o21a_1
X_5709_ _0576_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__buf_6
XFILLER_0_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8359_ clknet_leaf_61_hwclk sound4.osc.next_count\[17\] net78 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[17\] sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_96_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_hwclk
+ sky130_fd_sc_hd__clkbuf_16
Xhold171 sound1.sdiv.Q\[24\] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold160 sound2.count_m\[5\] vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 sound1.count_m\[4\] vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 sound2.count_m\[15\] vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_34_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_hwclk clknet_0_hwclk vssd1 vssd1 vccd1 vccd1 clknet_3_4__leaf_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _0676_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__nor2_8
X_5991_ _2400_ _2401_ _2397_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__a21o_1
X_4942_ _1129_ _1347_ _1343_ _1014_ _1427_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__o221a_1
X_7730_ clknet_leaf_64_hwclk _0015_ net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_7661_ _2053_ _3720_ vssd1 vssd1 vccd1 vccd1 _3722_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6612_ sound1.divisor_m\[9\] sound1.divisor_m\[8\] sound1.divisor_m\[7\] _2948_ vssd1
+ vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4873_ sound2.count\[14\] _1422_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3824_ _0481_ _0482_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__nand2_2
X_7592_ net774 _3674_ _2186_ vssd1 vssd1 vccd1 vccd1 _3675_ sky130_fd_sc_hd__mux2_1
X_6543_ _2913_ _2914_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6474_ _2865_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8213_ clknet_leaf_46_hwclk net568 net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5425_ _1935_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5356_ sound4.count\[4\] _1866_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__nand2_1
X_8144_ clknet_leaf_82_hwclk _0265_ net74 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_4307_ _0876_ _0877_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__nand2_1
X_5287_ _1146_ _1777_ _1792_ _1134_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__o221a_1
X_8075_ clknet_leaf_80_hwclk _0217_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_4238_ seq.clk_div.count\[8\] _0824_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__or2_1
X_7026_ _3286_ _3287_ vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4169_ net931 inputcont.INTERNAL_SYNCED_I\[0\] vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7928_ clknet_leaf_11_hwclk _0091_ net88 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7859_ clknet_leaf_96_hwclk seq.clk_div.next_count\[16\] net64 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5210_ net875 _1732_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6190_ sound2.sdiv.Q\[4\] _0578_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5141_ _1001_ _1570_ _1668_ _1671_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__o211a_1
X_5072_ _1556_ _1557_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4023_ _0588_ _0584_ _0585_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__or3b_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5974_ sound1.count_m\[2\] vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__inv_2
X_7713_ net748 net33 _0645_ vssd1 vssd1 vccd1 vccd1 _3756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ _1095_ _1343_ _1472_ _1473_ _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4856_ _1126_ _1347_ _1341_ _1166_ _1406_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7644_ _2069_ _2140_ vssd1 vssd1 vccd1 vccd1 _3710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7575_ net758 _3664_ _3419_ vssd1 vssd1 vccd1 vccd1 _3665_ sky130_fd_sc_hd__mux2_1
X_3807_ _0477_ _0478_ _0479_ _0485_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__and4b_1
X_6526_ net488 _2895_ sound1.sdiv.next_dived _2899_ vssd1 vssd1 vccd1 vccd1 _0109_
+ sky130_fd_sc_hd__a22o_1
X_4787_ _1337_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6457_ sound1.count\[16\] _2201_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6388_ _2439_ _2581_ _2805_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__mux2_1
X_5408_ _0954_ _1777_ _1792_ _0985_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__o22ai_1
X_8127_ clknet_leaf_84_hwclk _0248_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_5339_ _1844_ _1845_ _1849_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__or3_2
X_8058_ clknet_leaf_92_hwclk _0200_ net67 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_7009_ _3164_ _3271_ _3272_ _3174_ net238 vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _1274_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_5690_ sound4.sdiv.A\[23\] _2038_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4641_ _1210_ _0869_ _0965_ _1011_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7360_ sound3.divisor_m\[10\] _3515_ vssd1 vssd1 vccd1 vccd1 _3526_ sky130_fd_sc_hd__or2_1
X_4572_ _0981_ _1138_ _1139_ _0969_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7291_ sound3.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _3464_ sky130_fd_sc_hd__inv_2
Xhold715 pm.count\[0\] vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
X_6311_ _2703_ _2707_ _2741_ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__a21o_1
Xhold726 _0776_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 sound2.count\[8\] vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 sound2.count\[15\] vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 sound3.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__dlygate4sd3_1
X_6242_ sound4.sdiv.Q\[5\] _2290_ _2674_ _2292_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__o2bb2a_1
Xhold759 sound1.count\[5\] vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6173_ _2507_ _2573_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__and2_1
X_5124_ _1005_ _1578_ _1550_ _1017_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__o221a_2
X_5055_ _1057_ _1567_ _1565_ _1056_ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__o221a_1
X_4006_ net869 vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5957_ _2389_ _2390_ _2391_ _2392_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__and4b_1
XFILLER_0_48_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4908_ _1010_ _1456_ _1458_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7627_ _3697_ _2132_ vssd1 vssd1 vccd1 vccd1 _3698_ sky130_fd_sc_hd__or2b_1
X_5888_ sound4.count_m\[12\] vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4839_ _0954_ _1347_ _1345_ _1182_ _1389_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7558_ net893 _1859_ _3419_ vssd1 vssd1 vccd1 vccd1 _3655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7489_ _3437_ _3637_ _3639_ _3440_ net655 vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__a32o_1
X_6509_ net789 _2886_ _2864_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold31 _0355_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 sound3.sdiv.Q\[22\] vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 sound3.sdiv.Q\[24\] vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0263_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 _2001_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 sound3.count_m\[1\] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _0271_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 sound4.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_6 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6860_ _1412_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__inv_2
X_5811_ _2248_ _2252_ _2247_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__a21boi_1
X_6791_ net371 _2893_ _0867_ sound1.sdiv.Q\[17\] _2848_ vssd1 vssd1 vccd1 vccd1 _0159_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5742_ net305 _2182_ _2185_ net368 _2202_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5673_ _2155_ _2049_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7412_ _3570_ _3572_ vssd1 vssd1 vccd1 vccd1 _3573_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4624_ _1193_ _0967_ _0943_ _1158_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__o221a_1
X_7343_ sound3.sdiv.A\[8\] _3509_ vssd1 vssd1 vccd1 vccd1 _3511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4555_ _0959_ net59 vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__nor2_4
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold501 seq.player_3.state\[0\] vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 sound3.sdiv.A\[20\] vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 sound1.sdiv.A\[20\] vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 sound3.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold534 seq.player_4.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__dlygate4sd3_1
X_7274_ sound3.divisor_m\[1\] sound3.divisor_m\[0\] _3448_ vssd1 vssd1 vccd1 vccd1
+ _3449_ sky130_fd_sc_hd__o21a_1
Xhold567 pm.current_waveform\[0\] vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _1748_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
X_4486_ _0695_ _0970_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold556 seq.clk_div.count\[17\] vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6225_ _2620_ _2657_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__xnor2_1
Xhold589 sound2.count\[7\] vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
X_6156_ sound2.sdiv.Q\[0\] sound2.sdiv.Q\[1\] _0578_ _2499_ vssd1 vssd1 vccd1 vccd1
+ _2591_ sky130_fd_sc_hd__o211a_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _1204_ _1553_ _1580_ _1199_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _2521_ sound3.divisor_m\[14\] sound3.divisor_m\[13\] _2522_ vssd1 vssd1 vccd1
+ vccd1 _2523_ sky130_fd_sc_hd__a22o_1
X_5038_ _1563_ _1568_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6989_ _3164_ _3253_ _3254_ _3174_ net307 vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 beat_led[0] sky130_fd_sc_hd__clkbuf_4
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 multi[1] sky130_fd_sc_hd__clkbuf_4
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 note3[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4340_ seq.player_6.state\[0\] _0894_ _0896_ _0910_ vssd1 vssd1 vccd1 vccd1 _0911_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4271_ seq.clk_div.count\[16\] _0847_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6010_ sound2.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7961_ clknet_leaf_21_hwclk _0124_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7892_ clknet_leaf_4_hwclk net114 net71 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6912_ sound2.divisor_m\[2\] sound2.divisor_m\[1\] sound2.divisor_m\[0\] _3177_ vssd1
+ vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__o31a_1
XFILLER_0_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6843_ net889 _3136_ _2864_ vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3986_ net197 vssd1 vssd1 vccd1 vccd1 pm.next_count\[0\] sky130_fd_sc_hd__inv_2
X_6774_ net536 sound1.sdiv.next_dived _2436_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5725_ net401 _2182_ _2185_ sound4.sdiv.Q\[13\] _2193_ vssd1 vssd1 vccd1 vccd1 _0014_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5656_ _2070_ _2072_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4607_ _0954_ _0994_ _0992_ _1129_ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold320 _0378_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__dlygate4sd3_1
X_5587_ net493 vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold353 sound3.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__dlygate4sd3_1
X_7326_ _3491_ _3494_ vssd1 vssd1 vccd1 vccd1 _3496_ sky130_fd_sc_hd__nand2_1
X_4538_ _0677_ _1084_ _1090_ _0952_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__o22a_1
Xhold331 sound2.count_m\[14\] vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 sound2.count\[13\] vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__dlygate4sd3_1
X_7257_ _3435_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__clkbuf_1
Xhold375 sound3.count\[4\] vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _0207_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _0674_ _0977_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__nor2_2
Xhold364 sound4.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 sound3.count_m\[9\] vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ sound4.sdiv.Q\[2\] _2641_ _2582_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__a21o_1
X_7188_ sound3.count\[8\] _2863_ vssd1 vssd1 vccd1 vccd1 _3395_ sky130_fd_sc_hd__and2_1
X_6139_ _2374_ _2574_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3840_ inputcont.INTERNAL_SYNCED_I\[3\] _0502_ _0512_ _0513_ vssd1 vssd1 vccd1 vccd1
+ _0514_ sky130_fd_sc_hd__a211o_1
X_3771_ inputcont.INTERNAL_SYNCED_I\[8\] _0443_ _0444_ vssd1 vssd1 vccd1 vccd1 _0454_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5510_ net174 net154 vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6490_ _2005_ _1196_ _2874_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ sound4.count\[4\] _1944_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__nand2_1
X_8160_ clknet_leaf_31_hwclk _0281_ net91 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_5372_ _0679_ net59 _1784_ _1882_ _1778_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__o311a_1
XFILLER_0_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7111_ _3343_ _3361_ _3362_ _3352_ vssd1 vssd1 vccd1 vccd1 _3363_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8091_ clknet_leaf_77_hwclk _0233_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_4323_ select1.sequencer_on _0893_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7042_ _3299_ _3301_ vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__nor2_1
X_4254_ seq.clk_div.count\[12\] _0835_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_0_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_4185_ seq.clk_div.count\[18\] vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7944_ clknet_leaf_6_hwclk _0107_ net83 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7875_ clknet_leaf_96_hwclk net112 net68 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6826_ net426 _2857_ _3127_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6757_ sound1.sdiv.C\[1\] sound1.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5708_ net564 _2183_ sound4.sdiv.next_dived net632 vssd1 vssd1 vccd1 vccd1 _0007_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3969_ net33 _0632_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__nor2_2
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6688_ sound1.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5639_ sound4.divisor_m\[1\] _2121_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__xnor2_1
X_8358_ clknet_leaf_61_hwclk sound4.osc.next_count\[16\] net94 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7309_ _3468_ _3471_ _3479_ vssd1 vssd1 vccd1 vccd1 _3481_ sky130_fd_sc_hd__or3b_1
Xhold150 _0155_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _0174_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _0074_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _0166_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
X_8289_ clknet_leaf_63_hwclk _0389_ net78 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold183 _0184_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5990_ _2382_ _2425_ _2389_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _1020_ _1333_ _1345_ _1083_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__o221a_1
X_7660_ _3681_ _3720_ _3721_ _2184_ net266 vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__a32o_1
X_4872_ sound2.count\[14\] _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6611_ _2962_ _2963_ _2975_ _2966_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__o211a_1
X_3823_ _0479_ _0478_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7591_ _1817_ vssd1 vssd1 vccd1 vccd1 _3674_ sky130_fd_sc_hd__inv_2
X_6542_ _2910_ _2912_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6473_ net765 _2862_ _2864_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8212_ clknet_leaf_46_hwclk _0333_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5424_ _1861_ _1886_ _1934_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__or3_1
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8143_ clknet_leaf_82_hwclk _0264_ net74 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5355_ _0696_ _1792_ _1794_ _1140_ _1865_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4306_ seq.player_2.state\[0\] seq.player_2.state\[1\] seq.player_2.state\[2\] seq.player_2.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__or4_1
X_5286_ _1154_ _1794_ _1796_ _1042_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8074_ clknet_leaf_80_hwclk _0216_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_4237_ _0824_ _0825_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[7\] sky130_fd_sc_hd__nor2_1
X_7025_ _3282_ _3285_ vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4168_ _0766_ _0765_ _0768_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_2.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_4099_ net900 net848 seq.player_7.state\[3\] _0722_ _0700_ vssd1 vssd1 vccd1 vccd1
+ _0723_ sky130_fd_sc_hd__a311o_1
X_7927_ clknet_leaf_10_hwclk _0090_ net88 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7858_ clknet_leaf_96_hwclk seq.clk_div.next_count\[15\] net64 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6809_ sound2.count\[4\] _2855_ vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7789_ clknet_leaf_89_hwclk net119 net68 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5140_ _0973_ _1553_ _1574_ _0979_ _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__o221a_1
X_5071_ sound3.count\[4\] _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_80_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_4022_ _0594_ _0669_ _0596_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5973_ sound1.count_m\[3\] vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_95_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7712_ _3755_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__clkbuf_1
X_4924_ _1041_ _1323_ _1327_ _1096_ _1474_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4855_ _1159_ _1343_ _1333_ _0997_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__o22a_1
X_7643_ _3681_ _3708_ _3709_ _2184_ net272 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7574_ _1897_ vssd1 vssd1 vccd1 vccd1 _3664_ sky130_fd_sc_hd__inv_2
X_3806_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__buf_2
X_4786_ net38 _1325_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6525_ _2891_ _2898_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_6456_ net407 _2836_ _2853_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6387_ _2811_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_1
X_5407_ _1912_ _1914_ _1917_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__or3b_1
XFILLER_0_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8126_ clknet_leaf_61_hwclk _0247_ net94 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5338_ _1125_ _1796_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__o21ai_1
X_8057_ clknet_leaf_80_hwclk _0199_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[11\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_48_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_7008_ _3259_ _3262_ _3270_ vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__o21bai_2
X_5269_ net46 _1770_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__nor2_2
XFILLER_0_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _0909_ _0937_ _1138_ _0974_ _0688_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__o32a_1
XFILLER_0_56_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6310_ _2698_ _2702_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__and2_1
X_4571_ _1000_ _1140_ _1141_ _0976_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7290_ _3461_ _3462_ net450 _3463_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__a2bb2o_1
Xhold716 inputcont.u1.ff_intermediate\[7\] vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold705 sound3.count\[16\] vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 seq.player_1.next_state\[3\] vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold749 sound3.count\[12\] vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__dlygate4sd3_1
X_6241_ _2639_ _2673_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__xor2_1
Xhold738 seq.player_6.state\[1\] vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__dlygate4sd3_1
X_6172_ _2585_ _2606_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5123_ _1025_ _1028_ _1553_ _1650_ _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__o311a_1
X_5054_ _0959_ _1133_ _1553_ _1578_ _0983_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__o32a_1
X_4005_ net143 _0655_ pm.count\[8\] vssd1 vssd1 vccd1 vccd1 pm.next_count\[8\] sky130_fd_sc_hd__a21boi_1
X_5956_ sound1.divisor_m\[9\] sound1.count_m\[8\] vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__or2b_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5887_ _2322_ sound4.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__or2_1
X_4907_ _0688_ _1418_ _1317_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4838_ _1129_ _1341_ _1336_ _1175_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__o22a_1
X_7626_ _2133_ _2093_ vssd1 vssd1 vccd1 vccd1 _3697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7557_ net175 _2843_ _2206_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4769_ _0499_ _1319_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__nor2_2
X_7488_ _3622_ _3631_ _3638_ _3636_ vssd1 vssd1 vccd1 vccd1 _3639_ sky130_fd_sc_hd__a31o_1
X_6508_ _1219_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__inv_2
X_6439_ _1073_ _2843_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8109_ clknet_leaf_93_hwclk sound2.osc.next_count\[10\] net66 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[10\] sky130_fd_sc_hd__dfrtp_1
Xhold21 _0362_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 seq.encode.keys_sync\[1\] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 sound2.sdiv.Q\[9\] vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold54 _0364_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 sound2.sdiv.Q\[20\] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 rate_clk.next_count\[2\] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 sound3.count_m\[16\] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold76 sound4.sdiv.Q\[26\] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 inputcont.INTERNAL_SYNCED_I\[7\] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5810_ _2254_ _2255_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__nand2_1
X_6790_ sound1.sdiv.Q\[17\] _2893_ _0867_ net138 _2847_ vssd1 vssd1 vccd1 vccd1 _0158_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5741_ sound4.count\[14\] _2201_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7411_ sound3.divisor_m\[16\] _3571_ vssd1 vssd1 vccd1 vccd1 _3572_ sky130_fd_sc_hd__xnor2_1
X_5672_ _2046_ _2048_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4623_ _0992_ _1028_ _1020_ _0990_ _1130_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7342_ sound3.sdiv.A\[8\] _3509_ vssd1 vssd1 vccd1 vccd1 _3510_ sky130_fd_sc_hd__and2_1
Xhold502 wave_comb.u1.A\[10\] vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4554_ _1124_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__clkbuf_4
X_7273_ sound3.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _3448_ sky130_fd_sc_hd__inv_4
Xhold513 seq.encode.keys_edge_det\[1\] vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 seq.player_2.state\[0\] vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold524 sound4.count_m\[15\] vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 sound1.sdiv.A\[21\] vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 wave_comb.u1.Q\[1\] vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ sound1.sdiv.Q\[3\] _2656_ _2621_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__a21oi_1
X_4485_ _0678_ _1055_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__nand2_4
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold546 seq.player_7.state\[0\] vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold557 sound4.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6155_ _2279_ _2586_ _2589_ _2289_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__a2bb2o_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ sound3.count_m\[12\] vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__inv_2
X_5106_ _1200_ _1567_ _1550_ _0686_ _1636_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ net45 _1555_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6988_ _3233_ _3237_ _3251_ _3241_ _3250_ vssd1 vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__a311o_1
X_5939_ sound1.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7609_ _2120_ _2125_ vssd1 vssd1 vccd1 vccd1 _3685_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 multi[2] sky130_fd_sc_hd__buf_2
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 beat_led[1] sky130_fd_sc_hd__clkbuf_4
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 note3[2] sky130_fd_sc_hd__buf_2
XFILLER_0_101_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ net972 _0847_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7960_ clknet_leaf_21_hwclk _0123_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_6911_ sound2.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__inv_2
X_7891_ clknet_leaf_2_hwclk net111 net70 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6842_ _1404_ vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6773_ _0866_ _3114_ _2277_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3985_ _0646_ vssd1 vssd1 vccd1 vccd1 wave_comb.u1.next_dived sky130_fd_sc_hd__buf_4
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5724_ sound4.count\[6\] _2186_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5655_ _2079_ _2137_ _2077_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4606_ _0950_ _0996_ _1176_ _0981_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7325_ _3491_ _3494_ vssd1 vssd1 vccd1 vccd1 _3495_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold310 sound4.count\[0\] vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5586_ _2067_ _2068_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__nor2_1
Xhold321 sound3.sdiv.A\[23\] vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _0683_ _0981_ _0992_ _1052_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__o211a_1
Xhold332 _0183_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 rate_clk.count\[6\] vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold365 sound3.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 sound1.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__dlygate4sd3_1
X_7256_ net904 _1604_ _3419_ vssd1 vssd1 vccd1 vccd1 _3435_ sky130_fd_sc_hd__mux2_1
X_4468_ _1019_ _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__or2_4
Xhold354 seq.player_2.state\[3\] vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 seq.player_4.state\[3\] vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 _0277_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__dlygate4sd3_1
X_7187_ net320 _3132_ _3394_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__a21o_1
X_6207_ _0576_ _2370_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__and2_1
X_6138_ _2507_ _2573_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__xor2_1
X_4399_ _0686_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__nand2_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _2439_ _2504_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__xnor2_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3770_ _0441_ _0445_ _0447_ _0452_ _0453_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__o2111ai_4
XFILLER_0_42_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5440_ _1947_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5371_ _1057_ _1792_ _1794_ _1063_ _1881_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7110_ sound2.sdiv.A\[22\] sound2.sdiv.A\[21\] _3329_ vssd1 vssd1 vccd1 vccd1 _3362_
+ sky130_fd_sc_hd__o21ai_1
X_8090_ clknet_leaf_76_hwclk _0232_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_4322_ seq.beat\[3\] seq.encode.play _0874_ inputcont.INTERNAL_SYNCED_I\[5\] vssd1
+ vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7041_ sound2.divisor_m\[16\] _3300_ vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__xnor2_1
X_4253_ _0837_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
X_4184_ _0777_ _0778_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[1\] sky130_fd_sc_hd__nor2_1
X_7943_ clknet_leaf_15_hwclk _0106_ net83 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7874_ clknet_leaf_99_hwclk net109 net65 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6825_ net823 _2855_ vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6756_ net590 sound1.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3968_ _0630_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__or2_2
X_5707_ sound4.sdiv.Q\[6\] _2183_ sound4.sdiv.next_dived net600 vssd1 vssd1 vccd1
+ vccd1 _0006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6687_ net431 _2895_ sound1.sdiv.next_dived _3044_ vssd1 vssd1 vccd1 vccd1 _0125_
+ sky130_fd_sc_hd__a22o_1
X_3899_ _0554_ _0568_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__nand2_8
X_5638_ sound4.sdiv.A\[26\] sound4.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8357_ clknet_leaf_62_hwclk sound4.osc.next_count\[15\] net79 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[15\] sky130_fd_sc_hd__dfrtp_2
X_5569_ sound4.divisor_m\[16\] _2051_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7308_ _3468_ _3471_ _3479_ vssd1 vssd1 vccd1 vccd1 _3480_ sky130_fd_sc_hd__o21bai_2
Xhold162 sound4.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 sound2.count_m\[11\] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 sound2.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 sound3.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 sound1.count_m\[11\] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
X_8288_ clknet_leaf_63_hwclk _0388_ net78 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[2\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold195 sound2.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
X_7239_ _3424_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__clkbuf_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _1028_ _1341_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4871_ _0695_ _1417_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__o21ai_2
X_6610_ _2969_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3822_ _0443_ _0444_ inputcont.INTERNAL_SYNCED_I\[8\] vssd1 vssd1 vccd1 vccd1 _0500_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7590_ _3673_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__clkbuf_1
X_6541_ _2910_ _2912_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6472_ _2863_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8211_ clknet_leaf_46_hwclk _0332_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5423_ _1911_ _1918_ _1925_ _1933_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__or4b_1
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5354_ _1138_ _1769_ _1778_ _1864_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__o211a_1
X_8142_ clknet_leaf_81_hwclk net146 net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4305_ select1.sequencer_on _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__and2_1
X_8073_ clknet_leaf_80_hwclk _0215_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_5285_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__clkbuf_4
X_4236_ net678 _0822_ _0813_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7024_ _3282_ _3285_ vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__or2_1
X_4167_ net729 seq.player_2.state\[2\] _0762_ net458 vssd1 vssd1 vccd1 vccd1 _0768_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4098_ seq.player_7.state\[0\] _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__and2_1
X_7926_ clknet_leaf_32_hwclk _0089_ net87 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7857_ clknet_leaf_94_hwclk seq.clk_div.next_count\[14\] net66 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[14\] sky130_fd_sc_hd__dfrtp_1
X_6808_ net602 _2857_ _3118_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7788_ clknet_leaf_9_hwclk net495 net2 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_6739_ _0866_ _3089_ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout90 net92 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_6
XFILLER_0_83_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5070_ _1135_ _1550_ _1570_ _1140_ _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__o221a_1
X_4021_ _0668_ _0602_ _0592_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5972_ _2407_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7711_ net735 net32 _0645_ vssd1 vssd1 vccd1 vccd1 _3755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4923_ _1347_ _1336_ _0960_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7642_ _2138_ _3707_ vssd1 vssd1 vccd1 vccd1 _3709_ sky130_fd_sc_hd__or2b_1
X_4854_ _0677_ _1336_ _1345_ _1077_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7573_ _3663_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3805_ _0480_ _0481_ _0482_ _0483_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and4_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4785_ _1335_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__clkbuf_4
X_6524_ sound1.sdiv.A\[0\] _2897_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6455_ sound1.count\[15\] _2201_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6386_ net691 _2810_ _2808_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__mux2_1
X_5406_ sound4.count\[17\] _1222_ _1913_ _1915_ _1916_ vssd1 vssd1 vccd1 vccd1 _1917_
+ sky130_fd_sc_hd__o311a_1
X_8125_ clknet_leaf_61_hwclk _0246_ net94 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5337_ _1199_ _1800_ _1846_ _1847_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__o211a_1
X_5268_ _1778_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__buf_4
X_8056_ clknet_leaf_92_hwclk _0198_ net67 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_7007_ _3259_ _3262_ _3270_ vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__or3b_1
X_4219_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__buf_4
X_5199_ _1727_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7909_ clknet_leaf_11_hwclk net544 net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4570_ _1038_ _1034_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__nor2_2
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 sound4.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 rate_clk.count\[1\] vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 sound4.count\[11\] vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6240_ sound4.sdiv.Q\[3\] _2641_ _2642_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__a21o_1
Xhold739 seq.player_6.next_state\[3\] vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__dlygate4sd3_1
X_6171_ _2600_ _2605_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5122_ _1011_ _1559_ _1572_ _1020_ _1652_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5053_ sound3.count\[0\] _1583_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__xor2_1
X_4004_ _0657_ _0655_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[7\] sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_100_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5955_ sound1.count_m\[9\] sound1.divisor_m\[10\] vssd1 vssd1 vccd1 vccd1 _2391_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5886_ sound4.count_m\[16\] vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__inv_2
X_4906_ _1324_ _1333_ _1055_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7625_ _3695_ _3696_ net415 _2183_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a2bb2o_1
X_4837_ sound2.count\[10\] _1387_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7556_ net246 _2843_ _2205_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a21o_1
X_4768_ _0507_ _1312_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__nand2_1
X_7487_ _3630_ _3623_ _3627_ vssd1 vssd1 vccd1 vccd1 _3638_ sky130_fd_sc_hd__or3b_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6507_ _2885_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__clkbuf_1
X_4699_ net951 _1263_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6438_ net304 _2836_ _2844_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6369_ _2794_ _2796_ net52 vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__or3_1
X_8108_ clknet_leaf_93_hwclk sound2.osc.next_count\[9\] net66 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[9\] sky130_fd_sc_hd__dfrtp_1
Xhold22 seq.encode.inter_keys\[1\] vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 inputcont.u1.ff_intermediate\[3\] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 sound1.count_m\[18\] vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 _0261_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dlygate4sd3_1
X_8039_ clknet_leaf_92_hwclk _0181_ net67 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold33 _0250_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 _0284_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 sound3.count_m\[18\] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 sound1.sdiv.Q\[7\] vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_1
Xhold77 _0027_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_94_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5740_ _0575_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7410_ sound3.divisor_m\[15\] _3561_ _3448_ vssd1 vssd1 vccd1 vccd1 _3571_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_47_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5671_ _2053_ _2153_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__or2_1
X_4622_ _1107_ _1100_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__or2_2
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7341_ sound3.divisor_m\[9\] _3508_ vssd1 vssd1 vccd1 vccd1 _3509_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4553_ _0683_ _1034_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7272_ sound3.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _3447_ sky130_fd_sc_hd__inv_2
Xhold514 wave_comb.u1.A\[3\] vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 seq.player_2.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 sound2.sdiv.A\[21\] vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4484_ _0676_ _0695_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__or2_4
Xhold525 _0382_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 pm.current_waveform\[8\] vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _0579_ _2434_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__and2_1
Xhold558 sound4.sdiv.A\[20\] vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6154_ _2587_ _2588_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ sound3.count_m\[13\] vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__inv_2
X_5105_ _0683_ _1107_ _1570_ _1562_ _1198_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__o32a_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6987_ _3250_ _3252_ vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__nand2_1
X_5938_ _2289_ _2372_ _2373_ _2290_ sound4.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 _2374_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5869_ _2291_ _2305_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7608_ net456 _2183_ sound4.sdiv.next_dived _3684_ vssd1 vssd1 vccd1 vccd1 _0406_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7539_ net419 _3403_ _2187_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput34 net56 vssd1 vssd1 vccd1 vccd1 note1[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 beat_led[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 note3[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6910_ _3176_ _3179_ vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__or2_1
X_7890_ clknet_leaf_1_hwclk net546 net70 vssd1 vssd1 vccd1 vccd1 seq.encode.play sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6841_ _3135_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6772_ _3098_ _3100_ _3113_ _3096_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _0645_ _0571_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5723_ sound4.sdiv.Q\[13\] _2182_ _2185_ net405 _2192_ vssd1 vssd1 vccd1 vccd1 _0013_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5654_ _2083_ _2135_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__a21boi_1
X_4605_ _0996_ _1019_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7324_ sound3.divisor_m\[7\] _3493_ vssd1 vssd1 vccd1 vccd1 _3494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold300 sound1.sdiv.A\[8\] vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 sound4.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__dlygate4sd3_1
X_5585_ _2063_ _2065_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold322 sound2.count_m\[12\] vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 sound2.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 rate_clk.next_count\[6\] vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__dlygate4sd3_1
X_4536_ _0685_ _0684_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__nor2_8
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7255_ _3434_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
Xhold366 sound1.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 seq.player_2.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 seq.player_4.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__dlygate4sd3_1
X_4467_ _0676_ _0695_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__nor2_8
Xhold399 sound3.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__dlygate4sd3_1
X_7186_ _1642_ _2843_ vssd1 vssd1 vccd1 vccd1 _3394_ sky130_fd_sc_hd__nor2_1
X_6206_ sound4.sdiv.Q\[3\] _0576_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4398_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__buf_4
Xhold388 sound2.count_m\[9\] vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__dlygate4sd3_1
X_6137_ _2289_ _2571_ _2572_ _2301_ sound3.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 _2573_
+ sky130_fd_sc_hd__a32o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _2289_ _2502_ _2503_ _2295_ sound2.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 _2504_
+ sky130_fd_sc_hd__a32o_1
X_5019_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5370_ _1056_ _1777_ _1800_ _1053_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4321_ _0890_ _0891_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7040_ sound2.divisor_m\[15\] sound2.divisor_m\[14\] _3283_ _3177_ vssd1 vssd1 vccd1
+ vccd1 _3300_ sky130_fd_sc_hd__o31a_1
X_4252_ _0835_ _0813_ _0836_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__and3b_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4183_ net557 net140 _0719_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7942_ clknet_leaf_18_hwclk _0105_ net84 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7873_ clknet_leaf_96_hwclk net120 net68 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_6824_ net244 _2857_ _3126_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__a21o_1
X_6755_ _3102_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3967_ _0607_ _0629_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__and2_1
X_5706_ net600 _2183_ sound4.sdiv.next_dived net610 vssd1 vssd1 vccd1 vccd1 _0005_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6686_ _3042_ _3043_ vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3898_ sound4.sdiv.dived _0557_ _0560_ sound2.sdiv.dived _0567_ vssd1 vssd1 vccd1
+ vccd1 _0568_ sky130_fd_sc_hd__a221o_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5637_ _2117_ _2119_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8356_ clknet_leaf_85_hwclk sound4.osc.next_count\[14\] net79 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[14\] sky130_fd_sc_hd__dfrtp_1
X_5568_ _2036_ _2033_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__and2_1
X_7307_ _3477_ _3478_ vssd1 vssd1 vccd1 vccd1 _3479_ sky130_fd_sc_hd__nand2_1
X_4519_ _0967_ _1025_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__or2_1
Xhold152 sound4.sdiv.Q\[24\] vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__dlygate4sd3_1
X_8287_ clknet_leaf_62_hwclk _0387_ net78 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[1\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold141 _0180_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _0176_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold163 sound3.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__dlygate4sd3_1
X_7238_ net793 _1690_ _3419_ vssd1 vssd1 vccd1 vccd1 _3424_ sky130_fd_sc_hd__mux2_1
Xhold185 _0081_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 sound1.sdiv.Q\[23\] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _1779_ _1936_ _1992_ _1993_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__and4_1
Xhold196 sound3.count_m\[12\] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
X_7169_ net271 _3167_ _1311_ net273 _3133_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__a221o_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4870_ _1111_ _1325_ _1334_ _1058_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3821_ _0499_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__inv_2
X_6540_ sound1.divisor_m\[3\] _2911_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6471_ _0575_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__clkbuf_8
X_8210_ clknet_leaf_47_hwclk _0331_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_5422_ sound4.count\[1\] _1931_ _1909_ sound4.count\[11\] _1932_ vssd1 vssd1 vccd1
+ vccd1 _1933_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5353_ _1135_ _1784_ _1796_ _1141_ _1863_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__o221a_1
X_8141_ clknet_leaf_91_hwclk _0262_ net67 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4304_ _0702_ seq.encode.play _0874_ inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1
+ vccd1 vccd1 _0875_ sky130_fd_sc_hd__a31o_1
X_8072_ clknet_leaf_78_hwclk _0214_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5284_ _1782_ _1771_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__or2_1
X_4235_ net939 seq.clk_div.count\[7\] _0819_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__and3_1
X_7023_ _2441_ _3284_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__xnor2_1
X_4166_ _0766_ _0765_ _0767_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_2.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4097_ seq.encode.keys_edge_det\[8\] inputcont.INTERNAL_SYNCED_I\[6\] vssd1 vssd1
+ vccd1 vccd1 _0721_ sky130_fd_sc_hd__and2b_1
X_7925_ clknet_leaf_12_hwclk net160 net85 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7856_ clknet_leaf_94_hwclk seq.clk_div.next_count\[13\] net66 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[13\] sky130_fd_sc_hd__dfrtp_1
X_6807_ _1318_ _2843_ vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4999_ _1535_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_7787_ clknet_leaf_8_hwclk net123 net70 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_6738_ net54 _3087_ _3084_ _3085_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6669_ sound1.divisor_m\[15\] sound1.divisor_m\[14\] _3011_ vssd1 vssd1 vccd1 vccd1
+ _3028_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8339_ clknet_leaf_55_hwclk _0439_ net96 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.M\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout91 net92 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_8
Xfanout80 net82 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_6
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4020_ _0599_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5971_ sound1.count_m\[17\] _2405_ sound1.count_m\[16\] _2406_ vssd1 vssd1 vccd1
+ vccd1 _2407_ sky130_fd_sc_hd__o22a_1
X_7710_ _3754_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4922_ _1101_ _1333_ _1345_ _1097_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7641_ _3707_ _2138_ vssd1 vssd1 vccd1 vccd1 _3708_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4853_ _1398_ _1400_ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__and3_2
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7572_ net762 _1884_ _3419_ vssd1 vssd1 vccd1 vccd1 _3663_ sky130_fd_sc_hd__mux2_1
X_3804_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[3\]
+ inputcont.INTERNAL_SYNCED_I\[2\] inputcont.INTERNAL_SYNCED_I\[4\] vssd1 vssd1 vccd1
+ vccd1 _0483_ sky130_fd_sc_hd__o41ai_4
X_4784_ _1330_ _1334_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__or2_1
X_6523_ sound1.divisor_m\[1\] _2896_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6454_ net331 _2836_ _2852_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5405_ sound4.count\[18\] _1778_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6385_ _2294_ _2310_ _2805_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8124_ clknet_leaf_61_hwclk net609 net94 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_5336_ _1198_ _1769_ _1777_ _1189_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8055_ clknet_leaf_91_hwclk _0197_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_5267_ _1772_ _1773_ _1777_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__nand3_4
X_7006_ _3268_ _3269_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__nand2_1
X_4218_ _0719_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__and2_1
X_5198_ _1721_ _1725_ _1726_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__and3_1
X_4149_ seq.player_3.state\[0\] seq.player_3.state\[1\] _0753_ vssd1 vssd1 vccd1 vccd1
+ _0756_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7908_ clknet_leaf_11_hwclk net184 net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_7839_ clknet_leaf_47_hwclk _0062_ net101 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold707 sound3.count\[13\] vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 sound4.count\[3\] vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold729 seq.player_5.state\[1\] vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6170_ sound3.sdiv.Q\[3\] _2301_ _2603_ _2604_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__o2bb2a_1
X_5121_ _0997_ _1562_ _1565_ _0973_ _1651_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5052_ _1554_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__nand2_1
X_4003_ net143 vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5954_ sound1.count_m\[8\] sound1.divisor_m\[9\] vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5885_ _2313_ sound4.divisor_m\[4\] _2317_ _2319_ _2320_ vssd1 vssd1 vccd1 vccd1
+ _2321_ sky130_fd_sc_hd__a2111oi_1
X_4905_ _1450_ _1334_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7624_ _2099_ _2131_ _2185_ vssd1 vssd1 vccd1 vccd1 _3696_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4836_ _1107_ net59 _1322_ _1380_ _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__o311a_2
X_7555_ net442 _2843_ _2204_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6506_ net798 _2884_ _2864_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__mux2_1
X_4767_ net881 vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__inv_2
X_7486_ _3629_ _3630_ _3631_ _3636_ vssd1 vssd1 vccd1 vccd1 _3637_ sky130_fd_sc_hd__o211ai_1
X_4698_ _1265_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6437_ _1237_ _2843_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__nor2_1
X_6368_ _2762_ _2791_ _2792_ _2793_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__nor4_1
XFILLER_0_3_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8107_ clknet_leaf_95_hwclk sound2.osc.next_count\[8\] net66 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[8\] sky130_fd_sc_hd__dfrtp_2
X_5319_ sound4.count\[8\] _1829_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__and2_1
X_6299_ _2728_ _2729_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__xnor2_1
Xhold23 wave_comb.u1.Q\[10\] vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 inputcont.INTERNAL_OCTAVE_INPUT vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _0088_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 sound1.sdiv.Q\[16\] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 sound4.sdiv.Q\[11\] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dlygate4sd3_1
X_8038_ clknet_leaf_92_hwclk net245 net66 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold67 _0286_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 sound1.count_m\[7\] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _0149_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _2050_ _2052_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4621_ _0939_ _1014_ _1188_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7340_ sound3.divisor_m\[8\] _3448_ _3501_ vssd1 vssd1 vccd1 vccd1 _3508_ sky130_fd_sc_hd__a21o_1
X_4552_ _0679_ _0971_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7271_ _3442_ sound3.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _3446_ sky130_fd_sc_hd__or2b_1
Xhold504 sound2.sdiv.Q\[4\] vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ _0679_ _0950_ net59 _1053_ _0992_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o32a_1
Xhold515 sound2.count_m\[10\] vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold526 sound4.divisor_m\[9\] vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 pm.next_pwm_o vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 sound1.sdiv.A\[19\] vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold537 sound3.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ wave_comb.u1.next_start _2654_ _2655_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6153_ net392 _0579_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ sound3.divisor_m\[1\] _2517_ _2518_ _2519_ vssd1 vssd1 vccd1 vccd1 _2520_
+ sky130_fd_sc_hd__o211ai_1
X_5104_ _1181_ _1559_ _1578_ _1028_ _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__o221a_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _1560_ _1551_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__or2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6986_ _3233_ _3237_ _3251_ _3241_ vssd1 vssd1 vccd1 vccd1 _3252_ sky130_fd_sc_hd__a31o_1
X_5937_ sound4.sdiv.Q\[1\] _2181_ _2370_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__nand3_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5868_ _2303_ _2304_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__nor2_1
X_7607_ _2123_ _3682_ vssd1 vssd1 vccd1 vccd1 _3684_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5799_ wave_comb.u1.next_dived _2245_ _2246_ _0573_ net257 vssd1 vssd1 vccd1 vccd1
+ _0035_ sky130_fd_sc_hd__a32o_1
X_4819_ _1318_ _1352_ _1360_ sound2.count\[12\] _1369_ vssd1 vssd1 vccd1 vccd1 _1370_
+ sky130_fd_sc_hd__a221o_1
X_7538_ sound3.sdiv.Q\[27\] _3440_ _3437_ net132 vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__a22o_1
X_7469_ net982 _3595_ vssd1 vssd1 vccd1 vccd1 _3622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 beat_led[3] sky130_fd_sc_hd__clkbuf_4
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 note4[0] sky130_fd_sc_hd__buf_2
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 note1[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7__f_hwclk clknet_0_hwclk vssd1 vssd1 vccd1 vccd1 clknet_3_7__leaf_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6840_ net917 _1477_ _2864_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6771_ net987 sound1.divisor_m\[17\] sound1.sdiv.A\[26\] _3036_ vssd1 vssd1 vccd1
+ vccd1 _3113_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3983_ _0644_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5722_ sound4.count\[5\] _2186_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5653_ sound4.sdiv.A\[8\] _2082_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4604_ _1001_ _1028_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5584_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__inv_2
X_7323_ _3448_ _3492_ vssd1 vssd1 vccd1 vccd1 _3493_ sky130_fd_sc_hd__and2_1
X_4535_ sound1.count\[2\] _1032_ _1072_ sound1.count\[6\] _1105_ vssd1 vssd1 vccd1
+ vccd1 _1106_ sky130_fd_sc_hd__a221o_1
Xhold301 sound4.sdiv.Q\[12\] vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold334 sound3.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 sound3.sdiv.Q\[8\] vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold323 sound3.count\[13\] vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 sound3.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__dlygate4sd3_1
X_7254_ net767 _3433_ _3419_ vssd1 vssd1 vccd1 vccd1 _3434_ sky130_fd_sc_hd__mux2_1
X_4466_ _0992_ _1033_ _1035_ _0981_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__o221a_1
Xhold378 sound2.count_m\[13\] vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 sound2.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 sound2.count\[4\] vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7185_ net269 _3132_ _3393_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a21o_1
X_6205_ sound4.sdiv.Q\[4\] _0576_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4397_ _0918_ _0941_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__or2_1
Xhold389 sound4.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6136_ _2570_ _2275_ sound3.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _2500_ _2276_ _2499_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__or3b_1
X_5018_ _0540_ _1548_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__or2_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6969_ _3224_ _3228_ _3235_ vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_93_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4320_ seq.player_5.state\[0\] seq.player_5.state\[1\] seq.player_5.state\[2\] seq.player_5.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__or4_1
X_4251_ seq.clk_div.count\[11\] _0832_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4182_ net557 net948 vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7941_ clknet_leaf_18_hwclk _0104_ net84 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7872_ clknet_leaf_89_hwclk net115 net68 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6823_ net887 _2855_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__and2_1
X_6754_ _0867_ _2893_ net779 vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3966_ _0607_ _0629_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__nor2_2
X_6685_ _3031_ _3035_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__nand2_1
X_5705_ net610 _2183_ sound4.sdiv.next_dived net633 vssd1 vssd1 vccd1 vccd1 _0004_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3897_ sound3.sdiv.dived _0563_ _0566_ sound1.sdiv.dived vssd1 vssd1 vccd1 vccd1
+ _0567_ sky130_fd_sc_hd__a22o_1
X_5636_ sound4.divisor_m\[2\] _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5567_ sound4.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__inv_2
X_8355_ clknet_leaf_85_hwclk sound4.osc.next_count\[13\] net79 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[13\] sky130_fd_sc_hd__dfrtp_2
X_7306_ _3474_ _3476_ vssd1 vssd1 vccd1 vccd1 _3478_ sky130_fd_sc_hd__nand2_1
Xhold131 sound3.sdiv.A\[8\] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 wave_comb.u1.A\[7\] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 sound1.count_m\[5\] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _1075_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__nand2_1
X_8286_ clknet_leaf_60_hwclk _0386_ net94 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_5498_ sound4.count\[16\] _1988_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__or2_1
Xhold142 sound4.count_m\[17\] vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__dlygate4sd3_1
X_7237_ _3423_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__clkbuf_1
Xhold175 _0165_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _1018_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__or2_4
Xhold186 net827 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_1
XFILLER_0_0_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold164 sound2.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _0280_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7168_ net273 _3167_ _1311_ net453 _3131_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__a221o_1
X_6119_ _2551_ sound3.count_m\[0\] _2552_ _2553_ _2554_ vssd1 vssd1 vccd1 vccd1 _2555_
+ sky130_fd_sc_hd__o2111a_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _3350_ _3351_ _3352_ vssd1 vssd1 vccd1 vccd1 _3353_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3820_ _0472_ _0487_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__o21ba_4
XFILLER_0_55_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6470_ _1032_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5421_ sound4.count\[1\] _1931_ _1891_ sound4.count\[15\] vssd1 vssd1 vccd1 vccd1
+ _1932_ sky130_fd_sc_hd__o2bb2a_1
X_5352_ _1127_ _1777_ _1800_ _1126_ _1862_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__o221a_1
X_8140_ clknet_leaf_91_hwclk net148 net67 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8071_ clknet_leaf_78_hwclk _0213_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4303_ seq.beat\[0\] seq.beat\[2\] seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__nor3b_1
X_7022_ _3177_ _3283_ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__nand2_1
X_5283_ _1793_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4234_ _0822_ _0823_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[6\] sky130_fd_sc_hd__nor2_1
X_4165_ net775 _0764_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4096_ net860 _0716_ _0720_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_8.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_7924_ clknet_leaf_12_hwclk net334 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_7855_ clknet_leaf_94_hwclk seq.clk_div.next_count\[12\] net66 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[12\] sky130_fd_sc_hd__dfrtp_2
X_6806_ net645 _2857_ _3117_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4998_ _1533_ _1534_ _1504_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__and3b_1
X_7786_ clknet_leaf_9_hwclk net623 net70 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6737_ _3084_ _3085_ net54 _3087_ vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3949_ _0459_ _0481_ inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1 vccd1 vccd1 _0613_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6668_ sound1.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6599_ net404 _2895_ _2964_ _2965_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__a22o_1
X_5619_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8338_ clknet_leaf_57_hwclk _0438_ net96 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.M\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8269_ clknet_leaf_63_hwclk net178 net78 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout92 net103 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_8
Xfanout81 net82 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_8
Xfanout70 net72 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_8
XFILLER_0_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ sound1.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__inv_2
X_4921_ _1341_ _1322_ _0948_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4852_ _1005_ _1322_ _1339_ _0964_ _1402_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__o221a_1
X_7640_ _2139_ _2073_ vssd1 vssd1 vccd1 vccd1 _3707_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3803_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__o21ai_4
X_7571_ _3662_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__clkbuf_1
X_4783_ net41 _1313_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__nand2_2
X_6522_ sound1.sdiv.A\[26\] sound1.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6453_ sound1.count\[14\] _2201_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5404_ sound4.count\[18\] _1778_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6384_ _2809_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__clkbuf_1
X_8123_ clknet_leaf_61_hwclk net572 net94 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5335_ _1204_ _1786_ _1790_ _1014_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8054_ clknet_leaf_81_hwclk _0196_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_5266_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__buf_6
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _0786_ _0795_ _0801_ _0810_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__or4bb_1
X_7005_ _3265_ _3267_ vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__nand2_1
X_5197_ net862 sound3.count\[1\] sound3.count\[2\] vssd1 vssd1 vccd1 vccd1 _1726_
+ sky130_fd_sc_hd__nand3_1
X_4148_ net605 _0753_ _0755_ vssd1 vssd1 vccd1 vccd1 seq.player_3.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_4079_ _0709_ vssd1 vssd1 vccd1 vccd1 seq_power_on sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7907_ clknet_leaf_11_hwclk net311 net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7838_ clknet_leaf_47_hwclk _0061_ net101 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7769_ clknet_leaf_47_hwclk net144 net102 vssd1 vssd1 vccd1 vccd1 pm.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold708 sound4.sdiv.C\[5\] vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_1
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold719 sound2.count\[12\] vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5120_ _1016_ _1580_ _1570_ _1024_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__o22a_1
X_5051_ _0996_ _1025_ _1559_ _1577_ _1581_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__o311a_1
X_4002_ _0655_ net570 vssd1 vssd1 vccd1 vccd1 pm.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_79_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5953_ sound1.count_m\[15\] _2381_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5884_ sound4.count_m\[2\] sound4.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__and2b_1
X_4904_ sound2.count\[15\] _1454_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7623_ _2099_ _2131_ vssd1 vssd1 vccd1 vccd1 _3695_ sky130_fd_sc_hd__and2_1
X_4835_ _1317_ _1382_ _1385_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4766_ _1314_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__or2_4
X_7554_ net628 _2843_ _2203_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__a21o_1
X_6505_ _1215_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7485_ _3634_ _3635_ vssd1 vssd1 vccd1 vccd1 _3636_ sky130_fd_sc_hd__nand2_1
X_4697_ _1263_ _1264_ _1256_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6436_ _0554_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6367_ _2783_ _2786_ _2795_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5318_ _1778_ _1824_ _1828_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__and3_1
X_8106_ clknet_leaf_95_hwclk sound2.osc.next_count\[7\] net68 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_6298_ _2695_ _2697_ _2694_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__a21oi_1
Xhold13 seq.encode.keys_sync\[10\] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _1761_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
Xhold35 _0158_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _0056_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 _0012_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dlygate4sd3_1
X_8037_ clknet_leaf_92_hwclk net620 net66 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold68 sound3.sdiv.Q\[12\] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 sound1.count_m\[1\] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 seq.encode.keys_edge_det\[7\] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4620_ _0677_ _0958_ _1077_ _0981_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4551_ sound1.count\[13\] _1120_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7270_ _3437_ _3444_ _3445_ _3440_ net230 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold505 _0245_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 sound4.sdiv.A\[19\] vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ net60 _1001_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__nor2_4
Xhold516 _0179_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 sound3.sdiv.Q\[3\] vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 sound3.sdiv.Q\[7\] vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ net621 _0573_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6152_ sound1.sdiv.Q\[0\] sound1.sdiv.Q\[1\] _0579_ _2434_ vssd1 vssd1 vccd1 vccd1
+ _2587_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _1176_ _1562_ _1572_ _0954_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__o221a_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ sound3.divisor_m\[2\] sound3.count_m\[1\] vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__or2b_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _1564_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__buf_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6985_ _3240_ vssd1 vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _2181_ _2370_ _2371_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_118_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5867_ _2302_ _2300_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__and2b_1
X_7606_ _3681_ _3682_ net871 _2184_ net529 vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5798_ _2238_ _2243_ _2244_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__a21o_1
X_4818_ sound2.count\[12\] _1360_ _1368_ sound2.count\[7\] vssd1 vssd1 vccd1 vccd1
+ _1369_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7537_ net132 _3654_ _3643_ net352 _3406_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__a221o_1
X_4749_ _1256_ _1302_ _1303_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7468_ sound3.sdiv.A\[23\] _3595_ vssd1 vssd1 vccd1 vccd1 _3621_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 beat_led[4] sky130_fd_sc_hd__buf_2
X_6419_ net929 _2832_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__nand2_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 note4[1] sky130_fd_sc_hd__clkbuf_4
X_7399_ sound3.divisor_m\[14\] _3552_ vssd1 vssd1 vccd1 vccd1 _3561_ sky130_fd_sc_hd__or2_1
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 note1[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6770_ _3112_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
X_3982_ _0554_ _0568_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ sound4.sdiv.Q\[12\] _2182_ _2185_ net149 _2191_ vssd1 vssd1 vccd1 vccd1 _0012_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5652_ _2089_ _2134_ _2087_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8371_ clknet_leaf_53_hwclk wave_comb.u1.next_dived net103 vssd1 vssd1 vccd1 vccd1
+ wave_comb.u1.dived sky130_fd_sc_hd__dfrtp_1
X_4603_ _0695_ net60 net59 vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__a21o_2
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5583_ _2063_ _2065_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__or2_1
X_7322_ sound3.divisor_m\[6\] _3483_ vssd1 vssd1 vccd1 vccd1 _3492_ sky130_fd_sc_hd__or2_1
X_4534_ _1073_ _1089_ _1104_ sound1.count\[0\] vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__a22o_1
Xhold302 _0013_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 sound1.sdiv.Q\[8\] vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 sound3.count\[0\] vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 sound1.count\[12\] vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold346 sound3.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7253_ _1608_ vssd1 vssd1 vccd1 vccd1 _3433_ sky130_fd_sc_hd__inv_2
Xhold368 sound1.count\[0\] vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _0940_ _0944_ _1004_ _0974_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__a211o_1
Xhold357 sound2.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6204_ _2631_ _2637_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__xnor2_1
X_7184_ net875 _2863_ vssd1 vssd1 vccd1 vccd1 _3393_ sky130_fd_sc_hd__and2_1
X_4396_ _0966_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__clkbuf_4
Xhold379 _0182_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__dlygate4sd3_1
X_6135_ _2275_ _2570_ sound3.sdiv.Q\[1\] _0577_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__a2bb2o_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ sound2.sdiv.Q\[0\] _0578_ _2499_ _2501_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__a31o_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5017_ _0542_ _1547_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6968_ _3224_ _3228_ _3235_ vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5919_ _2346_ sound4.count_m\[0\] _2347_ _2348_ _2354_ vssd1 vssd1 vccd1 vccd1 _2355_
+ sky130_fd_sc_hd__o2111a_1
X_6899_ _0578_ vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__buf_6
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold880 sound2.count\[3\] vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4250_ seq.clk_div.count\[10\] seq.clk_div.count\[11\] _0829_ vssd1 vssd1 vccd1 vccd1
+ _0835_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4181_ _0700_ net140 vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[0\] sky130_fd_sc_hd__nor2_1
X_7940_ clknet_leaf_18_hwclk _0103_ net84 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7871_ clknet_leaf_97_hwclk net106 net65 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6822_ net619 _2857_ _3125_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6753_ net728 _2895_ sound1.sdiv.next_dived _3101_ vssd1 vssd1 vccd1 vccd1 _0134_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _0446_ _0628_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3896_ _0565_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__inv_2
X_6684_ _3040_ _3041_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__nand2_1
X_5704_ net633 _2183_ sound4.sdiv.next_dived net634 vssd1 vssd1 vccd1 vccd1 _0003_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5635_ sound4.divisor_m\[1\] sound4.divisor_m\[0\] _2036_ vssd1 vssd1 vccd1 vccd1
+ _2118_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold110 sound4.sdiv.Q\[25\] vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dlygate4sd3_1
X_5566_ _2046_ _2048_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8354_ clknet_leaf_84_hwclk sound4.osc.next_count\[12\] net79 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[12\] sky130_fd_sc_hd__dfrtp_2
X_7305_ _3474_ _3476_ vssd1 vssd1 vccd1 vccd1 _3477_ sky130_fd_sc_hd__or2_1
Xhold132 sound3.count_m\[5\] vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _0075_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4517_ net60 _0939_ _1077_ _1081_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__o311a_1
X_8285_ clknet_leaf_60_hwclk _0385_ net95 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold143 _0384_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ sound4.count\[16\] _1988_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold176 sound3.sdiv.Q\[0\] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7236_ net744 _3422_ _3419_ vssd1 vssd1 vccd1 vccd1 _3423_ sky130_fd_sc_hd__mux2_1
Xhold165 sound3.count_m\[6\] vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 sound3.sdiv.Q\[10\] vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _0675_ _0945_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__nor2_4
Xhold187 sound1.sdiv.Q\[12\] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 sound4.count_m\[4\] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
X_4379_ _0949_ _0909_ _0940_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__nand3_4
X_7167_ sound2.sdiv.Q\[23\] _3167_ _3349_ net145 _3130_ vssd1 vssd1 vccd1 vccd1 _0263_
+ sky130_fd_sc_hd__a221o_1
X_6118_ _2547_ sound3.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__or2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ sound2.sdiv.A\[20\] net961 _3329_ vssd1 vssd1 vccd1 vccd1 _3352_ sky130_fd_sc_hd__o21ai_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ sound2.count_m\[3\] _2484_ sound2.divisor_m\[1\] _2480_ vssd1 vssd1 vccd1
+ vccd1 _2485_ sky130_fd_sc_hd__a22o_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5420_ _0997_ _1781_ _1926_ _1930_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5351_ _1139_ _1786_ _1790_ _1134_ _1834_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__o221a_1
X_4302_ _0871_ _0872_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__nand2_1
X_8070_ clknet_leaf_83_hwclk _0212_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5282_ _1771_ _1775_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__or2_1
X_4233_ net689 _0819_ _0813_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_92_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_7021_ sound2.divisor_m\[13\] _3274_ vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__or2_1
X_4164_ seq.player_2.state\[2\] seq.player_2.state\[3\] vssd1 vssd1 vccd1 vccd1 _0766_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4095_ net727 net807 _0713_ net537 vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a31o_1
X_7923_ clknet_leaf_19_hwclk net465 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7854_ clknet_leaf_98_hwclk seq.clk_div.next_count\[11\] net65 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[11\] sky130_fd_sc_hd__dfrtp_1
X_7785_ clknet_leaf_44_hwclk net113 net99 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_MODE
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_30_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6805_ _1470_ _2843_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__nor2_1
X_6736_ sound1.sdiv.A\[22\] sound1.sdiv.A\[21\] sound1.sdiv.A\[20\] sound1.sdiv.A\[19\]
+ _3055_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__o41a_1
XFILLER_0_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ sound2.count\[12\] sound2.count\[13\] _1527_ sound2.count\[14\] vssd1 vssd1
+ vccd1 vccd1 _1534_ sky130_fd_sc_hd__a31o_1
X_3948_ inputcont.INTERNAL_SYNCED_I\[4\] vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6667_ _2890_ _3025_ _3026_ _2894_ net317 vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__a32o_1
X_3879_ _0549_ _0534_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__nand2_4
XFILLER_0_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6598_ _2962_ _2963_ _0866_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__a21oi_1
X_5618_ sound4.divisor_m\[5\] _2100_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8337_ clknet_leaf_57_hwclk _0437_ net96 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5549_ sound4.divisor_m\[12\] _2031_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8268_ clknet_leaf_63_hwclk net330 net78 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_8199_ clknet_leaf_43_hwclk net285 net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_7219_ _1641_ vssd1 vssd1 vccd1 vccd1 _3412_ sky130_fd_sc_hd__inv_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout82 net2 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_6
Xfanout71 net72 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_8
XFILLER_0_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_6
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4920_ _0996_ _1025_ _1339_ _1393_ _0977_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__o32a_1
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4851_ _0869_ _1343_ _1345_ _1001_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3802_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1
+ vccd1 vccd1 _0481_ sky130_fd_sc_hd__nand2_2
X_7570_ net777 _1810_ _3419_ vssd1 vssd1 vccd1 vccd1 _3662_ sky130_fd_sc_hd__mux2_1
X_4782_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__buf_4
X_6521_ _2893_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6452_ net384 _2836_ _2851_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5403_ _1222_ _1913_ sound4.count\[17\] vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6383_ net671 _2806_ _2808_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8122_ clknet_leaf_60_hwclk _0243_ net94 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5334_ _0686_ _1784_ _1781_ _1146_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__o22ai_1
X_8053_ clknet_leaf_81_hwclk _0195_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_5265_ _1765_ _1775_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__or2_1
X_5196_ sound3.count\[0\] sound3.count\[1\] sound3.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1725_ sky130_fd_sc_hd__a21o_1
X_4216_ _0804_ _0805_ _0808_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__and4_1
X_7004_ _3265_ _3267_ vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4147_ net824 seq.player_3.state\[2\] net890 _0754_ _0700_ vssd1 vssd1 vccd1 vccd1
+ _0755_ sky130_fd_sc_hd__a311o_1
X_4078_ net1 net19 vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__and2b_1
X_7906_ clknet_leaf_0_hwclk _0069_ net65 vssd1 vssd1 vccd1 vccd1 seq.beat\[3\] sky130_fd_sc_hd__dfrtp_4
X_7837_ clknet_leaf_52_hwclk _0060_ net101 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7768_ clknet_leaf_47_hwclk pm.next_count\[7\] net102 vssd1 vssd1 vccd1 vccd1 pm.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6719_ _3072_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__inv_2
X_7699_ _3747_ vssd1 vssd1 vccd1 vccd1 _3748_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold709 sound2.count\[6\] vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5050_ _0993_ _1012_ _1578_ _1580_ _0948_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__o32a_1
X_4001_ net569 _0652_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5952_ _2382_ _2384_ _2386_ _2387_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4903_ _0683_ _1316_ _1451_ _1453_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5883_ _2318_ sound4.divisor_m\[6\] sound4.divisor_m\[5\] _2312_ vssd1 vssd1 vccd1
+ vccd1 _2319_ sky130_fd_sc_hd__a22o_1
X_7622_ _3681_ _3693_ _3694_ _2184_ net383 vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__a32o_1
X_4834_ _1151_ _1323_ _1339_ _1095_ _1384_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4765_ _1314_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nor2_2
X_7553_ net506 _3403_ _2202_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6504_ _2883_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7484_ sound3.sdiv.A\[25\] _3595_ vssd1 vssd1 vccd1 vccd1 _3635_ sky130_fd_sc_hd__or2_1
X_4696_ sound1.count\[0\] net913 sound1.count\[2\] net944 vssd1 vssd1 vccd1 vccd1
+ _1264_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ net224 _2836_ _2842_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6366_ _2779_ _2782_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5317_ _1154_ _1784_ _1826_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__o211a_1
X_8105_ clknet_leaf_95_hwclk sound2.osc.next_count\[6\] net68 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[6\] sky130_fd_sc_hd__dfrtp_1
Xhold14 inputcont.INTERNAL_MODE vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dlygate4sd3_1
X_6297_ _2726_ _2727_ vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__nand2_1
X_8036_ clknet_leaf_93_hwclk _0178_ net66 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_5248_ _1721_ _1759_ _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__and3_1
Xhold47 sound1.sdiv.Q\[26\] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 seq.clk_div.count\[0\] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 rate_clk.count\[4\] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold69 _0352_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _0680_ _0959_ _1574_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__or3_1
Xhold58 seq.player_6.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4550_ sound1.count\[13\] _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold517 wave_comb.u1.Q\[4\] vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 sound4.sdiv.Q\[4\] vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__dlygate4sd3_1
X_4481_ _0944_ _0969_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold539 sound3.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ net679 _2653_ _0645_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__mux2_1
Xhold528 sound4.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6151_ sound1.sdiv.Q\[3\] _0579_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _0996_ _1550_ _1630_ _1632_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ sound3.count_m\[1\] sound3.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__or2b_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _1547_ _1563_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__or2_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6984_ _3248_ _3249_ vssd1 vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__nand2_1
X_5935_ sound4.sdiv.Q\[1\] _0576_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__nand2_1
X_5866_ _2300_ _2302_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7605_ sound4.divisor_m\[0\] net870 vssd1 vssd1 vccd1 vccd1 _3683_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4817_ _1362_ _1364_ _1367_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__and3_2
XFILLER_0_118_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5797_ _2238_ _2243_ _2244_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7536_ sound3.sdiv.Q\[25\] _3654_ _3643_ net157 _3405_ vssd1 vssd1 vccd1 vccd1 _0364_
+ sky130_fd_sc_hd__a221o_1
X_4748_ sound1.count\[16\] _1299_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__or2_1
X_7467_ net425 _3463_ sound3.sdiv.next_dived _3620_ vssd1 vssd1 vccd1 vccd1 _0329_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4679_ sound1.count\[4\] _1145_ _1249_ sound1.count\[12\] vssd1 vssd1 vccd1 vccd1
+ _1250_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6418_ seq.beat\[2\] _2832_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__or2_1
X_7398_ sound3.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _3560_ sky130_fd_sc_hd__inv_2
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 note1[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 note4[2] sky130_fd_sc_hd__clkbuf_4
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 beat_led[5] sky130_fd_sc_hd__clkbuf_4
X_6349_ _2772_ _2778_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8019_ clknet_leaf_17_hwclk _0161_ net83 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ net33 _0643_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__nor2_2
X_5720_ sound4.count\[4\] _2186_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _2093_ _2132_ _2133_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__a21boi_1
X_4602_ _1009_ _1051_ _1106_ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or4_1
X_8370_ clknet_leaf_72_hwclk rate_clk.next_count\[7\] net82 vssd1 vssd1 vccd1 vccd1
+ rate_clk.count\[7\] sky130_fd_sc_hd__dfrtp_4
X_5582_ sound4.divisor_m\[12\] _2064_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__xor2_1
XFILLER_0_130_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7321_ sound3.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 _3491_ sky130_fd_sc_hd__inv_2
X_4533_ _1094_ _1099_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__and3_2
Xhold325 sound1.sdiv.A\[18\] vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__dlygate4sd3_1
X_7252_ _3432_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
Xhold314 sound1.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 sound1.count_m\[15\] vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6203_ _2292_ _2634_ _2635_ _2636_ _2279_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__o32a_1
Xhold347 sound1.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _0150_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 sound4.sdiv.Q\[9\] vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold369 seq.encode.keys_edge_det\[10\] vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__dlygate4sd3_1
X_4464_ _0952_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__nor2_2
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7183_ net236 _3132_ _3392_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4395_ _0918_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6134_ _2516_ _2556_ _2569_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__o21a_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _2500_ sound2.sdiv.next_start vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__nor2_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _0546_ _1546_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _3233_ _3234_ vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5918_ _2350_ _2353_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6898_ sound2.divisor_m\[0\] sound2.sdiv.Q\[27\] _3171_ vssd1 vssd1 vccd1 vccd1 _3173_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _2181_ _2284_ _2285_ _2286_ _0645_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7519_ net416 _3654_ _3643_ net642 _3387_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold881 sound1.count\[7\] vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold870 _2832_ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4180_ _0774_ _0773_ net830 _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_1.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_7870_ clknet_leaf_8_hwclk net466 net70 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_6821_ sound2.count\[10\] _2855_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6752_ _3098_ _3100_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ _0626_ _0627_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3895_ sound1.sdiv.C\[4\] sound1.sdiv.C\[3\] sound1.sdiv.C\[2\] _0564_ net878 vssd1
+ vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__a311oi_4
X_6683_ sound1.sdiv.A\[16\] _3039_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__or2_1
X_5703_ sound4.sdiv.Q\[2\] _2183_ sound4.sdiv.next_dived net524 vssd1 vssd1 vccd1
+ vccd1 _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5634_ sound4.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8353_ clknet_leaf_85_hwclk sound4.osc.next_count\[11\] net79 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[11\] sky130_fd_sc_hd__dfrtp_2
X_7304_ sound3.divisor_m\[5\] _3475_ vssd1 vssd1 vccd1 vccd1 _3476_ sky130_fd_sc_hd__xnor2_1
Xhold100 sound3.sdiv.Q\[11\] vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5565_ sound4.divisor_m\[17\] _2047_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold122 sound3.count_m\[4\] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _0273_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 sound3.sdiv.Q\[13\] vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 sound1.sdiv.Q\[25\] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4516_ _1082_ _1084_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__and3_1
X_8284_ clknet_leaf_63_hwclk net247 net81 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_5496_ _1991_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
Xhold177 _0340_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
X_7235_ _1714_ vssd1 vssd1 vccd1 vccd1 _3422_ sky130_fd_sc_hd__inv_2
Xhold166 _0274_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _0350_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4447_ _0674_ _0964_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__nor2_4
Xhold199 _0371_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
X_7166_ net145 _3167_ _3349_ net370 _3129_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__a221o_1
Xhold188 sound2.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
X_6117_ _2509_ sound3.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__or2_1
X_4378_ _0926_ _0936_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__nor2_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ sound2.sdiv.A\[20\] _3329_ _3343_ vssd1 vssd1 vccd1 vccd1 _3351_ sky130_fd_sc_hd__o21bai_1
X_6048_ sound2.divisor_m\[4\] vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__inv_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7999_ clknet_leaf_40_hwclk _0141_ net98 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5350_ _1804_ _1822_ _1852_ _1860_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4301_ seq.player_1.state\[0\] seq.player_1.state\[1\] seq.player_1.state\[2\] seq.player_1.state\[3\]
+ _0698_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__o41a_1
X_5281_ _1791_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__buf_4
X_4232_ net689 _0819_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__and2_1
X_7020_ sound2.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4163_ seq.player_2.state\[2\] net458 _0764_ _0765_ _0700_ vssd1 vssd1 vccd1 vccd1
+ seq.player_2.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_4094_ net860 _0716_ _0718_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_8.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
X_7922_ clknet_leaf_17_hwclk net408 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7853_ clknet_leaf_98_hwclk seq.clk_div.next_count\[10\] net65 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[10\] sky130_fd_sc_hd__dfrtp_2
X_7784_ clknet_leaf_74_hwclk net116 net76 vssd1 vssd1 vccd1 vccd1 inputcont.u2.next_in
+ sky130_fd_sc_hd__dfrtp_1
X_4996_ sound2.count\[13\] sound2.count\[14\] _1530_ vssd1 vssd1 vccd1 vccd1 _1533_
+ sky130_fd_sc_hd__and3_1
X_6804_ net186 _2857_ _3116_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__a21o_1
X_6735_ _3069_ _3073_ _3078_ _3081_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__nor4b_1
X_3947_ inputcont.INTERNAL_SYNCED_I\[10\] _0610_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6666_ _3014_ _3018_ _3024_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3878_ _0545_ _0547_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__and3_2
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6597_ _2962_ _2963_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__or2_1
X_5617_ sound4.divisor_m\[4\] _2026_ _2036_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8336_ clknet_leaf_57_hwclk _0436_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5548_ sound4.divisor_m\[11\] sound4.divisor_m\[10\] _2030_ vssd1 vssd1 vccd1 vccd1
+ _2031_ sky130_fd_sc_hd__or3_1
X_8267_ clknet_leaf_67_hwclk net420 net95 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7218_ _3411_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__clkbuf_1
X_5479_ _1977_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__inv_2
X_8198_ clknet_leaf_28_hwclk _0319_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_7149_ sound2.sdiv.Q\[5\] _3168_ _3164_ net608 vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__a22o_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout83 net86 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_8
XFILLER_0_76_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout72 net2 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_4
XFILLER_0_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout94 net103 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_8
XFILLER_0_37_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4850_ _0978_ _0944_ _1333_ _1347_ _0997_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__o32a_1
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3801_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[2\]
+ inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__o31ai_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6520_ _2890_ _2891_ _2892_ _2894_ net499 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4781_ _1319_ _1331_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6451_ sound1.count\[13\] _2201_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6382_ _2807_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__clkbuf_4
X_5402_ _1772_ _1773_ _1777_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__and3_1
X_8121_ clknet_leaf_60_hwclk _0242_ net94 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5333_ _1011_ _1015_ _1842_ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8052_ clknet_leaf_81_hwclk _0194_ net74 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_5264_ _1766_ _1774_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__or2_1
X_5195_ _1724_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4215_ _0806_ seq.clk_div.count\[9\] seq.tempo_select.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0809_ sky130_fd_sc_hd__a21o_1
X_7003_ sound2.divisor_m\[12\] _3266_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__xnor2_1
X_4146_ seq.player_3.state\[0\] _0753_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__and2_1
X_4077_ _0708_ vssd1 vssd1 vccd1 vccd1 seq_play_on sky130_fd_sc_hd__clkbuf_1
X_7905_ clknet_leaf_0_hwclk _0068_ net65 vssd1 vssd1 vccd1 vccd1 seq.beat\[2\] sky130_fd_sc_hd__dfrtp_4
X_7836_ clknet_leaf_52_hwclk _0059_ net101 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7767_ clknet_leaf_47_hwclk pm.next_count\[6\] net102 vssd1 vssd1 vccd1 vccd1 pm.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4979_ net815 _1520_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6718_ sound1.sdiv.A\[20\] _3055_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__xor2_1
X_7698_ sound4.sdiv.C\[2\] sound4.sdiv.C\[1\] sound4.sdiv.C\[0\] vssd1 vssd1 vccd1
+ vccd1 _3747_ sky130_fd_sc_hd__and3_1
X_6649_ sound1.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8319_ clknet_leaf_71_hwclk _0419_ net82 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_91_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4000_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_44_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _2385_ sound1.divisor_m\[12\] sound1.count_m\[10\] _2378_ vssd1 vssd1 vccd1
+ vccd1 _2387_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4902_ _0688_ _1334_ _1452_ _1317_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_59_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ sound4.count_m\[5\] vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7621_ _2129_ _3692_ vssd1 vssd1 vccd1 vccd1 _3694_ sky130_fd_sc_hd__or2b_1
X_4833_ _1134_ _1343_ _1333_ _1146_ _1383_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4764_ _0698_ _0504_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__or2_2
X_7552_ net219 _3403_ _2200_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__a21o_1
X_7483_ net952 _3595_ vssd1 vssd1 vccd1 vccd1 _3634_ sky130_fd_sc_hd__nand2_1
X_6503_ net732 _2882_ _2864_ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6434_ net863 _2201_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__and2_1
X_4695_ sound1.count\[0\] sound1.count\[1\] sound1.count\[2\] sound1.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ _2762_ _2791_ _2792_ _2793_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__o22a_1
X_6296_ _2725_ _2717_ _2721_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__or3_1
X_5316_ _1166_ _1800_ _1796_ _0677_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8104_ clknet_leaf_89_hwclk sound2.osc.next_count\[5\] net68 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_5247_ net981 _1756_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__nand2_1
X_8035_ clknet_leaf_93_hwclk _0177_ net66 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold37 sound3.sdiv.Q\[9\] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 inputcont.u1.ff_intermediate\[11\] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _2003_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 _0168_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _1158_ _1578_ _1550_ _1004_ _1708_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__o221a_1
Xhold59 sound2.count_m\[18\] vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4129_ net753 _0740_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7819_ clknet_leaf_2_hwclk net481 net70 vssd1 vssd1 vccd1 vccd1 seq.player_4.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold518 _0050_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__dlygate4sd3_1
X_4480_ sound1.count\[2\] _1032_ _1050_ sound1.count\[11\] vssd1 vssd1 vccd1 vccd1
+ _1051_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold507 seq.player_6.state\[2\] vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold529 sound4.sdiv.Q\[3\] vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6150_ _2289_ _2583_ _2584_ _2290_ sound4.sdiv.Q\[3\] vssd1 vssd1 vccd1 vccd1 _2585_
+ sky130_fd_sc_hd__a32o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _1129_ _1580_ _1570_ _1182_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__o221a_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ sound3.count_m\[0\] vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__inv_2
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _0698_ _0540_ _1557_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__o21ai_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6983_ _3244_ _3247_ vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__nand2_1
X_5934_ _2314_ _2321_ _2356_ _2369_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5865_ _2275_ _2292_ _2301_ sound3.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_118_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7604_ sound4.divisor_m\[0\] net870 vssd1 vssd1 vccd1 vccd1 _3682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4816_ _1085_ _1322_ _1339_ _1078_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5796_ wave_comb.u1.A\[6\] _2224_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7535_ net157 _3654_ _3643_ net274 _3404_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4747_ net983 _1299_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7466_ _3618_ _3619_ vssd1 vssd1 vccd1 vccd1 _3620_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4678_ _1239_ _1241_ _1244_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__and4_2
X_7397_ _3437_ _3558_ _3559_ _3440_ net284 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6417_ _2831_ net974 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6348_ sound4.sdiv.Q\[8\] _2290_ _2369_ _2773_ _2777_ vssd1 vssd1 vccd1 vccd1 _2778_
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 note4[3] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 beat_led[6] sky130_fd_sc_hd__clkbuf_4
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 note2[0] sky130_fd_sc_hd__clkbuf_4
X_6279_ _2708_ _2710_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__xnor2_1
X_8018_ clknet_leaf_17_hwclk net377 net84 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _0630_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ net949 _2092_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ _1121_ _1122_ _1145_ sound1.count\[4\] _1171_ vssd1 vssd1 vccd1 vccd1 _1172_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _2036_ _2031_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__nand2_1
X_7320_ _3437_ _3489_ _3490_ _3440_ net309 vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a32o_1
X_4532_ _0981_ _1041_ _1101_ _0990_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__o221a_1
XFILLER_0_41_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold326 _0126_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__dlygate4sd3_1
X_7251_ net854 _3431_ _3419_ vssd1 vssd1 vccd1 vccd1 _3432_ sky130_fd_sc_hd__mux2_1
Xhold304 _0085_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 sound4.count_m\[0\] vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ _0685_ _0677_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__nor2_2
XFILLER_0_111_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold337 sound1.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ sound3.sdiv.Q\[4\] _0577_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__nand2_1
Xhold359 _0010_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 inputcont.INTERNAL_SYNCED_I\[5\] vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__dlygate4sd3_1
X_7182_ sound3.count\[5\] _2863_ vssd1 vssd1 vccd1 vccd1 _3392_ sky130_fd_sc_hd__and2_1
X_4394_ _0909_ _0955_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__nand2_1
X_6133_ _2544_ _2568_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__nor2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ net880 vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__inv_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _0699_ net45 vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__and2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _3229_ _3232_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__nand2_1
X_5917_ _2346_ sound4.count_m\[0\] _2351_ _2352_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6897_ _3165_ _3171_ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5848_ net29 net30 vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5779_ _2225_ _2222_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7518_ _0577_ vssd1 vssd1 vccd1 vccd1 _3654_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7449_ _3599_ _3602_ _3605_ vssd1 vssd1 vccd1 vccd1 _3606_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold871 sound3.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 wave_comb.u1.A\[4\] vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold860 sound2.sdiv.A\[21\] vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6820_ net492 _2857_ _3124_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__a21o_1
X_6751_ _3089_ _3092_ _3099_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3963_ _0456_ _0625_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__nand2_1
X_6682_ sound1.sdiv.A\[16\] _3039_ vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__nand2_1
X_3894_ sound1.sdiv.start vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__inv_2
X_5702_ sound4.sdiv.Q\[1\] _2183_ sound4.sdiv.next_dived net262 vssd1 vssd1 vccd1
+ vccd1 _0001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5633_ _2114_ _2115_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5564_ _2036_ _2034_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8352_ clknet_leaf_85_hwclk sound4.osc.next_count\[10\] net77 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7303_ sound3.divisor_m\[4\] _3465_ _3448_ vssd1 vssd1 vccd1 vccd1 _3475_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4515_ _0952_ _1000_ _1003_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 sound2.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold123 sound3.count_m\[2\] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _0167_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlygate4sd3_1
X_8283_ clknet_leaf_63_hwclk net443 net78 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_5495_ _1779_ _1936_ _1989_ _1990_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__and4_1
Xhold134 sound2.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7234_ _2843_ _1706_ _3421_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__o21ai_1
X_4446_ _0683_ _0947_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__nor2_2
Xhold156 sound4.count_m\[3\] vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 sound2.sdiv.Q\[25\] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 sound4.count_m\[12\] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold178 sound4.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ _0944_ _0947_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__or2_4
X_7165_ sound2.sdiv.Q\[21\] _3167_ _3349_ net147 _3128_ vssd1 vssd1 vccd1 vccd1 _0261_
+ sky130_fd_sc_hd__a221o_1
Xhold189 _0208_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
X_6116_ _2545_ sound3.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ net979 _3329_ vssd1 vssd1 vccd1 vccd1 _3350_ sky130_fd_sc_hd__xnor2_1
X_6047_ sound2.divisor_m\[1\] _2480_ _2481_ _2482_ vssd1 vssd1 vccd1 vccd1 _2483_
+ sky130_fd_sc_hd__o211ai_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ clknet_leaf_58_hwclk sound2.sdiv.next_dived net95 vssd1 vssd1 vccd1 vccd1
+ sound2.sdiv.dived sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6949_ _3206_ _3209_ _3217_ vssd1 vssd1 vccd1 vccd1 _3219_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold690 sound4.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4300_ _0702_ seq.encode.play _0870_ inputcont.INTERNAL_SYNCED_I\[0\] vssd1 vssd1
+ vccd1 vccd1 _0871_ sky130_fd_sc_hd__a31o_2
X_5280_ _1767_ _1773_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__or2_1
X_4231_ _0821_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4162_ net882 _0762_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__nor2_1
X_4093_ _0698_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__buf_6
X_7921_ clknet_leaf_18_hwclk net332 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7852_ clknet_leaf_98_hwclk seq.clk_div.next_count\[9\] net65 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[9\] sky130_fd_sc_hd__dfrtp_1
X_7783_ clknet_leaf_44_hwclk net118 net99 vssd1 vssd1 vccd1 vccd1 inputcont.u3.next_in
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4995_ net446 _1530_ _1532_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[13\] sky130_fd_sc_hd__a21oi_1
X_6803_ net925 _2855_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__and2_1
X_6734_ sound1.sdiv.A\[23\] _3055_ vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3946_ _0608_ _0609_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_0__f_hwclk clknet_0_hwclk vssd1 vssd1 vccd1 vccd1 clknet_3_0__leaf_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6665_ _3014_ _3018_ _3024_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3877_ _0518_ _0527_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6596_ _2946_ _2953_ _2951_ vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__o21a_1
X_5616_ _2097_ _2098_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8335_ clknet_leaf_57_hwclk _0435_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5547_ sound4.divisor_m\[9\] _2029_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__or2_1
X_8266_ clknet_leaf_40_hwclk net133 net100 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5478_ sound4.count\[12\] _1973_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__and2_1
X_7217_ net734 _3410_ _3142_ vssd1 vssd1 vccd1 vccd1 _3411_ sky130_fd_sc_hd__mux2_1
X_4429_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__buf_4
X_8197_ clknet_leaf_28_hwclk _0318_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7148_ sound2.sdiv.Q\[4\] _3168_ _3164_ net571 vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__a22o_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7079_ sound2.sdiv.A\[19\] _3329_ vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout73 net75 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_8
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout84 net86 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_6
Xfanout95 net97 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_6
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _0443_ _0463_ inputcont.INTERNAL_SYNCED_I\[6\] vssd1 vssd1 vccd1 vccd1 _0479_
+ sky130_fd_sc_hd__o21ai_4
X_4780_ _1315_ _1330_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6450_ net389 _2836_ _2850_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6381_ wave_comb.u1.dived _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5401_ sound4.count\[7\] _1897_ _1903_ sound4.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1912_ sky130_fd_sc_hd__a2bb2o_1
X_8120_ clknet_leaf_60_hwclk _0241_ net94 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5332_ _1200_ _1792_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8051_ clknet_leaf_81_hwclk _0193_ net74 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5263_ _0698_ _0673_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__nor2_1
X_5194_ _1721_ _1722_ _1723_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__and3_1
X_4214_ seq.tempo_select.state\[1\] _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__nand2_1
X_7002_ sound2.divisor_m\[11\] _3256_ _3177_ vssd1 vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__o21a_1
X_4145_ net915 inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4076_ net1 net18 vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__and2b_1
X_7904_ clknet_leaf_96_hwclk _0067_ net65 vssd1 vssd1 vccd1 vccd1 seq.beat\[1\] sky130_fd_sc_hd__dfrtp_4
X_7835_ clknet_leaf_52_hwclk _0058_ net101 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7766_ clknet_leaf_48_hwclk net510 net102 vssd1 vssd1 vccd1 vccd1 pm.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ net934 _1521_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[7\] sky130_fd_sc_hd__nor2_1
X_6717_ net616 _2895_ _3069_ _3071_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7697_ net562 sound4.sdiv.C\[0\] net586 vssd1 vssd1 vccd1 vccd1 _3746_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3929_ _0593_ net55 _0590_ _0521_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__o31a_1
X_6648_ _2890_ _3008_ _3009_ _2894_ net316 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6579_ sound1.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__inv_2
X_8318_ clknet_leaf_70_hwclk _0418_ net82 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_8249_ clknet_leaf_37_hwclk net142 net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5950_ _2383_ sound1.count_m\[12\] _2385_ sound1.divisor_m\[12\] vssd1 vssd1 vccd1
+ vccd1 _2386_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4901_ _1138_ _1324_ _1315_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__or3b_1
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7620_ _3692_ _2129_ vssd1 vssd1 vccd1 vccd1 _3693_ sky130_fd_sc_hd__or2b_1
X_5881_ _2315_ sound4.divisor_m\[8\] _2316_ sound4.divisor_m\[7\] vssd1 vssd1 vccd1
+ vccd1 _2317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4832_ _1012_ _1338_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__or2_1
X_4763_ _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__or2_2
X_7551_ net249 _3403_ _2199_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__a21o_1
X_7482_ net511 _3463_ sound3.sdiv.next_dived _3633_ vssd1 vssd1 vccd1 vccd1 _0331_
+ sky130_fd_sc_hd__a22o_1
X_6502_ _1235_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4694_ _1262_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6433_ net297 _2836_ _2841_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6364_ _2772_ _2778_ vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__nor2_1
X_6295_ _2717_ _2721_ _2725_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__o21ai_1
X_5315_ _0685_ _1769_ _1794_ _1077_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__o221a_1
X_8103_ clknet_leaf_95_hwclk sound2.osc.next_count\[4\] net68 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[4\] sky130_fd_sc_hd__dfrtp_2
X_5246_ sound3.count\[18\] _1756_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8034_ clknet_leaf_81_hwclk net234 net73 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold38 _0349_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 inputcont.u1.ff_intermediate\[4\] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 rate_clk.next_count\[5\] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 sound1.sdiv.Q\[15\] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _1014_ _1567_ _1570_ _1083_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__o22a_1
X_4128_ seq.player_5.state\[2\] net877 vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__nand2_1
X_4059_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7818_ clknet_leaf_1_hwclk net638 net70 vssd1 vssd1 vccd1 vccd1 seq.player_4.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7749_ clknet_leaf_54_hwclk _0034_ net101 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold508 seq.player_6.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold519 net838 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_2
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6080_ _2510_ _2512_ _2515_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__nand3b_1
X_5100_ _1026_ _1567_ _1574_ _1175_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__o22a_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__buf_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6982_ _3244_ _3247_ vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5933_ sound4.count_m\[17\] _2349_ sound4.count_m\[18\] _2368_ vssd1 vssd1 vccd1
+ vccd1 _2369_ sky130_fd_sc_hd__a211o_1
X_5864_ sound3.sdiv.next_start _2279_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__nor2_2
XFILLER_0_118_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7603_ _1764_ vssd1 vssd1 vccd1 vccd1 _3681_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4815_ _1083_ _1321_ _1341_ _1079_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__o221a_1
X_5795_ wave_comb.u1.next_dived _2242_ _2243_ _0573_ net514 vssd1 vssd1 vccd1 vccd1
+ _0034_ sky130_fd_sc_hd__a32o_1
X_7534_ sound3.sdiv.Q\[23\] _3654_ _3643_ net124 _3402_ vssd1 vssd1 vccd1 vccd1 _0362_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4746_ _1301_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
X_7465_ sound3.sdiv.A\[21\] _3595_ _3616_ vssd1 vssd1 vccd1 vccd1 _3619_ sky130_fd_sc_hd__a21oi_1
X_4677_ _0992_ _1245_ _1246_ _1247_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7396_ _3546_ _3549_ _3557_ vssd1 vssd1 vccd1 vccd1 _3559_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6416_ net973 seq.beat\[0\] _2830_ vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__and3_1
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 beat_led[7] sky130_fd_sc_hd__clkbuf_4
X_6347_ _2292_ _2776_ vssd1 vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__nor2_1
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 note2[1] sky130_fd_sc_hd__clkbuf_4
X_6278_ _2672_ _2675_ _2709_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_90_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5229_ net681 _1744_ _1721_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__o21ai_1
X_8017_ clknet_leaf_17_hwclk net372 net84 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600_ sound1.count\[10\] _1157_ _1170_ sound1.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _1171_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5580_ sound4.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__inv_2
X_4531_ _0977_ _0950_ _0996_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7250_ _1615_ vssd1 vssd1 vccd1 vccd1 _3431_ sky130_fd_sc_hd__inv_2
Xhold316 _0367_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__dlygate4sd3_1
X_4462_ _0679_ _0971_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__or2_2
XFILLER_0_4_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold305 sound4.count\[7\] vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ sound3.sdiv.Q\[3\] _0577_ _2633_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__a21oi_1
Xhold327 sound1.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 sound4.count_m\[16\] vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold349 sound2.sdiv.Q\[23\] vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7181_ net226 _3132_ _3391_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__a21o_1
X_4393_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__buf_8
X_6132_ _2552_ _2567_ _2546_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__a21oi_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _2459_ _2469_ _2487_ _2498_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__a31o_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _1545_ vssd1 vssd1 vccd1 vccd1 sound3.sdiv.next_dived sky130_fd_sc_hd__buf_4
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _3229_ _3232_ vssd1 vssd1 vccd1 vccd1 _3233_ sky130_fd_sc_hd__or2_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5916_ sound4.divisor_m\[2\] sound4.count_m\[1\] vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6896_ sound2.sdiv.A\[0\] _3170_ vssd1 vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5847_ _2181_ _2284_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5778_ _2227_ _2228_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7517_ net642 _3440_ _3437_ net649 vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__a22o_1
X_4729_ _1287_ _1288_ _1256_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7448_ sound3.sdiv.A\[18\] _3595_ _3600_ _3603_ _3604_ vssd1 vssd1 vccd1 vccd1 _3605_
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7379_ sound3.divisor_m\[12\] sound3.divisor_m\[11\] _3526_ vssd1 vssd1 vccd1 vccd1
+ _3543_ sky130_fd_sc_hd__or3_1
Xhold872 sound3.sdiv.A\[24\] vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold850 wave_comb.u1.A\[4\] vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 sound2.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold883 sound1.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6750_ sound1.sdiv.A\[24\] sound1.sdiv.A\[23\] _3055_ vssd1 vssd1 vccd1 vccd1 _3099_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3962_ _0456_ _0625_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__or2_1
X_5701_ _2182_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__clkbuf_8
X_3893_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__inv_2
X_6681_ _3038_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5632_ _2111_ _2113_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5563_ sound4.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8351_ clknet_leaf_86_hwclk sound4.osc.next_count\[9\] net77 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7302_ sound3.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 _3474_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4514_ _0959_ _0952_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold102 sound3.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 net820 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_2
X_5494_ sound4.count\[15\] _1984_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__or2_1
Xhold124 sound2.count_m\[0\] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 sound4.sdiv.Q\[15\] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__dlygate4sd3_1
X_8282_ clknet_leaf_64_hwclk net629 net80 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7233_ net641 _2843_ vssd1 vssd1 vccd1 vccd1 _3421_ sky130_fd_sc_hd__nand2_1
X_4445_ _1015_ _0869_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__nand2_2
Xhold157 _0370_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 sound4.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _0379_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold179 _0430_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
X_4376_ _0675_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nor2_4
X_7164_ net147 _3167_ _3349_ net166 _3127_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6115_ sound3.divisor_m\[1\] vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _1311_ vssd1 vssd1 vccd1 vccd1 _3349_ sky130_fd_sc_hd__buf_6
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ sound2.divisor_m\[2\] sound2.count_m\[1\] vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__or2b_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ clknet_leaf_5_hwclk sound1.osc.next_count\[18\] net72 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6948_ _3206_ _3209_ _3217_ vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__nand3_1
XFILLER_0_107_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6879_ _3159_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold680 sound2.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold691 sound1.divisor_m\[5\] vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _0819_ _0820_ _0813_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__and3b_1
X_4161_ seq.player_2.state\[0\] seq.player_2.state\[1\] _0761_ vssd1 vssd1 vccd1 vccd1
+ _0764_ sky130_fd_sc_hd__and3_1
X_4092_ net731 _0715_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__xor2_1
X_7920_ clknet_leaf_18_hwclk net385 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_7851_ clknet_leaf_98_hwclk seq.clk_div.next_count\[8\] net65 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[8\] sky130_fd_sc_hd__dfrtp_2
X_6802_ net228 _2857_ _3115_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__a21o_1
X_7782_ clknet_leaf_55_hwclk net128 net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_4994_ net446 _1530_ _1504_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__o21ai_1
X_6733_ sound1.sdiv.A\[23\] _3055_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3945_ inputcont.INTERNAL_SYNCED_I\[6\] inputcont.INTERNAL_SYNCED_I\[8\] vssd1 vssd1
+ vccd1 vccd1 _0609_ sky130_fd_sc_hd__nor2_1
X_6664_ _3022_ _3023_ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__nand2_1
X_5615_ sound4.sdiv.A\[5\] _2096_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__or2_1
X_3876_ _0520_ _0541_ net55 vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6595_ _2960_ _2961_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8334_ clknet_leaf_57_hwclk net587 net96 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5546_ sound4.divisor_m\[8\] sound4.divisor_m\[7\] _2028_ vssd1 vssd1 vccd1 vccd1
+ _2029_ sky130_fd_sc_hd__or3_1
X_8265_ clknet_leaf_38_hwclk net353 net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5477_ _1976_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7216_ _1655_ vssd1 vssd1 vccd1 vccd1 _3410_ sky130_fd_sc_hd__inv_2
X_4428_ _0940_ _0974_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8196_ clknet_leaf_27_hwclk _0317_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_7147_ net571 _3168_ sound2.sdiv.next_dived net598 vssd1 vssd1 vccd1 vccd1 _0243_
+ sky130_fd_sc_hd__a22o_1
X_4359_ _0928_ _0929_ _0892_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__o21a_1
X_7078_ net595 _3168_ sound2.sdiv.next_dived _3334_ vssd1 vssd1 vccd1 vccd1 _0226_
+ sky130_fd_sc_hd__a22o_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _2463_ sound2.divisor_m\[6\] sound2.divisor_m\[5\] _2464_ vssd1 vssd1 vccd1
+ vccd1 _2465_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout74 net75 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_8
Xfanout85 net86 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_4
Xfanout96 net97 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_4
XFILLER_0_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6380_ _2280_ _2274_ _2805_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__mux2_1
X_5400_ sound4.count\[15\] _1891_ _1897_ sound4.count\[7\] _1910_ vssd1 vssd1 vccd1
+ vccd1 _1911_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5331_ _1771_ _1775_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__nor2_1
X_8050_ clknet_leaf_89_hwclk _0192_ net68 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_7001_ sound2.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _3265_ sky130_fd_sc_hd__inv_2
X_5262_ _0698_ _0587_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__or2_4
X_5193_ net428 sound3.count\[1\] vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__nand2_1
X_4213_ seq.tempo_select.state\[0\] _0802_ seq.clk_div.count\[9\] _0806_ vssd1 vssd1
+ vccd1 vccd1 _0807_ sky130_fd_sc_hd__a211o_1
X_4144_ _0750_ _0749_ _0752_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_4.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_4075_ _0706_ _0707_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__nor2_1
X_7903_ clknet_leaf_96_hwclk _0066_ net64 vssd1 vssd1 vccd1 vccd1 seq.beat\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7834_ clknet_leaf_51_hwclk _0057_ net102 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7765_ clknet_leaf_50_hwclk pm.next_count\[4\] net102 vssd1 vssd1 vccd1 vccd1 pm.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6716_ _0866_ _3070_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ net693 _1518_ _1504_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7696_ _3681_ _3744_ _3745_ _2184_ net562 vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3928_ _0545_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__inv_2
X_6647_ _2996_ _3000_ _3007_ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3859_ _0520_ _0524_ _0528_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__a211o_1
X_6578_ _2942_ _2943_ _2940_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__o21a_1
X_5529_ _2012_ pm.current_waveform\[3\] vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8317_ clknet_leaf_71_hwclk _0417_ net82 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_8248_ clknet_leaf_41_hwclk _0348_ net98 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_8179_ clknet_leaf_29_hwclk _0300_ net91 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5880_ sound4.count_m\[6\] vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__inv_2
X_4900_ net59 _1449_ _1450_ _0944_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__a22o_1
X_4831_ _1053_ _1347_ _1341_ _0983_ _1381_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7550_ net423 _3403_ _2198_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__a21o_1
X_4762_ _0698_ _0507_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7481_ _3629_ _3632_ vssd1 vssd1 vccd1 vccd1 _3633_ sky130_fd_sc_hd__xnor2_1
X_6501_ _2881_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
X_4693_ _1256_ net914 _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6432_ sound1.count\[4\] _2201_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6363_ _2766_ _2771_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8102_ clknet_leaf_95_hwclk sound2.osc.next_count\[3\] net68 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_6294_ _2289_ _2723_ _2724_ _2293_ sound1.sdiv.Q\[7\] vssd1 vssd1 vccd1 vccd1 _2725_
+ sky130_fd_sc_hd__a32o_1
X_5314_ _0997_ _1777_ _1792_ _1159_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__o22a_1
X_5245_ _1758_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
X_8033_ clknet_leaf_81_hwclk net400 net73 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold28 sound3.sdiv.Q\[26\] vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 sound4.sdiv.Q\[20\] vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold39 pm.count\[7\] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ sound3.count\[8\] _1706_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4127_ seq.player_5.state\[2\] net541 _0740_ _0741_ _0700_ vssd1 vssd1 vccd1 vccd1
+ seq.player_5.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4058_ _0698_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__inv_4
XFILLER_0_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7817_ clknet_leaf_2_hwclk net835 net70 vssd1 vssd1 vccd1 vccd1 seq.player_5.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_7748_ clknet_leaf_53_hwclk _0033_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_7679_ _3733_ _3734_ net654 _2183_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_62_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold509 net955 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_1
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _1547_ _1560_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__or2_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ sound2.divisor_m\[10\] _3246_ vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__xnor2_1
X_5932_ _2323_ _2367_ _2350_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__a21oi_1
X_5863_ _2281_ _2299_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5794_ _2240_ _2241_ _2239_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__a21o_1
X_7602_ _3680_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _0680_ _1336_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__or2_1
X_7533_ net124 _3654_ _3643_ net397 _3401_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__a221o_1
X_4745_ _1299_ _1300_ _1256_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7464_ sound3.sdiv.A\[22\] _3595_ vssd1 vssd1 vccd1 vccd1 _3618_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4676_ _0967_ _1004_ _1133_ _1110_ _0976_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__o32a_1
X_7395_ _3546_ _3549_ _3557_ vssd1 vssd1 vccd1 vccd1 _3558_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6415_ net686 _2830_ net736 vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__a21oi_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 mode_out[0] sky130_fd_sc_hd__buf_2
X_6346_ _2774_ _2775_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6277_ _2668_ _2671_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__or2_1
X_8016_ clknet_leaf_17_hwclk net139 net83 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_5228_ net853 _1744_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__and2_1
X_5159_ _1684_ _1689_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap60 _0684_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_12
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4530_ _1100_ _0959_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__or2_4
XFILLER_0_13_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold306 sound3.count_m\[17\] vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _0990_ _0973_ _0939_ _1010_ _1031_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__o221a_1
Xhold317 sound2.sdiv.A\[23\] vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ sound3.sdiv.Q\[3\] _0577_ _2633_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__and3_1
Xhold328 sound1.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__dlygate4sd3_1
X_7180_ net803 _2863_ vssd1 vssd1 vccd1 vccd1 _3391_ sky130_fd_sc_hd__and2_1
Xhold339 _0383_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6131_ _2560_ _2541_ _2554_ _2566_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__a31o_1
X_4392_ _0676_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__or2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _2472_ _2497_ _2477_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__a21o_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _0575_ _0563_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__nor2_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6964_ sound2.divisor_m\[8\] _3231_ vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__xnor2_1
X_5915_ sound4.count_m\[1\] sound4.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__and2b_1
X_6895_ sound2.divisor_m\[1\] _3169_ vssd1 vssd1 vccd1 vccd1 _3170_ sky130_fd_sc_hd__xnor2_1
X_5846_ _2275_ _2282_ _2283_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5777_ wave_comb.u1.A\[3\] _2224_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__nand2_1
X_7516_ sound3.sdiv.Q\[6\] _3440_ _3437_ net603 vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__a22o_1
X_4728_ sound1.count\[9\] sound1.count\[10\] _1278_ net978 vssd1 vssd1 vccd1 vccd1
+ _1288_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7447_ sound3.sdiv.A\[18\] _3595_ _3589_ vssd1 vssd1 vccd1 vccd1 _3604_ sky130_fd_sc_hd__o21a_1
X_4659_ _0680_ _0950_ _0939_ net60 _0992_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7378_ sound3.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _3542_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold840 sound1.count\[3\] vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 sound2.sdiv.Q\[7\] vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 sound2.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 rate_clk.count\[6\] vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
X_6329_ _2472_ _2497_ _2477_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3961_ inputcont.INTERNAL_SYNCED_I\[9\] _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5700_ _0576_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__buf_6
XFILLER_0_57_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3892_ sound3.sdiv.C\[4\] sound3.sdiv.C\[3\] sound3.sdiv.C\[2\] _0561_ sound3.sdiv.C\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__a311oi_4
X_6680_ sound1.divisor_m\[17\] _3037_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5631_ _2111_ _2113_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5562_ sound4.sdiv.A\[21\] _2038_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__xnor2_1
X_8350_ clknet_leaf_85_hwclk sound4.osc.next_count\[8\] net79 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[8\] sky130_fd_sc_hd__dfrtp_1
X_7301_ _3471_ _3473_ net438 _3463_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__a2bb2o_1
X_4513_ _0950_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8281_ clknet_leaf_64_hwclk net507 net79 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold114 sound3.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7232_ _3420_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__clkbuf_1
Xhold103 sound1.sdiv.Q\[10\] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5493_ _1988_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold125 sound4.count_m\[8\] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 sound1.count_m\[9\] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 sound4.sdiv.Q\[0\] vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold136 _0016_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ _0695_ _0964_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__nand2_8
X_4375_ _0945_ net60 vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__nor2_8
X_7163_ net166 _3167_ _3349_ net344 _3126_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold169 sound2.sdiv.Q\[24\] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
X_6114_ _2544_ _2546_ _2548_ _2549_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7094_ _3164_ _3347_ _3348_ _3174_ net607 vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__a32o_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ sound2.count_m\[1\] sound2.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__or2b_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ clknet_leaf_4_hwclk sound1.osc.next_count\[17\] net71 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6947_ _3215_ _3216_ vssd1 vssd1 vccd1 vccd1 _3217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6878_ net784 _1422_ _3142_ vssd1 vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5829_ _2269_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_57_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold681 sound2.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold670 sound4.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 sound2.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4160_ net639 _0761_ _0763_ vssd1 vssd1 vccd1 vccd1 seq.player_2.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4091_ seq.player_8.state\[2\] net859 vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7850_ clknet_leaf_98_hwclk seq.clk_div.next_count\[7\] net65 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6801_ net899 _2855_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7781_ clknet_leaf_59_hwclk _0055_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _1530_ _1531_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[12\] sky130_fd_sc_hd__nor2_1
X_6732_ net670 _2895_ sound1.sdiv.next_dived _3083_ vssd1 vssd1 vccd1 vccd1 _0131_
+ sky130_fd_sc_hd__a22o_1
X_3944_ inputcont.INTERNAL_SYNCED_I\[6\] inputcont.INTERNAL_SYNCED_I\[8\] vssd1 vssd1
+ vccd1 vccd1 _0608_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6663_ _3019_ _3021_ vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3875_ _0546_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__inv_2
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5614_ sound4.sdiv.A\[5\] _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6594_ _2956_ _2959_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8333_ clknet_leaf_56_hwclk net563 net96 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5545_ sound4.divisor_m\[6\] _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__or2_1
X_8264_ clknet_leaf_38_hwclk net158 net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5476_ _1779_ _1936_ _1974_ _1975_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__and4_1
X_8195_ clknet_leaf_27_hwclk _0316_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_7215_ _3409_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__clkbuf_1
X_4427_ _0959_ _0992_ _0993_ _0994_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__o32a_1
X_7146_ net598 _3168_ sound2.sdiv.next_dived net635 vssd1 vssd1 vccd1 vccd1 _0242_
+ sky130_fd_sc_hd__a22o_1
X_4358_ select1.sequencer_on seq.player_6.state\[3\] _0893_ vssd1 vssd1 vccd1 vccd1
+ _0929_ sky130_fd_sc_hd__and3_1
X_7077_ _3332_ _3333_ vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__xnor2_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ net545 net111 vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__or2b_1
X_6028_ sound2.count_m\[4\] vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7979_ clknet_leaf_5_hwclk sound1.osc.next_count\[0\] net72 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[0\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_49_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout64 net65 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_8
Xfanout86 net103 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_4
Xfanout97 net103 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_8
XFILLER_0_52_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout75 net82 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5330_ sound4.count\[9\] _1840_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5261_ _1769_ _1770_ _1771_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__and3_1
X_4212_ seq.clk_div.count\[8\] vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__inv_2
X_7000_ net445 _3168_ sound2.sdiv.next_dived _3264_ vssd1 vssd1 vccd1 vccd1 _0218_
+ sky130_fd_sc_hd__a22o_1
X_5192_ sound3.count\[0\] sound3.count\[1\] vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__or2_1
X_4143_ net725 net906 _0746_ net480 vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__a31o_1
X_4074_ _0705_ _0707_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__nor2_1
X_7902_ clknet_leaf_40_hwclk sound1.sdiv.next_dived net98 vssd1 vssd1 vccd1 vccd1
+ sound1.sdiv.dived sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7833_ clknet_leaf_5_hwclk net831 net72 vssd1 vssd1 vccd1 vccd1 seq.player_1.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_7764_ clknet_leaf_47_hwclk net581 net102 vssd1 vssd1 vccd1 vccd1 pm.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6715_ _3068_ _3063_ _3065_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__and3_1
X_4976_ net933 sound2.count\[7\] _1515_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7695_ net562 sound4.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3745_ sky130_fd_sc_hd__or2_1
X_3927_ _0590_ _0591_ _0523_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__o21a_1
X_6646_ _2996_ _3000_ _3007_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3858_ _0529_ _0530_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__and3_1
X_3789_ net1 wave.mode\[0\] vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6577_ _2944_ _2945_ net467 _2895_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5528_ pm.count\[3\] vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__inv_2
X_8316_ clknet_leaf_71_hwclk _0416_ net80 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8247_ clknet_leaf_39_hwclk _0347_ net100 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_5459_ sound4.count\[7\] sound4.count\[8\] _1955_ vssd1 vssd1 vccd1 vccd1 _1962_
+ sky130_fd_sc_hd__and3_1
X_8178_ clknet_leaf_29_hwclk _0299_ net92 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_7129_ _3349_ _3375_ _3376_ _3174_ net550 vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__a32o_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4830_ _1042_ _1336_ _1345_ _1154_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__o22a_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _0699_ net41 vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__and2_1
X_7480_ _3630_ _3631_ vssd1 vssd1 vccd1 vccd1 _3632_ sky130_fd_sc_hd__and2b_1
X_6500_ net757 _1120_ _2864_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__mux2_1
X_4692_ net472 net913 sound1.count\[2\] vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6431_ net527 _2836_ _2840_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6362_ _2764_ _2765_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5313_ _1126_ _1781_ _1790_ _1165_ _1823_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8101_ clknet_leaf_89_hwclk sound2.osc.next_count\[2\] net68 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_6293_ sound1.sdiv.Q\[6\] _0579_ _2722_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__a21o_1
X_5244_ _1756_ _1757_ _1721_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8032_ clknet_leaf_91_hwclk net265 net74 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold29 _0366_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _1701_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__and2_1
Xhold18 _0021_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dlygate4sd3_1
X_4126_ net833 _0738_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4057_ select1.sequencer_on vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__buf_6
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7816_ clknet_leaf_2_hwclk seq.player_5.next_state\[2\] net70 vssd1 vssd1 vccd1 vccd1
+ seq.player_5.state\[2\] sky130_fd_sc_hd__dfrtp_4
X_7747_ clknet_leaf_54_hwclk _0032_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4959_ _1470_ _1506_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7678_ _2045_ _2171_ _3732_ _1763_ vssd1 vssd1 vccd1 vccd1 _3734_ sky130_fd_sc_hd__a31o_1
X_6629_ _2991_ _2992_ net451 _2895_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6980_ _3177_ _3245_ vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5931_ _2360_ net57 _2345_ _2366_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__a31o_1
X_5862_ _2297_ _2298_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__nor2_1
X_5793_ _2239_ _2240_ _2241_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7601_ net922 _1913_ _2186_ vssd1 vssd1 vccd1 vccd1 _3680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4813_ _0960_ _1333_ _1345_ _0952_ _1363_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7532_ sound3.sdiv.Q\[21\] _3654_ _3643_ net209 _3400_ vssd1 vssd1 vccd1 vccd1 _0360_
+ sky130_fd_sc_hd__a221o_1
X_4744_ sound1.count\[15\] _1296_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7463_ _3615_ _3617_ net576 _3463_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4675_ _0994_ _1025_ _1038_ _0954_ _0990_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__o32a_1
X_7394_ _3555_ _3556_ vssd1 vssd1 vccd1 vccd1 _3557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6414_ net686 _2830_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__xor2_1
X_6345_ sound4.sdiv.Q\[6\] _2641_ _2736_ vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__a21oi_1
X_6276_ _2703_ _2707_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5227_ _1746_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
X_8015_ clknet_leaf_15_hwclk _0157_ net83 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5158_ _1012_ _1578_ _1686_ _1688_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__o211a_1
X_5089_ _1605_ _1609_ _1616_ _1619_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__or4_1
X_4109_ _0456_ net161 vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap61 _0565_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold307 _0285_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__dlygate4sd3_1
X_4460_ _0981_ _0997_ _1023_ _1030_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold329 sound3.sdiv.Q\[16\] vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__dlygate4sd3_1
X_4391_ _0869_ _0939_ _0943_ _0948_ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold318 sound2.count\[0\] vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__dlygate4sd3_1
X_6130_ _2565_ _2539_ sound3.divisor_m\[16\] _2538_ vssd1 vssd1 vccd1 vccd1 _2566_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _2491_ _2496_ _2479_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__a21o_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _1544_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6963_ sound2.sdiv.A\[26\] _3230_ vssd1 vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5914_ sound4.count_m\[17\] _2349_ _2322_ sound4.divisor_m\[17\] vssd1 vssd1 vccd1
+ vccd1 _2350_ sky130_fd_sc_hd__a2bb2o_1
X_6894_ sound2.sdiv.A\[26\] sound2.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5845_ _2275_ _2279_ _2282_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__nor3_1
XFILLER_0_91_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5776_ wave_comb.u1.A\[3\] _2224_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__or2_1
X_7515_ sound3.sdiv.Q\[5\] _3463_ _3437_ net516 vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__a22o_1
X_4727_ sound1.count\[10\] sound1.count\[11\] _1281_ vssd1 vssd1 vccd1 vccd1 _1287_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7446_ _3573_ _3581_ _3582_ vssd1 vssd1 vccd1 vccd1 _3603_ sky130_fd_sc_hd__o21a_1
X_4658_ _0981_ _0994_ _0687_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold830 _1520_ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__dlygate4sd3_1
X_7377_ _3437_ _3540_ _3541_ _3440_ net211 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__a32o_1
Xhold863 pm.count\[3\] vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 sound3.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 sound1.count\[10\] vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
X_4589_ _0685_ _0981_ _0939_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__o22a_1
X_6328_ _2756_ _2757_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__xor2_1
Xhold874 sound1.count\[11\] vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6259_ sound1.sdiv.Q\[5\] _2690_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3960_ _0622_ _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3891_ sound3.sdiv.start vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5630_ sound4.divisor_m\[3\] _2112_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5561_ _2043_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7300_ _1545_ _3472_ vssd1 vssd1 vccd1 vccd1 _3473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5492_ sound4.count\[15\] _1984_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__and2_2
X_4512_ _0694_ _0996_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_4
XFILLER_0_14_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8280_ clknet_leaf_65_hwclk net220 net80 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold126 sound3.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7231_ net764 _1649_ _3419_ vssd1 vssd1 vccd1 vccd1 _3420_ sky130_fd_sc_hd__mux2_1
Xhold104 _0152_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold115 sound4.count_m\[13\] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold137 sound3.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _0079_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _0001_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _1013_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4374_ _0686_ _0680_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nor2_4
X_7162_ sound2.sdiv.Q\[18\] _3167_ _3349_ net338 _3125_ vssd1 vssd1 vccd1 vccd1 _0258_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6113_ _2514_ sound3.divisor_m\[6\] sound3.divisor_m\[5\] _2511_ vssd1 vssd1 vccd1
+ vccd1 _2549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7093_ _3336_ _3343_ _3346_ vssd1 vssd1 vccd1 vccd1 _3348_ sky130_fd_sc_hd__nand3_1
XFILLER_0_95_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ sound2.count_m\[0\] vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__inv_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7995_ clknet_leaf_4_hwclk sound1.osc.next_count\[16\] net71 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[16\] sky130_fd_sc_hd__dfrtp_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6946_ _3211_ _3214_ vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6877_ _3158_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5828_ _0569_ _2268_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5759_ _2207_ _2212_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7429_ sound3.divisor_m\[18\] _3587_ vssd1 vssd1 vccd1 vccd1 _3588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold660 sound3.divisor_m\[7\] vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 seq.player_2.state\[2\] vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 sound2.divisor_m\[10\] vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 sound2.divisor_m\[12\] vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4090_ seq.player_8.state\[2\] net537 _0715_ _0716_ _0700_ vssd1 vssd1 vccd1 vccd1
+ seq.player_8.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_6800_ sound1.sdiv.Q\[27\] _2894_ _2890_ net151 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7780_ clknet_leaf_59_hwclk _0054_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_4992_ net723 _1527_ _1504_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__o21ai_1
X_6731_ _3081_ _3082_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3943_ inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__inv_2
X_6662_ _3019_ _3021_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3874_ _0512_ _0544_ _0534_ _0545_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__o211a_2
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5613_ _2095_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6593_ _2956_ _2959_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__nor2_1
X_8332_ clknet_leaf_68_hwclk _0432_ net82 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5544_ sound4.divisor_m\[5\] sound4.divisor_m\[4\] _2026_ vssd1 vssd1 vccd1 vccd1
+ _2027_ sky130_fd_sc_hd__or3_1
X_8263_ clknet_leaf_37_hwclk _0363_ net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5475_ sound4.count\[9\] sound4.count\[10\] _1962_ sound4.count\[11\] vssd1 vssd1
+ vccd1 vccd1 _1975_ sky130_fd_sc_hd__a31o_1
X_8194_ clknet_leaf_27_hwclk _0315_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_7214_ net937 _3408_ _3142_ vssd1 vssd1 vccd1 vccd1 _3409_ sky130_fd_sc_hd__mux2_1
X_4426_ net60 _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__nor2_8
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7145_ net646 sound2.sdiv.next_dived _2501_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4357_ select1.sequencer_on _0896_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__and3_1
X_7076_ _3322_ _3325_ _3321_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__a21bo_1
X_4288_ net494 _0859_ _0862_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[21\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ sound2.count_m\[5\] vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__inv_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7978_ clknet_leaf_31_hwclk sound1.sdiv.next_start net90 vssd1 vssd1 vccd1 vccd1
+ sound1.sdiv.start sky130_fd_sc_hd__dfrtp_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _3187_ _3191_ _3199_ vssd1 vssd1 vccd1 vccd1 _3201_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout65 net2 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_6
Xfanout98 net100 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_8
Xfanout87 net88 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_8
XFILLER_0_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout76 net82 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__buf_8
XFILLER_0_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold490 inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_41_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5260_ _0698_ _0605_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__or2_2
X_4211_ _0789_ seq.clk_div.count\[14\] _0782_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__o21ai_1
X_5191_ net428 _1721_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[0\] sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_56_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_4142_ _0750_ _0749_ _0751_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_4.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
X_4073_ _0704_ _0707_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__nor2_1
X_7901_ clknet_leaf_95_hwclk net117 net66 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_7832_ clknet_leaf_5_hwclk seq.player_1.next_state\[2\] net71 vssd1 vssd1 vccd1 vccd1
+ seq.player_1.state\[2\] sky130_fd_sc_hd__dfrtp_2
X_7763_ clknet_leaf_50_hwclk net548 net102 vssd1 vssd1 vccd1 vccd1 pm.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_4975_ _1518_ _1519_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6714_ _3063_ _3065_ _3068_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _0515_ _0521_ _0519_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__o21ba_1
X_7694_ net562 sound4.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3744_ sky130_fd_sc_hd__nand2_1
X_6645_ _3005_ _3006_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3857_ _0525_ _0526_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6576_ _2942_ _2943_ _0866_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3788_ _0468_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_2
X_5527_ _0651_ pm.current_waveform\[4\] vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__and2_1
X_8315_ clknet_leaf_72_hwclk _0415_ net80 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_8246_ clknet_leaf_46_hwclk _0346_ net100 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5458_ _1961_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
X_8177_ clknet_3_5__leaf_hwclk _0298_ net91 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_4409_ _0918_ _0909_ _0949_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__or3b_1
X_5389_ _1017_ _1784_ _1781_ _1020_ _1899_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7128_ net550 sound2.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3376_ sky130_fd_sc_hd__or2_1
X_7059_ _3164_ _3316_ _3317_ _3174_ net295 vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a32o_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4760_ _1311_ vssd1 vssd1 vccd1 vccd1 sound2.sdiv.next_dived sky130_fd_sc_hd__buf_4
XFILLER_0_28_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4691_ sound1.count\[0\] net913 sound1.count\[2\] vssd1 vssd1 vccd1 vccd1 _1260_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6430_ sound1.count\[3\] _2201_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6361_ wave_comb.u1.next_start _2789_ _2790_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5312_ _1004_ _1038_ _1786_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8100_ clknet_leaf_89_hwclk sound2.osc.next_count\[1\] net69 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[1\] sky130_fd_sc_hd__dfrtp_1
X_6292_ sound1.sdiv.Q\[6\] _2722_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5243_ net845 sound3.count\[16\] _1750_ sound3.count\[17\] vssd1 vssd1 vccd1 vccd1
+ _1757_ sky130_fd_sc_hd__a31o_1
X_8031_ clknet_leaf_81_hwclk net374 net74 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold19 net817 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_1
X_5174_ _1591_ _1703_ _1587_ _1704_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__and4_1
X_4125_ seq.player_5.state\[0\] seq.player_5.state\[1\] _0737_ vssd1 vssd1 vccd1 vccd1
+ _0740_ sky130_fd_sc_hd__and3_1
X_4056_ _0682_ _0683_ _0694_ _0697_ vssd1 vssd1 vccd1 vccd1 oct.next_state\[2\] sky130_fd_sc_hd__a211o_1
XFILLER_0_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7815_ clknet_leaf_2_hwclk net542 net70 vssd1 vssd1 vccd1 vccd1 seq.player_5.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7746_ clknet_leaf_55_hwclk _0031_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4958_ _1507_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3909_ _0575_ net62 vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nor2_8
XFILLER_0_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7677_ _2171_ _3732_ _2045_ vssd1 vssd1 vccd1 vccd1 _3733_ sky130_fd_sc_hd__a21oi_1
X_4889_ _0696_ _1343_ _1436_ _1439_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6628_ _2989_ _2990_ _0866_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6559_ sound1.divisor_m\[5\] _2928_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8229_ clknet_leaf_32_hwclk sound3.osc.next_count\[10\] net87 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5930_ sound4.count_m\[15\] _2341_ _2365_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__a21oi_1
X_5861_ _2294_ _2296_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7600_ _2005_ _1018_ _1779_ _3679_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5792_ _2233_ _2234_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4812_ _1039_ _1347_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__or2_1
X_7531_ net209 _3654_ _3643_ net391 _3399_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__a221o_1
X_4743_ sound1.count\[15\] _1296_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7462_ _2863_ _0563_ _3616_ vssd1 vssd1 vccd1 vccd1 _3617_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4674_ _1018_ _0959_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__or2_2
X_6413_ _0811_ _2829_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7393_ _3551_ _3554_ vssd1 vssd1 vccd1 vccd1 _3556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6344_ sound4.sdiv.Q\[7\] _0576_ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6275_ _2289_ _2705_ _2706_ _2290_ sound4.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 _2707_
+ sky130_fd_sc_hd__a32o_1
X_5226_ _1744_ _1745_ _1721_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__and3b_1
X_8014_ clknet_leaf_13_hwclk _0156_ net85 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5157_ _1053_ _1572_ _1550_ _1125_ _1687_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__o221a_1
X_5088_ sound3.count\[18\] _1618_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__xnor2_1
X_4108_ net849 _0725_ _0728_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_7.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_4039_ _0674_ _0678_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__nor2_8
XFILLER_0_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ clknet_leaf_64_hwclk net402 net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap62 _0562_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold308 sound3.count_m\[8\] vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4390_ _0950_ _0954_ _0958_ _0960_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__o22a_1
Xhold319 sound4.count_m\[11\] vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _2493_ _2495_ _2459_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__o21ai_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _1504_ _1542_ _1543_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__and3_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6962_ sound2.divisor_m\[7\] _3221_ vssd1 vssd1 vccd1 vccd1 _3230_ sky130_fd_sc_hd__nor2_1
X_5913_ sound4.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__inv_2
X_6893_ _3164_ _3165_ _3166_ _3168_ net489 vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__a32o_1
X_5844_ _2276_ _2277_ _2281_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7514_ net516 _3463_ _3437_ net653 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5775_ net618 _0573_ wave_comb.u1.next_dived _2226_ vssd1 vssd1 vccd1 vccd1 _0031_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4726_ _1286_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_3__f_hwclk clknet_0_hwclk vssd1 vssd1 vccd1 vccd1 clknet_3_3__leaf_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_7445_ _3564_ _3568_ _3575_ _3583_ _3601_ vssd1 vssd1 vccd1 vccd1 _3602_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_114_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4657_ _1220_ _1221_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7376_ _3529_ _3532_ _3539_ vssd1 vssd1 vccd1 vccd1 _3541_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold820 sound4.divisor_m\[4\] vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6327_ sound2.sdiv.Q\[7\] _0578_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__nand2_1
Xhold842 sound1.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 sound1.count\[13\] vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
X_4588_ _1100_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__or2_2
Xhold864 sound1.count\[18\] vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold831 seq.clk_div.count\[1\] vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold875 sound2.sdiv.A\[21\] vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
X_6258_ sound1.sdiv.Q\[4\] _2656_ _2657_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__a21bo_1
X_6189_ _2279_ _2620_ _2622_ _2292_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__o22a_1
X_5209_ _1734_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3890_ _0559_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5560_ sound4.sdiv.A\[22\] _2038_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__xor2_2
XFILLER_0_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4511_ _0680_ _0976_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5491_ _1987_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7230_ _2863_ vssd1 vssd1 vccd1 vccd1 _3419_ sky130_fd_sc_hd__buf_8
Xhold105 sound3.sdiv.Q\[20\] vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ _0944_ _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold116 _0380_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _0307_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold149 sound1.sdiv.Q\[13\] vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 sound4.sdiv.Q\[18\] vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__dlygate4sd3_1
X_7161_ net338 _3167_ _3349_ net382 _3124_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4373_ _0674_ _0677_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__nor2_8
X_6112_ _2547_ sound3.divisor_m\[8\] _2513_ sound3.divisor_m\[7\] vssd1 vssd1 vccd1
+ vccd1 _2548_ sky130_fd_sc_hd__a22o_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7092_ _3336_ _3343_ _3346_ vssd1 vssd1 vccd1 vccd1 _3347_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ sound2.count_m\[16\] _2471_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__and2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7994_ clknet_leaf_4_hwclk sound1.osc.next_count\[15\] net71 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _3211_ _3214_ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__or2_1
X_6876_ net787 _3157_ _3142_ vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5827_ _0571_ _2267_ net865 vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5758_ wave_comb.u1.A\[0\] _2211_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4709_ _1272_ _1273_ _1256_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__and3b_1
XFILLER_0_32_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7428_ sound3.divisor_m\[17\] _3578_ _3448_ vssd1 vssd1 vccd1 vccd1 _3587_ sky130_fd_sc_hd__o21a_1
X_5689_ sound4.sdiv.A\[23\] _2038_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7359_ sound3.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _3525_ sky130_fd_sc_hd__inv_2
Xhold661 sound1.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 seq.player_2.next_state\[2\] vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 sound2.divisor_m\[9\] vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold694 sound1.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 sound2.divisor_m\[13\] vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6730_ sound1.sdiv.A\[21\] _3055_ _3079_ vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4991_ net823 _1527_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _0587_ _0606_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__nand2_8
XFILLER_0_46_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6661_ sound1.divisor_m\[15\] _3020_ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__xnor2_1
X_3873_ _0520_ _0524_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__nand2_1
X_6592_ sound1.divisor_m\[8\] _2958_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5612_ sound4.divisor_m\[6\] _2094_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8331_ clknet_leaf_68_hwclk net718 net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_5543_ sound4.divisor_m\[3\] sound4.divisor_m\[2\] sound4.divisor_m\[1\] sound4.divisor_m\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8262_ clknet_leaf_37_hwclk net125 net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_5474_ _1973_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__inv_2
X_8193_ clknet_leaf_29_hwclk _0314_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_7213_ _1673_ vssd1 vssd1 vccd1 vccd1 _3408_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4425_ _0995_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__clkbuf_16
X_7144_ sound2.sdiv.next_dived _3386_ _2276_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__a21bo_1
X_4356_ seq.player_7.state\[3\] _0897_ _0901_ seq.player_8.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _0927_ sky130_fd_sc_hd__a22o_1
X_7075_ _3330_ _3331_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__or2b_1
X_4287_ net494 _0859_ _0813_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__o21ai_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ sound2.count_m\[7\] _2460_ _2461_ sound2.divisor_m\[7\] vssd1 vssd1 vccd1
+ vccd1 _2462_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7977_ clknet_leaf_31_hwclk _0140_ net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ _3187_ _3191_ _3199_ vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_92_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6859_ _3146_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout99 net100 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_8
Xfanout88 net103 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout66 net69 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_6
Xfanout77 net79 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__buf_6
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold480 sound2.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 sound2.sdiv.A\[19\] vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4210_ seq.clk_div.count\[10\] _0779_ _0777_ _0803_ vssd1 vssd1 vccd1 vccd1 _0804_
+ sky130_fd_sc_hd__o211a_1
X_5190_ _1720_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4141_ net752 _0748_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__xor2_1
X_4072_ _0701_ _0707_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__nor2_1
X_7900_ clknet_leaf_0_hwclk net191 net64 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7831_ clknet_leaf_5_hwclk net566 net71 vssd1 vssd1 vccd1 vccd1 seq.player_1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_7762_ clknet_leaf_50_hwclk pm.next_count\[1\] net102 vssd1 vssd1 vccd1 vccd1 pm.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4974_ net715 _1515_ _1504_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__o21ai_1
X_6713_ _3066_ _3067_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__nand2_1
X_7693_ _3743_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__clkbuf_1
X_3925_ _0548_ _0543_ _0582_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__nand3_2
XFILLER_0_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6644_ _3001_ _3004_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3856_ inputcont.INTERNAL_SYNCED_I\[3\] _0502_ _0512_ vssd1 vssd1 vccd1 vccd1 _0530_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6575_ _2942_ _2943_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3787_ _0462_ _0467_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or2_1
X_5526_ _2009_ pm.current_waveform\[5\] vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__and2_1
X_8314_ clknet_leaf_71_hwclk _0414_ net80 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_8245_ clknet_leaf_46_hwclk net604 net100 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_5457_ _1779_ _1936_ _1959_ _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__and4_1
X_4408_ _0978_ _0971_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__or2_4
X_8176_ clknet_leaf_27_hwclk _0297_ net92 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_5388_ _1025_ _1794_ _1796_ _1027_ _1898_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4339_ seq.player_7.state\[0\] _0898_ _0901_ seq.player_8.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _0910_ sky130_fd_sc_hd__a22o_1
X_7127_ net550 sound2.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7058_ _3302_ _3306_ _3315_ vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6009_ sound2.count_m\[10\] _2443_ _2444_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _1259_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6360_ net667 _0572_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5311_ _1811_ _1812_ _1818_ _1821_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6291_ sound1.sdiv.Q\[5\] _2656_ _2690_ vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8030_ clknet_leaf_90_hwclk _0172_ net68 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5242_ sound3.count\[16\] sound3.count\[17\] _1753_ vssd1 vssd1 vccd1 vccd1 _1756_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_87_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5173_ _1025_ _1046_ _1559_ _1578_ _1165_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__o32a_1
X_4124_ net624 _0737_ _0739_ vssd1 vssd1 vccd1 vccd1 seq.player_5.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
Xinput1 cs vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_6
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4055_ _0682_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__nor2_1
X_7814_ clknet_leaf_2_hwclk net625 net70 vssd1 vssd1 vccd1 vccd1 seq.player_5.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7745_ clknet_leaf_55_hwclk _0030_ net95 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4957_ _1504_ _1505_ _1506_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__and3_1
X_7676_ _2042_ _2168_ vssd1 vssd1 vccd1 vccd1 _3732_ sky130_fd_sc_hd__or2b_1
X_3908_ _0576_ vssd1 vssd1 vccd1 vccd1 sound4.sdiv.next_start sky130_fd_sc_hd__inv_2
X_4888_ _1123_ _1339_ _1336_ _1141_ _1438_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6627_ _2989_ _2990_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3839_ _0480_ _0481_ _0482_ _0483_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6558_ sound1.divisor_m\[4\] _2919_ _2903_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6489_ net701 _2005_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__nor2_1
X_5509_ net154 vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[0\] sky130_fd_sc_hd__inv_2
X_8228_ clknet_leaf_33_hwclk sound3.osc.next_count\[9\] net87 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[9\] sky130_fd_sc_hd__dfrtp_1
X_8159_ clknet_leaf_31_hwclk net301 net91 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5860_ _2294_ _2296_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _1015_ _1323_ _1327_ _0946_ _1361_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5791_ net986 wave_comb.u1.A\[3\] _2224_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7530_ sound3.sdiv.Q\[19\] _3654_ _3643_ net342 _3398_ vssd1 vssd1 vccd1 vccd1 _0358_
+ sky130_fd_sc_hd__a221o_1
X_4742_ _1298_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7461_ _3613_ _3614_ _3612_ vssd1 vssd1 vccd1 vccd1 _3616_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4673_ _0985_ _0939_ _1242_ _0950_ _1243_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__o221a_1
X_6412_ _0719_ seq.encode.play vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__nand2_1
X_7392_ _3551_ _3554_ vssd1 vssd1 vccd1 vccd1 _3555_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6343_ net30 net29 vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6274_ sound4.sdiv.Q\[5\] _2704_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5225_ sound3.count\[9\] net802 _1738_ sound3.count\[11\] vssd1 vssd1 vccd1 vccd1
+ _1745_ sky130_fd_sc_hd__a31o_1
X_8013_ clknet_leaf_13_hwclk net254 net85 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5156_ _0983_ _1580_ _1565_ _1146_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__o22a_1
X_5087_ _0695_ _1617_ _1591_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__o21a_1
X_4107_ net726 net814 _0722_ net496 vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a31o_1
X_4038_ net930 inputcont.INTERNAL_OCTAVE_INPUT vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _2384_ _2424_ _2377_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__a21o_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7728_ clknet_leaf_64_hwclk net406 net78 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7659_ _3719_ _2154_ vssd1 vssd1 vccd1 vccd1 _3721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap52 net53 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xmax_cap63 _0559_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold309 _0276_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ sound2.count\[18\] _1539_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__nand2_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6961_ net965 vssd1 vssd1 vccd1 vccd1 _3229_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5912_ sound4.divisor_m\[3\] sound4.count_m\[2\] vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__or2b_1
X_6892_ _3167_ vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5843_ sound2.sdiv.Q\[0\] _0578_ _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7513_ sound3.sdiv.Q\[3\] _3463_ sound3.sdiv.next_dived net643 vssd1 vssd1 vccd1
+ vccd1 _0342_ sky130_fd_sc_hd__a22o_1
X_5774_ _2222_ _2225_ vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4725_ _1256_ _1284_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7444_ _3600_ vssd1 vssd1 vccd1 vccd1 _3601_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4656_ sound1.count\[11\] _1050_ _1224_ _1226_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7375_ _3529_ _3532_ _3539_ vssd1 vssd1 vccd1 vccd1 _3540_ sky130_fd_sc_hd__or3b_1
Xhold810 _1260_ vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 sound2.count\[1\] vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__dlygate4sd3_1
X_4587_ _0685_ _0982_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold843 wave_comb.u1.A\[7\] vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__dlygate4sd3_1
X_6326_ sound2.sdiv.Q\[6\] _2660_ _2718_ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__a21oi_1
Xhold854 _1297_ vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 _0816_ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 sound1.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 sound1.count\[0\] vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6257_ _2687_ _2688_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__nand2_1
X_6188_ _2586_ _2621_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__xor2_1
X_5208_ _1732_ _1733_ _1721_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__and3b_1
X_5139_ _0869_ _1567_ _1550_ _0954_ _1669_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4510_ _0990_ _0960_ _0994_ _1039_ _1080_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5490_ _1779_ _1936_ _1985_ _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__and4_1
Xhold106 _0360_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _0675_ _0970_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__nor2_8
Xhold117 sound2.sdiv.A\[8\] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold128 sound4.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlygate4sd3_1
X_7160_ sound2.sdiv.Q\[16\] _3167_ _3349_ net345 _3123_ vssd1 vssd1 vccd1 vccd1 _0256_
+ sky130_fd_sc_hd__a221o_1
Xhold139 _0018_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__dlygate4sd3_1
X_6111_ sound3.count_m\[7\] vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__inv_2
X_4372_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__buf_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7091_ _3345_ vssd1 vssd1 vccd1 vccd1 _3346_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ sound2.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__inv_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7993_ clknet_leaf_16_hwclk sound1.osc.next_count\[14\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[14\] sky130_fd_sc_hd__dfrtp_1
X_6944_ sound2.divisor_m\[6\] _3213_ vssd1 vssd1 vccd1 vccd1 _3214_ sky130_fd_sc_hd__xnor2_1
X_6875_ _1434_ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__inv_2
X_5826_ _0646_ _2266_ _2267_ _0573_ net614 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5757_ wave_comb.u1.M\[1\] _2210_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4708_ sound1.count\[6\] _1269_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7427_ sound3.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 _3586_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5688_ sound4.sdiv.A\[20\] sound4.sdiv.A\[19\] _2038_ vssd1 vssd1 vccd1 vccd1 _2171_
+ sky130_fd_sc_hd__o21ai_4
X_4639_ _0949_ _0988_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7358_ _3437_ _3523_ _3524_ _3440_ net206 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__a32o_1
Xhold640 sound3.divisor_m\[9\] vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 sound1.divisor_m\[11\] vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 sound4.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
X_7289_ _0577_ vssd1 vssd1 vccd1 vccd1 _3463_ sky130_fd_sc_hd__clkbuf_8
X_6309_ _2735_ _2739_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__xnor2_1
Xhold673 sound4.divisor_m\[5\] vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 sound2.divisor_m\[6\] vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 sound4.divisor_m\[11\] vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4990_ _1529_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3941_ _0588_ _0589_ _0598_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__o31a_4
XFILLER_0_128_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6660_ sound1.divisor_m\[14\] _3011_ _2903_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3872_ inputcont.INTERNAL_SYNCED_I\[3\] _0502_ _0543_ vssd1 vssd1 vccd1 vccd1 _0544_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6591_ sound1.sdiv.A\[26\] _2957_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5611_ _2036_ _2027_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__and2_1
X_5542_ net651 _2024_ _2025_ vssd1 vssd1 vccd1 vccd1 pm.next_pwm_o sky130_fd_sc_hd__o21a_1
X_8330_ clknet_leaf_68_hwclk net283 net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8261_ clknet_leaf_34_hwclk _0361_ net88 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_5473_ sound4.count\[10\] sound4.count\[11\] _1966_ vssd1 vssd1 vccd1 vccd1 _1973_
+ sky130_fd_sc_hd__and3_1
X_8192_ clknet_leaf_28_hwclk _0313_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7212_ _3407_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__clkbuf_1
X_4424_ _0686_ _0674_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__nor2_1
X_4355_ net36 _0925_ _0698_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__mux2_2
X_7143_ _3373_ _3385_ vssd1 vssd1 vccd1 vccd1 _3386_ sky130_fd_sc_hd__nand2_1
X_7074_ sound2.sdiv.A\[18\] _3329_ vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__nand2_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _0861_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[20\] sky130_fd_sc_hd__clkbuf_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ sound2.count_m\[6\] vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__inv_2
X_7976_ clknet_leaf_24_hwclk _0139_ net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _3197_ _3198_ vssd1 vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6858_ net745 _3145_ _3142_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout89 net103 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__buf_8
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5809_ wave_comb.u1.A\[8\] _2224_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__or2_1
Xfanout78 net79 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_6
Xfanout67 net69 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6789_ net138 _2893_ _0867_ net153 _2846_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold470 _0146_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 sound1.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 sound1.sdiv.C\[2\] vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ net906 seq.player_4.state\[3\] vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__nand2_1
X_4071_ seq.beat\[3\] net51 vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__nand2_8
X_7830_ clknet_leaf_7_hwclk net932 net71 vssd1 vssd1 vccd1 vccd1 seq.player_1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7761_ clknet_leaf_51_hwclk pm.next_count\[0\] net101 vssd1 vssd1 vccd1 vccd1 pm.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4973_ net715 _1515_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6712_ sound1.sdiv.A\[19\] _3055_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__nand2_1
X_7692_ _1764_ _2182_ net801 vssd1 vssd1 vccd1 vccd1 _3743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3924_ _0584_ _0585_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6643_ _3001_ _3004_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3855_ _0513_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6574_ _2932_ _2933_ _2930_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__o21a_1
X_3786_ inputcont.INTERNAL_SYNCED_I\[8\] _0448_ _0455_ _0466_ vssd1 vssd1 vccd1 vccd1
+ _0467_ sky130_fd_sc_hd__a211o_1
X_5525_ pm.count\[5\] vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__inv_2
X_8313_ clknet_leaf_71_hwclk _0413_ net80 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_8244_ clknet_leaf_47_hwclk net517 net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5456_ sound4.count\[7\] _1955_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__or2_1
X_4407_ _0685_ _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__nor2_4
X_8175_ clknet_leaf_29_hwclk _0296_ net91 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_5387_ _1024_ _1028_ _1786_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4338_ net35 _0908_ _0698_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__mux2_4
X_7126_ _3374_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_7057_ _3302_ _3306_ _3315_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__o21ai_1
X_4269_ _0849_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
X_6008_ sound2.divisor_m\[10\] sound2.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2444_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ clknet_leaf_21_hwclk _0122_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6290_ _2289_ _2719_ _2720_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__and3_1
X_5310_ sound4.count\[16\] _1820_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5241_ net367 _1753_ _1755_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[16\] sky130_fd_sc_hd__a21oi_1
X_5172_ _1159_ _1567_ _1565_ _0997_ _1702_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__o221a_1
X_4123_ seq.player_5.state\[1\] seq.player_5.state\[2\] seq.player_5.state\[3\] _0738_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__a311o_1
Xinput2 n_rst vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_8
X_4054_ _0695_ _0687_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__nand2_4
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7813_ clknet_leaf_100_hwclk net843 net64 vssd1 vssd1 vccd1 vccd1 seq.player_6.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_7744_ clknet_leaf_55_hwclk net366 net95 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4956_ sound2.count\[0\] sound2.count\[1\] vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3907_ _0575_ _0556_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__nor2_4
X_7675_ net688 _2184_ _3681_ _3731_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__a22o_1
X_4887_ _1138_ _1323_ _1341_ _1126_ _1437_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__o221a_1
X_6626_ _2970_ _2980_ _2976_ _2979_ _2974_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__o32a_1
XFILLER_0_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3838_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__buf_2
X_6557_ net980 vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5508_ _2000_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3769_ inputcont.INTERNAL_SYNCED_I\[5\] _0443_ inputcont.INTERNAL_SYNCED_I\[4\] inputcont.INTERNAL_SYNCED_I\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__or4b_2
XFILLER_0_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6488_ _2873_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8227_ clknet_leaf_33_hwclk sound3.osc.next_count\[8\] net87 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[8\] sky130_fd_sc_hd__dfrtp_1
X_5439_ _1779_ _1936_ _1945_ _1946_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__and4_1
X_8158_ clknet_leaf_31_hwclk net348 net91 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_7109_ _3346_ _3350_ _3355_ vssd1 vssd1 vccd1 vccd1 _3361_ sky130_fd_sc_hd__or3b_1
X_8089_ clknet_leaf_72_hwclk _0231_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4810_ _0684_ _1077_ _1343_ _1338_ _0971_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__o32a_1
X_5790_ _2237_ _2238_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4741_ _1296_ net958 _1256_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__and3b_1
X_7460_ _3612_ _3613_ _3614_ vssd1 vssd1 vccd1 vccd1 _3615_ sky130_fd_sc_hd__and3_1
X_4672_ _0958_ _0944_ _1004_ _1025_ _0981_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__o32a_1
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6411_ _2828_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7391_ sound3.divisor_m\[14\] _3553_ vssd1 vssd1 vccd1 vccd1 _3554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6342_ _2766_ _2771_ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6273_ sound4.sdiv.Q\[5\] _0576_ _2704_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__a21o_1
X_5224_ sound3.count\[10\] sound3.count\[11\] _1741_ vssd1 vssd1 vccd1 vccd1 _1744_
+ sky130_fd_sc_hd__and3_1
X_8012_ clknet_leaf_13_hwclk _0154_ net86 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5155_ _1134_ _1567_ _1570_ _1154_ _1685_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5086_ net60 _1603_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__nand2_1
X_4106_ net849 _0725_ _0727_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_7.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4037_ _0676_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__nor2_4
XFILLER_0_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _2387_ _2423_ _2386_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__a21bo_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7727_ clknet_leaf_64_hwclk net150 net78 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_4939_ _1189_ _1327_ _1365_ _0959_ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__o221a_1
X_7658_ _3719_ _2154_ vssd1 vssd1 vccd1 vccd1 _3720_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6609_ _0866_ _2972_ _2973_ sound1.sdiv.next_start _2974_ vssd1 vssd1 vccd1 vccd1
+ _0117_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_104_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7589_ net892 _1875_ _2186_ vssd1 vssd1 vccd1 vccd1 _3673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6960_ _3164_ _3227_ _3228_ _3174_ net205 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5911_ _2316_ sound4.divisor_m\[7\] _2318_ sound4.divisor_m\[6\] vssd1 vssd1 vccd1
+ vccd1 _2347_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6891_ _0578_ vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__buf_6
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5842_ _2279_ _2277_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5773_ wave_comb.u1.A\[2\] _2224_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7512_ net643 _3463_ sound3.sdiv.next_dived net658 vssd1 vssd1 vccd1 vccd1 _0341_
+ sky130_fd_sc_hd__a22o_1
X_4724_ sound1.count\[10\] _1281_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7443_ _3591_ _3596_ vssd1 vssd1 vccd1 vccd1 _3600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4655_ sound1.count\[17\] _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7374_ _3537_ _3538_ vssd1 vssd1 vccd1 vccd1 _3539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold800 sound3.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__dlygate4sd3_1
X_4586_ _1150_ _1153_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__and3_2
Xhold811 seq.encode.keys_edge_det\[4\] vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 sound3.divisor_m\[1\] vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__dlygate4sd3_1
X_6325_ _2292_ _2751_ _2754_ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__o21a_1
Xhold855 sound1.count\[17\] vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold844 seq.clk_div.count\[0\] vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 sound2.count\[18\] vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 sound3.count\[18\] vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 seq.clk_div.count\[20\] vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6256_ sound2.sdiv.Q\[5\] _2686_ _2292_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__a21oi_1
X_6187_ sound1.sdiv.Q\[0\] sound1.sdiv.Q\[1\] sound1.sdiv.Q\[2\] _0579_ _2434_ vssd1
+ vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__o311a_1
X_5207_ sound3.count\[4\] _1728_ sound3.count\[5\] vssd1 vssd1 vccd1 vccd1 _1733_
+ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_54_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5138_ _0959_ _0993_ _1580_ _1562_ _0985_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__o32a_1
X_5069_ _1126_ _1580_ _1598_ _1599_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold107 sound3.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dlygate4sd3_1
X_4440_ _0695_ _0678_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__or2_4
XFILLER_0_41_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold118 sound4.sdiv.Q\[8\] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold129 sound2.count_m\[7\] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlygate4sd3_1
X_6110_ sound3.count_m\[17\] _2543_ _2545_ sound3.divisor_m\[17\] vssd1 vssd1 vccd1
+ vccd1 _2546_ sky130_fd_sc_hd__a2bb2o_1
X_4371_ _0940_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ sound2.sdiv.A\[20\] _3329_ vssd1 vssd1 vccd1 vccd1 _3345_ sky130_fd_sc_hd__xor2_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ sound2.count_m\[17\] _2470_ sound2.count_m\[18\] vssd1 vssd1 vccd1 vccd1 _2477_
+ sky130_fd_sc_hd__a21o_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7992_ clknet_leaf_4_hwclk sound1.osc.next_count\[13\] net71 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[13\] sky130_fd_sc_hd__dfrtp_4
X_6943_ _3177_ _3212_ vssd1 vssd1 vccd1 vccd1 _3213_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6874_ _3156_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
X_5825_ wave_comb.u1.C\[2\] wave_comb.u1.C\[0\] wave_comb.u1.C\[1\] vssd1 vssd1 vccd1
+ vccd1 _2267_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5756_ wave_comb.u1.M\[0\] _2209_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4707_ sound1.count\[6\] _1269_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__and2_1
X_5687_ sound4.sdiv.A\[22\] sound4.sdiv.A\[21\] _2038_ vssd1 vssd1 vccd1 vccd1 _2170_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7426_ net457 _3463_ sound3.sdiv.next_dived _3585_ vssd1 vssd1 vccd1 vccd1 _0323_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4638_ sound1.count\[3\] _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 sound3.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7357_ _3503_ _3507_ _3521_ _3511_ _3520_ vssd1 vssd1 vccd1 vccd1 _3524_ sky130_fd_sc_hd__a311o_1
Xhold663 sound3.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 sound1.divisor_m\[7\] vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _0945_ _1038_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold641 sound2.divisor_m\[7\] vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__dlygate4sd3_1
X_7288_ _3454_ _3452_ _3460_ _0563_ _2005_ vssd1 vssd1 vccd1 vccd1 _3462_ sky130_fd_sc_hd__a311o_1
Xhold674 sound3.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 sound1.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ _2289_ _2737_ _2738_ _2290_ sound4.sdiv.Q\[7\] vssd1 vssd1 vccd1 vccd1 _2739_
+ sky130_fd_sc_hd__a32o_1
Xhold696 sound2.divisor_m\[5\] vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlygate4sd3_1
X_6239_ _2668_ _2671_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__xnor2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3940_ _0603_ _0595_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__or3b_2
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3871_ _0513_ _0531_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__nor2_1
X_6590_ sound1.divisor_m\[7\] _2948_ vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5610_ sound4.sdiv.A\[6\] _2092_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__or2_1
X_5541_ net651 _2024_ pm.count\[8\] vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8260_ clknet_leaf_34_hwclk net210 net91 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7211_ net945 _1583_ _3142_ vssd1 vssd1 vccd1 vccd1 _3407_ sky130_fd_sc_hd__mux2_1
X_5472_ _1972_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
X_8191_ clknet_leaf_28_hwclk _0312_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4423_ _0949_ _0909_ _0918_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nand3_4
XFILLER_0_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4354_ seq.player_1.state\[2\] _0871_ _0873_ _0924_ vssd1 vssd1 vccd1 vccd1 _0925_
+ sky130_fd_sc_hd__a22o_1
X_7142_ net868 _3327_ _3177_ vssd1 vssd1 vccd1 vccd1 _3385_ sky130_fd_sc_hd__o21ai_1
X_7073_ sound2.sdiv.A\[18\] _3329_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__nor2_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _0859_ _0813_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__and3b_1
X_6024_ sound2.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__inv_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7975_ clknet_leaf_24_hwclk _0138_ net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _3193_ _3196_ vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6857_ _1368_ vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__inv_2
X_5808_ wave_comb.u1.A\[8\] _2224_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__nand2_1
X_6788_ net153 _2893_ _0867_ net296 _2845_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__a221o_1
Xfanout79 net82 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout68 net69 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_6
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5739_ sound4.sdiv.Q\[21\] _2182_ _2185_ net121 _2200_ vssd1 vssd1 vccd1 vccd1 _0021_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7409_ sound3.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _3570_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold471 sound1.sdiv.A\[22\] vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 sound4.sdiv.Q\[7\] vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 sound1.sdiv.Q\[3\] vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 sound4.sdiv.C\[2\] vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4070_ _0703_ _0706_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__nor2_1
XFILLER_0_92_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7760_ clknet_leaf_51_hwclk wave_comb.u1.next_start net101 vssd1 vssd1 vccd1 vccd1
+ wave_comb.u1.start sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _1517_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6711_ sound1.sdiv.A\[19\] _3055_ vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7691_ _3681_ _2179_ _3742_ _2184_ net717 vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ _0581_ _0583_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6642_ sound1.divisor_m\[13\] _3003_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3854_ _0515_ _0518_ _0521_ _0523_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__o41a_1
XFILLER_0_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6573_ _2940_ _2941_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__nand2_1
X_8312_ clknet_leaf_70_hwclk _0412_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3785_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__inv_2
X_5524_ _2007_ pm.current_waveform\[6\] vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8243_ clknet_leaf_46_hwclk _0343_ net100 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5455_ sound4.count\[7\] _1955_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__nand2_1
X_8174_ clknet_leaf_30_hwclk _0295_ net91 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4406_ _0678_ _0964_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__nand2_8
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7125_ _1311_ _3167_ net770 vssd1 vssd1 vccd1 vccd1 _3374_ sky130_fd_sc_hd__mux2_1
X_5386_ _1892_ _1893_ _1896_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__and3_2
X_4337_ seq.player_1.state\[1\] _0871_ _0873_ _0907_ vssd1 vssd1 vccd1 vccd1 _0908_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7056_ _3313_ _3314_ vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__nor2_1
X_4268_ _0847_ _0813_ _0848_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__and3b_1
X_6007_ sound2.divisor_m\[11\] vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__inv_2
X_4199_ seq.tempo_select.state\[1\] _0791_ _0792_ seq.clk_div.count\[12\] vssd1 vssd1
+ vccd1 vccd1 _0793_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ clknet_leaf_21_hwclk _0121_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7889_ clknet_leaf_3_hwclk seq.encode.next_sequencer_on net71 vssd1 vssd1 vccd1 vccd1
+ select1.sequencer_on sky130_fd_sc_hd__dfrtp_4
X_6909_ _3164_ _3181_ _3182_ _3174_ net255 vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold290 sound2.count\[16\] vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ net367 _1753_ _1721_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5171_ _1004_ _1038_ _1553_ _1580_ _1166_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__o32a_1
X_4122_ seq.player_5.state\[0\] _0737_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__and2_1
X_4053_ _0674_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__buf_12
Xinput3 piano_keys[0] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7812_ clknet_leaf_100_hwclk seq.player_6.next_state\[2\] net64 vssd1 vssd1 vccd1
+ vccd1 seq.player_6.state\[2\] sky130_fd_sc_hd__dfrtp_2
X_7743_ clknet_leaf_55_hwclk net522 net95 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4955_ sound2.count\[0\] sound2.count\[1\] vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3906_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__buf_12
X_7674_ _2040_ _3730_ vssd1 vssd1 vccd1 vccd1 _3731_ sky130_fd_sc_hd__xor2_1
X_4886_ _1129_ _1347_ _1345_ _1140_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6625_ _2987_ _2988_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__or2_1
X_3837_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6556_ net470 _2895_ sound1.sdiv.next_dived _2926_ vssd1 vssd1 vccd1 vccd1 _0112_
+ sky130_fd_sc_hd__a22o_1
X_3768_ inputcont.INTERNAL_SYNCED_I\[8\] _0448_ _0451_ vssd1 vssd1 vccd1 vccd1 _0452_
+ sky130_fd_sc_hd__a21oi_1
X_5507_ _1779_ _1998_ _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6487_ net740 _2872_ _2864_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__mux2_1
X_8226_ clknet_leaf_11_hwclk sound3.osc.next_count\[7\] net88 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_5438_ sound4.count\[3\] _1940_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__or2_1
X_8157_ clknet_leaf_31_hwclk _0278_ net90 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_5369_ _1064_ _1781_ _1878_ _1879_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8088_ clknet_leaf_76_hwclk _0230_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_7108_ _3358_ _3359_ vssd1 vssd1 vccd1 vccd1 _3360_ sky130_fd_sc_hd__nand2_1
X_7039_ sound2.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4740_ sound1.count\[12\] net957 _1287_ sound1.count\[14\] vssd1 vssd1 vccd1 vccd1
+ _1297_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4671_ _1012_ _1028_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7390_ _3448_ _3552_ vssd1 vssd1 vccd1 vccd1 _3553_ sky130_fd_sc_hd__and2_1
X_6410_ net651 _2827_ _2808_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6341_ _2289_ _2769_ _2770_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6272_ sound4.sdiv.Q\[4\] _2641_ _2673_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5223_ net349 _1741_ _1743_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[10\] sky130_fd_sc_hd__a21oi_1
X_8011_ clknet_leaf_13_hwclk net189 net86 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_5154_ _1151_ _1562_ _1574_ _1042_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__o22a_1
X_4105_ net780 _0724_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__xor2_1
X_5085_ sound3.count\[15\] _1615_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4036_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__clkinv_8
XFILLER_0_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ sound1.count_m\[10\] _2378_ _2390_ _2391_ _2379_ vssd1 vssd1 vccd1 vccd1 _2423_
+ sky130_fd_sc_hd__a221o_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7726_ clknet_leaf_63_hwclk _0011_ net78 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4938_ _1077_ _1323_ _1339_ _1193_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4869_ _0964_ _1418_ _1419_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__or3b_1
X_7657_ _2145_ _2150_ _3715_ _2147_ vssd1 vssd1 vccd1 vccd1 _3719_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6608_ net432 vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7588_ _3672_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__clkbuf_1
X_6539_ sound1.divisor_m\[2\] sound1.divisor_m\[1\] sound1.divisor_m\[0\] _2903_ vssd1
+ vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8209_ clknet_leaf_47_hwclk _0330_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5910_ sound4.divisor_m\[1\] vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__inv_2
X_6890_ sound2.divisor_m\[0\] sound2.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3166_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5841_ _2278_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5772_ _2223_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__buf_4
X_7511_ sound3.sdiv.Q\[1\] _3463_ sound3.sdiv.next_dived net280 vssd1 vssd1 vccd1
+ vccd1 _0340_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4723_ net956 _1281_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7442_ sound3.sdiv.A\[19\] _3595_ vssd1 vssd1 vccd1 vccd1 _3599_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4654_ _0988_ _0955_ _0971_ _1069_ _1018_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7373_ _3534_ _3536_ vssd1 vssd1 vccd1 vccd1 _3538_ sky130_fd_sc_hd__nand2_1
X_4585_ _0967_ _1095_ _1042_ _0976_ _1155_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold801 sound2.count\[9\] vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 seq.player_3.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__dlygate4sd3_1
X_6324_ sound1.sdiv.Q\[8\] _2293_ _2752_ _2753_ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__o2bb2a_1
Xhold834 sound1.count\[7\] vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 sound4.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 sound2.count\[14\] vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 sound3.sdiv.A\[23\] vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 sound3.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ sound2.sdiv.Q\[5\] _0578_ _2686_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__a21o_1
Xhold856 sound4.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
X_5206_ sound3.count\[4\] sound3.count\[5\] _1728_ vssd1 vssd1 vccd1 vccd1 _1732_
+ sky130_fd_sc_hd__and3_1
X_6186_ sound1.sdiv.Q\[4\] _0579_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5137_ _0978_ _0944_ _1565_ _1572_ _0997_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__o32a_1
X_5068_ _1123_ _1559_ _1565_ _1127_ _1591_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4019_ _0587_ _0597_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7709_ net761 net31 _0645_ vssd1 vssd1 vccd1 vccd1 _3754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 sound3.count_m\[15\] vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold119 _0009_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ _0937_ _0909_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__or2b_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _2474_ sound2.divisor_m\[4\] _2475_ sound2.divisor_m\[3\] vssd1 vssd1 vccd1
+ vccd1 _2476_ sky130_fd_sc_hd__a22o_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7991_ clknet_leaf_16_hwclk sound1.osc.next_count\[12\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6942_ sound2.divisor_m\[5\] sound2.divisor_m\[4\] _3194_ vssd1 vssd1 vccd1 vccd1
+ _3212_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6873_ net797 _3155_ _3142_ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__mux2_1
X_5824_ wave_comb.u1.C\[0\] wave_comb.u1.C\[1\] net614 vssd1 vssd1 vccd1 vccd1 _2266_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5755_ wave_comb.u1.A\[10\] vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4706_ _1271_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
X_5686_ _2042_ _2044_ _2045_ _2168_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__or4b_2
XFILLER_0_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7425_ _3583_ _3584_ vssd1 vssd1 vccd1 vccd1 _3585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4637_ _0981_ _1198_ _0992_ _1199_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold620 sound2.count\[8\] vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7356_ _3520_ _3522_ vssd1 vssd1 vccd1 vccd1 _3523_ sky130_fd_sc_hd__nand2_1
Xhold642 sound3.divisor_m\[12\] vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold631 wave_comb.u1.M\[1\] vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 sound1.divisor_m\[13\] vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _0959_ _1028_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7287_ _3454_ _3452_ _3460_ vssd1 vssd1 vccd1 vccd1 _3461_ sky130_fd_sc_hd__a21oi_1
Xhold675 sound1.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
X_6307_ sound4.sdiv.Q\[6\] _2736_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__nand2_1
X_4499_ _0988_ _0955_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__a21o_4
Xhold697 sound4.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 seq.player_6.state\[3\] vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 sound4.divisor_m\[12\] vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
X_6238_ sound3.sdiv.Q\[5\] _2301_ _2670_ _2292_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__o2bb2a_1
X_6169_ sound3.sdiv.Q\[2\] _2602_ _2292_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__a21o_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3870_ _0542_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__inv_2
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5540_ _0657_ pm.current_waveform\[7\] _2023_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5471_ _1779_ _1936_ _1970_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7210_ net170 _3403_ _3406_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a21o_1
X_4422_ _0674_ _0680_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nor2_4
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8190_ clknet_leaf_43_hwclk _0311_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_4353_ seq.player_2.state\[2\] _0876_ _0878_ _0923_ vssd1 vssd1 vccd1 vccd1 _0924_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7141_ _3384_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
X_4284_ _0791_ _0858_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__nand2_1
X_7072_ _3328_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__buf_4
X_6023_ _2442_ _2445_ _2453_ _2458_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__and4bb_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7974_ clknet_leaf_24_hwclk _0137_ net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6925_ _3193_ _3196_ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6856_ _3144_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
X_3999_ pm.count\[6\] _0652_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5807_ net561 _0573_ wave_comb.u1.next_dived _2253_ vssd1 vssd1 vccd1 vccd1 _0036_
+ sky130_fd_sc_hd__a22o_1
X_6787_ sound1.sdiv.Q\[14\] _2893_ _0867_ net253 _2844_ vssd1 vssd1 vccd1 vccd1 _0155_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout69 net2 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_4
X_5738_ sound4.count\[13\] _2186_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5669_ _2057_ _2061_ _2141_ _2148_ _2151_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__a41o_1
XFILLER_0_130_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7408_ _3564_ _3568_ vssd1 vssd1 vccd1 vccd1 _3569_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold472 sound3.sdiv.A\[22\] vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__dlygate4sd3_1
X_7339_ _3437_ _3506_ _3507_ _3440_ net235 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a32o_1
Xhold461 seq.player_1.state\[3\] vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 seq.player_8.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 sound2.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _0434_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4971_ _1515_ _1516_ _1504_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__and3b_1
X_6710_ _3022_ _3026_ _3033_ _3042_ _3064_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__a2111o_1
X_7690_ _2178_ _2175_ _2176_ vssd1 vssd1 vccd1 vccd1 _3742_ sky130_fd_sc_hd__nand3_1
X_3922_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6641_ _2903_ _3002_ vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3853_ _0514_ _0525_ _0526_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__and3b_1
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6572_ _2936_ _2939_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__nand2_1
X_8311_ clknet_leaf_66_hwclk _0411_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3784_ inputcont.INTERNAL_SYNCED_I\[6\] _0443_ _0463_ inputcont.INTERNAL_SYNCED_I\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__or4b_1
XFILLER_0_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5523_ pm.count\[6\] vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8242_ clknet_leaf_47_hwclk net644 net101 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5454_ _1958_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_8173_ clknet_leaf_30_hwclk _0294_ net91 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4405_ _0975_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__clkbuf_4
X_5385_ _0960_ _1777_ _1894_ _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__o211a_1
X_4336_ seq.player_2.state\[1\] _0876_ _0878_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7124_ _3349_ _3371_ _3373_ _3174_ net713 vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__a32o_1
X_7055_ sound2.sdiv.A\[16\] _3311_ vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__nor2_1
X_4267_ seq.clk_div.count\[15\] _0844_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__or2_1
X_6006_ sound2.count_m\[14\] _2440_ sound2.count_m\[13\] _2441_ vssd1 vssd1 vccd1
+ vccd1 _2442_ sky130_fd_sc_hd__a22o_1
X_4198_ seq.tempo_select.state\[1\] seq.clk_div.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0792_ sky130_fd_sc_hd__nand2_1
X_7957_ clknet_leaf_21_hwclk _0120_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7888_ clknet_leaf_96_hwclk tempo_select_on net68 vssd1 vssd1 vccd1 vccd1 seq.encode.inter_keys\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_6908_ _3175_ _3172_ _3180_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__nand3_1
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6839_ net163 _3132_ _3134_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold280 sound1.count_m\[13\] vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 sound4.count_m\[7\] vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5170_ _0685_ _1562_ _1572_ _1126_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__o221a_1
X_4121_ _0612_ seq.encode.keys_edge_det\[6\] vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__nor2_1
X_4052_ _0676_ _0675_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__nor2_2
Xinput4 piano_keys[10] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
X_7811_ clknet_leaf_100_hwclk net612 net64 vssd1 vssd1 vccd1 vccd1 seq.player_6.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_7742_ clknet_leaf_58_hwclk net181 net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_4954_ net422 _1504_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3905_ rate_clk.count\[6\] rate_clk.count\[7\] _0552_ vssd1 vssd1 vccd1 vccd1 _0574_
+ sky130_fd_sc_hd__and3_1
X_7673_ sound4.sdiv.A\[19\] _2038_ _3728_ vssd1 vssd1 vccd1 vccd1 _3730_ sky130_fd_sc_hd__a21oi_1
X_4885_ _1135_ _1321_ _1333_ _1127_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6624_ _2983_ _2986_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__and2_1
X_3836_ _0471_ _0487_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__nand2_1
X_6555_ _2924_ _2925_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3767_ _0449_ inputcont.INTERNAL_SYNCED_I\[2\] inputcont.INTERNAL_SYNCED_I\[4\] _0450_
+ inputcont.INTERNAL_SYNCED_I\[0\] vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_6__f_hwclk clknet_0_hwclk vssd1 vssd1 vccd1 vccd1 clknet_3_6__leaf_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5506_ sound4.count\[16\] sound4.count\[17\] sound4.count\[18\] _1988_ vssd1 vssd1
+ vccd1 vccd1 _1999_ sky130_fd_sc_hd__nand4_1
X_8225_ clknet_leaf_35_hwclk sound3.osc.next_count\[6\] net87 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[6\] sky130_fd_sc_hd__dfrtp_2
X_6486_ _1170_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5437_ _1944_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__inv_2
X_8156_ clknet_leaf_31_hwclk net502 net90 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_5368_ _0677_ _1038_ _1796_ _1769_ _1059_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__o32a_1
X_5299_ _0954_ _1781_ _1805_ _1809_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__o211ai_4
X_8087_ clknet_leaf_77_hwclk _0229_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_7107_ sound2.sdiv.A\[23\] _3329_ vssd1 vssd1 vccd1 vccd1 _3359_ sky130_fd_sc_hd__nand2_1
X_4319_ select1.sequencer_on _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__and2_1
X_7038_ _3164_ _3297_ _3298_ _3174_ net308 vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4670_ _0969_ _1101_ _1240_ _0943_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6340_ _2569_ _2753_ sound3.sdiv.Q\[8\] _2301_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6271_ _2698_ _2702_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5222_ net349 _1741_ _1721_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__o21ai_1
X_8010_ clknet_leaf_10_hwclk net208 net85 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_5153_ _1095_ _1559_ _1553_ _1127_ _1591_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__o221a_1
X_4104_ net848 seq.player_7.state\[3\] vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__nand2_1
X_5084_ _1610_ _1612_ _1614_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__and3_2
XFILLER_0_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4035_ _0675_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__nor2_4
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5986_ _2408_ _2411_ _2412_ _2421_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__nor4_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7725_ clknet_leaf_63_hwclk net463 net78 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _1001_ _1480_ _1482_ _1487_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__o211a_2
X_7656_ net468 _2183_ sound4.sdiv.next_dived _3718_ vssd1 vssd1 vccd1 vccd1 _0420_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4868_ _0695_ _0499_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__or2_1
X_6607_ _2966_ _2964_ _2971_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3819_ _0492_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__or2_1
X_7587_ net790 _1924_ _2186_ vssd1 vssd1 vccd1 vccd1 _3672_ sky130_fd_sc_hd__mux2_1
X_4799_ _1014_ _1338_ _1339_ _0688_ _1349_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__o221a_1
X_6538_ sound1.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__inv_2
X_6469_ _2861_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8208_ clknet_leaf_48_hwclk _0329_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8139_ clknet_leaf_92_hwclk _0260_ net67 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5840_ wave.mode\[0\] net1 wave.mode\[1\] vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__or3b_1
XFILLER_0_76_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5771_ wave_comb.u1.M\[0\] wave_comb.u1.M\[1\] wave_comb.u1.M\[2\] _2209_ vssd1 vssd1
+ vccd1 vccd1 _2223_ sky130_fd_sc_hd__o31a_1
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7510_ _2275_ _3653_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4722_ _1283_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7441_ net647 _3463_ sound3.sdiv.next_dived _3598_ vssd1 vssd1 vccd1 vccd1 _0325_
+ sky130_fd_sc_hd__a22o_1
X_4653_ sound1.count\[18\] _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7372_ _3534_ _3536_ vssd1 vssd1 vccd1 vccd1 _3537_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4584_ _0950_ _1125_ _1154_ _1000_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold802 seq.player_4.state\[2\] vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__dlygate4sd3_1
X_6323_ net1 wave.mode\[1\] wave.mode\[0\] vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__or3b_2
Xhold824 sound3.count\[14\] vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 seq.clk_div.count\[6\] vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold846 sound2.sdiv.A\[24\] vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 sound2.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6254_ sound2.sdiv.Q\[4\] _2660_ _2661_ vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__a21bo_1
Xhold879 sound1.count\[16\] vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold857 sound2.sdiv.A\[19\] vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold868 seq.clk_div.count\[16\] vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
X_5205_ net479 _1728_ _1731_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[4\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6185_ _2617_ _2599_ _2618_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5136_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__inv_2
X_5067_ _1134_ _1578_ _1553_ _1139_ _1597_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4018_ _0662_ _0666_ vssd1 vssd1 vccd1 vccd1 seq.tempo_select.next_state\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5969_ sound1.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7708_ _3753_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7639_ _1763_ _3705_ _3706_ sound4.sdiv.next_start _2070_ vssd1 vssd1 vccd1 vccd1
+ _0415_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold109 _0283_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7990_ clknet_leaf_16_hwclk sound1.osc.next_count\[11\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[11\] sky130_fd_sc_hd__dfrtp_2
X_6941_ net977 vssd1 vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6872_ _1360_ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5823_ _0646_ _2264_ _2265_ _0573_ net588 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5754_ wave_comb.u1.next_dived _2207_ _2208_ _0573_ net521 vssd1 vssd1 vccd1 vccd1
+ _0028_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4705_ _1269_ _1270_ _1256_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__and3b_1
X_5685_ sound4.sdiv.A\[18\] _2038_ _2158_ _2166_ _2167_ vssd1 vssd1 vccd1 vccd1 _2168_
+ sky130_fd_sc_hd__a221o_1
X_7424_ _3569_ _3575_ _3573_ vssd1 vssd1 vccd1 vccd1 _3584_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_114_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4636_ _0958_ _1027_ _1203_ _1206_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7355_ _3503_ _3507_ _3521_ _3511_ vssd1 vssd1 vccd1 vccd1 _3522_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold610 sound1.sdiv.C\[3\] vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold621 seq.player_4.state\[1\] vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 sound3.divisor_m\[13\] vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ sound4.sdiv.Q\[6\] _0576_ _2736_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__a21o_1
X_4567_ _0685_ _0678_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__nand2_4
Xhold654 sound4.divisor_m\[7\] vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold632 seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
X_7286_ _3458_ _3459_ vssd1 vssd1 vccd1 vccd1 _3460_ sky130_fd_sc_hd__or2_1
X_4498_ _0949_ _0937_ _0974_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__nand3b_1
Xhold665 sound4.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 seq.player_7.state\[2\] vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 sound2.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6237_ _2636_ _2669_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__xor2_1
Xhold698 sound3.count\[10\] vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__dlygate4sd3_1
X_6168_ sound3.sdiv.Q\[2\] _0577_ _2602_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__a21oi_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _1010_ _1567_ _1574_ _1027_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__o22a_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ sound3.divisor_m\[11\] sound3.count_m\[10\] vssd1 vssd1 vccd1 vccd1 _2535_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5470_ sound4.count\[10\] _1966_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4421_ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7140_ net733 _0554_ vssd1 vssd1 vccd1 vccd1 _3384_ sky130_fd_sc_hd__and2_1
X_4352_ seq.player_3.state\[2\] _0881_ _0883_ _0922_ vssd1 vssd1 vccd1 vccd1 _0923_
+ sky130_fd_sc_hd__a22o_1
X_4283_ _0791_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__nor2_1
X_7071_ sound2.sdiv.A\[26\] _3327_ vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6022_ _2454_ _2455_ _2456_ _2457_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__and4b_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7973_ clknet_leaf_24_hwclk net591 net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ _2484_ _3195_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6855_ net799 _1378_ _3142_ vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3998_ _0652_ net509 vssd1 vssd1 vccd1 vccd1 pm.next_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_107_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5806_ _2249_ _2252_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__xnor2_1
X_6786_ net253 _2893_ _2890_ net291 _2842_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5737_ net121 _2182_ _2185_ net318 _2199_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7407_ _3437_ _3567_ _3568_ _3440_ net267 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5668_ _2145_ _2150_ _2147_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4619_ _0950_ _1004_ _1189_ _0969_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5599_ _2081_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__inv_2
X_7338_ _3495_ _3499_ _3505_ vssd1 vssd1 vccd1 vccd1 _3507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold440 _0072_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 sound4.sdiv.A\[24\] vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 seq.player_1.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7269_ sound3.divisor_m\[0\] sound3.sdiv.Q\[27\] _3443_ vssd1 vssd1 vccd1 vccd1 _3445_
+ sky130_fd_sc_hd__a21o_1
Xhold495 sound3.sdiv.C\[2\] vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 wave_comb.u1.C\[1\] vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 wave_comb.u1.A\[9\] vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ net984 sound2.count\[4\] _1508_ sound2.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _1516_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3921_ _0581_ _0583_ _0584_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__and4b_1
X_6640_ sound1.divisor_m\[12\] sound1.divisor_m\[11\] _2984_ vssd1 vssd1 vccd1 vccd1
+ _3002_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3852_ _0478_ _0485_ _0479_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6571_ _2936_ _2939_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__or2_1
X_8310_ clknet_leaf_68_hwclk _0410_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5522_ _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[7\] sky130_fd_sc_hd__nor2_1
X_3783_ inputcont.INTERNAL_SYNCED_I\[3\] _0460_ _0462_ _0464_ vssd1 vssd1 vccd1 vccd1
+ net36 sky130_fd_sc_hd__a211o_1
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8241_ clknet_leaf_47_hwclk _0341_ net101 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5453_ _1779_ _1936_ _1956_ _1957_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__and4_1
X_8172_ clknet_leaf_35_hwclk _0293_ net87 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_4404_ _0918_ _0974_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__or2_1
X_5384_ _1015_ _1769_ _1784_ _1083_ _1833_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7123_ _3359_ _3367_ _3372_ _3370_ vssd1 vssd1 vccd1 vccd1 _3373_ sky130_fd_sc_hd__a31o_1
X_4335_ seq.player_3.state\[1\] _0881_ _0883_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_
+ sky130_fd_sc_hd__a22o_1
X_4266_ seq.clk_div.count\[14\] seq.clk_div.count\[15\] _0841_ vssd1 vssd1 vccd1 vccd1
+ _0847_ sky130_fd_sc_hd__and3_1
X_7054_ _3312_ vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__inv_2
X_6005_ sound2.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__inv_2
X_4197_ net970 vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7956_ clknet_leaf_21_hwclk _0119_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7887_ clknet_leaf_49_hwclk net15 net102 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_6907_ _3175_ _3172_ _3180_ vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6838_ net926 _2855_ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6769_ net730 _2843_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 _0173_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _0083_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _0374_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_67_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4120_ _0734_ _0733_ _0736_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_6.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_4051_ _0693_ vssd1 vssd1 vccd1 vccd1 oct.next_state\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 piano_keys[11] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7810_ clknet_leaf_0_hwclk net162 net64 vssd1 vssd1 vccd1 vccd1 seq.player_6.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7741_ clknet_leaf_58_hwclk _0026_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4953_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__buf_4
X_3904_ _0573_ vssd1 vssd1 vccd1 vccd1 wave_comb.u1.next_start sky130_fd_sc_hd__inv_2
XFILLER_0_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7672_ net662 _2183_ _3681_ _3729_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__a22o_1
X_6623_ _2983_ _2986_ vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__nor2_1
X_4884_ _1134_ _1338_ _1322_ _1041_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3835_ _0509_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_4
X_6554_ _2909_ _2915_ _2913_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__o21ai_1
X_3766_ _0443_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
X_6485_ _2871_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
X_5505_ sound4.count\[16\] sound4.count\[17\] _1988_ sound4.count\[18\] vssd1 vssd1
+ vccd1 vccd1 _1998_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8224_ clknet_leaf_35_hwclk sound3.osc.next_count\[5\] net87 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5436_ sound4.count\[3\] _1940_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8155_ clknet_leaf_31_hwclk net413 net90 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_5367_ _0959_ _1133_ _1786_ _1790_ _0983_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__o32a_1
X_5298_ _0996_ _1784_ _1806_ _1808_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__o211a_1
X_8086_ clknet_leaf_78_hwclk _0228_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_7106_ sound2.sdiv.A\[23\] _3329_ vssd1 vssd1 vccd1 vccd1 _3358_ sky130_fd_sc_hd__or2_1
X_4318_ seq.beat\[3\] seq.encode.play _0870_ inputcont.INTERNAL_SYNCED_I\[4\] vssd1
+ vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__a31o_1
X_7037_ _3286_ _3290_ _3296_ vssd1 vssd1 vccd1 vccd1 _3298_ sky130_fd_sc_hd__a21o_1
X_4249_ _0834_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ clknet_leaf_17_hwclk _0102_ net83 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6270_ _2289_ _2700_ _2701_ _2301_ sound3.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 _2702_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5221_ _1741_ _1742_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[9\] sky130_fd_sc_hd__nor2_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5152_ sound3.count\[12\] _1681_ _1655_ sound3.count\[2\] _1682_ vssd1 vssd1 vccd1
+ vccd1 _1683_ sky130_fd_sc_hd__o221a_1
X_4103_ seq.player_7.state\[2\] net496 _0724_ _0725_ _0700_ vssd1 vssd1 vccd1 vccd1
+ seq.player_7.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_5083_ _1011_ _1559_ _1613_ _1590_ _1591_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4034_ _0676_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__nand2_8
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5985_ sound1.count_m\[2\] _2413_ _2414_ _2418_ _2420_ vssd1 vssd1 vccd1 vccd1 _2421_
+ sky130_fd_sc_hd__a2111o_1
X_7724_ clknet_leaf_63_hwclk net223 net78 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4936_ _1004_ _1483_ _1484_ _1486_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__o211a_1
XANTENNA_10 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4867_ _1314_ _1315_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__or2_1
X_7655_ _3717_ _2148_ vssd1 vssd1 vccd1 vccd1 _3718_ sky130_fd_sc_hd__xor2_1
X_6606_ _2966_ _2964_ _2971_ vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3818_ _0474_ _0491_ _0494_ _0495_ _0496_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__a221o_1
X_7586_ _3671_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6537_ _2901_ _2906_ _2908_ vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4798_ _1199_ _1341_ _1343_ _1200_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__o221a_1
XFILLER_0_120_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6468_ net897 _1008_ _2005_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__mux2_1
X_8207_ clknet_leaf_45_hwclk _0328_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6399_ _2819_ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__inv_2
X_5419_ _0973_ _1786_ _1928_ _1929_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8138_ clknet_leaf_93_hwclk _0259_ net67 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_8069_ clknet_leaf_77_hwclk _0211_ net74 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap56 net34 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_4
XFILLER_0_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _2216_ _2218_ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _1281_ _1282_ _1256_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7440_ _3596_ _3597_ vssd1 vssd1 vccd1 vccd1 _3598_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4652_ _1222_ _1216_ _1070_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7371_ sound3.divisor_m\[12\] _3535_ vssd1 vssd1 vccd1 vccd1 _3536_ sky130_fd_sc_hd__xnor2_1
X_4583_ _1018_ _0978_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__or2_4
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold803 seq.player_4.next_state\[3\] vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 sound3.count\[2\] vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__dlygate4sd3_1
X_6322_ _2407_ _2432_ _2412_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__a21oi_2
Xhold825 seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 seq.player_6.state\[2\] vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6253_ sound2.sdiv.Q\[6\] _2295_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__nand2_1
Xhold847 sound1.count\[4\] vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 sound2.count\[8\] vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
X_5204_ net479 _1728_ _1721_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__o21ai_1
X_6184_ _2590_ _2595_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__nand2_1
X_5135_ _1591_ _1660_ _1665_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5066_ _1129_ _1572_ _1574_ _1141_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__o221a_1
X_4017_ net847 _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__nand2_1
X_5968_ _2397_ _2400_ _2401_ _2403_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7707_ net739 _0554_ vssd1 vssd1 vccd1 vccd1 _3753_ sky130_fd_sc_hd__and2_1
X_4919_ net903 vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5899_ _2333_ sound4.divisor_m\[10\] sound4.divisor_m\[9\] _2334_ vssd1 vssd1 vccd1
+ vccd1 _2335_ sky130_fd_sc_hd__a22o_1
X_7638_ _2079_ _2137_ vssd1 vssd1 vccd1 vccd1 _3706_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7569_ _3661_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6940_ _3164_ _3209_ _3210_ _3174_ net299 vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6871_ _3154_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
X_5822_ wave_comb.u1.C\[0\] wave_comb.u1.C\[1\] vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5753_ wave_comb.u1.M\[0\] wave_comb.u1.Q\[11\] vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4704_ sound1.count\[4\] _1263_ net863 vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5684_ sound4.sdiv.A\[18\] _2038_ _2162_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__o21a_1
X_7423_ _3581_ _3582_ vssd1 vssd1 vccd1 vccd1 _3583_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4635_ _0688_ _0967_ _0969_ _1204_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7354_ _3510_ vssd1 vssd1 vccd1 vccd1 _3521_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold600 sound4.sdiv.C\[3\] vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _0696_ _0939_ _1003_ _1041_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold611 sound2.count\[6\] vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold633 sound1.divisor_m\[12\] vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 wave_comb.u1.M\[2\] vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ sound4.sdiv.Q\[5\] _2641_ _2704_ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold622 seq.player_7.state\[1\] vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlygate4sd3_1
X_7285_ _3455_ _3457_ vssd1 vssd1 vccd1 vccd1 _3459_ sky130_fd_sc_hd__and2_1
Xhold677 sound3.divisor_m\[6\] vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _0677_ _0976_ _1038_ _1054_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__o311a_1
Xhold688 seq.player_1.state\[2\] vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 sound2.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 sound2.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
X_6236_ sound3.sdiv.Q\[3\] _2632_ _2633_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__a21o_1
Xhold699 sound3.count\[4\] vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__dlygate4sd3_1
X_6167_ _2570_ _2601_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__nor2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5118_ _1643_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nand2_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ sound3.divisor_m\[10\] sound3.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2534_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4420_ _0988_ _0937_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4351_ seq.player_4.state\[2\] _0886_ _0888_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4282_ net677 _0855_ net856 _0813_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[19\]
+ sky130_fd_sc_hd__o211a_1
X_7070_ _3308_ _2471_ _2470_ vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__and3b_1
X_6021_ sound2.divisor_m\[9\] sound2.count_m\[8\] vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__or2b_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7972_ clknet_leaf_24_hwclk _0135_ net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6923_ _3177_ _3194_ vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__nand2_1
X_6854_ _3143_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3997_ pm.count\[4\] _0649_ net508 vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__a21oi_1
X_5805_ _2250_ _2251_ _2240_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__or3b_1
X_6785_ sound1.sdiv.Q\[12\] _2893_ _2890_ net188 _2841_ vssd1 vssd1 vccd1 vccd1 _0153_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5736_ net873 _2186_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5667_ _2149_ _2056_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7406_ _3555_ _3559_ _3566_ vssd1 vssd1 vccd1 vccd1 _3568_ sky130_fd_sc_hd__a21o_1
X_4618_ _1001_ _1040_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nor2_4
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5598_ sound4.divisor_m\[9\] _2080_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__xnor2_1
X_7337_ _3495_ _3499_ _3505_ vssd1 vssd1 vccd1 vccd1 _3506_ sky130_fd_sc_hd__nand3_1
Xhold463 sound3.sdiv.C\[1\] vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkdlybuf4s25_1
X_4549_ _1107_ _1108_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold452 seq.clk_div.count\[2\] vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 inputcont.INTERNAL_SYNCED_I\[6\] vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 seq.encode.keys_edge_det\[0\] vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__dlygate4sd3_1
X_7268_ _3438_ _3443_ vssd1 vssd1 vccd1 vccd1 _3444_ sky130_fd_sc_hd__or2b_1
Xhold485 _0040_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 sound4.sdiv.Q\[5\] vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 sound2.sdiv.C\[2\] vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__dlygate4sd3_1
X_6219_ _2650_ _2652_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__xnor2_1
X_7199_ net341 _3132_ _3400_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__a21o_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _0529_ _0549_ _0582_ _0525_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3851_ _0478_ _0485_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__or2_2
XFILLER_0_128_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6570_ sound1.divisor_m\[6\] _2938_ vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3782_ inputcont.INTERNAL_SYNCED_I\[6\] _0463_ _0450_ vssd1 vssd1 vccd1 vccd1 _0464_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5521_ net722 _0553_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__nor2_1
X_8240_ clknet_leaf_47_hwclk net281 net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5452_ sound4.count\[6\] _1951_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__or2_1
X_8171_ clknet_leaf_30_hwclk _0292_ net91 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_4403_ _0909_ _0936_ _0926_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__or3b_4
X_5383_ _1079_ _1800_ _1794_ _0952_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__o22a_1
X_7122_ _3360_ _3363_ _3366_ vssd1 vssd1 vccd1 vccd1 _3372_ sky130_fd_sc_hd__or3_1
X_4334_ seq.player_4.state\[1\] _0886_ _0888_ _0904_ vssd1 vssd1 vccd1 vccd1 _0905_
+ sky130_fd_sc_hd__a22o_1
X_7053_ sound2.sdiv.A\[16\] _3311_ vssd1 vssd1 vccd1 vccd1 _3312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6004_ sound2.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__inv_2
X_4265_ _0846_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4196_ _0789_ seq.clk_div.count\[14\] seq.tempo_select.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0790_ sky130_fd_sc_hd__a21oi_1
X_7955_ clknet_leaf_19_hwclk _0118_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7886_ clknet_leaf_94_hwclk net14 net66 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6906_ _3176_ _3179_ vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6837_ net477 _3132_ _3133_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6768_ _3111_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6699_ _3054_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5719_ net149 _2182_ _2185_ net328 _2190_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8369_ clknet_leaf_72_hwclk net448 net76 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold271 sound3.sdiv.Q\[17\] vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _0163_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 sound3.sdiv.Q\[21\] vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 sound2.sdiv.Q\[12\] vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4050_ _0679_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__or2_1
Xinput6 piano_keys[12] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_7740_ clknet_leaf_60_hwclk _0025_ net94 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_4952_ _1317_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__and2_1
X_3903_ _0572_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__clkbuf_8
X_7671_ _3727_ _3728_ vssd1 vssd1 vccd1 vccd1 _3729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4883_ _1317_ _1426_ _1431_ _1433_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__and4_2
XFILLER_0_117_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6622_ sound1.divisor_m\[11\] _2985_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__xnor2_1
X_3834_ net1 wave.mode\[1\] vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6553_ _2922_ _2923_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3765_ inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
X_6484_ net756 _1089_ _2864_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__mux2_1
X_5504_ _1997_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
X_8223_ clknet_leaf_35_hwclk sound3.osc.next_count\[4\] net88 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[4\] sky130_fd_sc_hd__dfrtp_2
X_5435_ _1943_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8154_ clknet_leaf_31_hwclk _0275_ net90 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5366_ sound4.count\[13\] _1875_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__or2_1
X_5297_ _1182_ _1794_ _1796_ _1175_ _1807_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__o221a_1
X_8085_ clknet_leaf_75_hwclk _0227_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_7105_ net421 _3168_ sound2.sdiv.next_dived _3357_ vssd1 vssd1 vccd1 vccd1 _0230_
+ sky130_fd_sc_hd__a22o_1
X_4317_ _0886_ _0887_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__nand2_1
X_7036_ _3286_ _3290_ _3296_ vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__nand3_1
X_4248_ _0832_ _0813_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4179_ net829 seq.player_1.state\[2\] _0770_ net565 vssd1 vssd1 vccd1 vccd1 _0776_
+ sky130_fd_sc_hd__a31o_1
X_7938_ clknet_leaf_19_hwclk _0101_ net85 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7869_ clknet_leaf_7_hwclk net105 net72 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5220_ net674 _1738_ _1721_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__o21ai_1
X_5151_ sound3.count\[1\] _1673_ _1666_ sound3.count\[13\] vssd1 vssd1 vccd1 vccd1
+ _1682_ sky130_fd_sc_hd__o2bb2a_1
X_5082_ _1138_ _1551_ _1568_ _0688_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__o22a_1
X_4102_ net900 _0722_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nor2_1
X_4033_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__buf_12
XFILLER_0_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ sound1.count_m\[3\] _2419_ sound1.divisor_m\[1\] _2415_ vssd1 vssd1 vccd1
+ vccd1 _2420_ sky130_fd_sc_hd__a22o_1
X_7723_ clknet_leaf_60_hwclk _0008_ net94 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _0947_ _1325_ _1485_ _1033_ _1341_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__o32a_1
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4866_ _0680_ _1321_ _1415_ _1416_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__o211a_1
X_7654_ _2150_ _3715_ vssd1 vssd1 vccd1 vccd1 _3717_ sky130_fd_sc_hd__nand2_1
X_6605_ _2969_ _2970_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3817_ inputcont.INTERNAL_SYNCED_I\[2\] _0459_ _0481_ vssd1 vssd1 vccd1 vccd1 _0496_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_34_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7585_ net788 _3670_ _2186_ vssd1 vssd1 vccd1 vccd1 _3671_ sky130_fd_sc_hd__mux2_1
X_4797_ _0683_ _1107_ _1345_ _1347_ _1146_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__o32a_1
X_6536_ _2902_ _2905_ vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6467_ _2860_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
X_8206_ clknet_leaf_45_hwclk _0327_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6398_ _2659_ _2682_ _2805_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__mux2_1
X_5418_ _0959_ _0993_ _1800_ _1792_ _0869_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__o32a_1
X_5349_ sound4.count\[0\] _1859_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8137_ clknet_leaf_93_hwclk net339 net67 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_66_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_8068_ clknet_leaf_77_hwclk _0210_ net74 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_7019_ _3164_ _3280_ _3281_ _3174_ net294 vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ sound1.count\[9\] _1278_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4651_ _0685_ net60 vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__nand2_2
Xinput20 tempo_select vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7370_ sound3.divisor_m\[11\] _3526_ _3448_ vssd1 vssd1 vccd1 vccd1 _3535_ sky130_fd_sc_hd__o21a_1
X_4582_ _0939_ _1134_ _1151_ _0981_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold837 wave_comb.u1.A\[5\] vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__dlygate4sd3_1
X_6321_ _2749_ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__xor2_1
Xhold804 sound4.count\[17\] vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 inputcont.u2.next_in vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold815 _0734_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold848 sound3.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__dlygate4sd3_1
X_6252_ _2678_ _2679_ _2683_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__o21ai_1
Xhold859 sound4.sdiv.Q\[0\] vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6183_ _2590_ _2595_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__nor2_1
X_5203_ _1730_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5134_ _0952_ _1025_ _1559_ _1661_ _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__o311a_1
X_5065_ _1138_ _1562_ _1567_ _0696_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__o22a_1
X_4016_ seq.tempo_select.state\[1\] seq.tempo_select.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _0665_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5967_ sound1.divisor_m\[5\] _2399_ _2402_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7706_ _3752_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4918_ _1466_ _1468_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5898_ sound4.count_m\[8\] vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__inv_2
X_7637_ _2079_ _2137_ vssd1 vssd1 vccd1 vccd1 _3705_ sky130_fd_sc_hd__nor2_1
X_4849_ _0985_ _1323_ _1338_ _0948_ _1399_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__o221a_1
X_7568_ net924 _1866_ _3419_ vssd1 vssd1 vccd1 vccd1 _3661_ sky130_fd_sc_hd__mux2_1
X_7499_ _3643_ _3644_ _3646_ _3440_ net599 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__a32o_1
X_6519_ _2893_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__buf_6
XFILLER_0_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6870_ net742 _3153_ _3142_ vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__mux2_1
X_5821_ wave_comb.u1.C\[0\] net588 vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__nand2_1
X_5752_ wave_comb.u1.M\[0\] wave_comb.u1.Q\[11\] vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ sound1.count\[4\] sound1.count\[5\] _1263_ vssd1 vssd1 vccd1 vccd1 _1269_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_57_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5683_ _2164_ _2165_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7422_ _3577_ _3580_ vssd1 vssd1 vccd1 vccd1 _3582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4634_ _0683_ _1107_ _1000_ _0943_ _1014_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__o32a_1
XFILLER_0_71_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7353_ _3518_ _3519_ vssd1 vssd1 vccd1 vccd1 _3520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4565_ _0943_ _1134_ _1135_ _0950_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold612 seq.beat\[3\] vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold601 sound2.sdiv.C\[3\] vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold645 sound3.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _2730_ _2734_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__xor2_1
Xhold634 sound2.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 seq.player_8.state\[1\] vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__dlygate4sd3_1
X_7284_ _3455_ _3457_ vssd1 vssd1 vccd1 vccd1 _3458_ sky130_fd_sc_hd__nor2_1
Xhold678 sound1.divisor_m\[10\] vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4496_ _0990_ _1056_ _1061_ _1066_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__o211a_1
Xhold656 seq.player_6.state\[2\] vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold667 sound4.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 sound3.divisor_m\[10\] vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
X_6235_ _2666_ _2667_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6166_ sound3.sdiv.Q\[0\] sound3.sdiv.Q\[1\] _0577_ vssd1 vssd1 vccd1 vccd1 _2601_
+ sky130_fd_sc_hd__o21ai_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _2531_ sound3.divisor_m\[10\] sound3.divisor_m\[9\] _2532_ vssd1 vssd1 vccd1
+ vccd1 _2533_ sky130_fd_sc_hd__a22o_1
X_5117_ _0971_ _1578_ _1645_ _1647_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__o211a_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5048_ _1551_ _1563_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6999_ _3262_ _3263_ vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4350_ seq.player_5.state\[2\] _0890_ _0892_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4281_ net855 seq.clk_div.count\[19\] _0853_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__nand3_1
X_6020_ sound2.count_m\[9\] sound2.divisor_m\[10\] vssd1 vssd1 vccd1 vccd1 _2456_
+ sky130_fd_sc_hd__or2b_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7971_ clknet_leaf_24_hwclk _0134_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6922_ sound2.divisor_m\[3\] sound2.divisor_m\[2\] sound2.divisor_m\[1\] sound2.divisor_m\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3194_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6853_ net800 _3141_ _3142_ vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5804_ wave_comb.u1.A\[6\] wave_comb.u1.A\[5\] _2224_ vssd1 vssd1 vccd1 vccd1 _2251_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3996_ net508 pm.count\[4\] _0649_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__and3_1
X_6784_ net188 _2893_ _2890_ net207 _2840_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5735_ net318 _2182_ _2185_ net242 _2198_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5666_ sound4.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__inv_2
X_7405_ _3555_ _3559_ _3566_ vssd1 vssd1 vccd1 vccd1 _3567_ sky130_fd_sc_hd__nand3_1
X_4617_ _0676_ _1003_ _1083_ _1000_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold420 sound4.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__dlygate4sd3_1
X_5597_ _2036_ _2029_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7336_ _3503_ _3504_ vssd1 vssd1 vccd1 vccd1 _3505_ sky130_fd_sc_hd__nand2_1
Xhold431 pm.count\[1\] vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__dlygate4sd3_1
X_4548_ _0676_ _1003_ _1034_ _1109_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__o311a_1
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold453 seq.clk_div.count\[1\] vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 seq.encode.next_play vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _0334_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__dlygate4sd3_1
X_7267_ sound3.sdiv.A\[0\] _3442_ vssd1 vssd1 vccd1 vccd1 _3443_ sky130_fd_sc_hd__xnor2_1
Xhold475 pm.count\[3\] vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold486 sound1.sdiv.C\[1\] vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _1037_ _1045_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__and3_2
X_6218_ _2610_ _2612_ _2651_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__a21bo_1
Xhold497 _0006_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__dlygate4sd3_1
X_7198_ _1658_ _2843_ vssd1 vssd1 vccd1 vccd1 _3400_ sky130_fd_sc_hd__nor2_1
X_6149_ sound4.sdiv.Q\[2\] _0576_ _2582_ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__a21o_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _0473_ _0486_ _0521_ _0523_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__nor4_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3781_ inputcont.INTERNAL_SYNCED_I\[5\] inputcont.INTERNAL_SYNCED_I\[4\] vssd1 vssd1
+ vccd1 vccd1 _0463_ sky130_fd_sc_hd__or2_2
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5520_ _0575_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__buf_12
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5451_ _1955_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8170_ clknet_leaf_36_hwclk _0291_ net93 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_4402_ _0971_ _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__or2_4
XFILLER_0_10_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5382_ _0684_ _1077_ _1792_ _1781_ _1039_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__o32a_1
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7121_ _3365_ _3366_ _3367_ _3370_ vssd1 vssd1 vccd1 vccd1 _3371_ sky130_fd_sc_hd__o211ai_1
X_4333_ seq.player_5.state\[1\] _0890_ _0892_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_
+ sky130_fd_sc_hd__a22o_1
X_4264_ _0844_ _0813_ _0845_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__and3b_1
X_7052_ _3310_ vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__inv_2
X_6003_ _2289_ _2437_ _2438_ _2293_ sound1.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 _2439_
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4195_ seq.clk_div.count\[2\] vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__inv_2
X_7954_ clknet_leaf_20_hwclk _0117_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6905_ sound2.divisor_m\[2\] _3178_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__xnor2_1
X_7885_ clknet_leaf_99_hwclk net13 net65 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6836_ net840 _2855_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__and2_1
X_6767_ _2843_ _3110_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5718_ net822 _2186_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__and2_1
X_3979_ _0640_ _0641_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__xnor2_2
X_6698_ sound1.divisor_m\[18\] sound1.divisor_m\[17\] _3036_ _2903_ vssd1 vssd1 vccd1
+ vccd1 _3054_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5649_ _2099_ _2131_ _2097_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8368_ clknet_leaf_72_hwclk net131 net76 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7319_ _3477_ _3480_ _3488_ vssd1 vssd1 vccd1 vccd1 _3490_ sky130_fd_sc_hd__a21o_1
Xhold261 wave_comb.u1.A\[1\] vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold250 sound4.count_m\[6\] vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 sound1.sdiv.Q\[19\] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 sound2.count_m\[8\] vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _0253_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__dlygate4sd3_1
X_8299_ clknet_leaf_66_hwclk _0399_ net80 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 piano_keys[13] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_4951_ _1370_ _1414_ _1443_ _1501_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3902_ _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__and2_1
X_7670_ _2041_ _2168_ vssd1 vssd1 vccd1 vccd1 _3728_ sky130_fd_sc_hd__and2b_1
X_4882_ _0952_ _1025_ _1339_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__o31a_1
X_6621_ _2903_ _2984_ vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__and2_1
X_3833_ _0508_ _0477_ _0505_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__a21o_2
XFILLER_0_116_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6552_ _2918_ _2921_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3764_ _0443_ _0444_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6483_ _2870_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
X_5503_ _1779_ _1936_ _1995_ _1996_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8222_ clknet_leaf_35_hwclk sound3.osc.next_count\[3\] net87 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_5434_ _1779_ _1936_ _1941_ _1942_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8153_ clknet_leaf_33_hwclk net270 net90 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7104_ _3355_ _3356_ vssd1 vssd1 vccd1 vccd1 _3357_ sky130_fd_sc_hd__xnor2_1
X_5365_ sound4.count\[13\] _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5296_ _1129_ _1800_ _1792_ _1026_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__o22a_1
X_8084_ clknet_leaf_75_hwclk _0226_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_4316_ seq.player_4.state\[0\] seq.player_4.state\[1\] seq.player_4.state\[2\] seq.player_4.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__or4_1
X_7035_ _3294_ _3295_ vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__nand2_1
X_4247_ seq.clk_div.count\[10\] _0829_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__or2_1
X_4178_ net921 _0773_ _0775_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_1.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7937_ clknet_leaf_19_hwclk _0100_ net84 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ clknet_leaf_4_hwclk net126 net71 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_sync\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6819_ net905 _2855_ vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7799_ clknet_leaf_8_hwclk oct.next_state\[0\] net71 vssd1 vssd1 vccd1 vccd1 oct.state\[0\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_107_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _1675_ _1677_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__and3_1
X_5081_ _1611_ _1565_ _1213_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__a21o_1
X_4101_ seq.player_7.state\[0\] seq.player_7.state\[1\] _0721_ vssd1 vssd1 vccd1 vccd1
+ _0724_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4032_ oct.state\[1\] vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__buf_12
X_5983_ sound1.divisor_m\[4\] vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7722_ clknet_leaf_58_hwclk _0007_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4934_ _0977_ _1419_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4865_ _1347_ _1323_ _0687_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__a21o_1
X_7653_ _3681_ _3715_ _3716_ _2184_ net380 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__a32o_1
XANTENNA_12 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6604_ net943 _2968_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3816_ _0480_ _0481_ _0482_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__and3_1
X_4796_ _1346_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__buf_4
X_7584_ _1909_ vssd1 vssd1 vccd1 vccd1 _3670_ sky130_fd_sc_hd__inv_2
X_6535_ net485 _2895_ sound1.sdiv.next_dived _2907_ vssd1 vssd1 vccd1 vccd1 _0110_
+ sky130_fd_sc_hd__a22o_1
X_8205_ clknet_leaf_45_hwclk _0326_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_6466_ net874 _2859_ _2005_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6397_ _2818_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
X_5417_ _0985_ _1769_ _1796_ _0979_ _1927_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5348_ _1041_ _1769_ _1777_ _1101_ _1858_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__o221ai_4
X_8136_ clknet_leaf_93_hwclk _0257_ net66 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8067_ clknet_leaf_83_hwclk _0209_ net74 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_7018_ _3268_ _3272_ _3279_ vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__nand3_1
X_5279_ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4650_ sound1.count\[15\] _1215_ _1219_ sound1.count\[16\] vssd1 vssd1 vccd1 vccd1
+ _1221_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 piano_keys[2] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6320_ sound1.sdiv.Q\[7\] _0579_ vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__nand2_1
X_4581_ _1107_ _1003_ net59 vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold816 seq.player_1.state\[3\] vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 seq.encode.keys_edge_det\[2\] vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold805 seq.player_4.state\[1\] vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 sound1.sdiv.C\[4\] vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _2676_ _2677_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__or2b_1
Xhold838 sound2.sdiv.C\[4\] vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__dlygate4sd3_1
X_6182_ wave_comb.u1.next_start _2615_ _2616_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__a21o_1
X_5202_ _1728_ _1729_ _1721_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5133_ _1016_ _1553_ _1567_ _0997_ _1663_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__o221a_1
X_5064_ sound3.count\[6\] _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4015_ seq.tempo_select.state\[1\] net846 vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ sound1.divisor_m\[8\] sound1.count_m\[7\] vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7705_ _2843_ _3751_ vssd1 vssd1 vccd1 vccd1 _3752_ sky130_fd_sc_hd__and2_1
X_5897_ sound4.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__inv_2
X_4917_ _1014_ _1322_ _1467_ _0499_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4848_ _0954_ _1321_ _1327_ _0973_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__o22a_1
X_7636_ _3681_ _3703_ _3704_ _2184_ net360 vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7567_ _3660_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__clkbuf_1
X_4779_ _0698_ _0499_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__or2_1
X_7498_ _3645_ vssd1 vssd1 vccd1 vccd1 _3646_ sky130_fd_sc_hd__inv_2
X_6518_ _0579_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__buf_6
X_6449_ net417 _2201_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8119_ clknet_leaf_60_hwclk _0240_ net94 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_50_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5820_ _2263_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5751_ sound4.sdiv.Q\[27\] _2183_ sound4.sdiv.next_dived net180 vssd1 vssd1 vccd1
+ vccd1 _0027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4702_ _1268_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[4\] sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_65_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7421_ _3577_ _3580_ vssd1 vssd1 vccd1 vccd1 _3581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5682_ sound4.sdiv.A\[18\] _2037_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4633_ _0978_ _0996_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__or2_2
XFILLER_0_130_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7352_ _3514_ _3517_ vssd1 vssd1 vccd1 vccd1 _3519_ sky130_fd_sc_hd__nand2_1
X_4564_ _1107_ net59 vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold602 _3381_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__dlygate4sd3_1
X_7283_ sound3.divisor_m\[3\] _3456_ vssd1 vssd1 vccd1 vccd1 _3457_ sky130_fd_sc_hd__xnor2_1
Xhold624 sound1.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ sound3.sdiv.Q\[7\] _2301_ _2732_ _2733_ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold635 sound4.sdiv.C\[5\] vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold613 sound4.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold679 wave_comb.u1.C\[0\] vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _2619_ _2629_ _2628_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__a21o_1
Xhold646 sound1.divisor_m\[4\] vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 wave_comb.u1.M\[0\] vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ _1000_ _1063_ _1064_ _0994_ _1065_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__o221a_1
Xhold668 sound2.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
X_6165_ _2596_ _2599_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ sound3.count_m\[8\] vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5116_ _1083_ _1550_ _1565_ _0960_ _1646_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__o221a_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _0540_ _1552_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__nand2_4
Xclkbuf_leaf_18_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_6998_ _3248_ _3254_ _3261_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5949_ sound1.count_m\[11\] vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7619_ _2130_ _2103_ vssd1 vssd1 vccd1 vccd1 _3692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4280_ _0857_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7970_ clknet_leaf_24_hwclk _0133_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_6921_ sound2.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__inv_2
X_6852_ _2863_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__buf_8
X_5803_ _2239_ _2241_ _2244_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__nor3_1
XFILLER_0_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3995_ _0651_ _0649_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[4\] sky130_fd_sc_hd__xnor2_1
X_6783_ net207 _2894_ _2890_ net336 _2839_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5734_ net832 _2186_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5665_ _2146_ _2147_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__nor2_1
X_7404_ _3564_ _3565_ vssd1 vssd1 vccd1 vccd1 _3566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4616_ sound1.count\[5\] _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7335_ _3500_ _3502_ vssd1 vssd1 vccd1 vccd1 _3504_ sky130_fd_sc_hd__nand2_1
Xhold410 wave_comb.u1.A\[6\] vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlygate4sd3_1
X_5596_ _2077_ _2078_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__nand2_1
Xhold443 pm.count\[2\] vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 sound1.sdiv.Q\[0\] vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _0002_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _0958_ _1110_ _1115_ _1117_ _1070_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__o2111a_1
Xhold454 seq.clk_div.next_count\[1\] vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 pm.count\[6\] vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__dlygate4sd3_1
X_7266_ sound3.divisor_m\[1\] _3441_ vssd1 vssd1 vccd1 vccd1 _3442_ sky130_fd_sc_hd__xnor2_1
Xhold476 _0650_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _0136_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _1001_ _1047_ _1048_ _0947_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__o22a_1
X_7197_ net300 _3132_ _3399_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a21o_1
X_6217_ _2607_ _2609_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold498 sound2.count_m\[3\] vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__dlygate4sd3_1
X_6148_ sound4.sdiv.Q\[2\] _2582_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__nand2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _2513_ sound3.divisor_m\[7\] _2514_ sound3.divisor_m\[6\] vssd1 vssd1 vccd1
+ vccd1 _2515_ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3780_ _0447_ _0461_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5450_ sound4.count\[6\] _1951_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__and2_1
X_4401_ _0675_ _0687_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5381_ _0946_ _1786_ _1790_ _0971_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7120_ net868 _3329_ vssd1 vssd1 vccd1 vccd1 _3370_ sky130_fd_sc_hd__xnor2_1
X_4332_ seq.player_6.state\[1\] _0894_ _0896_ _0902_ vssd1 vssd1 vccd1 vccd1 _0903_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4263_ seq.clk_div.count\[14\] _0841_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__or2_1
X_7051_ sound2.divisor_m\[17\] _3309_ vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__xnor2_1
X_6002_ _2435_ _2277_ _2434_ vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__or3b_1
X_4194_ seq.clk_div.count\[6\] seq.clk_div.count\[12\] seq.clk_div.count\[16\] _0779_
+ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__or4_1
X_7953_ clknet_leaf_20_hwclk _0116_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6904_ sound2.divisor_m\[1\] sound2.divisor_m\[0\] _3177_ vssd1 vssd1 vccd1 vccd1
+ _3178_ sky130_fd_sc_hd__o21a_1
X_7884_ clknet_leaf_92_hwclk net12 net66 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6835_ _0554_ vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__buf_6
XFILLER_0_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6766_ sound1.sdiv.C\[3\] _0565_ _3106_ net953 vssd1 vssd1 vccd1 vccd1 _3110_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3978_ _0446_ _0628_ _0626_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__o21a_1
X_5717_ net328 _2182_ _2185_ net462 _2189_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a221o_1
X_6697_ _2890_ _3052_ _3053_ _2894_ net429 vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5648_ _2103_ _2129_ _2130_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8367_ clknet_leaf_73_hwclk rate_clk.next_count\[4\] net76 vssd1 vssd1 vccd1 vccd1
+ rate_clk.count\[4\] sky130_fd_sc_hd__dfrtp_1
X_5579_ _2060_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__inv_2
X_7318_ _3477_ _3480_ _3488_ vssd1 vssd1 vccd1 vccd1 _3489_ sky130_fd_sc_hd__nand3_1
Xhold262 _0029_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 sound2.sdiv.Q\[18\] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd3_1
X_8298_ clknet_leaf_72_hwclk _0398_ net80 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[12\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold251 _0373_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__dlygate4sd3_1
X_7249_ _3430_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__clkbuf_1
Xhold284 sound1.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _0160_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 sound2.count_m\[6\] vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput8 piano_keys[14] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4950_ _1444_ _1461_ _1479_ _1500_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__or4_1
X_3901_ wave_comb.u1.C\[3\] wave_comb.u1.C\[2\] _0570_ wave_comb.u1.C\[5\] wave_comb.u1.C\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__a2111o_4
X_4881_ _0687_ _1001_ _1338_ _1336_ _1112_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__o32a_1
XFILLER_0_47_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6620_ sound1.divisor_m\[10\] _2977_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__or2_1
X_3832_ _0479_ _0478_ _0485_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__and3_1
X_6551_ _2918_ _2921_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__nor2_1
X_5502_ sound4.count\[15\] sound4.count\[16\] _1984_ sound4.count\[17\] vssd1 vssd1
+ vccd1 vccd1 _1996_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3763_ _0446_ inputcont.INTERNAL_SYNCED_I\[11\] inputcont.INTERNAL_SYNCED_I\[10\]
+ _0445_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or4_2
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6482_ net773 _1071_ _2864_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8221_ clknet_leaf_37_hwclk sound3.osc.next_count\[2\] net93 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[2\] sky130_fd_sc_hd__dfrtp_4
X_5433_ sound4.count\[0\] sound4.count\[1\] sound4.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1942_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8152_ clknet_leaf_30_hwclk net237 net90 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5364_ _1778_ _1874_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7103_ net964 _3329_ _3354_ vssd1 vssd1 vccd1 vccd1 _3356_ sky130_fd_sc_hd__a21boi_1
X_4315_ select1.sequencer_on _0885_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__and2_1
X_5295_ _1176_ _1769_ _1777_ _1174_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__o22a_1
X_8083_ clknet_leaf_75_hwclk _0225_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_7034_ _3291_ _3293_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__nand2_1
X_4246_ seq.clk_div.count\[8\] seq.clk_div.count\[9\] seq.clk_div.count\[10\] _0824_
+ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__and4_1
X_4177_ net792 _0772_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7936_ clknet_leaf_19_hwclk _0099_ net85 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7867_ clknet_leaf_3_hwclk net107 net70 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_sync\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6818_ net398 _2857_ _3123_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7798_ clknet_leaf_43_hwclk net8 net99 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6749_ _3096_ _3097_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5080_ _0542_ _1551_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__or2_1
X_4100_ net650 _0721_ net901 vssd1 vssd1 vccd1 vccd1 seq.player_7.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_4031_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__inv_6
X_5982_ sound1.divisor_m\[1\] _2415_ _2416_ _2417_ vssd1 vssd1 vccd1 vccd1 _2418_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7721_ clknet_leaf_58_hwclk net601 net94 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_4933_ _1041_ _1343_ _1333_ _1129_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7652_ _2061_ _2141_ _2057_ vssd1 vssd1 vccd1 vccd1 _3716_ sky130_fd_sc_hd__a21o_1
X_4864_ _0684_ _1343_ _1333_ _0686_ _1341_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__o221a_1
X_6603_ sound1.sdiv.A\[8\] _2968_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3815_ _0483_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__nand2_1
X_4795_ net38 _1315_ _1319_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__or3_1
X_7583_ _3669_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6534_ _2901_ _2906_ vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6465_ _1104_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8204_ clknet_leaf_44_hwclk _0325_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_5416_ _0978_ _0944_ _1777_ _1794_ _1001_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__o32a_1
XFILLER_0_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6396_ net700 _2817_ _2808_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5347_ _0948_ _1800_ _1853_ _1857_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8135_ clknet_leaf_93_hwclk net346 net67 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_8066_ clknet_leaf_84_hwclk net293 net74 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5278_ net46 _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__or2_1
X_7017_ _3268_ _3272_ _3279_ vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__a21o_1
X_4229_ seq.clk_div.count\[4\] _0815_ seq.clk_div.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0820_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap59 _1040_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_8
X_7919_ clknet_leaf_18_hwclk net390 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4580_ _0696_ _1055_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nand2_2
Xinput11 piano_keys[3] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold817 _0774_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 seq.player_1.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold806 seq.player_4.next_state\[2\] vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 sound1.sdiv.A\[8\] vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__dlygate4sd3_1
X_6250_ wave_comb.u1.next_start _2681_ _2682_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6181_ net679 _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__and3_1
X_5201_ sound3.count\[0\] sound3.count\[1\] sound3.count\[2\] sound3.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5132_ _1113_ _1570_ _1574_ _1112_ _1662_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__o221a_1
X_5063_ _1586_ _1593_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__nand2_1
X_4014_ net474 _0663_ vssd1 vssd1 vccd1 vccd1 seq.tempo_select.next_state\[0\] sky130_fd_sc_hd__nand2_1
X_5965_ _2396_ sound1.divisor_m\[7\] _2398_ sound1.divisor_m\[6\] vssd1 vssd1 vccd1
+ vccd1 _2401_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7704_ sound4.sdiv.C\[3\] _0556_ _3747_ net898 vssd1 vssd1 vccd1 vccd1 _3751_ sky130_fd_sc_hd__a31o_1
X_4916_ _1025_ _1028_ _1325_ _1418_ _1011_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__o32a_1
X_5896_ sound4.count_m\[14\] _2331_ sound4.count_m\[13\] _2142_ vssd1 vssd1 vccd1
+ vccd1 _2332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4847_ _0959_ _0993_ _1341_ _1336_ _0979_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__o32a_1
X_7635_ _2135_ _3702_ vssd1 vssd1 vccd1 vccd1 _3704_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7566_ net794 _1850_ _3419_ vssd1 vssd1 vccd1 vccd1 _3660_ sky130_fd_sc_hd__mux2_1
X_4778_ _0686_ _1321_ _1322_ _1134_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__o221a_1
X_7497_ sound3.sdiv.C\[2\] sound3.sdiv.C\[1\] sound3.sdiv.C\[0\] vssd1 vssd1 vccd1
+ vccd1 _3645_ sky130_fd_sc_hd__and3_1
X_6517_ sound1.divisor_m\[0\] sound1.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6448_ net288 _2836_ _2849_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__a21o_1
X_6379_ net33 _2804_ _0700_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__o21a_4
X_8118_ clknet_leaf_40_hwclk sound3.sdiv.next_dived net98 vssd1 vssd1 vccd1 vccd1
+ sound3.sdiv.dived sky130_fd_sc_hd__dfrtp_1
X_8049_ clknet_leaf_90_hwclk _0191_ net68 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5750_ net180 _2182_ _2185_ net214 _2206_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4701_ _1256_ _1266_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__and3_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _2162_ _2163_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__or2b_1
X_7420_ sound3.divisor_m\[17\] _3579_ vssd1 vssd1 vccd1 vccd1 _3580_ sky130_fd_sc_hd__xnor2_1
X_4632_ _1003_ _1134_ _1125_ _0976_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7351_ _3514_ _3517_ vssd1 vssd1 vccd1 vccd1 _3518_ sky130_fd_sc_hd__or2_1
Xhold603 pm.current_waveform\[7\] vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlygate4sd3_1
X_4563_ _1107_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__nor2_4
XFILLER_0_130_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7282_ sound3.divisor_m\[2\] sound3.divisor_m\[1\] sound3.divisor_m\[0\] _3448_ vssd1
+ vssd1 vccd1 vccd1 _3456_ sky130_fd_sc_hd__o31a_1
X_6302_ sound3.sdiv.Q\[6\] _2731_ _2292_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__a21o_1
Xhold636 sound1.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _0979_ _1003_ _0943_ _0983_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__o22a_1
Xhold614 _0431_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 seq.player_2.state\[1\] vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold647 sound3.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold669 sound1.divisor_m\[6\] vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ _2664_ _2665_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__and2b_1
Xhold658 sound4.divisor_m\[6\] vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6164_ _2597_ _2506_ _2598_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__a21oi_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ sound3.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5115_ _1078_ _1559_ _1572_ _1039_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__o22a_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5046_ _1041_ _1562_ _1565_ _1101_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6997_ _3248_ _3254_ _3261_ vssd1 vssd1 vccd1 vccd1 _3262_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5948_ sound1.count_m\[13\] _2376_ _2383_ sound1.count_m\[12\] vssd1 vssd1 vccd1
+ vccd1 _2384_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5879_ sound4.count_m\[7\] vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7618_ _3681_ _3690_ _3691_ _2184_ net232 vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7549_ net518 _3403_ _2197_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6920_ net437 _3168_ sound2.sdiv.next_dived _3192_ vssd1 vssd1 vccd1 vccd1 _0210_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6851_ _1396_ vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__inv_2
X_5802_ _2247_ _2248_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3994_ net692 vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__inv_2
X_6782_ net336 _2894_ _2890_ net439 _2838_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5733_ net242 _2182_ _2185_ sound4.sdiv.Q\[17\] _2197_ vssd1 vssd1 vccd1 vccd1 _0018_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5664_ sound4.sdiv.A\[14\] _2144_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__nor2_1
X_7403_ _3560_ _3563_ vssd1 vssd1 vccd1 vccd1 _3565_ sky130_fd_sc_hd__nand2_1
X_4615_ _1026_ _0939_ _1174_ _0990_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5595_ sound4.sdiv.A\[9\] _2076_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__or2_1
X_7334_ _3500_ _3502_ vssd1 vssd1 vccd1 vccd1 _3503_ sky130_fd_sc_hd__or2_2
Xhold400 _0306_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 wave_comb.u1.A\[5\] vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _0990_ _1064_ _1116_ _0994_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold444 pm.next_count\[2\] vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 seq.clk_div.count\[4\] vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold433 seq.player_8.state\[3\] vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 _0656_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 pm.next_count\[3\] vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__dlygate4sd3_1
X_7265_ sound3.sdiv.A\[26\] sound3.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 _3441_ sky130_fd_sc_hd__and2b_1
Xhold455 sound1.count_m\[10\] vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _0990_ _0996_ net59 _0969_ _0943_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__o221a_1
Xhold499 sound3.sdiv.Q\[5\] vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__dlygate4sd3_1
X_6216_ _2648_ _2649_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__or2b_1
X_7196_ net853 _2863_ vssd1 vssd1 vccd1 vccd1 _3399_ sky130_fd_sc_hd__and2_1
Xhold488 sound4.sdiv.A\[23\] vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__dlygate4sd3_1
X_6147_ sound4.sdiv.Q\[0\] sound4.sdiv.Q\[1\] _0576_ _2370_ vssd1 vssd1 vccd1 vccd1
+ _2582_ sky130_fd_sc_hd__o211a_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ sound3.count_m\[5\] vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__inv_2
X_5029_ _0698_ _0540_ net43 vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__or3_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_64_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4400_ _0674_ _0970_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__nor2_8
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5380_ _1778_ _1887_ _1890_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__and3_2
X_4331_ seq.player_7.state\[1\] _0898_ _0901_ seq.player_8.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _0902_ sky130_fd_sc_hd__a22o_1
X_4262_ seq.clk_div.count\[13\] seq.clk_div.count\[14\] _0838_ vssd1 vssd1 vccd1 vccd1
+ _0844_ sky130_fd_sc_hd__and3_1
X_7050_ _3177_ _3308_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__and2_1
X_6001_ sound1.sdiv.Q\[0\] _0579_ _2434_ _2436_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4193_ seq.tempo_select.state\[0\] seq.clk_div.count\[4\] vssd1 vssd1 vccd1 vccd1
+ _0787_ sky130_fd_sc_hd__nand2_1
X_7952_ clknet_leaf_20_hwclk _0115_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6903_ sound2.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7883_ clknet_leaf_94_hwclk net11 net66 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6834_ net358 _2857_ _3131_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6765_ _2005_ _3108_ _3109_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__nor3_1
XFILLER_0_92_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3977_ _0638_ _0639_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5716_ sound4.count\[2\] _2186_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6696_ _3050_ _3051_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5647_ sound4.sdiv.A\[4\] _2102_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8366_ clknet_leaf_73_hwclk rate_clk.next_count\[3\] net76 vssd1 vssd1 vccd1 vccd1
+ rate_clk.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_5578_ _2058_ _2060_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__nand2_1
X_7317_ _3486_ _3487_ vssd1 vssd1 vccd1 vccd1 _3488_ sky130_fd_sc_hd__nand2_1
Xhold230 _0087_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 sound1.sdiv.Q\[20\] vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _0674_ _0687_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__nor2_1
Xhold241 sound2.sdiv.Q\[15\] vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__dlygate4sd3_1
X_8297_ clknet_leaf_72_hwclk _0397_ net80 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_7248_ net749 _1628_ _3419_ vssd1 vssd1 vccd1 vccd1 _3430_ sky130_fd_sc_hd__mux2_1
Xhold263 sound3.count\[16\] vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 sound1.count_m\[12\] vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 sound2.count\[10\] vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _0175_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7179_ net200 _3132_ _3390_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a21o_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 piano_keys[1] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3900_ wave_comb.u1.start vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__inv_2
X_4880_ _1034_ _1427_ _1428_ _1430_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3831_ _0507_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__inv_2
X_6550_ _2419_ _2920_ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3762_ inputcont.INTERNAL_SYNCED_I\[12\] vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5501_ sound4.count\[16\] sound4.count\[17\] _1988_ vssd1 vssd1 vccd1 vccd1 _1995_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_27_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6481_ _2869_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8220_ clknet_leaf_35_hwclk sound3.osc.next_count\[1\] net93 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[1\] sky130_fd_sc_hd__dfrtp_4
X_5432_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__inv_2
X_8151_ clknet_leaf_30_hwclk _0272_ net90 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5363_ _1107_ _1869_ _1872_ _1873_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7102_ sound2.sdiv.A\[22\] _3329_ vssd1 vssd1 vccd1 vccd1 _3355_ sky130_fd_sc_hd__xor2_1
X_4314_ _0702_ seq.encode.play _0884_ inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1
+ vccd1 vccd1 _0885_ sky130_fd_sc_hd__a31o_1
X_5294_ _1180_ _1786_ _1790_ _1028_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__o22a_1
X_8082_ clknet_leaf_79_hwclk _0224_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7033_ _3291_ _3293_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__or2_1
X_4245_ _0831_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_4176_ seq.player_1.state\[2\] net920 vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7935_ clknet_leaf_10_hwclk _0098_ net83 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7866_ clknet_leaf_93_hwclk seq.tempo_select.next_state\[1\] net66 vssd1 vssd1 vccd1
+ vccd1 seq.tempo_select.state\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6817_ net808 _2855_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__and2_1
X_7797_ clknet_leaf_74_hwclk net7 net76 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6748_ sound1.sdiv.A\[25\] _3055_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6679_ _2903_ _3036_ vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8349_ clknet_leaf_85_hwclk sound4.osc.next_count\[7\] net77 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4030_ oct.state\[2\] vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__buf_12
X_5981_ sound1.divisor_m\[2\] sound1.count_m\[1\] vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7720_ clknet_leaf_58_hwclk _0005_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4932_ _0944_ _1336_ _1345_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7651_ _2057_ _2061_ _2141_ vssd1 vssd1 vccd1 vccd1 _3715_ sky130_fd_sc_hd__nand3_1
X_6602_ sound1.divisor_m\[9\] _2967_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__xnor2_1
X_4863_ _1379_ _1388_ _1397_ _1413_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__or4_1
X_3814_ _0479_ _0478_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__or2b_1
X_4794_ _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__buf_4
X_7582_ net884 _1803_ _3419_ vssd1 vssd1 vccd1 vccd1 _3669_ sky130_fd_sc_hd__mux2_1
X_6533_ _2902_ _2905_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6464_ net159 _2857_ _2858_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__a21o_1
X_8203_ clknet_leaf_45_hwclk _0324_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_113_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5415_ _0954_ _1784_ _1790_ _0948_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__o22a_1
X_6395_ _2816_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5346_ _1095_ _1792_ _1855_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8134_ clknet_leaf_91_hwclk net326 net67 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8065_ clknet_leaf_83_hwclk net490 net74 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5277_ _0673_ _1773_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__or2_1
X_7016_ _3277_ _3278_ vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__nand2_1
X_4228_ seq.clk_div.count\[4\] seq.clk_div.count\[5\] _0815_ vssd1 vssd1 vccd1 vccd1
+ _0819_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4159_ seq.player_2.state\[1\] seq.player_2.state\[2\] seq.player_2.state\[3\] _0762_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__a311o_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ clknet_leaf_17_hwclk net289 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7849_ clknet_leaf_99_hwclk seq.clk_div.next_count\[6\] net65 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 piano_keys[4] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold807 sound3.count\[1\] vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold818 sound4.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold829 sound2.count\[6\] vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6180_ _2613_ _2614_ net695 _0569_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__a2bb2o_1
X_5200_ net862 sound3.count\[1\] sound3.count\[2\] sound3.count\[3\] vssd1 vssd1 vccd1
+ vccd1 _1728_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5131_ _1064_ _1565_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5062_ _1038_ _1587_ _1589_ _1592_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__o211a_1
X_4013_ _0661_ net473 seq.tempo_select.state\[0\] vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5964_ _2398_ sound1.divisor_m\[6\] sound1.divisor_m\[5\] _2399_ vssd1 vssd1 vccd1
+ vccd1 _2400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7703_ _2005_ _3749_ _3750_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4915_ _1025_ _1345_ _1462_ _1465_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__o211a_1
X_5895_ sound4.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ sound2.count\[7\] _1368_ _1396_ sound2.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _1397_ sky130_fd_sc_hd__a2bb2o_1
X_7634_ _3702_ _2135_ vssd1 vssd1 vccd1 vccd1 _3703_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7565_ _3659_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6516_ sound1.divisor_m\[0\] sound1.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4777_ _1198_ _1323_ _1327_ _1204_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7496_ net567 net806 net599 vssd1 vssd1 vccd1 vccd1 _3644_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6447_ sound1.count\[11\] _2201_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6378_ _0632_ _0643_ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8117_ clknet_leaf_82_hwclk sound2.osc.next_count\[18\] net74 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[18\] sky130_fd_sc_hd__dfrtp_1
X_5329_ _0959_ _1833_ _1834_ _1835_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__o2111a_1
X_8048_ clknet_leaf_90_hwclk _0190_ net68 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4700_ sound1.count\[4\] _1263_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__or2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _2159_ _2161_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4631_ _0939_ _1200_ _1189_ _0990_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7350_ sound3.divisor_m\[10\] _3516_ vssd1 vssd1 vccd1 vccd1 _3517_ sky130_fd_sc_hd__xnor2_1
X_4562_ _0674_ _0681_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__nor2_4
XFILLER_0_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7281_ sound3.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _3455_ sky130_fd_sc_hd__inv_2
Xhold626 sound1.sdiv.C\[5\] vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 pm.current_waveform\[6\] vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
X_6301_ sound3.sdiv.Q\[6\] _0577_ _2731_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__a21oi_1
Xhold604 wave_comb.u1.Q\[7\] vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4493_ _0674_ _0684_ _0683_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a21oi_4
Xhold637 sound3.divisor_m\[5\] vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _2659_ _2663_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold648 seq.player_4.state\[2\] vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 seq.player_3.state\[2\] vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6163_ _2439_ _2504_ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__and2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ sound3.divisor_m\[14\] _2521_ _2529_ sound3.count_m\[14\] vssd1 vssd1 vccd1
+ vccd1 _2530_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5114_ _1015_ _1562_ _1570_ _0952_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__o221a_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _1095_ _1567_ _1570_ _1097_ _1575_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__o221a_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6996_ _3259_ _3260_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5947_ sound1.divisor_m\[13\] vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__inv_2
X_7617_ _2110_ _2128_ vssd1 vssd1 vccd1 vccd1 _3691_ sky130_fd_sc_hd__or2_1
X_5878_ sound4.divisor_m\[5\] _2312_ _2313_ sound4.divisor_m\[4\] vssd1 vssd1 vccd1
+ vccd1 _2314_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4829_ _1125_ _1321_ _1327_ _1127_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__o22a_1
X_7548_ net455 _3403_ _2196_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__a21o_1
X_7479_ net976 _3595_ vssd1 vssd1 vccd1 vccd1 _3631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1 net816 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_1
X_6850_ _3140_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ wave_comb.u1.A\[7\] _2224_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__or2_1
X_6781_ sound1.sdiv.Q\[8\] _2894_ _2890_ net192 _2837_ vssd1 vssd1 vccd1 vccd1 _0149_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3993_ _0649_ net580 vssd1 vssd1 vccd1 vccd1 pm.next_count\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_85_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5732_ sound4.count\[10\] _2186_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5663_ _2145_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__inv_2
X_7402_ _3560_ _3563_ vssd1 vssd1 vccd1 vccd1 _3564_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4614_ _0958_ _1141_ _1179_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5594_ net960 _2076_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__nand2_1
X_7333_ sound3.divisor_m\[8\] _3501_ vssd1 vssd1 vccd1 vccd1 _3502_ sky130_fd_sc_hd__xnor2_1
X_4545_ _0695_ net60 net59 vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold401 sound4.sdiv.A\[8\] vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold412 sound3.sdiv.Q\[4\] vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 sound3.count_m\[10\] vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 sound1.count_m\[3\] vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold434 seq.player_8.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7264_ _3437_ _3438_ _3439_ _3440_ net503 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a32o_1
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold478 wave_comb.u1.A\[4\] vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 _0080_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 sound2.sdiv.Q\[3\] vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _0950_ _0996_ _1046_ _0994_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7195_ net347 _3132_ _3398_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6215_ _2645_ _2647_ vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__nand2_1
Xhold489 wave_comb.u1.A\[2\] vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6146_ wave_comb.u1.next_start _2580_ _2581_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__a21o_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ sound3.count_m\[6\] vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__inv_2
X_5028_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__buf_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6979_ sound2.divisor_m\[9\] sound2.divisor_m\[8\] sound2.divisor_m\[7\] _3221_ vssd1
+ vssd1 vccd1 vccd1 _3245_ sky130_fd_sc_hd__or4_1
XFILLER_0_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_hwclk hwclk vssd1 vssd1 vccd1 vccd1 clknet_0_hwclk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4330_ select1.sequencer_on _0897_ _0899_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__a31oi_2
X_4261_ _0843_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
X_6000_ _2435_ sound1.sdiv.next_start vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4192_ seq.tempo_select.state\[0\] _0781_ _0784_ _0785_ vssd1 vssd1 vccd1 vccd1 _0786_
+ sky130_fd_sc_hd__o22ai_1
X_7951_ clknet_leaf_32_hwclk _0114_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7882_ clknet_leaf_99_hwclk net10 net65 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6902_ sound2.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__inv_2
X_6833_ net394 _2855_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6764_ _0565_ _3106_ net714 vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3976_ inputcont.INTERNAL_SYNCED_I\[9\] _0624_ _0622_ vssd1 vssd1 vccd1 vccd1 _0639_
+ sky130_fd_sc_hd__a21oi_1
X_6695_ _3050_ _3051_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5715_ sound4.sdiv.Q\[9\] _2184_ _2185_ net222 _2188_ vssd1 vssd1 vccd1 vccd1 _0009_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5646_ _2110_ _2128_ _2107_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold220 sound3.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8365_ clknet_leaf_73_hwclk net169 net76 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5577_ sound4.divisor_m\[13\] _2059_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__xnor2_2
X_7316_ _3482_ _3485_ vssd1 vssd1 vccd1 vccd1 _3487_ sky130_fd_sc_hd__nand2_1
Xhold231 sound1.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _0162_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ _0939_ _1095_ _1056_ _0958_ _1098_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__o221a_1
Xhold242 _0256_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8296_ clknet_leaf_64_hwclk _0396_ net79 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_7247_ _3429_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__clkbuf_1
Xhold286 _0082_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _1000_ _1025_ _1027_ _0976_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__o221a_1
Xhold275 sound2.sdiv.Q\[13\] vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 sound4.sdiv.Q\[21\] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 sound4.sdiv.Q\[14\] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__dlygate4sd3_1
X_7178_ sound3.count\[3\] _2863_ vssd1 vssd1 vccd1 vccd1 _3390_ sky130_fd_sc_hd__and2_1
X_6129_ _2564_ _2530_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__or2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3830_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3761_ inputcont.INTERNAL_SYNCED_I\[9\] inputcont.INTERNAL_SYNCED_I\[8\] _0443_ _0444_
+ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__or4_4
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5500_ _1994_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6480_ net795 _1186_ _2864_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5431_ sound4.count\[0\] sound4.count\[1\] sound4.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1940_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8150_ clknet_leaf_34_hwclk net201 net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5362_ _0677_ _1083_ _1784_ _1777_ _1064_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__o32a_1
XFILLER_0_112_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8081_ clknet_leaf_78_hwclk _0223_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_7101_ _3349_ _3353_ _3354_ _3174_ net476 vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__a32o_1
X_4313_ seq.beat\[0\] seq.beat\[2\] seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__and3b_1
X_7032_ sound2.divisor_m\[15\] _3292_ vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__xnor2_1
X_5293_ sound4.count\[10\] _1803_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__xor2_1
X_4244_ _0829_ _0813_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__and3b_1
XFILLER_0_93_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4175_ seq.player_1.state\[2\] net565 _0772_ _0773_ _0700_ vssd1 vssd1 vccd1 vccd1
+ seq.player_1.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
XFILLER_0_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7934_ clknet_leaf_19_hwclk _0097_ net85 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7865_ clknet_leaf_95_hwclk net475 net66 vssd1 vssd1 vccd1 vccd1 seq.tempo_select.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_7796_ clknet_leaf_55_hwclk net6 net96 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_6816_ net233 _2857_ _3122_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6747_ net699 _3055_ vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3959_ inputcont.INTERNAL_SYNCED_I\[7\] _0621_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6678_ sound1.divisor_m\[16\] _3028_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5629_ sound4.divisor_m\[2\] sound4.divisor_m\[1\] sound4.divisor_m\[0\] _2036_ vssd1
+ vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8348_ clknet_leaf_87_hwclk sound4.osc.next_count\[6\] net77 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[6\] sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_78_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_8279_ clknet_leaf_65_hwclk net250 net79 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_16_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5980_ sound1.count_m\[1\] sound1.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4931_ _1035_ _1323_ _1322_ _1039_ _1481_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4862_ sound2.count\[1\] _1404_ _1412_ sound2.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _1413_ sky130_fd_sc_hd__a2bb2o_1
X_7650_ net661 _2183_ sound4.sdiv.next_dived _3714_ vssd1 vssd1 vccd1 vccd1 _0418_
+ sky130_fd_sc_hd__a22o_1
X_6601_ _2395_ _2957_ sound1.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3813_ inputcont.INTERNAL_SYNCED_I\[10\] _0445_ _0488_ _0491_ vssd1 vssd1 vccd1 vccd1
+ _0492_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4793_ _1331_ _1334_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__or2_1
X_7581_ _2005_ _1840_ _3668_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__a21oi_1
X_6532_ sound1.divisor_m\[2\] _2904_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6463_ sound1.count\[18\] _2855_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8202_ clknet_leaf_43_hwclk _0323_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5414_ sound4.count\[12\] _1924_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__xor2_1
X_6394_ _2623_ _2655_ _2805_ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8133_ clknet_leaf_91_hwclk _0254_ net67 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5345_ _0993_ _1012_ _1790_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8064_ clknet_leaf_82_hwclk _0206_ net74 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_5276_ _1125_ _1784_ _1786_ _1127_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__o22a_1
X_7015_ _3273_ _3276_ vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__nand2_1
X_4227_ net526 _0815_ _0818_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[4\] sky130_fd_sc_hd__a21oi_1
X_4158_ seq.player_2.state\[0\] _0761_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__and2_1
X_4089_ net885 _0713_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__nor2_1
X_7917_ clknet_leaf_17_hwclk net560 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7848_ clknet_leaf_99_hwclk seq.clk_div.next_count\[5\] net65 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_7779_ clknet_leaf_59_hwclk _0053_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 piano_keys[5] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold819 sound3.sdiv.C\[4\] vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold808 inputcont.u1.ff_intermediate\[1\] vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5130_ _0687_ _1001_ _1578_ _1572_ _1116_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__o32a_1
X_5061_ _1026_ _1559_ _1572_ _1064_ _1591_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__o221a_1
X_4012_ _0661_ net473 net846 vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5963_ sound1.count_m\[4\] vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__inv_2
X_7702_ _0556_ _3747_ net704 vssd1 vssd1 vccd1 vccd1 _3750_ sky130_fd_sc_hd__a21oi_1
X_4914_ _1005_ _1338_ _1336_ _1027_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__o221a_1
X_5894_ sound4.divisor_m\[13\] _2324_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4845_ _1390_ _1392_ _1395_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7633_ _2136_ _2083_ vssd1 vssd1 vccd1 vccd1 _3702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7564_ net766 _3658_ _3419_ vssd1 vssd1 vccd1 vccd1 _3659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4776_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6515_ _0867_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__buf_6
XFILLER_0_90_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7495_ _1545_ vssd1 vssd1 vccd1 vccd1 _3643_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6446_ net559 _2836_ _2848_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__a21o_1
X_6377_ wave_comb.u1.Q\[11\] _0573_ wave_comb.u1.next_dived net127 vssd1 vssd1 vccd1
+ vccd1 _0056_ sky130_fd_sc_hd__a22o_1
X_8116_ clknet_leaf_82_hwclk sound2.osc.next_count\[17\] net74 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[17\] sky130_fd_sc_hd__dfrtp_2
X_5328_ _1077_ _1769_ _1836_ _1838_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8047_ clknet_leaf_90_hwclk _0189_ net2 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_5259_ _0673_ _1765_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4630_ _0686_ _0950_ _0994_ _1146_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6300_ sound3.sdiv.Q\[5\] _2632_ _2699_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__a21o_1
X_4561_ _0967_ _1123_ _1125_ _0958_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__o221a_1
X_7280_ _3447_ _3450_ vssd1 vssd1 vccd1 vccd1 _3454_ sky130_fd_sc_hd__or2_1
Xhold616 sound3.sdiv.C\[3\] vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold605 sound1.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _0964_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__nand2_2
Xhold627 seq.player_8.state\[2\] vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6231_ _2659_ _2663_ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__nor2_1
Xhold638 sound2.divisor_m\[11\] vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 seq.player_5.state\[2\] vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__dlygate4sd3_1
X_6162_ _2439_ _2504_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5113_ _1079_ _1580_ _1574_ _0680_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ sound3.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__inv_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5044_ _1572_ _1574_ _0960_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__a21o_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6995_ _3255_ _3258_ vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5946_ sound1.count_m\[15\] _2381_ sound1.count_m\[14\] _2375_ vssd1 vssd1 vccd1
+ vccd1 _2382_ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5877_ sound4.count_m\[3\] vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__inv_2
X_7616_ _3689_ vssd1 vssd1 vccd1 vccd1 _3690_ sky130_fd_sc_hd__inv_2
X_4828_ sound2.count\[6\] _1378_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4759_ _0575_ _0560_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__nor2_4
X_7547_ net229 _3403_ _2195_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a21o_1
X_7478_ sound3.sdiv.A\[24\] _3595_ vssd1 vssd1 vccd1 vccd1 _3630_ sky130_fd_sc_hd__nor2_1
X_6429_ net543 _2836_ _2839_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2 inputcont.u1.ff_intermediate\[2\] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3992_ net579 _0647_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__nor2_1
X_5800_ net947 _2224_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__nand2_1
X_6780_ net192 _2894_ _2890_ net585 vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5731_ net350 _2182_ _2185_ sound4.sdiv.Q\[16\] _2196_ vssd1 vssd1 vccd1 vccd1 _0017_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5662_ sound4.sdiv.A\[14\] _2144_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__nand2_1
X_7401_ sound3.divisor_m\[15\] _3562_ vssd1 vssd1 vccd1 vccd1 _3563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4613_ _0969_ _1180_ _1181_ _0967_ _1183_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5593_ _2075_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__inv_2
X_7332_ sound3.divisor_m\[7\] _3492_ _3448_ vssd1 vssd1 vccd1 vccd1 _3501_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4544_ _0976_ _1112_ _1113_ _1000_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold402 sound4.count_m\[14\] vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _0344_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__dlygate4sd3_1
X_7263_ _0577_ vssd1 vssd1 vccd1 vccd1 _3440_ sky130_fd_sc_hd__clkbuf_8
Xhold424 _0073_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold435 seq.player_3.state\[3\] vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6214_ _2645_ _2647_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__nor2_1
Xhold457 wave_comb.u1.A\[8\] vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _0244_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _0674_ _0945_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__nor2_4
Xhold446 sound2.sdiv.C\[1\] vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_1
Xhold479 sound1.sdiv.A\[24\] vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7194_ sound3.count\[11\] _2863_ vssd1 vssd1 vccd1 vccd1 _3398_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6145_ wave_comb.u1.Q\[2\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ sound3.divisor_m\[5\] _2511_ _2508_ sound3.divisor_m\[4\] vssd1 vssd1 vccd1
+ vccd1 _2512_ sky130_fd_sc_hd__o22a_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _1556_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__or2_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6978_ sound2.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5929_ _2364_ _2332_ _2342_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _0841_ _0813_ _0842_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4191_ seq.tempo_select.state\[0\] seq.tempo_select.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7950_ clknet_leaf_24_hwclk _0113_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6901_ _3170_ sound2.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__or2b_1
X_7881_ clknet_leaf_71_hwclk net9 net80 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6832_ net286 _2857_ _3130_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6763_ net714 _0565_ _3106_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3975_ _0633_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__xnor2_1
X_6694_ _3041_ _3043_ _3040_ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__a21boi_1
X_5714_ sound4.count\[1\] _2186_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5645_ _2116_ _2127_ _2114_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 sound4.count_m\[5\] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8364_ clknet_leaf_76_hwclk rate_clk.next_count\[1\] net76 vssd1 vssd1 vccd1 vccd1
+ rate_clk.count\[1\] sky130_fd_sc_hd__dfrtp_1
X_5576_ _2036_ _2032_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__and2_1
X_7315_ _3482_ _3485_ vssd1 vssd1 vccd1 vccd1 _3486_ sky130_fd_sc_hd__or2_1
Xhold243 sound3.count_m\[11\] vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 sound1.sdiv.Q\[9\] vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ _0969_ _1096_ _1097_ _1000_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__o22a_1
Xhold221 sound2.sdiv.Q\[14\] vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlygate4sd3_1
X_8295_ clknet_leaf_72_hwclk _0395_ net80 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_7246_ net747 _1667_ _3419_ vssd1 vssd1 vccd1 vccd1 _3429_ sky130_fd_sc_hd__mux2_1
Xhold287 sound3.sdiv.Q\[19\] vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ _0969_ _1025_ _1028_ _1005_ _0943_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__o32a_1
Xhold254 sound2.count_m\[16\] vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold265 _0022_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 sound4.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
X_7177_ net227 _3132_ _3389_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__a21o_1
Xhold298 _0014_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__dlygate4sd3_1
X_6128_ _2562_ _2527_ _2528_ _2563_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__o31a_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ _0959_ _0944_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__or2_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _2474_ sound2.divisor_m\[4\] _2476_ _2494_ _2469_ vssd1 vssd1 vccd1 vccd1
+ _2495_ sky130_fd_sc_hd__o221a_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ inputcont.INTERNAL_SYNCED_I\[5\] inputcont.INTERNAL_SYNCED_I\[4\] inputcont.INTERNAL_SYNCED_I\[7\]
+ inputcont.INTERNAL_SYNCED_I\[6\] vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__or4_4
XFILLER_0_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5430_ _1939_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ _0997_ _1792_ _1796_ _1112_ _1871_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__o221a_1
XFILLER_0_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8080_ clknet_leaf_75_hwclk _0222_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7100_ _3351_ _3352_ _3350_ vssd1 vssd1 vccd1 vccd1 _3354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4312_ _0881_ _0882_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__nand2_1
X_5292_ _1053_ _1781_ _1787_ _1802_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_10_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7031_ sound2.divisor_m\[14\] _3283_ _3177_ vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__o21a_1
X_4243_ seq.clk_div.count\[8\] _0824_ seq.clk_div.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _0830_ sky130_fd_sc_hd__a21o_1
X_4174_ net829 _0770_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__nor2_1
X_7933_ clknet_leaf_19_hwclk _0096_ net85 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7864_ clknet_leaf_94_hwclk seq.clk_div.next_count\[21\] net66 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7795_ clknet_leaf_92_hwclk net5 net66 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_6815_ sound2.count\[7\] _2855_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__and2_1
X_6746_ net441 _2895_ sound1.sdiv.next_dived _3095_ vssd1 vssd1 vccd1 vccd1 _0133_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3958_ inputcont.INTERNAL_SYNCED_I\[7\] _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6677_ _2890_ _3034_ _3035_ _2894_ net388 vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__a32o_1
X_3889_ sound2.sdiv.C\[4\] sound2.sdiv.C\[3\] sound2.sdiv.C\[2\] _0558_ sound2.sdiv.C\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__a311oi_4
X_5628_ sound4.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5559_ _2040_ _2041_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8347_ clknet_leaf_87_hwclk sound4.osc.next_count\[5\] net78 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_8278_ clknet_leaf_84_hwclk net424 net80 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_7229_ _3418_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_2__f_hwclk clknet_0_hwclk vssd1 vssd1 vccd1 vccd1 clknet_3_2__leaf_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _1043_ _1339_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4861_ _1405_ _1408_ _1411_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__and3_2
X_6600_ _2960_ vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3812_ _0490_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__clkbuf_4
X_4792_ _1342_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__buf_4
X_7580_ net630 _2005_ vssd1 vssd1 vccd1 vccd1 _3668_ sky130_fd_sc_hd__nor2_1
X_6531_ sound1.divisor_m\[1\] sound1.divisor_m\[0\] _2903_ vssd1 vssd1 vccd1 vccd1
+ _2904_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6462_ _0554_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__buf_6
X_8201_ clknet_leaf_43_hwclk _0322_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_6393_ _2815_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
X_5413_ _1079_ _1842_ _1919_ _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__a211o_2
XFILLER_0_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8132_ clknet_leaf_91_hwclk net387 net69 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_5344_ _0977_ _0996_ _1784_ _1854_ _0960_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__o32a_1
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8063_ clknet_leaf_83_hwclk _0205_ net74 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_5275_ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__buf_4
X_7014_ _3273_ _3276_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__or2_1
X_4226_ net526 _0815_ _0813_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__o21ai_1
X_4157_ _0449_ seq.encode.keys_edge_det\[3\] vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4088_ seq.player_8.state\[0\] seq.player_8.state\[1\] _0712_ vssd1 vssd1 vccd1 vccd1
+ _0715_ sky130_fd_sc_hd__and3_1
X_7916_ clknet_leaf_17_hwclk net252 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7847_ clknet_leaf_97_hwclk seq.clk_div.next_count\[4\] net65 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7778_ clknet_leaf_59_hwclk net676 net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6729_ sound1.sdiv.A\[22\] _3055_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput14 piano_keys[6] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_1
Xhold809 sound1.count\[1\] vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5060_ _1556_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__or2_4
X_4011_ net117 vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ sound1.count_m\[5\] vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7701_ net704 _0556_ _3747_ vssd1 vssd1 vccd1 vccd1 _3749_ sky130_fd_sc_hd__and3_1
X_4913_ _0997_ _1323_ _1343_ _1010_ _1463_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_77_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5893_ _2326_ sound4.divisor_m\[12\] vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4844_ _0985_ _1322_ _1339_ _1181_ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7632_ _3700_ _3701_ net505 _2183_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_62_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7563_ _1903_ vssd1 vssd1 vccd1 vccd1 _3658_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4775_ _0499_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__or2_1
X_6514_ _2889_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7494_ _3437_ _3641_ _3642_ _3440_ net567 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6445_ sound1.count\[10\] _2201_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6376_ _0645_ _2801_ _2802_ _2803_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_15_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_8115_ clknet_leaf_90_hwclk sound2.osc.next_count\[16\] net74 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[16\] sky130_fd_sc_hd__dfrtp_1
X_5327_ _1020_ _1777_ _1792_ _1014_ _1837_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8046_ clknet_leaf_89_hwclk _0188_ net68 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_5258_ _1768_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__buf_4
X_5189_ _1621_ _1719_ _1591_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__o21a_1
X_4209_ seq.clk_div.count\[7\] seq.clk_div.count\[11\] _0802_ seq.clk_div.count\[21\]
+ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4560_ _0992_ _1126_ _1127_ _0990_ _1130_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold617 _3648_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold606 sound3.count\[15\] vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4491_ _0676_ _0685_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nand2_4
Xhold639 sound3.sdiv.C\[5\] vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 sound1.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ sound2.sdiv.Q\[5\] _2295_ _2662_ _2292_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6161_ _2590_ _2595_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ net60 _1077_ _1567_ _1553_ _0946_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__o32a_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ sound3.divisor_m\[13\] _2522_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5043_ _1573_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__clkbuf_4
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6994_ _3255_ _3258_ vssd1 vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__nor2_1
X_5945_ sound1.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5876_ sound4.count_m\[4\] vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7615_ _2110_ _2128_ vssd1 vssd1 vccd1 vccd1 _3689_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4827_ _0983_ _1338_ _1371_ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_105_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4758_ _1310_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7546_ net395 _3403_ _2194_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__a21o_1
X_7477_ _3621_ _3627_ _3622_ vssd1 vssd1 vccd1 vccd1 _3629_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4689_ _1256_ _1257_ _1258_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6428_ sound1.count\[2\] _2201_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__and2_1
Xsass_synth_104 vssd1 vssd1 vccd1 vccd1 sass_synth_104/HI multi[3] sky130_fd_sc_hd__conb_1
X_6359_ net708 _0569_ _2787_ _2788_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8029_ clknet_3_1__leaf_hwclk _0171_ net77 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 seq.encode.inter_keys\[0\] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3991_ net967 _0647_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5730_ net836 _2186_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7400_ _3448_ _3561_ vssd1 vssd1 vccd1 vccd1 _3562_ sky130_fd_sc_hd__and2_1
X_5661_ sound4.divisor_m\[15\] _2143_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__xnor2_1
X_4612_ _1182_ _1000_ _1003_ _0985_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__o22a_1
X_5592_ sound4.divisor_m\[10\] _2074_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__xnor2_1
X_7331_ net971 vssd1 vssd1 vccd1 vccd1 _3500_ sky130_fd_sc_hd__inv_2
X_4543_ _0687_ _1001_ _0943_ _0997_ _0939_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o32a_1
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7262_ sound3.divisor_m\[0\] sound3.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3439_ sky130_fd_sc_hd__or2_1
Xhold425 sound4.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold414 sound4.count_m\[10\] vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 _0381_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 seq.player_3.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6213_ _2585_ _2606_ _2646_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__a21oi_1
Xhold469 sound1.sdiv.Q\[4\] vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 sound4.sdiv.C\[1\] vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_1
X_4474_ _1003_ _1039_ _1041_ _0939_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__o221a_1
Xhold447 _0235_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7193_ net549 _3132_ _3397_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__a21o_1
X_6144_ net683 _0569_ _2578_ _2579_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__a22o_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ sound3.count_m\[4\] vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _0698_ _0542_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _3164_ _3242_ _3243_ _3174_ net319 vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5928_ _2362_ _2329_ _2330_ _2363_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5859_ _2276_ _2292_ _2295_ sound2.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7529_ net342 _3654_ _3643_ net375 _3397_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4190_ seq.clk_div.count\[19\] _0782_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__a21oi_1
X_7880_ clknet_3_5__leaf_hwclk net3 net92 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6900_ _3164_ _3172_ _3173_ _3174_ net292 vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6831_ sound2.count\[15\] _2855_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6762_ _2890_ _3105_ _3107_ _2894_ net596 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3974_ _0634_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__xnor2_1
X_6693_ _3048_ _3049_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__nand2_1
X_5713_ net222 _2184_ _2185_ net564 _2187_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5644_ _2120_ _2125_ _2126_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8363_ clknet_leaf_76_hwclk rate_clk.next_count\[0\] net76 vssd1 vssd1 vccd1 vccd1
+ rate_clk.count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7314_ sound3.divisor_m\[6\] _3484_ vssd1 vssd1 vccd1 vccd1 _3485_ sky130_fd_sc_hd__xnor2_1
Xhold200 sound1.count_m\[6\] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold211 _0372_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlygate4sd3_1
X_5575_ sound4.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold244 _0279_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _0151_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__dlygate4sd3_1
X_4526_ _0952_ _0972_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__nor2_2
Xhold222 _0255_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlygate4sd3_1
X_8294_ clknet_leaf_66_hwclk _0394_ net80 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_7245_ _3428_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__clkbuf_1
X_4457_ _0695_ _0946_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__nor2_8
Xhold266 sound2.sdiv.Q\[21\] vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _0185_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 sound2.sdiv.Q\[10\] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 sound3.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 sound1.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__dlygate4sd3_1
X_7176_ net940 _2863_ vssd1 vssd1 vccd1 vccd1 _3389_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6127_ _2523_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__inv_2
X_4388_ _0951_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__buf_8
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _2481_ _2483_ _2475_ sound2.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2494_
+ sky130_fd_sc_hd__o2bb2a_1
X_5009_ sound2.count\[18\] _1539_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__or2_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5360_ _1016_ _1786_ _1781_ _1116_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5291_ _1012_ _1790_ _1798_ _1801_ _1778_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4311_ seq.player_3.state\[0\] seq.player_3.state\[1\] seq.player_3.state\[2\] seq.player_3.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__or4_1
X_7030_ sound2.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__inv_2
X_4242_ seq.clk_div.count\[8\] seq.clk_div.count\[9\] _0824_ vssd1 vssd1 vccd1 vccd1
+ _0829_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4173_ seq.player_1.state\[0\] seq.player_1.state\[1\] _0769_ vssd1 vssd1 vccd1 vccd1
+ _0772_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7932_ clknet_leaf_20_hwclk _0095_ net85 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7863_ clknet_leaf_94_hwclk seq.clk_div.next_count\[20\] net66 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6814_ net399 _2857_ _3121_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__a21o_1
X_7794_ clknet_leaf_71_hwclk net4 net80 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_6745_ _3091_ _3094_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3957_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6676_ _3022_ _3026_ _3033_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__a21o_1
X_3888_ sound2.sdiv.start vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5627_ _2109_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5558_ sound4.sdiv.A\[19\] _2038_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__xnor2_1
X_8346_ clknet_leaf_87_hwclk sound4.osc.next_count\[4\] net78 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4509_ _0956_ _1078_ _1079_ _0992_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8277_ clknet_leaf_72_hwclk net519 net80 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7228_ net781 _1594_ _3142_ vssd1 vssd1 vccd1 vccd1 _3418_ sky130_fd_sc_hd__mux2_1
X_5489_ sound4.count\[12\] sound4.count\[13\] _1973_ sound4.count\[14\] vssd1 vssd1
+ vccd1 vccd1 _1986_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7159_ sound2.sdiv.Q\[15\] _3167_ _3349_ net325 _3122_ vssd1 vssd1 vccd1 vccd1 _0255_
+ sky130_fd_sc_hd__a221o_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4860_ _1317_ _1409_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__and3_1
X_3811_ _0479_ _0478_ _0485_ _0489_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__and4_1
X_6530_ sound1.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4791_ net39 _1330_ _1324_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6461_ net333 _2836_ _2856_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8200_ clknet_leaf_43_hwclk _0321_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6392_ net694 _2814_ _2808_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5412_ _1025_ _1920_ _1922_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__o21ai_1
X_8131_ clknet_leaf_91_hwclk net199 net69 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_5343_ _1780_ _1832_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__nor2_1
X_8062_ clknet_leaf_81_hwclk _0204_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_5274_ _0719_ _0587_ _0672_ _0673_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__or4_1
X_7013_ sound2.divisor_m\[13\] _3275_ vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__xnor2_1
X_4225_ _0817_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_4156_ _0758_ _0757_ net825 _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_3.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4087_ net553 _0712_ _0714_ vssd1 vssd1 vccd1 vccd1 seq.player_8.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_7915_ clknet_leaf_17_hwclk net313 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_7846_ clknet_leaf_97_hwclk seq.clk_div.next_count\[3\] net65 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7777_ clknet_leaf_59_hwclk _0051_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4989_ _1527_ _1528_ _1504_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6728_ _3079_ _3080_ net575 _2895_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_34_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6659_ sound1.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8329_ clknet_leaf_56_hwclk _0429_ net96 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 piano_keys[7] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4010_ net498 _0659_ vssd1 vssd1 vccd1 vccd1 wave.next_state\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_74_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5961_ sound1.count_m\[7\] _2395_ _2396_ sound1.divisor_m\[7\] vssd1 vssd1 vccd1
+ vccd1 _2397_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7700_ _3681_ _3746_ _3748_ _2184_ net586 vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__a32o_1
X_4912_ _1020_ _1347_ _1333_ _0973_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5892_ _2326_ sound4.divisor_m\[12\] _2327_ sound4.divisor_m\[11\] vssd1 vssd1 vccd1
+ vccd1 _2328_ sky130_fd_sc_hd__a22o_1
X_7631_ _2089_ _2134_ _1764_ vssd1 vssd1 vccd1 vccd1 _3701_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4843_ _1026_ _1343_ _1333_ _1174_ _1393_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7562_ _3657_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4774_ _0504_ _1324_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7493_ sound3.sdiv.C\[1\] sound3.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3642_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6513_ net864 _1223_ _2864_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6444_ net251 _2836_ _2847_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6375_ _2796_ net52 vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8114_ clknet_leaf_90_hwclk sound2.osc.next_count\[15\] net69 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[15\] sky130_fd_sc_hd__dfrtp_2
X_5326_ _1158_ _1790_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__or2_1
X_8045_ clknet_leaf_86_hwclk net164 net77 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_5257_ _1765_ _1767_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__or2_1
X_4208_ seq.clk_div.count\[13\] vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__inv_2
X_5188_ _1629_ _1657_ _1692_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4139_ seq.player_4.state\[2\] net480 _0748_ _0749_ _0700_ vssd1 vssd1 vccd1 vccd1
+ seq.player_4.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7829_ clknet_leaf_5_hwclk net883 net71 vssd1 vssd1 vccd1 vccd1 seq.player_2.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold607 pm.current_waveform\[2\] vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4490_ _0939_ _1057_ _1058_ _0958_ _1060_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold618 rate_clk.count\[7\] vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold629 sound2.sdiv.C\[5\] vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__dlygate4sd3_1
X_6160_ _2292_ _2592_ _2593_ _2594_ _2279_ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__o32ai_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5111_ net858 vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _2524_ sound3.divisor_m\[12\] vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__nor2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _1560_ _1568_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__or2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6993_ sound2.divisor_m\[11\] _3257_ vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__xnor2_1
X_5944_ sound1.count_m\[10\] _2378_ _2379_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5875_ _2306_ _2307_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7614_ _3681_ _3687_ _3688_ _2184_ net190 vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4826_ _0676_ _1372_ _1373_ _1375_ _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_118_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7545_ net354 _3403_ _2193_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__a21o_1
X_4757_ _1256_ _1308_ _1309_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7476_ net530 _3463_ sound3.sdiv.next_dived _3628_ vssd1 vssd1 vccd1 vccd1 _0330_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4688_ net969 sound1.count\[1\] vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6427_ net183 _2836_ _2838_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6358_ _2783_ _2786_ _0569_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__a21oi_1
X_5309_ _1010_ _1772_ _1778_ _1819_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__o211a_1
X_6289_ sound2.sdiv.Q\[6\] _0578_ _2718_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__a21o_1
X_8028_ clknet_leaf_82_hwclk net187 net74 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_76_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 inputcont.u1.ff_intermediate\[13\] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3990_ _0647_ _0648_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[2\] sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_14_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _2142_ _2054_ sound4.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4611_ _0959_ _0944_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5591_ _2036_ _2030_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__and2_1
X_7330_ _3437_ _3498_ _3499_ _3440_ net241 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__a32o_1
X_4542_ _1015_ _1062_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nand2_2
XFILLER_0_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold426 sound3.sdiv.A\[24\] vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold404 pm.count\[5\] vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__dlygate4sd3_1
X_7261_ sound3.divisor_m\[0\] sound3.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3438_ sky130_fd_sc_hd__nand2_1
X_4473_ _0958_ _1042_ _1043_ _0967_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__o22a_1
Xhold415 _0377_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _2605_ _2600_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__and2b_1
Xhold459 _0433_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 sound2.sdiv.Q\[8\] vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 seq.player_5.state\[3\] vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7192_ net349 _2863_ vssd1 vssd1 vccd1 vccd1 _3397_ sky130_fd_sc_hd__and2_1
X_6143_ _2311_ _2577_ _0569_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _2508_ sound3.divisor_m\[4\] _2509_ sound3.divisor_m\[3\] vssd1 vssd1 vccd1
+ vccd1 _2510_ sky130_fd_sc_hd__a22o_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _1555_ _1546_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__or2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6976_ _3233_ _3237_ _3240_ _3241_ vssd1 vssd1 vccd1 vccd1 _3243_ sky130_fd_sc_hd__a211o_1
X_5927_ _2325_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5858_ sound2.sdiv.next_start _2279_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5789_ net941 _2224_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__nand2_1
X_4809_ _1354_ _1356_ _1359_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__and3_2
X_7528_ net375 _3654_ _3643_ net433 _3396_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7459_ sound3.sdiv.A\[20\] sound3.sdiv.A\[19\] _3595_ vssd1 vssd1 vccd1 vccd1 _3614_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6830_ net435 _2857_ _3129_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__a21o_1
X_6761_ _3106_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5712_ sound4.count\[0\] _2186_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__and2_1
X_3973_ inputcont.INTERNAL_SYNCED_I\[11\] _0635_ _0619_ vssd1 vssd1 vccd1 vccd1 _0636_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6692_ _3045_ _3047_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__nand2_1
X_5643_ _2117_ _2119_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8362_ clknet_leaf_46_hwclk wave.next_state\[1\] net100 vssd1 vssd1 vccd1 vccd1 wave.mode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5574_ sound4.sdiv.A\[13\] _2056_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__xnor2_1
X_7313_ _3448_ _3483_ vssd1 vssd1 vccd1 vccd1 _3484_ sky130_fd_sc_hd__and2_1
X_4525_ _0983_ _0978_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__or2_2
Xhold201 sound4.sdiv.Q\[22\] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 sound1.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlygate4sd3_1
X_8293_ clknet_leaf_66_hwclk _0393_ net81 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[7\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold234 sound2.sdiv.Q\[17\] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 sound2.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7244_ net746 _3427_ _3419_ vssd1 vssd1 vccd1 vccd1 _3428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold245 sound3.count\[10\] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 sound1.sdiv.Q\[18\] vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _0964_ _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nand2_2
Xhold278 sound2.sdiv.Q\[16\] vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 sound4.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__dlygate4sd3_1
X_7175_ net179 _3132_ _3388_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__a21o_1
Xhold289 _0144_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__dlygate4sd3_1
X_4387_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__buf_4
X_6126_ _2533_ _2561_ _2526_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__a21oi_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _2467_ _2492_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__and2_1
X_5008_ _1541_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6959_ _3215_ _3219_ _3226_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold790 sound4.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5290_ _1151_ _1769_ _1800_ _0983_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4310_ select1.sequencer_on _0880_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4241_ _0828_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_4172_ net648 _0769_ _0771_ vssd1 vssd1 vccd1 vccd1 seq.player_1.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_7931_ clknet_leaf_12_hwclk _0094_ net85 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7862_ clknet_leaf_95_hwclk net857 net68 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_7793_ clknet_leaf_23_hwclk net17 net89 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6813_ net813 _2855_ vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6744_ _3092_ _3093_ vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3956_ _0611_ _0618_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6675_ _3022_ _3026_ _3033_ vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__nand3_1
XFILLER_0_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3887_ _0556_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__inv_2
X_5626_ _2107_ _2108_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5557_ sound4.sdiv.A\[20\] _2038_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__xnor2_1
X_8345_ clknet_leaf_62_hwclk sound4.osc.next_count\[3\] net78 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[3\] sky130_fd_sc_hd__dfrtp_2
X_4508_ _0970_ _0869_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nand2_4
XFILLER_0_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8276_ clknet_leaf_65_hwclk _0376_ net80 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_5488_ _1984_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__inv_2
X_7227_ _3417_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__clkbuf_1
X_4439_ _0685_ _0681_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__nand2_8
X_7158_ net325 _3167_ _3349_ net379 _3121_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__a221o_1
X_6109_ sound3.count_m\[16\] vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__inv_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _3342_ _3344_ net656 _3168_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_96_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ inputcont.INTERNAL_SYNCED_I\[6\] _0443_ _0463_ inputcont.INTERNAL_SYNCED_I\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__o31ai_2
X_4790_ _1340_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6460_ sound1.count\[17\] _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6391_ _2590_ _2616_ _2805_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5411_ _1245_ _1800_ _1796_ _1110_ _1921_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5342_ _1096_ _1786_ _1794_ _1097_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8130_ clknet_leaf_90_hwclk _0251_ net69 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_8061_ clknet_leaf_80_hwclk _0203_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_7012_ _3177_ _3274_ vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__and2_1
X_5273_ _1783_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__buf_4
X_4224_ _0815_ net936 _0813_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__and3b_1
X_4155_ net824 seq.player_3.state\[2\] _0754_ net539 vssd1 vssd1 vccd1 vccd1 _0760_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4086_ seq.player_8.state\[1\] seq.player_8.state\[2\] seq.player_8.state\[3\] _0713_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a311o_1
X_7914_ clknet_leaf_19_hwclk _0077_ net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7845_ clknet_leaf_97_hwclk seq.clk_div.next_count\[2\] net64 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_7776_ clknet_leaf_53_hwclk net622 net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4988_ sound2.count\[10\] _1524_ net887 vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6727_ _3078_ _3076_ _3077_ _0866_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3939_ _0587_ _0597_ _0596_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__and3_1
X_6658_ _2890_ _3017_ _3018_ _2894_ net418 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5609_ _2091_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__inv_2
X_6589_ sound1.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__inv_2
X_8328_ clknet_leaf_56_hwclk _0428_ net96 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_8259_ clknet_leaf_30_hwclk _0359_ net91 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 piano_keys[8] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5960_ sound1.count_m\[6\] vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__inv_2
X_4911_ _1017_ _1321_ _1341_ _1016_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__o22a_1
X_5891_ sound4.count_m\[10\] vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7630_ _2089_ _2134_ vssd1 vssd1 vccd1 vccd1 _3700_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4842_ _0996_ _1321_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7561_ net879 _3656_ _3419_ vssd1 vssd1 vccd1 vccd1 _3657_ sky130_fd_sc_hd__mux2_1
X_4773_ _0698_ _0507_ net41 vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__or3_2
X_7492_ net567 sound3.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6512_ _2888_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6443_ sound1.count\[9\] _2201_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6374_ _0569_ _2794_ vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8113_ clknet_leaf_91_hwclk sound2.osc.next_count\[14\] net69 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[14\] sky130_fd_sc_hd__dfrtp_1
X_5325_ _1028_ _1800_ _1794_ _1083_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8044_ clknet_leaf_86_hwclk net478 net77 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_5256_ _0673_ _1766_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__nand2_1
X_4207_ _0796_ _0797_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__o21ai_1
X_5187_ sound3.count\[11\] _1699_ _1707_ _1716_ _1717_ vssd1 vssd1 vccd1 vccd1 _1718_
+ sky130_fd_sc_hd__a2111o_1
X_4138_ net909 _0746_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__nor2_1
X_4069_ seq.beat\[0\] seq.beat\[2\] seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7828_ clknet_leaf_4_hwclk net776 net71 vssd1 vssd1 vccd1 vccd1 seq.player_2.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7759_ clknet_leaf_51_hwclk _0044_ net101 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold608 sound2.count\[9\] vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold619 sound2.count\[12\] vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6090_ _2524_ sound3.divisor_m\[12\] _2525_ sound3.divisor_m\[11\] vssd1 vssd1 vccd1
+ vccd1 _2526_ sky130_fd_sc_hd__a22o_1
X_5110_ _0688_ _1559_ _1578_ _1014_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__o221a_2
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _1571_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__buf_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6992_ _3177_ _3256_ vssd1 vssd1 vccd1 vccd1 _3257_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5943_ sound1.divisor_m\[10\] sound1.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2379_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5874_ wave_comb.u1.next_start _2309_ _2310_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7613_ _2116_ _2127_ vssd1 vssd1 vccd1 vccd1 _3688_ sky130_fd_sc_hd__nand2_1
X_4825_ _0677_ _1038_ _1336_ _1339_ _1026_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__o32a_1
XFILLER_0_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7544_ net314 _3403_ _2192_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__a21o_1
X_4756_ net968 _1305_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nand2_1
X_7475_ _3623_ _3627_ vssd1 vssd1 vccd1 vccd1 _3628_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4687_ sound1.count\[0\] sound1.count\[1\] vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6426_ sound1.count\[1\] _2201_ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6357_ _2783_ _2786_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__or2_1
X_5308_ _1773_ _1777_ _1055_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__a21o_1
X_6288_ sound2.sdiv.Q\[6\] _2718_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__nand2_1
X_5239_ _1753_ _1754_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[15\] sky130_fd_sc_hd__nor2_1
X_8027_ clknet_leaf_86_hwclk _0169_ net77 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 inputcont.u1.ff_intermediate\[5\] vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4610_ _0952_ _1004_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5590_ _2070_ _2072_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__nand2_1
X_4541_ _1015_ _1111_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__nand2_4
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold427 wave.mode\[0\] vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 _0653_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__dlygate4sd3_1
X_7260_ _1545_ vssd1 vssd1 vccd1 vccd1 _3437_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4472_ _0679_ _0944_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold416 sound2.sdiv.A\[24\] vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7191_ net501 _3132_ _3396_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__a21o_1
X_6211_ _2638_ _2644_ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__xnor2_1
Xhold449 seq.player_8.state\[0\] vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 seq.player_5.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__dlygate4sd3_1
X_6142_ _2311_ _2577_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__or2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ sound3.count_m\[2\] vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__inv_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _0698_ _0546_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__nor2_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _3240_ _3241_ _3233_ _3237_ vssd1 vssd1 vccd1 vccd1 _3242_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_76_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5926_ _2335_ _2361_ _2328_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5857_ _2277_ _2292_ _2293_ sound1.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5788_ wave_comb.u1.A\[5\] _2224_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4808_ _1242_ _1321_ _1327_ _1101_ _1358_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7527_ sound3.sdiv.Q\[16\] _3654_ _3643_ net134 _3395_ vssd1 vssd1 vccd1 vccd1 _0355_
+ sky130_fd_sc_hd__a221o_1
X_4739_ sound1.count\[13\] sound1.count\[14\] _1290_ vssd1 vssd1 vccd1 vccd1 _1296_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7458_ sound3.sdiv.A\[20\] _3595_ _3607_ vssd1 vssd1 vccd1 vccd1 _3613_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6409_ _2826_ vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__inv_2
X_7389_ sound3.divisor_m\[13\] _3543_ vssd1 vssd1 vccd1 vccd1 _3552_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6760_ sound1.sdiv.C\[2\] sound1.sdiv.C\[1\] sound1.sdiv.C\[0\] vssd1 vssd1 vccd1
+ vccd1 _3106_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5711_ _0575_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__clkbuf_8
X_3972_ _0617_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6691_ _3045_ _3047_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5642_ sound4.divisor_m\[0\] sound4.sdiv.Q\[27\] _2123_ _2124_ vssd1 vssd1 vccd1
+ vccd1 _2125_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_5_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8361_ clknet_leaf_44_hwclk wave.next_state\[0\] net100 vssd1 vssd1 vccd1 vccd1 wave.mode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5573_ sound4.divisor_m\[14\] _2055_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__xnor2_1
X_7312_ sound3.divisor_m\[5\] sound3.divisor_m\[4\] _3465_ vssd1 vssd1 vccd1 vccd1
+ _3483_ sky130_fd_sc_hd__or3_1
X_4524_ _0685_ _0677_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nand2_4
XFILLER_0_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold202 _0023_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold213 sound1.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 sound4.sdiv.Q\[10\] vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd3_1
X_8292_ clknet_leaf_64_hwclk _0392_ net78 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[6\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold235 _0258_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlygate4sd3_1
X_7243_ _1681_ vssd1 vssd1 vccd1 vccd1 _3427_ sky130_fd_sc_hd__inv_2
Xhold268 _0159_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 sound1.sdiv.Q\[22\] vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ _0695_ _0677_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__nand2_4
Xhold246 sound4.sdiv.Q\[17\] vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7174_ net911 _2863_ vssd1 vssd1 vccd1 vccd1 _3388_ sky130_fd_sc_hd__and2_1
X_4386_ _0909_ _0956_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__or2_1
Xhold279 sound4.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6125_ _2534_ _2535_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__nor2_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _2465_ _2466_ _2462_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__a21o_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5007_ _1539_ _1540_ _1504_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__and3b_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6958_ _3215_ _3219_ _3226_ vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__nand3_1
XFILLER_0_119_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5909_ _2315_ sound4.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_75_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_6889_ sound2.divisor_m\[0\] sound2.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_hwclk
+ sky130_fd_sc_hd__clkbuf_16
Xhold791 inputcont.u1.ff_intermediate\[12\] vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold780 sound4.divisor_m\[10\] vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _0813_ _0826_ _0827_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4171_ net829 seq.player_1.state\[2\] seq.player_1.state\[3\] _0770_ _0700_ vssd1
+ vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__a311o_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7930_ clknet_leaf_12_hwclk _0093_ net87 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_7861_ clknet_leaf_95_hwclk seq.clk_div.next_count\[18\] net68 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6812_ net264 _2857_ _3120_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__a21o_1
X_7792_ clknet_leaf_49_hwclk net16 net102 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6743_ sound1.sdiv.A\[24\] _3055_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3955_ _0611_ _0618_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__nor2_1
X_6674_ _3031_ _3032_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3886_ sound4.sdiv.C\[4\] sound4.sdiv.C\[3\] sound4.sdiv.C\[2\] _0555_ net812 vssd1
+ vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5625_ _2104_ _2106_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5556_ net810 _2038_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__nand2_1
X_8344_ clknet_leaf_62_hwclk sound4.osc.next_count\[2\] net79 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4507_ _0695_ _0680_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nand2_2
X_8275_ clknet_leaf_65_hwclk _0375_ net77 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_5487_ sound4.count\[13\] sound4.count\[14\] _1977_ vssd1 vssd1 vccd1 vccd1 _1984_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_130_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7226_ net741 _3416_ _3142_ vssd1 vssd1 vccd1 vccd1 _3417_ sky130_fd_sc_hd__mux2_1
X_4438_ sound1.count\[1\] _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ _0699_ net34 _0917_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__a21bo_2
X_7157_ net379 _3167_ _3349_ net386 _3120_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__a221o_1
X_6108_ sound3.count_m\[17\] _2543_ sound3.count_m\[18\] vssd1 vssd1 vccd1 vccd1 _2544_
+ sky130_fd_sc_hd__a21o_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _1311_ _3343_ vssd1 vssd1 vccd1 vccd1 _3344_ sky130_fd_sc_hd__nand2_1
X_6039_ sound2.count_m\[2\] vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6390_ _2813_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
X_5410_ _1101_ _1786_ _1790_ _1240_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5341_ _1830_ _1831_ _1841_ _1851_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8060_ clknet_leaf_81_hwclk _0202_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7011_ sound2.divisor_m\[12\] sound2.divisor_m\[11\] _3256_ vssd1 vssd1 vccd1 vccd1
+ _3274_ sky130_fd_sc_hd__or3_1
X_5272_ _1782_ _1770_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__or2_1
X_4223_ net935 seq.clk_div.count\[0\] seq.clk_div.count\[2\] seq.clk_div.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4154_ net891 _0757_ _0759_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_3.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4085_ seq.player_8.state\[0\] _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__and2_1
X_7913_ clknet_leaf_13_hwclk _0076_ net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_7844_ clknet_leaf_97_hwclk net558 net64 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_7775_ clknet_leaf_52_hwclk _0049_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6726_ _3076_ _3077_ _3078_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4987_ sound2.count\[10\] sound2.count\[11\] _1524_ vssd1 vssd1 vccd1 vccd1 _1527_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3938_ _0599_ _0602_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nor2_1
X_6657_ _3005_ _3008_ _3016_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3869_ _0520_ _0541_ _0512_ _0532_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__a211oi_4
X_6588_ _2954_ _2955_ net454 _2895_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5608_ sound4.divisor_m\[7\] _2090_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__xnor2_1
X_5539_ _0657_ pm.current_waveform\[7\] _2008_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_
+ sky130_fd_sc_hd__o22a_1
X_8327_ clknet_leaf_55_hwclk _0427_ net96 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8258_ clknet_leaf_31_hwclk net343 net91 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_8189_ clknet_leaf_42_hwclk _0310_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_7209_ sound3.count\[18\] _2863_ vssd1 vssd1 vccd1 vccd1 _3406_ sky130_fd_sc_hd__and2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 piano_keys[9] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4910_ sound2.count\[18\] _1445_ _1448_ _1455_ _1460_ vssd1 vssd1 vccd1 vccd1 _1461_
+ sky130_fd_sc_hd__a2111o_1
X_5890_ sound4.count_m\[11\] vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4841_ _1176_ _1323_ _1338_ _1028_ _1391_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7560_ _1931_ vssd1 vssd1 vccd1 vccd1 _3656_ sky130_fd_sc_hd__inv_2
X_4772_ _0504_ _1320_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__nand2_8
X_7491_ _3640_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6511_ net946 _1225_ _2864_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6442_ net312 _2836_ _2846_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6373_ net698 net127 _0571_ vssd1 vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__mux2_1
X_8112_ clknet_leaf_91_hwclk sound2.osc.next_count\[13\] net67 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5324_ _1004_ _1784_ _1786_ _1189_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__o22a_1
X_8043_ clknet_leaf_82_hwclk net359 net74 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_5255_ _0699_ net46 vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__and2_1
X_4206_ _0782_ _0798_ _0799_ seq.clk_div.count\[21\] seq.clk_div.count\[20\] vssd1
+ vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5186_ sound3.count\[3\] _1641_ _1681_ sound3.count\[12\] vssd1 vssd1 vccd1 vccd1
+ _1717_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_98_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ seq.player_4.state\[0\] seq.player_4.state\[1\] _0745_ vssd1 vssd1 vccd1 vccd1
+ _0748_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ _0703_ _0705_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__nor2_2
X_7827_ clknet_leaf_4_hwclk net459 net71 vssd1 vssd1 vccd1 vccd1 seq.player_2.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7758_ clknet_leaf_51_hwclk _0043_ net101 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6709_ _3050_ _3058_ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__or2_1
X_7689_ _3681_ _3740_ _3741_ _2184_ net282 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold609 sound2.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ net42 _1548_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__or2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6991_ sound2.divisor_m\[10\] _3245_ vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__or2_1
X_5942_ sound1.divisor_m\[11\] vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__inv_2
X_5873_ wave_comb.u1.Q\[1\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__and3_1
X_7612_ _2116_ _2127_ vssd1 vssd1 vccd1 vccd1 _3687_ sky130_fd_sc_hd__or2_1
X_4824_ _1053_ _1341_ _1345_ _1063_ _1374_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4755_ sound1.count\[18\] _1305_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7543_ net302 _3403_ _2191_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7474_ _3607_ _3618_ _3625_ _3626_ vssd1 vssd1 vccd1 vccd1 _3627_ sky130_fd_sc_hd__a31o_1
X_4686_ net472 _1256_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6425_ net310 _2836_ _2837_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6356_ _2784_ _2745_ _2785_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__a21o_1
X_5307_ sound4.count\[14\] _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__xnor2_1
X_8026_ clknet_leaf_11_hwclk net152 net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_6287_ sound2.sdiv.Q\[5\] _2660_ _2686_ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__a21o_1
X_5238_ net710 _1750_ _1721_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__o21ai_1
X_5169_ _1154_ _1550_ _1570_ _1077_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__o22a_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6 seq.encode.inter_keys\[10\] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4540_ _0685_ _0970_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__nand2_4
XFILLER_0_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold406 pm.next_count\[5\] vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold417 wave_comb.u1.A\[0\] vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__dlygate4sd3_1
X_4471_ _0944_ _0947_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 _0660_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__dlygate4sd3_1
X_7190_ sound3.count\[9\] _2863_ vssd1 vssd1 vccd1 vccd1 _3396_ sky130_fd_sc_hd__and2_1
Xhold439 sound1.count_m\[2\] vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _2639_ _2279_ _2292_ _2643_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6141_ _2575_ _2576_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ sound3.count_m\[3\] vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__inv_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _0977_ _0996_ _1550_ _1553_ _1096_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__o32a_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6974_ sound2.sdiv.A\[8\] _3239_ vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _2336_ _2337_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5856_ sound1.sdiv.next_start _2279_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4807_ _1110_ _1336_ _1345_ _1238_ _1357_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__o221a_1
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5787_ wave_comb.u1.next_dived _2235_ _2236_ _0573_ net515 vssd1 vssd1 vccd1 vccd1
+ _0033_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7526_ net134 _3654_ _3643_ net165 _3394_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__a221o_1
X_4738_ _1295_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7457_ sound3.sdiv.A\[21\] _3595_ vssd1 vssd1 vccd1 vccd1 _3612_ sky130_fd_sc_hd__xnor2_1
X_4669_ _0683_ _0959_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__or2_2
X_6408_ _2755_ _2790_ _2805_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7388_ sound3.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _3551_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6339_ _2767_ _2768_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8009_ clknet_leaf_11_hwclk net337 net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5__f_hwclk clknet_0_hwclk vssd1 vssd1 vccd1 vccd1 clknet_3_5__leaf_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3971_ inputcont.INTERNAL_SYNCED_I\[4\] _0512_ _0615_ _0502_ vssd1 vssd1 vccd1 vccd1
+ _0634_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5710_ _1764_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__buf_6
X_6690_ sound1.divisor_m\[18\] _3046_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5641_ _2122_ sound4.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8360_ clknet_leaf_61_hwclk sound4.osc.next_count\[18\] net94 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5572_ sound4.sdiv.A\[26\] _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7311_ sound3.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _3482_ sky130_fd_sc_hd__inv_2
X_4523_ _0996_ _1090_ _1091_ _1092_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o2111a_1
X_8291_ clknet_leaf_66_hwclk _0391_ net81 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7242_ _3426_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
Xhold225 sound4.count_m\[1\] vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 sound2.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold214 sound4.sdiv.Q\[19\] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold236 sound1.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _0164_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__buf_6
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold269 sound2.count_m\[4\] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _0017_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__dlygate4sd3_1
X_7173_ net533 _3132_ _3387_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__a21o_1
X_4385_ _0940_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__nand2_1
X_6124_ _2559_ _2515_ _2548_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__a21o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _2447_ _2490_ _2454_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__a21o_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ sound2.count\[15\] sound2.count\[16\] _1533_ sound2.count\[17\] vssd1 vssd1
+ vccd1 vccd1 _1540_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_9_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6957_ _3224_ _3225_ vssd1 vssd1 vccd1 vccd1 _3226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6888_ _1311_ vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__buf_6
X_5908_ _2325_ _2328_ _2339_ _2343_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5839_ net536 _0579_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7509_ _3634_ _3639_ _3652_ _0563_ _2005_ vssd1 vssd1 vccd1 vccd1 _3653_ sky130_fd_sc_hd__a311o_1
XFILLER_0_91_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold770 sound1.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 seq.player_8.state\[1\] vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 sound1.count\[6\] vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4170_ seq.player_1.state\[0\] _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__and2_1
X_7860_ clknet_leaf_96_hwclk seq.clk_div.next_count\[17\] net68 vssd1 vssd1 vccd1
+ vccd1 seq.clk_div.count\[17\] sky130_fd_sc_hd__dfrtp_1
X_6811_ sound2.count\[5\] _2855_ vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7791_ clknet_leaf_74_hwclk net108 net76 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_OCTAVE_INPUT
+ sky130_fd_sc_hd__dfrtp_1
X_6742_ sound1.sdiv.A\[24\] _3055_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3954_ inputcont.INTERNAL_SYNCED_I\[11\] _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6673_ _3027_ _3030_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__nand2_1
X_3885_ sound4.sdiv.start vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5624_ _2104_ _2106_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8343_ clknet_leaf_62_hwclk sound4.osc.next_count\[1\] net79 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5555_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4506_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5486_ _1983_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
X_8274_ clknet_leaf_64_hwclk net396 net80 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_7225_ _1635_ vssd1 vssd1 vccd1 vccd1 _3416_ sky130_fd_sc_hd__inv_2
X_4437_ _0962_ _0987_ _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7156_ sound2.sdiv.Q\[12\] _3167_ _3349_ net198 _3119_ vssd1 vssd1 vccd1 vccd1 _0252_
+ sky130_fd_sc_hd__a221o_1
X_6107_ net852 vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__inv_2
X_4368_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__clkbuf_8
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _3339_ _3341_ _3337_ vssd1 vssd1 vccd1 vccd1 _3343_ sky130_fd_sc_hd__a21o_1
X_4299_ seq.beat\[1\] seq.beat\[0\] seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nor3_1
X_6038_ sound2.count_m\[3\] vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7989_ clknet_leaf_16_hwclk sound1.osc.next_count\[10\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[10\] sky130_fd_sc_hd__dfrtp_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5340_ sound4.count\[3\] _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5271_ _1766_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7010_ sound2.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__inv_2
X_4222_ seq.clk_div.count\[2\] seq.clk_div.count\[3\] _0777_ vssd1 vssd1 vccd1 vccd1
+ _0815_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_74_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4153_ net763 _0756_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4084_ seq.encode.keys_edge_det\[9\] inputcont.INTERNAL_SYNCED_I\[7\] vssd1 vssd1
+ vccd1 vccd1 _0712_ sky130_fd_sc_hd__and2b_1
X_7912_ clknet_leaf_13_hwclk net225 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_89_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7843_ clknet_leaf_97_hwclk seq.clk_div.next_count\[0\] net64 vssd1 vssd1 vccd1 vccd1
+ seq.clk_div.count\[0\] sky130_fd_sc_hd__dfrtp_1
X_7774_ clknet_leaf_52_hwclk _0048_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4986_ net378 _1524_ _1526_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[10\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6725_ sound1.sdiv.A\[21\] _3055_ vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_12_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_3937_ _0600_ _0590_ _0601_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6656_ _3005_ _3008_ _3016_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__nand3_1
X_3868_ _0521_ _0523_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_27_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_6587_ _2946_ _2953_ _0866_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__a21o_1
X_5607_ _2036_ _2028_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__and2_1
X_3799_ inputcont.INTERNAL_SYNCED_I\[4\] _0443_ inputcont.INTERNAL_SYNCED_I\[5\] vssd1
+ vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__o21ai_4
X_5538_ _2007_ pm.current_waveform\[6\] _2010_ _2021_ vssd1 vssd1 vccd1 vccd1 _2022_
+ sky130_fd_sc_hd__o22a_1
X_8326_ clknet_leaf_56_hwclk _0426_ net96 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_8257_ clknet_leaf_31_hwclk _0357_ net90 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7208_ net410 _3403_ _3405_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__a21o_1
X_5469_ sound4.count\[10\] _1966_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__nand2_1
X_8188_ clknet_leaf_43_hwclk _0309_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_7139_ _3383_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 seq_play vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4840_ _1180_ _1327_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6510_ _2887_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4771_ _0499_ _1316_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__nand2_4
X_7490_ _1545_ _0577_ net778 vssd1 vssd1 vccd1 vccd1 _3640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6441_ net886 _2201_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6372_ _0645_ _2798_ _2799_ net668 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8111_ clknet_leaf_91_hwclk sound2.osc.next_count\[12\] net67 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5323_ net46 _1129_ _1770_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__or3_1
X_8042_ clknet_leaf_81_hwclk net287 net73 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_5254_ _0698_ _0606_ net48 vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__or3_2
X_5185_ _1642_ _1649_ _1714_ sound3.count\[9\] _1715_ vssd1 vssd1 vccd1 vccd1 _1716_
+ sky130_fd_sc_hd__o221ai_1
X_4205_ seq.clk_div.count\[11\] seq.clk_div.count\[19\] vssd1 vssd1 vccd1 vccd1 _0799_
+ sky130_fd_sc_hd__nand2_1
X_4136_ net637 _0745_ _0747_ vssd1 vssd1 vccd1 vccd1 seq.player_4.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_4067_ seq.beat\[1\] seq.beat\[0\] seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__or3b_4
Xwire53 _2797_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7826_ clknet_leaf_5_hwclk net640 net71 vssd1 vssd1 vccd1 vccd1 seq.player_2.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7757_ clknet_leaf_53_hwclk _0042_ net101 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4969_ sound2.count\[4\] sound2.count\[5\] _1511_ vssd1 vssd1 vccd1 vccd1 _1515_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_19_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6708_ _3050_ _3061_ _3058_ _3062_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__o31a_1
X_7688_ _2173_ _2174_ _3739_ vssd1 vssd1 vccd1 vccd1 _3741_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6639_ sound1.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8309_ clknet_leaf_68_hwclk _0409_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6990_ sound2.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__inv_2
X_5941_ sound1.count_m\[14\] _2375_ sound1.count_m\[13\] _2376_ vssd1 vssd1 vccd1
+ vccd1 _2377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5872_ net486 _2308_ _0645_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7611_ _3681_ _3685_ _3686_ _2184_ net321 vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__a32o_1
X_4823_ _1057_ _1343_ _1333_ _1056_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4754_ _1307_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7542_ net260 _3403_ _2190_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7473_ sound3.sdiv.A\[22\] sound3.sdiv.A\[21\] sound3.sdiv.A\[20\] sound3.sdiv.A\[19\]
+ _3595_ vssd1 vssd1 vccd1 vccd1 _3626_ sky130_fd_sc_hd__o41a_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4685_ _1173_ _1255_ _1070_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__o21a_4
XFILLER_0_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6424_ sound1.count\[0\] _2201_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__and2_1
X_6355_ _2740_ _2742_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6286_ sound2.sdiv.Q\[7\] _0578_ _2286_ vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__and3_1
X_5306_ _1062_ _1777_ _1813_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__o211a_1
X_5237_ net845 _1750_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__and2_1
X_8025_ clknet_leaf_14_hwclk net216 net88 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_5168_ _1043_ _1559_ _1580_ _1033_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__o221a_2
X_5099_ _1180_ _1553_ _1565_ _1174_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__o22a_1
X_4119_ net842 net760 _0730_ net768 vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7809_ clknet_leaf_0_hwclk net850 net64 vssd1 vssd1 vccd1 vccd1 seq.player_7.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7 seq.encode.keys_sync\[0\] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold407 sound3.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 _0028_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__dlygate4sd3_1
X_4470_ _1019_ net59 vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__nor2_8
Xhold429 sound3.count_m\[0\] vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6140_ _2291_ _2305_ _2303_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _2505_ _2506_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__xnor2_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ net42 _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__nand2_4
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6973_ sound2.sdiv.A\[8\] _3239_ vssd1 vssd1 vccd1 vccd1 _3240_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5924_ _2347_ _2359_ _2317_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__a21o_1
X_5855_ net29 net30 vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__nand2_8
XFILLER_0_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4806_ _1004_ _1133_ _1339_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5786_ _2228_ _2233_ _2234_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7525_ net165 _3654_ _3643_ net248 _3393_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__a221o_1
X_4737_ _1256_ _1293_ _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7456_ net665 _3463_ sound3.sdiv.next_dived _3611_ vssd1 vssd1 vccd1 vccd1 _0327_
+ sky130_fd_sc_hd__a22o_1
X_4668_ _1004_ _1003_ _1028_ _1238_ _1000_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__o32a_1
XFILLER_0_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6407_ _2825_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkbuf_1
X_7387_ _3437_ _3549_ _3550_ _3440_ net218 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4599_ _1070_ _1161_ _1163_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__and4_2
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6338_ sound3.sdiv.Q\[7\] _0577_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__nand2_1
X_6269_ sound3.sdiv.Q\[5\] _0577_ _2699_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__a21o_1
X_8008_ clknet_leaf_11_hwclk net440 net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3970_ inputcont.INTERNAL_SYNCED_I\[10\] _0610_ _0608_ vssd1 vssd1 vccd1 vccd1 _0633_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5640_ sound4.sdiv.A\[0\] _2122_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5571_ sound4.divisor_m\[13\] _2032_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__nor2_1
X_7310_ _3437_ _3480_ _3481_ _3440_ net277 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__a32o_1
X_4522_ _0992_ _1003_ _0948_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__a21o_1
X_8290_ clknet_leaf_62_hwclk _0390_ net78 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_7241_ net844 _3425_ _3419_ vssd1 vssd1 vccd1 vccd1 _3426_ sky130_fd_sc_hd__mux2_1
Xhold226 _0368_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _0685_ _0681_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__nor2_1
Xhold204 sound2.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 sound2.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold237 sound3.count_m\[13\] vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 sound3.sdiv.Q\[25\] vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 sound1.sdiv.Q\[21\] vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7172_ net862 _2855_ vssd1 vssd1 vccd1 vccd1 _3387_ sky130_fd_sc_hd__and2_1
X_4384_ _0926_ _0936_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__nor2b_2
X_6123_ _2558_ _2512_ _2549_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__a21o_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _2449_ _2489_ _2442_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__a21o_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ sound2.count\[16\] sound2.count\[17\] _1536_ vssd1 vssd1 vccd1 vccd1 _1539_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _3220_ _3223_ vssd1 vssd1 vccd1 vccd1 _3225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5907_ _2340_ sound4.divisor_m\[16\] sound4.divisor_m\[9\] _2334_ _2342_ vssd1 vssd1
+ vccd1 vccd1 _2343_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6887_ _2843_ _1445_ _3163_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__o21ai_1
X_5838_ sound2.sdiv.Q\[0\] _0578_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5769_ _2219_ _2215_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7508_ sound3.divisor_m\[18\] sound3.divisor_m\[17\] sound3.sdiv.A\[26\] _3578_ vssd1
+ vssd1 vccd1 vccd1 _3652_ sky130_fd_sc_hd__or4_1
XFILLER_0_106_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7439_ _3590_ _3592_ _3589_ vssd1 vssd1 vccd1 vccd1 _3597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold771 sound3.count\[6\] vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 sound1.count\[8\] vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 sound1.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 sound1.divisor_m\[1\] vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6810_ net373 _2857_ _3119_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__a21o_1
X_7790_ clknet_leaf_7_hwclk net444 net71 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6741_ sound1.sdiv.A\[23\] _3055_ _3089_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3953_ _0615_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6672_ _3027_ _3030_ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__or2_1
X_3884_ rate_clk.count\[7\] _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__nand2_8
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5623_ sound4.divisor_m\[4\] _2105_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8342_ clknet_leaf_60_hwclk sound4.osc.next_count\[0\] net94 vssd1 vssd1 vccd1 vccd1
+ sound4.count\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5554_ sound4.divisor_m\[18\] _2035_ _2036_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4505_ _0679_ _1046_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__or2_1
X_5485_ _1779_ _1936_ _1981_ _1982_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__and4_1
X_8273_ clknet_leaf_64_hwclk net355 net81 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_7224_ _3415_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
X_4436_ _0990_ _0978_ _0944_ _0998_ _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__o311a_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4367_ _0909_ _0918_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__or3_1
X_7155_ net198 _3167_ _3349_ net381 _3118_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__a221o_1
X_6106_ _2541_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _3337_ _3339_ _3341_ vssd1 vssd1 vccd1 vccd1 _3342_ sky130_fd_sc_hd__and3_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__clkbuf_8
X_6037_ _2472_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__inv_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7988_ clknet_leaf_15_hwclk sound1.osc.next_count\[9\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[9\] sky130_fd_sc_hd__dfrtp_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6939_ _3197_ _3200_ _3208_ vssd1 vssd1 vccd1 vccd1 _3210_ sky130_fd_sc_hd__or3b_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold590 pm.current_waveform\[3\] vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5270_ _1780_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__clkinv_4
X_4221_ net556 _0777_ _0814_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[2\] sky130_fd_sc_hd__a21oi_1
X_4152_ seq.player_3.state\[2\] net890 vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__nand2_1
X_4083_ _0711_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7911_ clknet_leaf_12_hwclk net298 net84 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_7842_ clknet_leaf_47_hwclk _0065_ net101 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7773_ clknet_leaf_52_hwclk net684 net101 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4985_ net378 _1524_ _1504_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__o21ai_1
X_6724_ sound1.sdiv.A\[20\] sound1.sdiv.A\[19\] _3055_ vssd1 vssd1 vccd1 vccd1 _3077_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3936_ _0473_ _0486_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__nor2_1
X_6655_ _3014_ _3015_ vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__nand2_1
X_3867_ _0540_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__inv_2
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6586_ _2946_ _2953_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3798_ inputcont.INTERNAL_SYNCED_I\[10\] _0445_ _0474_ _0475_ _0476_ vssd1 vssd1
+ vccd1 vccd1 _0477_ sky130_fd_sc_hd__a2111o_1
X_5606_ _2087_ _2088_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__nand2_1
X_5537_ _2009_ pm.current_waveform\[5\] _2011_ _2020_ vssd1 vssd1 vccd1 vccd1 _2021_
+ sky130_fd_sc_hd__o22a_1
X_8325_ clknet_leaf_69_hwclk _0425_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8256_ clknet_leaf_31_hwclk net434 net90 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7207_ sound3.count\[17\] _2863_ vssd1 vssd1 vccd1 vccd1 _3405_ sky130_fd_sc_hd__and2_1
X_5468_ _1969_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_8187_ clknet_leaf_43_hwclk _0308_ net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4419_ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__clkbuf_8
X_5399_ sound4.count\[2\] _1903_ _1909_ sound4.count\[11\] vssd1 vssd1 vccd1 vccd1
+ _1910_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7138_ _2843_ _3382_ vssd1 vssd1 vccd1 vccd1 _3383_ sky130_fd_sc_hd__and2_1
X_7069_ net513 _3168_ sound2.sdiv.next_dived _3326_ vssd1 vssd1 vccd1 vccd1 _0225_
+ sky130_fd_sc_hd__a22o_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 seq_power vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ net39 _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nand2_4
XFILLER_0_99_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6440_ net182 _2836_ _2845_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6371_ wave_comb.u1.Q\[9\] _0573_ _0646_ net667 vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8110_ clknet_leaf_93_hwclk sound2.osc.next_count\[11\] net67 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[11\] sky130_fd_sc_hd__dfrtp_1
X_5322_ _0677_ _1832_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__nand2_1
X_8041_ clknet_leaf_91_hwclk net436 net67 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_5253_ _1764_ vssd1 vssd1 vccd1 vccd1 sound4.sdiv.next_dived sky130_fd_sc_hd__buf_4
X_5184_ sound3.count\[9\] _1714_ _1699_ sound3.count\[11\] vssd1 vssd1 vccd1 vccd1
+ _1715_ sky130_fd_sc_hd__o2bb2a_1
X_4204_ seq.clk_div.count\[3\] seq.clk_div.count\[17\] _0785_ seq.clk_div.count\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__or4bb_1
X_4135_ seq.player_4.state\[1\] seq.player_4.state\[2\] seq.player_4.state\[3\] _0746_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__a311o_1
X_4066_ _0703_ _0704_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__nor2_1
XFILLER_0_64_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire54 _3086_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_1
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7825_ clknet_leaf_3_hwclk net826 net71 vssd1 vssd1 vccd1 vccd1 seq.player_3.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7756_ clknet_leaf_51_hwclk net615 net101 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4968_ net471 _1511_ _1514_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[4\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6707_ _3048_ _3056_ _3057_ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__o21a_1
X_7687_ _2173_ _2174_ _3739_ vssd1 vssd1 vccd1 vccd1 _3740_ sky130_fd_sc_hd__or3_1
X_3919_ _0529_ _0525_ _0549_ _0582_ _0526_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__a41o_1
XFILLER_0_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4899_ _0499_ _1315_ _1319_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__a21oi_1
X_6638_ _2890_ _2999_ _3000_ _2894_ net340 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6569_ _2903_ _2937_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__and2_1
X_8308_ clknet_leaf_67_hwclk _0408_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_8239_ clknet_leaf_46_hwclk _0339_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5940_ sound1.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5871_ _2306_ _2307_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__xnor2_1
X_7610_ _2120_ _2125_ vssd1 vssd1 vccd1 vccd1 _3686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4822_ _1064_ _1347_ _1322_ _0979_ _1317_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__o221a_1
X_4753_ _1305_ _1306_ _1256_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__and3b_1
X_7541_ net177 _3403_ _2189_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7472_ _3624_ _3612_ vssd1 vssd1 vccd1 vccd1 _3625_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6423_ _0554_ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__clkbuf_8
X_4684_ _1187_ _1197_ _1209_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6354_ _2742_ _2740_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__or2b_1
X_6285_ wave_comb.u1.next_start _2714_ _2715_ _2716_ vssd1 vssd1 vccd1 vccd1 _0051_
+ sky130_fd_sc_hd__a31o_1
X_5305_ _1814_ _1815_ _0695_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__a21o_1
X_5236_ _1752_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_8024_ clknet_leaf_13_hwclk net276 net86 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5167_ _1004_ _1693_ _1694_ _1001_ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__o221a_1
X_5098_ sound3.count\[14\] _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__xor2_1
X_4118_ net919 _0733_ _0735_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_6.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
X_4049_ _0682_ _0683_ _0687_ _0689_ _0681_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__o32a_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7808_ clknet_leaf_97_hwclk seq.player_7.next_state\[2\] net65 vssd1 vssd1 vccd1
+ vccd1 seq.player_7.state\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7739_ clknet_leaf_60_hwclk net828 net94 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 inputcont.u1.ff_intermediate\[6\] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold408 sound4.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold419 sound3.count\[7\] vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _2281_ _2299_ _2297_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__a21o_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _0542_ _1551_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__nor2_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6972_ sound2.divisor_m\[9\] _3238_ vssd1 vssd1 vccd1 vccd1 _3239_ sky130_fd_sc_hd__xnor2_1
X_5923_ _2314_ _2358_ _2319_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5854_ _2181_ _2289_ _2290_ sound4.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4805_ _1025_ _1323_ _1338_ _1240_ _1355_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7524_ sound3.sdiv.Q\[13\] _3654_ _3643_ net172 _3392_ vssd1 vssd1 vccd1 vccd1 _0352_
+ sky130_fd_sc_hd__a221o_1
X_5785_ _2228_ _2233_ _2234_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4736_ sound1.count\[13\] _1290_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__or2_1
X_7455_ _3609_ _3610_ vssd1 vssd1 vccd1 vccd1 _3611_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4667_ _0681_ _0944_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nor2_1
X_7386_ _3537_ _3541_ _3548_ vssd1 vssd1 vccd1 vccd1 _3550_ sky130_fd_sc_hd__nand3_1
X_6406_ net707 _2824_ _2808_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6337_ sound3.sdiv.Q\[6\] _2632_ _2731_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4598_ _1003_ _1164_ _1165_ _0943_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__o221a_1
X_6268_ sound3.sdiv.Q\[5\] _2699_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6199_ sound3.sdiv.Q\[2\] _2632_ _2602_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__a21o_1
X_5219_ net674 _1738_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__and2_1
X_8007_ clknet_leaf_11_hwclk net193 net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5570_ _2050_ _2052_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__nor2_1
X_4521_ _0993_ _0943_ _1012_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold205 sound3.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
X_7240_ _1699_ vssd1 vssd1 vccd1 vccd1 _3425_ sky130_fd_sc_hd__inv_2
Xhold216 sound3.count_m\[7\] vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ _1011_ _0967_ _1003_ _1014_ _1022_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__o221a_1
Xhold238 sound3.sdiv.Q\[18\] vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _0365_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 sound1.count_m\[14\] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4383_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7171_ sound2.sdiv.Q\[27\] _3168_ _3164_ net155 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__a22o_1
X_6122_ _2553_ _2557_ _2510_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _2452_ _2488_ _2451_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__a21bo_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ net394 _1536_ _1538_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[16\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6955_ _3220_ _3223_ vssd1 vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5906_ sound4.count_m\[15\] _2341_ sound4.count_m\[14\] _2331_ vssd1 vssd1 vccd1
+ vccd1 _2342_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6886_ _2470_ _2005_ vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__or2_1
X_5837_ net280 _0577_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5768_ net593 _0573_ wave_comb.u1.next_dived _2220_ vssd1 vssd1 vccd1 vccd1 _0030_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7507_ _3651_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__clkbuf_1
X_4719_ sound1.count\[9\] _1278_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__and2_1
X_7438_ sound3.sdiv.A\[18\] _3595_ vssd1 vssd1 vccd1 vccd1 _3596_ sky130_fd_sc_hd__xnor2_1
X_5699_ _1763_ _2180_ _2181_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7369_ sound3.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _3534_ sky130_fd_sc_hd__inv_2
Xhold750 sound3.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 wave_comb.u1.C\[3\] vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold772 sound2.divisor_m\[4\] vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 sound4.sdiv.C\[4\] vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold783 sound2.count\[11\] vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6740_ net583 _2895_ _3088_ _3090_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__a22o_1
X_3952_ _0612_ _0614_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__and2_1
X_6671_ sound1.divisor_m\[16\] _3029_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3883_ net966 _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__and2_2
XFILLER_0_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5622_ _2036_ _2026_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__nand2_1
X_8341_ clknet_leaf_57_hwclk sound4.sdiv.next_start net96 vssd1 vssd1 vccd1 vccd1
+ sound4.sdiv.start sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5553_ sound4.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4504_ _0688_ _0958_ _0943_ _0971_ _1074_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8272_ clknet_leaf_64_hwclk net315 net81 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5484_ sound4.count\[13\] _1977_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7223_ net866 _3414_ _3142_ vssd1 vssd1 vccd1 vccd1 _3415_ sky130_fd_sc_hd__mux2_1
X_4435_ _1000_ _1001_ _1003_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o22a_1
X_4366_ _0926_ _0936_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7154_ sound2.sdiv.Q\[10\] _3167_ _3349_ net136 _3117_ vssd1 vssd1 vccd1 vccd1 _0250_
+ sky130_fd_sc_hd__a221o_1
X_6105_ _2523_ _2526_ _2537_ _2540_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _3321_ _3330_ _3331_ _3340_ vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__o211a_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _0674_ _0677_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__or2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ sound2.count_m\[17\] _2470_ sound2.count_m\[16\] _2471_ vssd1 vssd1 vccd1
+ vccd1 _2472_ sky130_fd_sc_hd__o22a_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7987_ clknet_leaf_15_hwclk sound1.osc.next_count\[8\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[8\] sky130_fd_sc_hd__dfrtp_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _3197_ _3200_ _3208_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__o21bai_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6869_ _1488_ vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold580 _0047_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 wave_comb.u1.Q\[2\] vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4220_ net556 _0777_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o21ai_1
X_4151_ seq.player_3.state\[2\] net539 _0756_ _0757_ _0700_ vssd1 vssd1 vccd1 vccd1
+ seq.player_3.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_4082_ net1 pm.pwm_o vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7910_ clknet_leaf_12_hwclk net528 net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_7841_ clknet_leaf_47_hwclk _0064_ net101 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_7772_ clknet_leaf_51_hwclk net487 net102 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4984_ _1524_ _1525_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[9\] sky130_fd_sc_hd__nor2_1
X_6723_ sound1.sdiv.A\[20\] _3055_ _3069_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3935_ _0547_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__inv_2
X_6654_ _3010_ _3013_ vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3866_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__clkbuf_4
X_5605_ sound4.sdiv.A\[7\] _2086_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__or2_1
X_6585_ _2951_ _2952_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3797_ inputcont.INTERNAL_SYNCED_I\[6\] _0443_ _0463_ inputcont.INTERNAL_SYNCED_I\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__o31a_1
X_5536_ _0651_ pm.current_waveform\[4\] _2013_ _2019_ vssd1 vssd1 vccd1 vccd1 _2020_
+ sky130_fd_sc_hd__o22a_1
X_8324_ clknet_leaf_69_hwclk _0424_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_8255_ clknet_leaf_31_hwclk net135 net90 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_5467_ _1779_ _1936_ _1967_ _1968_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__and4_1
X_7206_ net202 _3403_ _3404_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4418_ _0926_ _0936_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__or3_1
X_8186_ clknet_leaf_44_hwclk net231 net99 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5398_ _1035_ _1769_ _1792_ _1041_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__o221a_2
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7137_ net705 _0559_ _3378_ net942 vssd1 vssd1 vccd1 vccd1 _3382_ sky130_fd_sc_hd__a31o_1
X_4349_ seq.player_6.state\[2\] _0894_ _0896_ _0919_ vssd1 vssd1 vccd1 vccd1 _0920_
+ sky130_fd_sc_hd__a22o_1
X_7068_ _3323_ _3325_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__xnor2_1
X_6019_ sound2.count_m\[8\] sound2.divisor_m\[9\] vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__or2b_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6370_ _2794_ net53 _2796_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5321_ _1782_ _1771_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8040_ clknet_leaf_92_hwclk net483 net67 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_5252_ _1763_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__inv_2
X_5183_ _1709_ _1711_ _1713_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__and3_2
X_4203_ seq.clk_div.count\[20\] _0664_ _0665_ seq.clk_div.count\[21\] vssd1 vssd1
+ vccd1 vccd1 _0797_ sky130_fd_sc_hd__o22a_1
X_4134_ seq.player_4.state\[0\] _0745_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__and2_1
X_4065_ seq.beat\[0\] seq.beat\[2\] seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__or3b_4
Xwire55 _0537_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
X_7824_ clknet_leaf_3_hwclk seq.player_3.next_state\[2\] net71 vssd1 vssd1 vccd1 vccd1
+ seq.player_3.state\[2\] sky130_fd_sc_hd__dfrtp_2
X_7755_ clknet_leaf_51_hwclk net589 net101 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ net471 _1511_ _1504_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__o21ai_1
X_6706_ _3031_ _3040_ _3041_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__a21bo_1
X_7686_ sound4.sdiv.A\[24\] _2038_ vssd1 vssd1 vccd1 vccd1 _3739_ sky130_fd_sc_hd__xor2_1
X_3918_ _0549_ _0582_ _0529_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__a21o_1
X_4898_ _1333_ _1325_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6637_ _2987_ _2991_ _2998_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__o21bai_2
X_3849_ _0488_ _0491_ _0441_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__a211oi_4
X_6568_ sound1.divisor_m\[5\] sound1.divisor_m\[4\] _2919_ vssd1 vssd1 vccd1 vccd1
+ _2937_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8307_ clknet_leaf_68_hwclk net322 net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5519_ _0553_ _2004_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6499_ _2880_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8238_ clknet_leaf_58_hwclk sound4.sdiv.next_dived net95 vssd1 vssd1 vccd1 vccd1
+ sound4.sdiv.dived sky130_fd_sc_hd__dfrtp_1
X_8169_ clknet_leaf_30_hwclk _0290_ net91 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[3\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_7_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5870_ _2181_ _2286_ _2284_ _2283_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4821_ _0944_ _1327_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4752_ sound1.count\[15\] sound1.count\[16\] _1296_ net959 vssd1 vssd1 vccd1 vccd1
+ _1306_ sky130_fd_sc_hd__a31o_1
X_7540_ net329 _3403_ _2188_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7471_ _3609_ vssd1 vssd1 vccd1 vccd1 _3624_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4683_ _1228_ _1236_ _1251_ _1253_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__or4b_1
XFILLER_0_70_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6422_ net716 _2834_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6353_ _2779_ _2782_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6284_ net675 _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__and3_1
X_5304_ _0680_ _1784_ _1792_ _0684_ _1800_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__o221a_1
X_5235_ _1750_ _1751_ _1721_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__and3b_1
X_8023_ clknet_leaf_15_hwclk net279 net86 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5166_ _1041_ _1567_ _1565_ _1129_ _1696_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__o221a_1
X_5097_ _1624_ _1627_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__nand2_2
X_4117_ net611 _0732_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__xor2_1
X_4048_ _0691_ vssd1 vssd1 vccd1 vccd1 oct.next_state\[0\] sky130_fd_sc_hd__clkbuf_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5999_ net666 vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7807_ clknet_leaf_100_hwclk net497 net64 vssd1 vssd1 vccd1 vccd1 seq.player_7.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_7738_ clknet_leaf_64_hwclk net306 net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7669_ _2168_ _2041_ vssd1 vssd1 vccd1 vccd1 _3727_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold9 inputcont.u1.ff_intermediate\[14\] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 sound2.sdiv.A\[18\] vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _0698_ _0546_ net45 vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__or3_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6971_ _2460_ _3230_ sound2.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _3238_ sky130_fd_sc_hd__a21o_1
X_5922_ _2313_ sound4.divisor_m\[4\] _2348_ _2357_ _2320_ vssd1 vssd1 vccd1 vccd1
+ _2358_ sky130_fd_sc_hd__a221o_1
X_5853_ sound4.sdiv.next_start _2279_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5784_ net954 _2224_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__xnor2_1
X_4804_ _1004_ _1028_ _1322_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7523_ net172 _3654_ _3643_ net204 _3391_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__a221o_1
X_4735_ sound1.count\[13\] _1290_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7454_ sound3.sdiv.A\[19\] _3595_ _3607_ vssd1 vssd1 vccd1 vccd1 _3610_ sky130_fd_sc_hd__a21oi_1
X_4666_ net896 vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__inv_2
X_7385_ _3537_ _3541_ _3548_ vssd1 vssd1 vccd1 vccd1 _3549_ sky130_fd_sc_hd__a21o_1
X_6405_ _2725_ _2748_ _2805_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__mux2_1
X_4597_ _0990_ _0997_ _0992_ _1166_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6336_ _2764_ _2765_ vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6267_ sound3.sdiv.Q\[4\] _2632_ _2669_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__a21o_1
X_6198_ sound3.sdiv.next_start _2570_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__nor2_1
X_5218_ _1740_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_8006_ clknet_leaf_36_hwclk _0148_ net93 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_72_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5149_ _1101_ _1553_ _1678_ _1679_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_87_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4520_ _0976_ _0994_ _0960_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold206 sound1.count_m\[0\] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _0979_ _0958_ _0992_ _1016_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__o221a_1
Xhold217 sound4.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold239 _0358_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _0084_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7170_ net155 _3167_ _1311_ net271 _3134_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6121_ _2518_ _2520_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__nand2_1
X_4382_ _0951_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__or2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ sound2.count_m\[10\] _2443_ _2455_ _2456_ _2444_ vssd1 vssd1 vccd1 vccd1 _2488_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ net394 _1536_ _1504_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__o21ai_1
X_6954_ sound2.divisor_m\[7\] _3222_ vssd1 vssd1 vccd1 vccd1 _3223_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5905_ net867 vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6885_ _3162_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5836_ net486 _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5767_ _2215_ _2219_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7506_ net743 _0554_ vssd1 vssd1 vccd1 vccd1 _3651_ sky130_fd_sc_hd__and2_1
X_4718_ _1280_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_5698_ net963 _0576_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__and2_2
X_7437_ _3594_ vssd1 vssd1 vccd1 vccd1 _3595_ sky130_fd_sc_hd__buf_6
X_4649_ sound1.count\[15\] _1215_ _1219_ sound1.count\[16\] vssd1 vssd1 vccd1 vccd1
+ _1220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7368_ _3532_ _3533_ net469 _3463_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__a2bb2o_1
Xhold740 sound3.divisor_m\[11\] vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold762 sound3.divisor_m\[4\] vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 seq.clk_div.count\[18\] vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 seq.player_5.state\[3\] vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7299_ _3458_ _3461_ _3470_ vssd1 vssd1 vccd1 vccd1 _3472_ sky130_fd_sc_hd__or3b_1
Xhold784 sound1.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__dlygate4sd3_1
X_6319_ sound1.sdiv.Q\[6\] _2656_ _2722_ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__a21o_1
Xhold795 sound2.count\[0\] vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _0612_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__nor2_1
X_6670_ _2903_ _3028_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__and2_1
X_3882_ rate_clk.count\[5\] net129 _0551_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__and3_1
X_5621_ sound4.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__inv_2
X_8340_ clknet_leaf_53_hwclk _0440_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.M\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5552_ sound4.divisor_m\[17\] _2034_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4503_ _1015_ _0981_ _0969_ _0946_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__o22a_1
X_8271_ clknet_leaf_64_hwclk net303 net81 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5483_ sound4.count\[13\] _1977_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7222_ _1601_ vssd1 vssd1 vccd1 vccd1 _3414_ sky130_fd_sc_hd__inv_2
X_4434_ _0944_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__nor2_2
X_4365_ _0699_ net37 _0934_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7153_ net136 _3174_ _3349_ net552 _3116_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__a221o_1
X_6104_ _2538_ sound3.divisor_m\[16\] sound3.divisor_m\[9\] _2532_ _2539_ vssd1 vssd1
+ vccd1 vccd1 _2540_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7084_ _3323_ _3330_ _3331_ _3324_ vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__or4bb_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _0867_ vssd1 vssd1 vccd1 vccd1 sound1.sdiv.next_dived sky130_fd_sc_hd__buf_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ sound2.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__inv_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7986_ clknet_leaf_15_hwclk sound1.osc.next_count\[7\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[7\] sky130_fd_sc_hd__dfrtp_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6937_ _3206_ _3207_ vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__nand2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6868_ _3152_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5819_ _0646_ _0573_ net783 vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6799_ net151 _2893_ _0867_ net215 _2858_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold570 sound3.count\[9\] vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 wave_comb.u1.C\[5\] vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4150_ net824 _0754_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__nor2_1
X_4081_ _0710_ vssd1 vssd1 vccd1 vccd1 tempo_select_on sky130_fd_sc_hd__clkbuf_1
X_7840_ clknet_leaf_47_hwclk _0063_ net101 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7771_ clknet_leaf_53_hwclk _0045_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4983_ net712 _1522_ _1504_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6722_ _3074_ _3075_ net672 _2895_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3934_ _0514_ _0533_ _0510_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6653_ _3010_ _3013_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__or2_1
X_3865_ _0534_ _0535_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5604_ sound4.sdiv.A\[7\] _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__nand2_1
X_6584_ _2947_ _2950_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3796_ inputcont.INTERNAL_SYNCED_I\[8\] _0443_ _0444_ inputcont.INTERNAL_SYNCED_I\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__o31a_2
XFILLER_0_42_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5535_ _2012_ pm.current_waveform\[3\] pm.current_waveform\[2\] _2014_ _2018_ vssd1
+ vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__o221a_1
X_8323_ clknet_leaf_69_hwclk _0423_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8254_ clknet_leaf_32_hwclk _0354_ net87 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5466_ sound4.count\[9\] _1962_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7205_ net809 _2863_ vssd1 vssd1 vccd1 vccd1 _3404_ sky130_fd_sc_hd__and2_1
X_4417_ _0909_ _0940_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__or2_2
X_8185_ clknet_leaf_42_hwclk net504 net98 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5397_ _1129_ _1777_ _1905_ _1906_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__o2111a_1
X_4348_ seq.player_7.state\[2\] _0898_ _0901_ seq.player_8.state\[2\] vssd1 vssd1
+ vccd1 vccd1 _0919_ sky130_fd_sc_hd__a22o_1
X_7136_ _2005_ _3380_ net706 vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__nor3_1
X_7067_ _3306_ _3315_ _3324_ vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__a21o_1
X_4279_ _0855_ _0813_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__and3b_1
X_6018_ sound2.count_m\[15\] _2446_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__and2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7969_ clknet_leaf_23_hwclk _0132_ net103 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5320_ sound4.count\[8\] _1829_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__nor2_1
X_5251_ _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__buf_2
X_4202_ seq.clk_div.count\[7\] vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__inv_2
X_5182_ _1189_ _1553_ _1580_ _1028_ _1712_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__o221a_1
X_4133_ _0607_ seq.encode.keys_edge_det\[5\] vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__nor2_1
X_4064_ _0701_ _0703_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__nor2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7823_ clknet_leaf_3_hwclk net540 net70 vssd1 vssd1 vccd1 vccd1 seq.player_3.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_7754_ clknet_leaf_51_hwclk _0039_ net101 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6705_ net663 _2895_ sound1.sdiv.next_dived _3060_ vssd1 vssd1 vccd1 vccd1 _0127_
+ sky130_fd_sc_hd__a22o_1
X_4966_ _1513_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7685_ _1763_ _2174_ _3737_ _3738_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_61_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3917_ _0510_ _0513_ _0533_ _0530_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__o31a_2
X_4897_ sound2.count\[18\] _1445_ _1447_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6636_ _2987_ _2991_ _2998_ vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__or3b_1
X_3848_ inputcont.INTERNAL_SYNCED_I\[9\] _0454_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6567_ sound1.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3779_ inputcont.INTERNAL_SYNCED_I\[10\] _0445_ inputcont.INTERNAL_SYNCED_I\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__or3b_1
X_8306_ clknet_leaf_56_hwclk _0406_ net96 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5518_ net447 _0552_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6498_ net737 _2879_ _2864_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__mux2_1
X_8237_ clknet_leaf_36_hwclk sound3.osc.next_count\[18\] net93 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[18\] sky130_fd_sc_hd__dfrtp_1
X_5449_ _1954_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
X_8168_ clknet_leaf_42_hwclk _0289_ net98 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_7119_ net584 _3168_ sound2.sdiv.next_dived _3369_ vssd1 vssd1 vccd1 vccd1 _0232_
+ sky130_fd_sc_hd__a22o_1
X_8099_ clknet_leaf_89_hwclk sound2.osc.next_count\[0\] net69 vssd1 vssd1 vccd1 vccd1
+ sound2.count\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_97_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4820_ _0679_ net59 _1321_ _1323_ _1059_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__o32a_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ sound1.count\[16\] sound1.count\[17\] _1299_ vssd1 vssd1 vccd1 vccd1 _1305_
+ sky130_fd_sc_hd__and3_1
X_7470_ _3621_ _3622_ vssd1 vssd1 vccd1 vccd1 _3623_ sky130_fd_sc_hd__nand2_1
X_4682_ _1073_ _1089_ _1104_ sound1.count\[0\] _1252_ vssd1 vssd1 vccd1 vccd1 _1253_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6421_ _2835_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6352_ _2780_ _2739_ _2781_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6283_ net697 _0645_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__or2_1
X_5303_ _1769_ _1781_ _0687_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__a21o_1
X_5234_ sound3.count\[12\] sound3.count\[13\] _1744_ sound3.count\[14\] vssd1 vssd1
+ vccd1 vccd1 _1751_ sky130_fd_sc_hd__a31o_1
X_8022_ clknet_leaf_17_hwclk net362 net83 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_5165_ _0947_ _1611_ _1695_ _1035_ _1562_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__o32a_1
X_4116_ net918 seq.player_6.state\[3\] vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5096_ _1095_ _1550_ _1626_ _0695_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4047_ _0679_ _0690_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7806_ clknet_leaf_0_hwclk net902 net64 vssd1 vssd1 vccd1 vccd1 seq.player_7.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5998_ _2394_ _2404_ _2422_ _2433_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__a31o_2
XFILLER_0_93_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4949_ _1497_ _1499_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__nand2_1
X_7737_ clknet_leaf_64_hwclk net369 net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7668_ net631 _2183_ _3681_ _3726_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6619_ sound1.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7599_ net894 _0554_ vssd1 vssd1 vccd1 vccd1 _3679_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6970_ _3164_ _3236_ _3237_ _3174_ net221 vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _2351_ _2353_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5852_ _2288_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5783_ _2229_ _2231_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__or2b_1
X_4803_ _1245_ _1341_ _1343_ _0985_ _1353_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__o221a_1
X_7522_ net204 _3654_ _3643_ net258 _3390_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4734_ _1292_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7453_ sound3.sdiv.A\[20\] _3595_ vssd1 vssd1 vccd1 vccd1 _3609_ sky130_fd_sc_hd__xor2_2
X_4665_ sound1.count\[14\] _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7384_ _3546_ _3547_ vssd1 vssd1 vccd1 vccd1 _3548_ sky130_fd_sc_hd__nand2_1
X_6404_ _2823_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_6_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_4596_ _0994_ _1126_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6335_ _2728_ _2729_ _2726_ vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6266_ _2696_ _2697_ vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__xor2_1
X_8005_ clknet_leaf_38_hwclk _0147_ net93 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6197_ _2619_ _2630_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__xnor2_2
X_5217_ _1738_ _1739_ _1721_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__and3b_1
X_5148_ _1240_ _1578_ _1550_ _1242_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__o22a_1
X_5079_ _1562_ _1548_ _0869_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold207 _0070_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
X_4450_ _0950_ _1017_ _1020_ _0994_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold229 sound1.count_m\[17\] vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 _0407_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlygate4sd3_1
X_4381_ _0674_ _0684_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__nor2_8
X_6120_ _2520_ _2542_ _2550_ _2555_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__or4b_1
XFILLER_0_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _2473_ _2476_ _2477_ _2486_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__nor4_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _1536_ _1537_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[15\] sky130_fd_sc_hd__nor2_1
X_6953_ _3177_ _3221_ vssd1 vssd1 vccd1 vccd1 _3222_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6884_ net796 _1446_ _3142_ vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__mux2_1
X_5904_ sound4.count_m\[15\] vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__inv_2
X_5835_ net577 _2224_ _2261_ _2272_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5766_ _2216_ _2218_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7505_ _3650_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__clkbuf_1
X_4717_ _1278_ _1279_ _1256_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__and3b_1
X_5697_ sound4.divisor_m\[18\] sound4.sdiv.A\[26\] _2035_ _2039_ _2179_ vssd1 vssd1
+ vccd1 vccd1 _2180_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7436_ sound3.divisor_m\[18\] sound3.divisor_m\[17\] _3578_ _3448_ vssd1 vssd1 vccd1
+ vccd1 _3594_ sky130_fd_sc_hd__o31a_1
X_4648_ _0688_ _1216_ _1070_ _1217_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_4_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold730 _0744_ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__dlygate4sd3_1
X_7367_ _3518_ _3524_ _3531_ _0563_ _2005_ vssd1 vssd1 vccd1 vccd1 _3533_ sky130_fd_sc_hd__a311o_1
Xhold741 sound3.count\[15\] vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
X_4579_ _0680_ _0959_ _0958_ _1149_ _1070_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__o311a_1
Xhold752 _0858_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold763 sound4.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__dlygate4sd3_1
X_7298_ _3458_ _3461_ _3470_ vssd1 vssd1 vccd1 vccd1 _3471_ sky130_fd_sc_hd__o21ba_1
Xhold774 sound1.sdiv.C\[5\] vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6318_ wave_comb.u1.next_start _2747_ _2748_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a21o_1
Xhold796 seq.player_7.state\[1\] vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 sound2.divisor_m\[1\] vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__dlygate4sd3_1
X_6249_ wave_comb.u1.Q\[5\] _0572_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 sound4.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlygate4sd3_1
X_3950_ _0496_ _0613_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3881_ net176 _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5620_ sound4.sdiv.A\[4\] _2102_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_71_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5551_ sound4.divisor_m\[16\] _2033_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__or2_1
X_4502_ net938 vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__inv_2
X_8270_ clknet_leaf_63_hwclk net261 net78 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_7221_ _3413_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__clkbuf_1
X_5482_ _1980_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4433_ _0972_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__buf_6
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4364_ _0698_ seq.player_1.state\[3\] _0871_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__and3_1
X_7152_ net552 _3174_ _3349_ net613 _3115_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__a221o_1
X_6103_ _2538_ sound3.divisor_m\[16\] sound3.count_m\[14\] _2529_ vssd1 vssd1 vccd1
+ vccd1 _2539_ sky130_fd_sc_hd__o2bb2a_1
X_4295_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__inv_6
X_7083_ _3294_ _3298_ _3323_ _3338_ _3332_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ net791 vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__inv_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7985_ clknet_leaf_15_hwclk sound1.osc.next_count\[6\] net86 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[6\] sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_24_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _3203_ _3205_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__nand2_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6867_ net786 _3151_ _3142_ vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5818_ _2261_ _2262_ net606 _0573_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__a2bb2o_1
X_6798_ net215 _2893_ _0867_ net275 _2856_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_hwclk clknet_3_7__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5749_ net839 _2201_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7419_ _3448_ _3578_ vssd1 vssd1 vccd1 vccd1 _3579_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold571 wave_comb.u1.Q\[6\] vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 sound4.sdiv.A\[18\] vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold593 wave_comb.u1.Q\[5\] vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 seq.beat\[0\] vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4080_ net1 net20 vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__and2b_1
X_7770_ clknet_leaf_48_hwclk net652 net102 vssd1 vssd1 vccd1 vccd1 pm.pwm_o sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ net962 sound2.count\[9\] _1520_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6721_ _3067_ _3069_ _3073_ _0866_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3933_ _0595_ _0596_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6652_ _2376_ _3012_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3864_ _0530_ _0536_ net55 _0512_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5603_ _2085_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6583_ _2947_ _2950_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__or2_1
X_8322_ clknet_leaf_69_hwclk _0422_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_3795_ _0443_ _0444_ inputcont.INTERNAL_SYNCED_I\[8\] vssd1 vssd1 vccd1 vccd1 _0474_
+ sky130_fd_sc_hd__o21a_1
X_5534_ pm.next_count\[0\] pm.current_waveform\[0\] _2016_ _2017_ vssd1 vssd1 vccd1
+ vccd1 _2018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8253_ clknet_leaf_34_hwclk _0353_ net88 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5465_ _1966_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8184_ clknet_leaf_40_hwclk _0305_ net98 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4416_ _0964_ _0967_ _0969_ _0973_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__o221a_1
X_7204_ _0554_ vssd1 vssd1 vccd1 vccd1 _3403_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7135_ _0559_ _3378_ net705 vssd1 vssd1 vccd1 vccd1 _3381_ sky130_fd_sc_hd__a21oi_1
X_5396_ _1125_ _1780_ _1800_ _1033_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__o2bb2a_1
X_4347_ _0699_ net34 _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__a21boi_4
X_7066_ _3302_ _3313_ _3314_ vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__o21ba_1
X_4278_ seq.clk_div.count\[18\] _0853_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6017_ _2447_ _2449_ _2451_ _2452_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__and4_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ clknet_leaf_23_hwclk _0131_ net103 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7899_ clknet_leaf_0_hwclk net534 net64 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6919_ _3190_ _3191_ vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold390 seq.clk_div.count\[21\] vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5250_ _0575_ _0557_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__or2_1
X_4201_ _0787_ _0788_ _0790_ _0793_ _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__o32a_1
X_5181_ _1077_ _1562_ _1565_ _1020_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__o22a_1
X_4132_ _0742_ _0741_ net834 _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_5.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_4063_ _0702_ net51 vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__nand2_4
Xwire57 net58 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
X_7822_ clknet_leaf_8_hwclk net916 net70 vssd1 vssd1 vccd1 vccd1 seq.player_3.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7753_ clknet_leaf_53_hwclk _0038_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4965_ _1511_ _1512_ _1504_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__and3b_1
X_6704_ _3058_ _3059_ vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3916_ _0512_ _0533_ _0580_ _0502_ inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1 vccd1
+ vccd1 _0581_ sky130_fd_sc_hd__o311a_1
XFILLER_0_104_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7684_ net555 _2182_ vssd1 vssd1 vccd1 vccd1 _3738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4896_ sound2.count\[17\] _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6635_ _2996_ _2997_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3847_ _0500_ _0491_ _0475_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6566_ _2890_ _2934_ _2935_ _2894_ net335 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ inputcont.INTERNAL_SYNCED_I\[2\] _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8305_ clknet_leaf_58_hwclk _0405_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5517_ _0552_ net130 vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_30_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6497_ _1249_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__inv_2
X_8236_ clknet_leaf_38_hwclk sound3.osc.next_count\[17\] net93 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5448_ _1779_ _1936_ _1952_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__and4_1
X_8167_ clknet_leaf_40_hwclk _0288_ net98 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[1\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout100 net103 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_8
X_5379_ _1775_ _1888_ _1889_ _1774_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__o2bb2a_1
X_8098_ clknet_leaf_60_hwclk sound2.sdiv.next_start net95 vssd1 vssd1 vccd1 vccd1
+ sound2.sdiv.start sky130_fd_sc_hd__dfrtp_1
X_7118_ _3365_ _3368_ vssd1 vssd1 vccd1 vccd1 _3369_ sky130_fd_sc_hd__xnor2_1
X_7049_ sound2.divisor_m\[16\] sound2.divisor_m\[15\] sound2.divisor_m\[14\] _3283_
+ vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__or4_2
XFILLER_0_97_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _1304_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4681_ sound1.count\[12\] _1249_ _1170_ sound1.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _1252_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6420_ _2833_ _2834_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6351_ _2730_ _2734_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5302_ _1058_ _1771_ _1788_ _1111_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__o22a_1
X_6282_ _2712_ _2713_ _0569_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5233_ sound3.count\[13\] sound3.count\[14\] _1747_ vssd1 vssd1 vccd1 vccd1 _1750_
+ sky130_fd_sc_hd__and3_1
X_8021_ clknet_leaf_17_hwclk net364 net83 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5164_ _0540_ _1213_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__nor2_1
X_4115_ net611 seq.player_6.state\[3\] _0732_ _0733_ _0700_ vssd1 vssd1 vccd1 vccd1
+ seq.player_6.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_5095_ net60 _1567_ _1625_ _0687_ _1580_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__o221a_1
X_4046_ _0681_ _0682_ _0683_ net60 _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__o32a_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7805_ clknet_leaf_100_hwclk net861 net64 vssd1 vssd1 vccd1 vccd1 seq.player_8.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _2407_ _2432_ _2412_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4948_ sound2.count\[8\] _1412_ _1469_ _1470_ _1498_ vssd1 vssd1 vccd1 vccd1 _1499_
+ sky130_fd_sc_hd__o221a_1
X_7736_ clknet_leaf_64_hwclk net122 net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7667_ _3725_ _2165_ vssd1 vssd1 vccd1 vccd1 _3726_ sky130_fd_sc_hd__xnor2_1
X_4879_ _0997_ _1343_ _1333_ _1064_ _1429_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__o221a_1
X_6618_ _2890_ _2981_ _2982_ _2894_ net323 vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7598_ _2843_ _1820_ _3678_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__o21ai_1
X_6549_ _2903_ _2919_ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__nand2_1
X_8219_ clknet_leaf_36_hwclk sound3.osc.next_count\[0\] net94 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[0\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5920_ _2323_ net57 _2345_ _2355_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5851_ net29 net30 vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5782_ net582 _0573_ wave_comb.u1.next_dived _2232_ vssd1 vssd1 vccd1 vccd1 _0032_
+ sky130_fd_sc_hd__a22o_1
X_4802_ _1025_ _1038_ _1347_ _1333_ _0954_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__o32a_1
X_7521_ sound3.sdiv.Q\[10\] _3654_ _3643_ net141 _3389_ vssd1 vssd1 vccd1 vccd1 _0349_
+ sky130_fd_sc_hd__a221o_1
X_4733_ _1290_ _1291_ _1256_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7452_ net627 _3463_ sound3.sdiv.next_dived _3608_ vssd1 vssd1 vccd1 vccd1 _0326_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6403_ net719 _2822_ _2808_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__mux2_1
X_4664_ _0958_ _1112_ _1231_ _1234_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7383_ _3542_ _3545_ vssd1 vssd1 vccd1 vccd1 _3547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4595_ _1107_ _0996_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6334_ _2762_ _2763_ vssd1 vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__or2_1
X_6265_ _2665_ _2667_ _2664_ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8004_ clknet_leaf_38_hwclk net574 net93 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_5216_ sound3.count\[6\] sound3.count\[7\] _1732_ sound3.count\[8\] vssd1 vssd1 vccd1
+ vccd1 _1739_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6196_ _2628_ _2629_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__and2b_1
X_5147_ _1038_ _1562_ _1625_ _1025_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__a211o_1
X_5078_ sound3.count\[16\] _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__xnor2_1
X_4029_ _0606_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__inv_2
XFILLER_0_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7719_ clknet_leaf_58_hwclk _0004_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 sound1.count_m\[8\] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold219 sound1.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__dlygate4sd3_1
X_4380_ _0686_ _0675_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ sound2.count_m\[2\] _2478_ _2479_ _2483_ _2485_ vssd1 vssd1 vccd1 vccd1 _2486_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_56_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ net687 _1533_ _1504_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6952_ sound2.divisor_m\[6\] _3212_ vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6883_ _3161_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
X_5903_ _2329_ _2330_ _2332_ _2338_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__or4_1
X_5834_ wave_comb.u1.M\[0\] wave_comb.u1.M\[1\] wave_comb.u1.M\[2\] wave_comb.u1.A\[10\]
+ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__nor4_1
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5765_ wave_comb.u1.M\[2\] _2217_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7504_ _2843_ _3649_ vssd1 vssd1 vccd1 vccd1 _3650_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4716_ sound1.count\[6\] sound1.count\[7\] _1269_ net886 vssd1 vssd1 vccd1 vccd1
+ _1279_ sky130_fd_sc_hd__a31o_1
X_5696_ _2175_ _2176_ _2178_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7435_ net680 _3463_ sound3.sdiv.next_dived _3593_ vssd1 vssd1 vccd1 vccd1 _0324_
+ sky130_fd_sc_hd__a22o_1
X_4647_ _0974_ _1210_ _1010_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__a21o_1
X_7366_ _3518_ _3524_ _3531_ vssd1 vssd1 vccd1 vccd1 _3532_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold720 seq.player_3.state\[1\] vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__dlygate4sd3_1
X_6317_ wave_comb.u1.Q\[7\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__and3_1
X_4578_ _0943_ _1012_ _1127_ _0969_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold742 seq.tempo_select.state\[0\] vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 seq.clk_div.next_count\[19\] vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 sound2.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 seq.player_5.next_state\[3\] vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7297_ _3468_ _3469_ vssd1 vssd1 vccd1 vccd1 _3470_ sky130_fd_sc_hd__or2_1
Xhold775 sound4.divisor_m\[1\] vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 seq.player_3.state\[3\] vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _0723_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__dlygate4sd3_1
X_6248_ net621 _2680_ _0645_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__mux2_1
X_6179_ _2610_ _2612_ _0569_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold91 sound3.count_m\[14\] vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 _0071_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3880_ net821 net185 net167 vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5550_ sound4.divisor_m\[15\] sound4.divisor_m\[14\] sound4.divisor_m\[13\] _2032_
+ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__or4_1
X_4501_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__inv_2
X_5481_ _1779_ _1936_ _1978_ _1979_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7220_ net751 _3412_ _3142_ vssd1 vssd1 vccd1 vccd1 _3413_ sky130_fd_sc_hd__mux2_1
X_4432_ _1002_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__buf_4
XFILLER_0_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7151_ net613 _3168_ _3164_ net636 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__a22o_1
X_4363_ seq.player_2.state\[3\] _0878_ _0932_ _0933_ _0873_ vssd1 vssd1 vccd1 vccd1
+ _0934_ sky130_fd_sc_hd__o221a_1
X_6102_ sound3.count_m\[15\] vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__inv_2
X_4294_ _0865_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__clkbuf_8
X_7082_ _3304_ _3313_ _3314_ vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__or3_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _2462_ _2465_ _2466_ _2468_ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__and4bb_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7984_ clknet_leaf_15_hwclk sound1.osc.next_count\[5\] net86 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6935_ _3203_ _3205_ vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6866_ _1387_ vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5817_ _2254_ _2260_ _2259_ _0573_ _0645_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__a311o_1
X_6797_ net275 _2893_ _0867_ net278 _2854_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5748_ net214 _2182_ _2185_ net256 _2205_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5679_ _2159_ _2161_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__nor2_1
X_7418_ sound3.divisor_m\[16\] sound3.divisor_m\[15\] _3561_ vssd1 vssd1 vccd1 vccd1
+ _3578_ sky130_fd_sc_hd__or3_2
Xhold561 sound3.sdiv.A\[21\] vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__dlygate4sd3_1
X_7349_ _3448_ _3515_ vssd1 vssd1 vccd1 vccd1 _3516_ sky130_fd_sc_hd__and2_1
Xhold572 _0052_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 sound4.sdiv.A\[22\] vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 wave_comb.u1.Q\[9\] vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 sound2.count\[15\] vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _1522_ _1523_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[8\] sky130_fd_sc_hd__nor2_1
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6720_ _3067_ _3069_ _3073_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _0545_ _0543_ _0582_ _0489_ _0508_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a311o_1
XFILLER_0_46_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6651_ _2903_ _3011_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__nand2_1
X_3863_ _0500_ _0491_ _0519_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__nor3_1
XFILLER_0_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6582_ sound1.divisor_m\[7\] _2949_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5602_ sound4.divisor_m\[8\] _2084_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__xnor2_1
X_5533_ _2014_ pm.current_waveform\[2\] pm.current_waveform\[1\] _2015_ vssd1 vssd1
+ vccd1 vccd1 _2017_ sky130_fd_sc_hd__a22o_1
X_8321_ clknet_leaf_69_hwclk _0421_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3794_ inputcont.INTERNAL_SYNCED_I\[11\] _0461_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8252_ clknet_leaf_34_hwclk net173 net88 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_5464_ sound4.count\[9\] _1962_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7203_ net212 _3132_ _3402_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__a21o_1
X_8183_ clknet_leaf_36_hwclk _0304_ net94 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4415_ _0976_ _0979_ _0981_ _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5395_ net46 net59 _1788_ _0947_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4346_ _0698_ _0916_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand2_1
X_7134_ net705 _0559_ _3378_ vssd1 vssd1 vccd1 vccd1 _3380_ sky130_fd_sc_hd__and3_1
X_7065_ _3321_ _3322_ vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__nand2_1
X_4277_ seq.clk_div.count\[17\] net855 _0850_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__and3_1
X_6016_ _2450_ sound2.divisor_m\[12\] sound2.count_m\[10\] _2443_ vssd1 vssd1 vccd1
+ vccd1 _2452_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7967_ clknet_leaf_22_hwclk _0130_ net103 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6918_ _3183_ _3181_ _3189_ vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__a21oi_1
X_7898_ clknet_leaf_2_hwclk net452 net70 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6849_ net876 _1441_ _2864_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold380 sound4.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold391 net837 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_70_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_85_hwclk clknet_3_3__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_4200_ seq.tempo_select.state\[0\] seq.clk_div.count\[4\] seq.clk_div.count\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__or3b_1
X_5180_ _1193_ _1559_ _1572_ _1129_ _1710_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__o221a_1
X_4131_ net833 seq.player_5.state\[2\] _0738_ net541 vssd1 vssd1 vccd1 vccd1 _0744_
+ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_38_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_4062_ seq.beat\[3\] vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire58 _2344_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_7821_ clknet_leaf_3_hwclk net907 net70 vssd1 vssd1 vccd1 vccd1 seq.player_4.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_7752_ clknet_leaf_53_hwclk _0037_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ net984 _1508_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__or2_1
X_6703_ _3050_ _3051_ _3048_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__o21ai_1
X_3915_ _0510_ _0514_ _0533_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__nor3_1
X_7683_ _2173_ _2172_ _2169_ _2170_ _2171_ vssd1 vssd1 vccd1 vccd1 _3737_ sky130_fd_sc_hd__o2111a_1
X_4895_ _1018_ _1314_ _1316_ _0971_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6634_ _2993_ _2995_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3846_ _0515_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nor2_2
X_6565_ _2932_ _2933_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__nand2_1
X_3777_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1
+ vccd1 vccd1 _0459_ sky130_fd_sc_hd__or2_1
X_6496_ _2878_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__clkbuf_1
X_8304_ clknet_leaf_63_hwclk _0404_ net78 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_5516_ net129 _0551_ rate_clk.count\[5\] vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__a21oi_1
X_8235_ clknet_leaf_37_hwclk sound3.osc.next_count\[16\] net93 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[16\] sky130_fd_sc_hd__dfrtp_2
X_5447_ sound4.count\[3\] sound4.count\[4\] _1940_ sound4.count\[5\] vssd1 vssd1 vccd1
+ vccd1 _1953_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout101 net102 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_6
X_8166_ clknet_leaf_36_hwclk _0287_ net94 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_5378_ _0688_ _1771_ _1773_ _1138_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7117_ _3366_ _3367_ vssd1 vssd1 vccd1 vccd1 _3368_ sky130_fd_sc_hd__and2b_1
X_4329_ seq.beat\[3\] seq.encode.play _0884_ inputcont.INTERNAL_SYNCED_I\[7\] vssd1
+ vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__a31oi_1
X_8097_ clknet_leaf_72_hwclk _0239_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_7048_ net449 _3168_ sound2.sdiv.next_dived _3307_ vssd1 vssd1 vccd1 vccd1 _0223_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4680_ _1237_ _1071_ _1157_ sound1.count\[10\] _1250_ vssd1 vssd1 vccd1 vccd1 _1251_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6350_ _2730_ _2734_ vssd1 vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__nand2_1
X_5301_ sound4.count\[5\] _1810_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6281_ _2684_ _2711_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5232_ net427 _1747_ _1749_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[13\] sky130_fd_sc_hd__a21oi_1
X_8020_ clknet_leaf_17_hwclk net357 net83 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5163_ _1046_ _1572_ _1550_ _0996_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__o22a_1
X_4114_ net842 _0730_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__nor2_1
X_5094_ _1562_ _1572_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__and2_1
X_4045_ _0682_ _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7804_ clknet_leaf_100_hwclk seq.player_8.next_state\[2\] net64 vssd1 vssd1 vccd1
+ vccd1 seq.player_8.state\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _2426_ _2431_ _2414_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4947_ sound2.count\[11\] _1488_ _1495_ sound2.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _1498_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7735_ clknet_leaf_84_hwclk _0020_ net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7666_ _2158_ _2163_ _2162_ vssd1 vssd1 vccd1 vccd1 _3725_ sky130_fd_sc_hd__a21o_1
X_4878_ _1116_ _1347_ _1345_ _1113_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__o22a_1
X_6617_ _2970_ _2980_ _2976_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3829_ _0479_ _0478_ _0480_ _0483_ _0502_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__a41o_1
XFILLER_0_61_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7597_ _2341_ _2005_ vssd1 vssd1 vccd1 vccd1 _3678_ sky130_fd_sc_hd__or2_1
X_6548_ sound1.divisor_m\[3\] sound1.divisor_m\[2\] sound1.divisor_m\[1\] sound1.divisor_m\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6479_ _2868_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8218_ clknet_leaf_46_hwclk sound3.sdiv.next_start net100 vssd1 vssd1 vccd1 vccd1
+ sound3.sdiv.start sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8149_ clknet_leaf_37_hwclk _0270_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5850_ wave_comb.u1.next_dived _2273_ _2274_ _2287_ vssd1 vssd1 vccd1 vccd1 _0045_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5781_ _2229_ _2231_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4801_ _1329_ _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__nand2_1
X_7520_ net141 _3654_ _3643_ net416 _3388_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__a221o_1
X_4732_ sound1.count\[12\] _1287_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7451_ _3606_ _3607_ vssd1 vssd1 vccd1 vccd1 _3608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4663_ _0990_ _1062_ _1232_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6402_ _2693_ _2716_ _2805_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7382_ _3542_ _3545_ vssd1 vssd1 vccd1 vccd1 _3546_ sky130_fd_sc_hd__or2_1
X_4594_ _0952_ _1019_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nor2_2
X_6333_ _2755_ _2761_ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6264_ _2694_ _2695_ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__and2b_1
X_8003_ clknet_leaf_38_hwclk _0145_ net103 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5215_ sound3.count\[7\] sound3.count\[8\] _1735_ vssd1 vssd1 vccd1 vccd1 _1738_
+ sky130_fd_sc_hd__and3_1
X_6195_ _2623_ _2627_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5146_ _1245_ _1580_ _1574_ _1110_ _1676_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__o221a_1
X_5077_ _0688_ _1559_ _1591_ _1606_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__o2111a_2
X_4028_ _0587_ _0605_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__nand2_2
XFILLER_0_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5979_ sound1.count_m\[0\] vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__inv_2
X_7718_ clknet_leaf_57_hwclk _0003_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7649_ _3712_ _3713_ vssd1 vssd1 vccd1 vccd1 _3714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold209 _0078_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ net841 _1533_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__and2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6951_ sound2.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 _3220_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6882_ net785 _1459_ _3142_ vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__mux2_1
X_5902_ _2335_ _2336_ _2337_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__or3_1
X_5833_ _2271_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7503_ sound3.sdiv.C\[3\] _0562_ _3645_ net923 vssd1 vssd1 vccd1 vccd1 _3649_ sky130_fd_sc_hd__a31o_1
X_5764_ wave_comb.u1.M\[0\] wave_comb.u1.M\[1\] _2209_ vssd1 vssd1 vccd1 vccd1 _2217_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4715_ sound1.count\[7\] sound1.count\[8\] _1272_ vssd1 vssd1 vccd1 vccd1 _1278_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5695_ _2039_ _2177_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__nand2_1
X_7434_ _3591_ _3592_ vssd1 vssd1 vccd1 vccd1 _3593_ sky130_fd_sc_hd__xnor2_1
X_4646_ _0990_ _0937_ _1055_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7365_ _3529_ _3530_ vssd1 vssd1 vccd1 vccd1 _3531_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4577_ _0983_ _0992_ _1146_ _0990_ _1147_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold710 seq.player_7.state\[2\] vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold721 _0760_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ net675 _2746_ _0645_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__mux2_1
Xhold754 sound3.count\[7\] vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold743 _0664_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 sound4.count\[9\] vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 inputcont.u3.next_in vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__dlygate4sd3_1
X_7296_ _3464_ _3467_ vssd1 vssd1 vccd1 vccd1 _3469_ sky130_fd_sc_hd__and2_1
Xhold776 sound2.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _0758_ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__dlygate4sd3_1
X_6247_ _2678_ _2679_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__xor2_1
Xhold798 seq.player_7.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__dlygate4sd3_1
X_6178_ _2610_ _2612_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5129_ _0677_ _1083_ _1550_ _1659_ _1107_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__o32a_1
XFILLER_0_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold92 _0282_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 rate_clk.count\[0\] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 rate_clk.count\[1\] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4500_ _0676_ _1052_ _1068_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5480_ sound4.count\[12\] _1973_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4431_ _0940_ _0965_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _0699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7150_ net636 _3168_ _3164_ net659 vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__a22o_1
X_4362_ _0876_ _0877_ _0881_ seq.player_3.state\[3\] vssd1 vssd1 vccd1 vccd1 _0933_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6101_ _2527_ _2528_ _2530_ _2536_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__or4_1
X_4293_ _0575_ _0566_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7081_ _3335_ _3336_ vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__nand2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ sound2.divisor_m\[5\] _2464_ _2467_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__o21a_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7983_ clknet_leaf_15_hwclk sound1.osc.next_count\[4\] net86 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_107_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6934_ sound2.divisor_m\[5\] _3204_ vssd1 vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__xnor2_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6865_ _3150_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
X_5816_ _2254_ _2259_ _2260_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__a21oi_1
X_6796_ net278 _2893_ _0867_ net361 _2853_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5747_ net908 _2201_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7417_ sound3.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 _3577_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5678_ sound4.divisor_m\[18\] _2160_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4629_ _1165_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__inv_2
Xhold551 sound3.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__dlygate4sd3_1
X_7348_ sound3.divisor_m\[9\] sound3.divisor_m\[8\] sound3.divisor_m\[7\] _3492_ vssd1
+ vssd1 vccd1 vccd1 _3515_ sky130_fd_sc_hd__or4_1
Xhold540 _0342_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 sound1.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__dlygate4sd3_1
X_7279_ _3437_ _3452_ _3453_ _3440_ net324 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__a32o_1
Xhold595 sound1.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 sound4.sdiv.A\[21\] vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 seq.clk_div.count\[19\] vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4980_ net724 _1520_ _1504_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3931_ _0515_ _0590_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6650_ sound1.divisor_m\[13\] _3002_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__or2_1
X_3862_ _0525_ _0517_ _0513_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6581_ _2903_ _2948_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5601_ sound4.divisor_m\[7\] _2028_ _2036_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__o21a_1
X_5532_ _2015_ pm.current_waveform\[1\] vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3793_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8320_ clknet_leaf_70_hwclk _0420_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8251_ clknet_leaf_37_hwclk _0351_ net88 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5463_ _1965_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_8182_ clknet_leaf_42_hwclk _0303_ net98 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_7202_ sound3.count\[15\] _2863_ vssd1 vssd1 vccd1 vccd1 _3402_ sky130_fd_sc_hd__and2_1
X_4414_ _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__buf_4
X_5394_ _1001_ _0996_ _1784_ _1904_ _1004_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__o32a_1
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4345_ seq.player_1.state\[0\] _0871_ _0873_ _0915_ vssd1 vssd1 vccd1 vccd1 _0916_
+ sky130_fd_sc_hd__a22o_1
X_7133_ _3349_ _3377_ _3379_ _3174_ net578 vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7064_ sound2.sdiv.A\[17\] _3320_ vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__or2_1
X_4276_ net660 _0850_ _0854_ _0813_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[17\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6015_ _2448_ sound2.count_m\[12\] _2450_ sound2.divisor_m\[12\] vssd1 vssd1 vccd1
+ vccd1 _2451_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7966_ clknet_leaf_22_hwclk _0129_ net103 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6917_ _3183_ _3181_ _3189_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__and3_1
X_7897_ clknet_leaf_1_hwclk net669 net72 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6848_ _3139_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6779_ net585 _2894_ _2890_ net626 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_4_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_hwclk
+ sky130_fd_sc_hd__clkbuf_16
Xhold381 sound1.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 _0662_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 seq.player_7.state\[3\] vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4130_ _0742_ _0741_ _0743_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_5.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4061_ seq.beat\[1\] seq.beat\[0\] seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__or3_4
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7820_ clknet_leaf_3_hwclk net910 net70 vssd1 vssd1 vccd1 vccd1 seq.player_4.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_7751_ clknet_leaf_55_hwclk _0036_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4963_ net881 _1508_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6702_ _3056_ _3057_ vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__or2b_1
X_3914_ _0579_ vssd1 vssd1 vccd1 vccd1 sound1.sdiv.next_start sky130_fd_sc_hd__inv_2
X_7682_ net592 _2184_ _3681_ _3736_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6633_ _2993_ _2995_ vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4894_ _0695_ _0964_ _1418_ _1317_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__o31a_1
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3845_ _0514_ _0516_ _0517_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__or4_2
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6564_ _2932_ _2933_ vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3776_ _0455_ _0458_ _0453_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__nand3b_2
X_6495_ net755 _2877_ _2864_ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__mux2_1
X_8303_ clknet_leaf_62_hwclk _0403_ net78 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_5515_ net129 _0551_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[4\] sky130_fd_sc_hd__xor2_1
X_8234_ clknet_leaf_36_hwclk sound3.osc.next_count\[15\] net93 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5446_ _1951_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout102 net103 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_8
X_8165_ clknet_leaf_38_hwclk net171 net98 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_5377_ _0869_ _1765_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__nor2_1
X_7116_ net950 _3329_ vssd1 vssd1 vccd1 vccd1 _3367_ sky130_fd_sc_hd__nand2_1
X_4328_ seq.player_7.state\[0\] seq.player_7.state\[1\] seq.player_7.state\[2\] seq.player_7.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__or4_1
X_8096_ clknet_leaf_72_hwclk _0238_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_7047_ _3305_ _3306_ vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__nor2_1
X_4259_ seq.clk_div.count\[13\] _0838_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__or2_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ clknet_leaf_31_hwclk _0112_ net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5300_ sound4.count\[5\] _1810_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6280_ _2684_ _2711_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5231_ net427 _1747_ _1721_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5162_ _0944_ _1574_ _1570_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__o21a_1
X_5093_ _1062_ _1565_ _1617_ _1622_ _1623_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__o221a_1
X_4113_ seq.player_6.state\[0\] seq.player_6.state\[1\] _0729_ vssd1 vssd1 vccd1 vccd1
+ _0732_ sky130_fd_sc_hd__and3_1
X_4044_ _0685_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__nand2_8
XFILLER_0_79_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7803_ clknet_leaf_100_hwclk net538 net64 vssd1 vssd1 vccd1 vccd1 seq.player_8.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5995_ _2428_ _2430_ _2394_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__o21ai_1
X_7734_ clknet_leaf_84_hwclk _0019_ net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_4946_ _1318_ _1352_ _1396_ sound2.count\[5\] _1496_ vssd1 vssd1 vccd1 vccd1 _1497_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7665_ net664 _2183_ _3681_ _3724_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__a22o_1
X_4877_ _0677_ _1083_ _1321_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6616_ _2970_ _2976_ _2980_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__o21ai_1
X_3828_ _0472_ _0473_ _0486_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__a21boi_1
X_7596_ _3677_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6547_ sound1.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3759_ _0442_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__clkbuf_8
X_6478_ net750 _2867_ _2864_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8217_ clknet_leaf_39_hwclk _0338_ net100 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5429_ _1779_ _1936_ _1937_ _1938_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__and4_1
X_8148_ clknet_leaf_41_hwclk _0269_ net98 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_84_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_8079_ clknet_leaf_75_hwclk _0221_ net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_99_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_hwclk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_22_hwclk clknet_3_5__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_37_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4800_ _1189_ _1333_ _1336_ _1125_ _1350_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__o221a_1
X_5780_ wave_comb.u1.A\[2\] _2224_ _2230_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ sound1.count\[12\] _1287_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7450_ _3602_ _3605_ _3599_ vssd1 vssd1 vccd1 vccd1 _3607_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4662_ _0974_ _1058_ _1111_ _0941_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6401_ _2821_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7381_ sound3.divisor_m\[13\] _3544_ vssd1 vssd1 vccd1 vccd1 _3545_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4593_ _0683_ _0947_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6332_ _2755_ _2761_ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__nor2_1
X_6263_ _2693_ _2685_ _2689_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8002_ clknet_leaf_38_hwclk net393 net93 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5214_ net523 _1735_ _1737_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[7\] sky130_fd_sc_hd__a21oi_1
X_6194_ _2623_ _2627_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5145_ _0985_ _1567_ _1570_ _1238_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5076_ _1551_ _1565_ _1055_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__a21o_1
X_4027_ _0673_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__inv_2
XFILLER_0_79_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5978_ sound1.count_m\[16\] _2406_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7717_ clknet_leaf_57_hwclk net525 net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_4929_ _1046_ _1347_ _1393_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7648_ _2058_ _2060_ vssd1 vssd1 vccd1 vccd1 _3713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7579_ _3667_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1__f_hwclk clknet_0_hwclk vssd1 vssd1 vccd1 vccd1 clknet_3_1__leaf_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6950_ _3164_ _3218_ _3219_ _3174_ net268 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__a32o_1
X_5901_ sound4.divisor_m\[11\] sound4.count_m\[10\] vssd1 vssd1 vccd1 vccd1 _2337_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6881_ _3160_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5832_ net696 _0569_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__and2_1
X_5763_ wave_comb.u1.A\[1\] vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7502_ _2005_ _3647_ net721 vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__nor3_1
XFILLER_0_72_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4714_ _1277_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5694_ sound4.sdiv.A\[25\] _2038_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__or2_1
X_7433_ _3582_ _3584_ _3581_ vssd1 vssd1 vccd1 vccd1 _3592_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4645_ _0988_ _0955_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7364_ _3525_ _3528_ vssd1 vssd1 vccd1 vccd1 _3530_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4576_ _0994_ _1053_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__or2_1
Xhold711 sound2.count\[8\] vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold700 sound2.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6315_ _2743_ _2745_ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__xnor2_1
Xhold722 seq.player_3.next_state\[3\] vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 seq.player_7.state\[2\] vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 seq.player_8.state\[3\] vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 inputcont.u1.ff_intermediate\[10\] vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__dlygate4sd3_1
X_7295_ _3464_ _3467_ vssd1 vssd1 vccd1 vccd1 _3468_ sky130_fd_sc_hd__nor2_1
Xhold766 sound4.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 sound2.count\[3\] vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 sound4.divisor_m\[13\] vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _2649_ _2652_ _2648_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__a21oi_1
Xhold799 sound2.count\[2\] vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__dlygate4sd3_1
X_6177_ _2311_ _2577_ _2611_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__o21ai_1
X_5128_ _0683_ _1562_ _1580_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__o21a_1
X_5059_ _1557_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold71 sound4.count_m\[18\] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 sound2.count_m\[1\] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 _0187_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 net819 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_1
XFILLER_0_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_2 _0699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _0685_ _0680_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__nor2_8
X_6100_ _2533_ _2534_ _2535_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4361_ seq.player_4.state\[3\] _0888_ _0930_ _0931_ _0883_ vssd1 vssd1 vccd1 vccd1
+ _0932_ sky130_fd_sc_hd__o221a_1
X_4292_ _0700_ _0864_ vssd1 vssd1 vccd1 vccd1 seq.encode.next_sequencer_on sky130_fd_sc_hd__xnor2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7080_ net961 _3329_ vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ sound2.divisor_m\[8\] sound2.count_m\[7\] vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__or2b_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7982_ clknet_leaf_14_hwclk sound1.osc.next_count\[3\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6933_ sound2.divisor_m\[4\] _3194_ _3177_ vssd1 vssd1 vccd1 vccd1 _3204_ sky130_fd_sc_hd__o21a_1
X_6864_ net754 _3149_ _3142_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__mux2_1
X_5815_ wave_comb.u1.A\[9\] _2224_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6795_ net361 _2893_ _0867_ net363 _2852_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5746_ net256 _2182_ _2185_ net290 _2204_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5677_ _2036_ _2035_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7416_ net460 _3463_ sound3.sdiv.next_dived _3576_ vssd1 vssd1 vccd1 vccd1 _0322_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4628_ _0970_ _1078_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold530 sound4.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7347_ net975 vssd1 vssd1 vccd1 vccd1 _3514_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold563 wave_comb.u1.Q\[8\] vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _0994_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__or2_1
Xhold552 sound2.sdiv.A\[20\] vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold541 sound2.count_m\[2\] vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__dlygate4sd3_1
X_7278_ _3446_ _3444_ _3451_ vssd1 vssd1 vccd1 vccd1 _3453_ sky130_fd_sc_hd__nand3_1
Xhold596 pm.current_waveform\[4\] vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 seq.clk_div.count\[6\] vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 seq.clk_div.count\[7\] vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlygate4sd3_1
X_6229_ _2624_ _2661_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__xnor2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 pwm_o sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3930_ _0592_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__or2_2
XFILLER_0_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3861_ _0515_ _0519_ _0521_ _0523_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__or4b_1
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6580_ sound1.divisor_m\[6\] _2937_ vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5600_ sound4.sdiv.A\[8\] _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__or2_1
X_3792_ _0467_ _0470_ inputcont.INTERNAL_SYNCED_I\[12\] vssd1 vssd1 vccd1 vccd1 _0471_
+ sky130_fd_sc_hd__o21a_1
X_5531_ pm.count\[1\] vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8250_ clknet_leaf_37_hwclk net259 net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7201_ net195 _3132_ _3401_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a21o_1
X_5462_ _1779_ _1936_ _1963_ _1964_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__and4_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8181_ clknet_leaf_42_hwclk _0302_ net98 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_4413_ _0983_ _0951_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5393_ _0869_ _1832_ _1842_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__a21oi_1
X_4344_ seq.player_2.state\[0\] _0876_ _0878_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_
+ sky130_fd_sc_hd__a22o_1
X_7132_ _3378_ vssd1 vssd1 vccd1 vccd1 _3379_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7063_ sound2.sdiv.A\[17\] _3320_ vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__nand2_1
X_6014_ sound2.count_m\[11\] vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__inv_2
X_4275_ _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7965_ clknet_leaf_22_hwclk _0128_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _3187_ _3188_ vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__or2_1
X_7896_ clknet_leaf_7_hwclk net673 net72 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6847_ net872 _1352_ _2864_ vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6778_ sound1.sdiv.Q\[5\] _2894_ sound1.sdiv.next_dived net573 vssd1 vssd1 vccd1
+ vccd1 _0146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5729_ sound4.sdiv.Q\[16\] _2182_ _2185_ net239 _2195_ vssd1 vssd1 vccd1 vccd1 _0016_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 sound1.count_m\[16\] vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 seq.tempo_select.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 wave_comb.u1.Q\[0\] vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 seq.player_7.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4060_ _0700_ net1 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__nor2_4
XFILLER_0_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7750_ clknet_leaf_54_hwclk _0035_ net97 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4962_ _1510_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_6701_ sound1.sdiv.A\[18\] _3055_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__nand2_1
X_3913_ _0575_ net61 vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__nor2_8
X_7681_ _2043_ _3735_ vssd1 vssd1 vccd1 vccd1 _3736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4893_ sound2.count\[13\] _1434_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6632_ sound1.divisor_m\[12\] _2994_ vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3844_ _0479_ _0478_ _0485_ _0489_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6563_ _2923_ _2925_ _2922_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3775_ _0456_ inputcont.INTERNAL_SYNCED_I\[4\] _0443_ _0457_ inputcont.INTERNAL_SYNCED_I\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__o32a_1
X_6494_ _1050_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5514_ _0551_ _2002_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[3\] sky130_fd_sc_hd__nor2_1
X_8302_ clknet_leaf_65_hwclk _0402_ net80 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8233_ clknet_leaf_33_hwclk sound3.osc.next_count\[14\] net88 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[14\] sky130_fd_sc_hd__dfrtp_1
X_5445_ sound4.count\[4\] sound4.count\[5\] _1944_ vssd1 vssd1 vccd1 vccd1 _1951_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_112_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8164_ clknet_leaf_38_hwclk net411 net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout103 net2 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7115_ sound2.sdiv.A\[24\] _3329_ vssd1 vssd1 vccd1 vccd1 _3366_ sky130_fd_sc_hd__nor2_1
X_5376_ _1777_ _1788_ _1213_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__a21o_1
X_8095_ clknet_leaf_76_hwclk _0237_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4327_ select1.sequencer_on _0897_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7046_ _3294_ _3298_ _3304_ vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__a21oi_2
X_4258_ seq.clk_div.count\[11\] seq.clk_div.count\[12\] seq.clk_div.count\[13\] _0832_
+ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__and4_1
X_4189_ seq.clk_div.count\[5\] seq.clk_div.count\[15\] seq.clk_div.count\[17\] seq.clk_div.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__or4bb_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ clknet_leaf_31_hwclk _0111_ net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7879_ clknet_leaf_21_hwclk seq_power_on net89 vssd1 vssd1 vccd1 vccd1 seq.encode.inter_keys\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 sound2.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5230_ _1747_ net682 vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[12\] sky130_fd_sc_hd__nor2_1
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5161_ _1658_ _1667_ _1674_ _1683_ _1691_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__o2111ai_1
X_5092_ _1111_ _1611_ _1568_ _1058_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__o22a_1
X_4112_ seq.player_6.state\[0\] _0729_ _0731_ vssd1 vssd1 vccd1 vccd1 seq.player_6.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_4043_ _0686_ _0677_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__nor2_8
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5994_ _2409_ sound1.divisor_m\[4\] _2411_ _2429_ _2404_ vssd1 vssd1 vccd1 vccd1
+ _2430_ sky130_fd_sc_hd__o221a_1
X_7802_ clknet_leaf_0_hwclk net554 net64 vssd1 vssd1 vccd1 vccd1 seq.player_8.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4945_ sound2.count\[11\] _1488_ _1495_ sound2.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _1496_ sky130_fd_sc_hd__o22a_1
X_7733_ clknet_leaf_84_hwclk net243 net74 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_3_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7664_ _2158_ _2164_ vssd1 vssd1 vccd1 vccd1 _3724_ sky130_fd_sc_hd__xnor2_1
X_4876_ _0676_ _1322_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__or2_1
X_6615_ _2974_ _2979_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3827_ _0504_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__inv_2
X_7595_ net771 _3676_ _2186_ vssd1 vssd1 vccd1 vccd1 _3677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6546_ net491 _2895_ _2916_ _2917_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a22o_1
X_3758_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[3\]
+ inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6477_ _1145_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8216_ clknet_leaf_39_hwclk _0337_ net98 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5428_ sound4.count\[0\] sound4.count\[1\] vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__or2_1
X_8147_ clknet_leaf_40_hwclk _0268_ net98 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5359_ _0687_ _1001_ _1790_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8078_ clknet_leaf_79_hwclk _0220_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_7029_ _3164_ _3289_ _3290_ _3174_ net327 vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _1289_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4661_ _0685_ _0940_ _0965_ _0964_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__a211o_1
X_7380_ _3448_ _3543_ vssd1 vssd1 vccd1 vccd1 _3544_ sky130_fd_sc_hd__and2_1
X_6400_ net703 _2820_ _2808_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6331_ _2289_ _2758_ _2760_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__a21oi_1
X_4592_ _0677_ _0976_ _1046_ _1090_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6262_ _2685_ _2689_ _2693_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8001_ clknet_leaf_40_hwclk _0143_ net98 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5213_ net523 _1735_ _1721_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__o21ai_1
X_6193_ _2279_ _2624_ _2626_ _2292_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__o22a_1
X_5144_ _1004_ _1133_ _1559_ _1565_ _0954_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__o32a_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5075_ _1562_ _1548_ _1568_ _1010_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4026_ _0604_ _0595_ _0589_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5977_ sound1.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7716_ clknet_leaf_59_hwclk net263 net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_4928_ sound2.count\[1\] _1404_ _1469_ _1470_ _1478_ vssd1 vssd1 vccd1 vccd1 _1479_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7647_ _2066_ _3710_ vssd1 vssd1 vccd1 vccd1 _3712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4859_ _1004_ _1038_ _1327_ _1321_ _1154_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__o32a_1
XFILLER_0_50_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7578_ net769 _3666_ _3419_ vssd1 vssd1 vccd1 vccd1 _3667_ sky130_fd_sc_hd__mux2_1
X_6529_ sound1.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5900_ sound4.divisor_m\[10\] sound4.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2336_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6880_ net738 _1454_ _3142_ vssd1 vssd1 vccd1 vccd1 _3160_ sky130_fd_sc_hd__mux2_1
X_5831_ _2270_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5762_ wave_comb.u1.A\[0\] _2211_ _2213_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_83_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_7501_ _0562_ _3645_ net720 vssd1 vssd1 vccd1 vccd1 _3648_ sky130_fd_sc_hd__a21oi_1
X_4713_ _1256_ _1275_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5693_ net555 net592 _2038_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__o21ai_1
X_7432_ _3589_ _3590_ vssd1 vssd1 vccd1 vccd1 _3591_ sky130_fd_sc_hd__or2b_1
X_4644_ _0958_ _1058_ _1212_ _1214_ _1070_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_21_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7363_ _3525_ _3528_ vssd1 vssd1 vccd1 vccd1 _3529_ sky130_fd_sc_hd__nor2_1
Xhold701 wave.mode\[0\] vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold712 inputcont.u1.ff_intermediate\[0\] vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ _0683_ _0694_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_98_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7294_ sound3.divisor_m\[4\] _3466_ vssd1 vssd1 vccd1 vccd1 _3467_ sky130_fd_sc_hd__xor2_1
Xhold734 inputcont.u1.ff_intermediate\[8\] vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__dlygate4sd3_1
X_6314_ _2684_ _2711_ _2744_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__a21o_1
Xhold723 sound4.sdiv.Q\[23\] vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 _0726_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__dlygate4sd3_1
X_6245_ _2676_ _2677_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__xor2_1
Xhold767 _3683_ vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 seq.player_2.state\[1\] vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 _0717_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_21_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_hwclk
+ sky130_fd_sc_hd__clkbuf_16
Xhold789 sound4.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__dlygate4sd3_1
X_6176_ _2575_ _2576_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__or2_1
X_5127_ net811 vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_36_hwclk clknet_3_6__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5058_ _1059_ _1562_ _1570_ _1063_ _1588_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__o221a_1
X_4009_ _0659_ net532 vssd1 vssd1 vccd1 vccd1 wave.next_state\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold50 net818 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_1
Xhold61 sound3.sdiv.Q\[14\] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 rate_clk.count\[3\] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold83 _0170_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 sound2.sdiv.Q\[11\] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _0699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4360_ _0886_ _0887_ _0890_ seq.player_5.state\[3\] vssd1 vssd1 vccd1 vccd1 _0931_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4291_ net617 net114 vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__and2b_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _2461_ sound2.divisor_m\[7\] _2463_ sound2.divisor_m\[6\] vssd1 vssd1 vccd1
+ vccd1 _2466_ sky130_fd_sc_hd__o22a_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7981_ clknet_leaf_14_hwclk sound1.osc.next_count\[2\] net83 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6932_ sound2.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6863_ _1495_ vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__inv_2
X_5814_ wave_comb.u1.A\[8\] _2224_ _2257_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_76_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6794_ sound1.sdiv.Q\[21\] _2893_ _0867_ net356 _2851_ vssd1 vssd1 vccd1 vccd1 _0162_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5745_ sound4.count\[16\] _2201_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5676_ sound4.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__inv_2
X_7415_ _3569_ _3575_ vssd1 vssd1 vccd1 vccd1 _3576_ sky130_fd_sc_hd__xor2_1
X_4627_ _0685_ _0964_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__nand2_2
XFILLER_0_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold520 seq.player_5.state\[0\] vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__dlygate4sd3_1
X_7346_ _3437_ _3512_ _3513_ _3440_ net403 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold542 sound2.sdiv.Q\[0\] vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 sound2.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 inputcont.INTERNAL_SYNCED_I\[0\] vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4558_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__buf_4
X_7277_ _3446_ _3444_ _3451_ vssd1 vssd1 vccd1 vccd1 _3452_ sky130_fd_sc_hd__a21o_1
Xhold586 wave_comb.u1.C\[4\] vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 wave_comb.u1.Q\[3\] vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _2800_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 sound1.divisor_m\[9\] vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _0956_ _1026_ _1059_ _0981_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6228_ sound2.sdiv.Q\[3\] _2660_ _2625_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__a21oi_1
X_6159_ sound2.sdiv.Q\[3\] _0578_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__nand2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 note2[2] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 seq_led_on sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3860_ _0510_ _0514_ _0533_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__or3_2
X_3791_ _0464_ _0443_ _0461_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or3b_1
XFILLER_0_128_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5530_ pm.count\[2\] vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__inv_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5461_ sound4.count\[6\] sound4.count\[7\] _1951_ sound4.count\[8\] vssd1 vssd1 vccd1
+ vccd1 _1964_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7200_ net928 _2863_ vssd1 vssd1 vccd1 vccd1 _3401_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4412_ _0674_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__nor2_8
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8180_ clknet_leaf_29_hwclk _0301_ net91 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_5392_ _0993_ _1837_ _1900_ _1902_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__o211a_1
X_7131_ sound2.sdiv.C\[2\] sound2.sdiv.C\[1\] sound2.sdiv.C\[0\] vssd1 vssd1 vccd1
+ vccd1 _3378_ sky130_fd_sc_hd__and3_1
X_4343_ seq.player_3.state\[0\] _0881_ _0883_ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_
+ sky130_fd_sc_hd__a22o_1
X_7062_ _3319_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__inv_2
X_4274_ seq.clk_div.count\[15\] seq.clk_div.count\[16\] seq.clk_div.count\[17\] _0844_
+ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6013_ sound2.count_m\[13\] _2441_ _2448_ sound2.count_m\[12\] vssd1 vssd1 vccd1
+ vccd1 _2449_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7964_ clknet_leaf_23_hwclk _0127_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6915_ _3184_ _3186_ vssd1 vssd1 vccd1 vccd1 _3188_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7895_ clknet_leaf_1_hwclk net685 net70 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6846_ _3138_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6777_ net573 _2894_ sound1.sdiv.next_dived net597 vssd1 vssd1 vccd1 vccd1 _0145_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3989_ net535 net197 net547 vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__a21oi_1
X_5728_ net851 _2186_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5659_ sound4.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7329_ _3486_ _3490_ _3497_ vssd1 vssd1 vccd1 vccd1 _3499_ sky130_fd_sc_hd__a21o_1
Xhold350 sound1.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _0086_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold394 wave.mode\[1\] vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold383 _0046_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 sound2.sdiv.A\[22\] vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _1508_ _1504_ _1509_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__and3b_1
X_6700_ sound1.sdiv.A\[18\] _3055_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3912_ _0578_ vssd1 vssd1 vccd1 vccd1 sound2.sdiv.next_start sky130_fd_sc_hd__inv_2
X_7680_ sound4.sdiv.A\[21\] _2038_ _3733_ vssd1 vssd1 vccd1 vccd1 _3735_ sky130_fd_sc_hd__a21oi_1
X_4892_ _1423_ _1424_ _1434_ sound2.count\[13\] _1442_ vssd1 vssd1 vccd1 vccd1 _1443_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6631_ sound1.divisor_m\[11\] _2984_ _2903_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3843_ _0478_ _0485_ _0479_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6562_ _2930_ _2931_ vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3774_ inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1
+ vccd1 vccd1 _0457_ sky130_fd_sc_hd__nor2_1
X_8301_ clknet_leaf_66_hwclk _0401_ net80 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6493_ _2876_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__clkbuf_1
X_5513_ net176 _0550_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8232_ clknet_leaf_35_hwclk sound3.osc.next_count\[13\] net88 vssd1 vssd1 vccd1 vccd1
+ sound3.count\[13\] sky130_fd_sc_hd__dfrtp_1
X_5444_ _1950_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[4\] sky130_fd_sc_hd__clkbuf_1
X_8163_ clknet_leaf_41_hwclk net203 net98 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7114_ _3360_ _3363_ _3359_ vssd1 vssd1 vccd1 vccd1 _3365_ sky130_fd_sc_hd__o21a_1
X_5375_ _1867_ _1868_ _1876_ _1877_ _1885_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__a221o_1
X_4326_ seq.beat\[3\] seq.encode.play _0879_ inputcont.INTERNAL_SYNCED_I\[6\] vssd1
+ vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__a31o_1
X_8094_ clknet_leaf_77_hwclk _0236_ net76 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7045_ _3294_ _3298_ _3304_ vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__and3_1
X_4257_ _0840_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
X_4188_ seq.tempo_select.state\[1\] seq.tempo_select.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _0782_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7947_ clknet_leaf_31_hwclk _0110_ net90 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ clknet_leaf_3_hwclk seq_play_on net70 vssd1 vssd1 vccd1 vccd1 seq.encode.inter_keys\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6829_ net927 _2855_ vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold180 sound3.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold191 sound2.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5160_ sound3.count\[10\] _1690_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__xnor2_1
X_5091_ _0695_ _0540_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__nor2_1
X_4111_ seq.player_6.state\[1\] seq.player_6.state\[2\] seq.player_6.state\[3\] _0730_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__a311o_1
X_4042_ _0676_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__inv_6
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5993_ _2416_ _2418_ _2410_ sound1.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2429_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7801_ clknet_leaf_7_hwclk oct.next_state\[2\] net71 vssd1 vssd1 vccd1 vccd1 oct.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7732_ clknet_leaf_84_hwclk net351 net77 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_4944_ _1490_ _1492_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7663_ net484 _2183_ sound4.sdiv.next_dived _3723_ vssd1 vssd1 vccd1 vccd1 _0422_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4875_ _1341_ _1372_ _1425_ _1107_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6614_ sound1.divisor_m\[10\] _2978_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3826_ _0500_ _0475_ _0491_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__a31oi_4
X_7594_ _1891_ vssd1 vssd1 vccd1 vccd1 _3676_ sky130_fd_sc_hd__inv_2
X_6545_ _2909_ _2915_ _0866_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3757_ inputcont.INTERNAL_SYNCED_I\[10\] vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8215_ clknet_leaf_46_hwclk _0336_ net98 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6476_ _2005_ _1208_ _2866_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5427_ net414 sound4.count\[1\] vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8146_ clknet_leaf_83_hwclk net156 net75 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_5358_ _0683_ _1769_ _1794_ _0996_ _1800_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__o221a_1
X_8077_ clknet_leaf_79_hwclk _0219_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_4309_ _0702_ seq.encode.play _0879_ inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1
+ vccd1 vccd1 _0880_ sky130_fd_sc_hd__a31o_1
X_7028_ _3277_ _3280_ _3288_ vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__a21o_1
X_5289_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4660_ _1229_ _1230_ _0695_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6330_ _2759_ _2753_ sound2.sdiv.Q\[8\] _2295_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__a2bb2o_1
X_4591_ _0969_ _1004_ _1038_ _1077_ _1000_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__o32a_1
XFILLER_0_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6261_ _2289_ _2691_ _2692_ _2293_ sound1.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 _2693_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8000_ clknet_leaf_39_hwclk _0142_ net98 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5212_ _1735_ _1736_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[6\] sky130_fd_sc_hd__nor2_1
X_6192_ _2594_ _2625_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__xor2_1
X_5143_ sound3.count\[1\] _1673_ _1635_ sound3.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _1674_ sky130_fd_sc_hd__o22a_1
X_5074_ sound3.count\[17\] _1604_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__xor2_1
X_4025_ _0667_ _0670_ _0672_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__o21ai_4
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5976_ sound1.count_m\[17\] _2405_ sound1.count_m\[18\] vssd1 vssd1 vccd1 vccd1 _2412_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7715_ clknet_leaf_57_hwclk _0000_ net95 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4927_ sound2.count\[0\] _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4858_ _1025_ _1046_ _1339_ _1322_ _1164_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__o32a_1
X_7646_ _3681_ _3710_ _3711_ _2184_ net512 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3809_ _0474_ _0475_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4789_ _1331_ _1324_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__or2_1
X_7577_ _1829_ vssd1 vssd1 vccd1 vccd1 _3666_ sky130_fd_sc_hd__inv_2
X_6528_ sound1.divisor_m\[0\] sound1.sdiv.Q\[27\] _2898_ _2900_ vssd1 vssd1 vccd1
+ vccd1 _2901_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6459_ _0575_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__buf_6
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8129_ clknet_leaf_90_hwclk net137 net2 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_hwclk clknet_3_1__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_hwclk
+ sky130_fd_sc_hd__clkbuf_16
X_5830_ net690 _0569_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5761_ wave_comb.u1.next_dived _2213_ _2214_ _0573_ net365 vssd1 vssd1 vccd1 vccd1
+ _0029_ sky130_fd_sc_hd__a32o_1
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7500_ net720 _0562_ _3645_ vssd1 vssd1 vccd1 vccd1 _3647_ sky130_fd_sc_hd__and3_1
X_4712_ sound1.count\[7\] _1272_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7431_ _3586_ _3588_ vssd1 vssd1 vccd1 vccd1 _3590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5692_ sound4.sdiv.A\[24\] _2038_ _2174_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4643_ _0990_ _0941_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7362_ sound3.divisor_m\[11\] _3527_ vssd1 vssd1 vccd1 vccd1 _3528_ sky130_fd_sc_hd__xnor2_1
Xhold702 sound3.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__dlygate4sd3_1
X_4574_ _1070_ _1132_ _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7293_ _3448_ _3465_ vssd1 vssd1 vccd1 vccd1 _3466_ sky130_fd_sc_hd__nand2_1
Xhold713 inputcont.u1.ff_intermediate\[9\] vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ _2710_ _2708_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__and2b_1
Xhold735 sound4.count\[18\] vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 _0024_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 seq.player_7.next_state\[3\] vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ _2631_ _2637_ _2638_ _2644_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__o22ai_2
Xhold779 seq.player_2.next_state\[3\] vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 seq.player_8.next_state\[3\] vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 sound2.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6175_ _2607_ _2609_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5126_ sound3.count\[5\] _1635_ _1641_ sound3.count\[3\] _1656_ vssd1 vssd1 vccd1
+ vccd1 _1657_ sky130_fd_sc_hd__a221o_1
X_5057_ _0679_ net59 _1550_ _1580_ _1053_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__o32a_1
X_4008_ net118 _0658_ net531 vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5959_ sound1.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7629_ _3681_ _3698_ _3699_ _2184_ net194 vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold40 pm.next_count\[8\] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold73 sound4.count_m\[2\] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 sound2.sdiv.Q\[19\] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 sound2.sdiv.Q\[26\] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold84 sound1.sdiv.Q\[11\] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _0252_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_4 _1011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ seq.encode.play _0863_ vssd1 vssd1 vccd1 vccd1 seq.encode.next_play sky130_fd_sc_hd__xnor2_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7980_ clknet_leaf_6_hwclk sound1.osc.next_count\[1\] net72 vssd1 vssd1 vccd1 vccd1
+ sound1.count\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6931_ _3200_ _3202_ net461 _3168_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6862_ _3148_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5813_ net577 _0573_ wave_comb.u1.next_dived _2258_ vssd1 vssd1 vccd1 vccd1 _0037_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6793_ net356 _2893_ _0867_ net376 _2850_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5744_ net290 _2182_ _2185_ net305 _2203_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__a221o_1
X_5675_ _2049_ _2053_ _2152_ _2157_ _2155_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__a221o_1
X_7414_ _3573_ _3574_ vssd1 vssd1 vccd1 vccd1 _3575_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4626_ sound1.count\[9\] _1196_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7345_ _3503_ _3507_ _3510_ _3511_ vssd1 vssd1 vccd1 vccd1 _3513_ sky130_fd_sc_hd__a211o_1
Xhold510 wave_comb.u1.C\[2\] vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold543 sound3.sdiv.A\[19\] vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 sound3.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 sound2.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold521 seq.player_5.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _0995_ _0947_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__or2_1
Xhold576 sound3.sdiv.A\[18\] vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
X_7276_ _3447_ _3450_ vssd1 vssd1 vccd1 vccd1 _3451_ sky130_fd_sc_hd__xnor2_1
Xhold587 pm.current_waveform\[1\] vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ _1018_ _0959_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold565 inputcont.INTERNAL_SYNCED_I\[4\] vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 sound3.count\[6\] vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ _0578_ _2499_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__and2_1
X_6158_ sound2.sdiv.Q\[2\] _0578_ _2591_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__a21oi_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _1146_ _1572_ _1574_ _1125_ _1639_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__o221a_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ sound3.count_m\[10\] vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 mode_out[1] sky130_fd_sc_hd__buf_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 note2[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_hwclk clknet_3_2__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_97_hwclk clknet_3_0__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3790_ _0469_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5460_ _1962_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_35_hwclk clknet_3_4__leaf_hwclk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_hwclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4411_ _0676_ _0680_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5391_ _0997_ _1769_ _1792_ _1010_ _1901_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7130_ net550 net804 net578 vssd1 vssd1 vccd1 vccd1 _3377_ sky130_fd_sc_hd__a21o_1
X_4342_ seq.player_4.state\[0\] _0886_ _0888_ _0912_ vssd1 vssd1 vccd1 vccd1 _0913_
+ sky130_fd_sc_hd__a22o_1
X_7061_ sound2.divisor_m\[18\] _3318_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__xnor2_1
X_4273_ _0852_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6012_ sound2.divisor_m\[13\] vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__inv_2
.ends

