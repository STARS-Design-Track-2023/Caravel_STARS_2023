magic
tech sky130A
magscale 1 2
timestamp 1693931981
<< viali >>
rect 1501 35241 1535 35275
rect 27169 35241 27203 35275
rect 16865 35105 16899 35139
rect 8125 35037 8159 35071
rect 8217 35037 8251 35071
rect 13829 35037 13863 35071
rect 16405 35037 16439 35071
rect 17141 35037 17175 35071
rect 20085 35037 20119 35071
rect 21925 35037 21959 35071
rect 33149 35037 33183 35071
rect 1777 34969 1811 35003
rect 22477 34969 22511 35003
rect 27077 34969 27111 35003
rect 7941 34901 7975 34935
rect 8401 34901 8435 34935
rect 13645 34901 13679 34935
rect 15761 34901 15795 34935
rect 20269 34901 20303 34935
rect 32965 34901 32999 34935
rect 26065 34697 26099 34731
rect 7941 34629 7975 34663
rect 9873 34629 9907 34663
rect 12633 34629 12667 34663
rect 22109 34629 22143 34663
rect 32413 34629 32447 34663
rect 14197 34561 14231 34595
rect 16037 34561 16071 34595
rect 17325 34561 17359 34595
rect 19625 34561 19659 34595
rect 19901 34561 19935 34595
rect 21833 34561 21867 34595
rect 24317 34561 24351 34595
rect 3617 34493 3651 34527
rect 6377 34493 6411 34527
rect 7665 34493 7699 34527
rect 9597 34493 9631 34527
rect 11345 34493 11379 34527
rect 12357 34493 12391 34527
rect 14473 34493 14507 34527
rect 15945 34493 15979 34527
rect 16313 34493 16347 34527
rect 16773 34493 16807 34527
rect 17601 34493 17635 34527
rect 20177 34493 20211 34527
rect 22385 34493 22419 34527
rect 22661 34493 22695 34527
rect 24593 34493 24627 34527
rect 32137 34493 32171 34527
rect 17049 34425 17083 34459
rect 19809 34425 19843 34459
rect 3880 34357 3914 34391
rect 5365 34357 5399 34391
rect 7021 34357 7055 34391
rect 9413 34357 9447 34391
rect 14105 34357 14139 34391
rect 17233 34357 17267 34391
rect 19073 34357 19107 34391
rect 21649 34357 21683 34391
rect 24133 34357 24167 34391
rect 33885 34357 33919 34391
rect 4353 34153 4387 34187
rect 4629 34153 4663 34187
rect 7849 34153 7883 34187
rect 8033 34153 8067 34187
rect 14933 34153 14967 34187
rect 17049 34153 17083 34187
rect 17877 34153 17911 34187
rect 19717 34153 19751 34187
rect 22937 34153 22971 34187
rect 7113 34017 7147 34051
rect 15301 34017 15335 34051
rect 18797 34017 18831 34051
rect 20269 34017 20303 34051
rect 23949 34017 23983 34051
rect 33793 34017 33827 34051
rect 3985 33949 4019 33983
rect 4813 33949 4847 33983
rect 7481 33949 7515 33983
rect 8493 33949 8527 33983
rect 14289 33949 14323 33983
rect 18061 33949 18095 33983
rect 20545 33949 20579 33983
rect 23121 33949 23155 33983
rect 24501 33949 24535 33983
rect 26801 33949 26835 33983
rect 6837 33881 6871 33915
rect 7849 33881 7883 33915
rect 8125 33881 8159 33915
rect 8309 33881 8343 33915
rect 15577 33881 15611 33915
rect 18705 33881 18739 33915
rect 20085 33881 20119 33915
rect 26525 33881 26559 33915
rect 26985 33881 27019 33915
rect 27813 33881 27847 33915
rect 4353 33813 4387 33847
rect 4537 33813 4571 33847
rect 5365 33813 5399 33847
rect 18245 33813 18279 33847
rect 18613 33813 18647 33847
rect 20177 33813 20211 33847
rect 20637 33813 20671 33847
rect 23397 33813 23431 33847
rect 23765 33813 23799 33847
rect 23857 33813 23891 33847
rect 24593 33813 24627 33847
rect 25053 33813 25087 33847
rect 34345 33813 34379 33847
rect 5641 33609 5675 33643
rect 6377 33609 6411 33643
rect 18337 33609 18371 33643
rect 20545 33609 20579 33643
rect 24961 33609 24995 33643
rect 26617 33609 26651 33643
rect 5349 33541 5383 33575
rect 5549 33541 5583 33575
rect 17417 33541 17451 33575
rect 17877 33541 17911 33575
rect 18705 33541 18739 33575
rect 6561 33473 6595 33507
rect 6837 33473 6871 33507
rect 7021 33473 7055 33507
rect 7297 33473 7331 33507
rect 7481 33473 7515 33507
rect 8861 33473 8895 33507
rect 16681 33473 16715 33507
rect 17509 33473 17543 33507
rect 18797 33473 18831 33507
rect 19165 33473 19199 33507
rect 19349 33473 19383 33507
rect 20085 33473 20119 33507
rect 20269 33473 20303 33507
rect 20821 33473 20855 33507
rect 21005 33473 21039 33507
rect 25513 33473 25547 33507
rect 5825 33405 5859 33439
rect 5917 33405 5951 33439
rect 6009 33405 6043 33439
rect 6101 33405 6135 33439
rect 7113 33405 7147 33439
rect 17233 33405 17267 33439
rect 17785 33405 17819 33439
rect 18981 33405 19015 33439
rect 19625 33405 19659 33439
rect 20637 33405 20671 33439
rect 21833 33405 21867 33439
rect 22109 33405 22143 33439
rect 25973 33405 26007 33439
rect 5181 33269 5215 33303
rect 5365 33269 5399 33303
rect 9045 33269 9079 33303
rect 17693 33269 17727 33303
rect 19533 33269 19567 33303
rect 21189 33269 21223 33303
rect 23581 33269 23615 33303
rect 6653 33065 6687 33099
rect 8493 33065 8527 33099
rect 8677 33065 8711 33099
rect 19809 33065 19843 33099
rect 22017 33065 22051 33099
rect 25329 33065 25363 33099
rect 15025 32997 15059 33031
rect 1685 32929 1719 32963
rect 15117 32929 15151 32963
rect 15393 32929 15427 32963
rect 16865 32929 16899 32963
rect 17233 32929 17267 32963
rect 23121 32929 23155 32963
rect 34345 32929 34379 32963
rect 1409 32861 1443 32895
rect 4261 32861 4295 32895
rect 6193 32861 6227 32895
rect 6285 32861 6319 32895
rect 6377 32861 6411 32895
rect 6469 32861 6503 32895
rect 8125 32861 8159 32895
rect 8953 32861 8987 32895
rect 12817 32861 12851 32895
rect 13001 32861 13035 32895
rect 14749 32861 14783 32895
rect 14841 32861 14875 32895
rect 19257 32861 19291 32895
rect 19717 32861 19751 32895
rect 19901 32861 19935 32895
rect 22201 32861 22235 32895
rect 22937 32861 22971 32895
rect 24777 32861 24811 32895
rect 25145 32861 25179 32895
rect 26985 32861 27019 32895
rect 4077 32793 4111 32827
rect 9229 32793 9263 32827
rect 15025 32793 15059 32827
rect 19441 32793 19475 32827
rect 24961 32793 24995 32827
rect 25053 32793 25087 32827
rect 34069 32793 34103 32827
rect 3893 32725 3927 32759
rect 8493 32725 8527 32759
rect 10701 32725 10735 32759
rect 17877 32725 17911 32759
rect 19625 32725 19659 32759
rect 22477 32725 22511 32759
rect 22845 32725 22879 32759
rect 26341 32725 26375 32759
rect 32597 32725 32631 32759
rect 3893 32521 3927 32555
rect 8033 32521 8067 32555
rect 8953 32521 8987 32555
rect 15393 32521 15427 32555
rect 17049 32521 17083 32555
rect 24225 32521 24259 32555
rect 26709 32521 26743 32555
rect 6720 32453 6754 32487
rect 8201 32453 8235 32487
rect 8401 32453 8435 32487
rect 14473 32453 14507 32487
rect 14933 32453 14967 32487
rect 19441 32453 19475 32487
rect 23857 32453 23891 32487
rect 28457 32453 28491 32487
rect 4445 32385 4479 32419
rect 4629 32385 4663 32419
rect 6837 32385 6871 32419
rect 9413 32385 9447 32419
rect 12449 32385 12483 32419
rect 14841 32385 14875 32419
rect 15117 32385 15151 32419
rect 15577 32385 15611 32419
rect 15669 32385 15703 32419
rect 17233 32385 17267 32419
rect 17509 32385 17543 32419
rect 17601 32385 17635 32419
rect 17785 32385 17819 32419
rect 20361 32385 20395 32419
rect 20545 32385 20579 32419
rect 20913 32385 20947 32419
rect 21281 32385 21315 32419
rect 21465 32385 21499 32419
rect 21649 32385 21683 32419
rect 23581 32385 23615 32419
rect 23765 32385 23799 32419
rect 23949 32385 23983 32419
rect 26525 32385 26559 32419
rect 28733 32385 28767 32419
rect 30573 32385 30607 32419
rect 1869 32317 1903 32351
rect 2145 32317 2179 32351
rect 4261 32317 4295 32351
rect 6929 32317 6963 32351
rect 7205 32317 7239 32351
rect 9137 32317 9171 32351
rect 9229 32317 9263 32351
rect 9321 32317 9355 32351
rect 12725 32317 12759 32351
rect 15301 32317 15335 32351
rect 15393 32317 15427 32351
rect 17417 32317 17451 32351
rect 20453 32317 20487 32351
rect 20821 32317 20855 32351
rect 21005 32317 21039 32351
rect 21097 32317 21131 32351
rect 25697 32317 25731 32351
rect 25973 32317 26007 32351
rect 28825 32317 28859 32351
rect 30297 32317 30331 32351
rect 3617 32181 3651 32215
rect 3709 32181 3743 32215
rect 3893 32181 3927 32215
rect 4813 32181 4847 32215
rect 6561 32181 6595 32215
rect 8217 32181 8251 32215
rect 14197 32181 14231 32215
rect 14289 32181 14323 32215
rect 14473 32181 14507 32215
rect 19349 32181 19383 32215
rect 20637 32181 20671 32215
rect 24133 32181 24167 32215
rect 26985 32181 27019 32215
rect 2329 31977 2363 32011
rect 3893 31977 3927 32011
rect 4537 31977 4571 32011
rect 4997 31977 5031 32011
rect 5825 31977 5859 32011
rect 8125 31977 8159 32011
rect 9505 31977 9539 32011
rect 9965 31977 9999 32011
rect 13093 31977 13127 32011
rect 14105 31977 14139 32011
rect 17785 31977 17819 32011
rect 19901 31977 19935 32011
rect 23765 31977 23799 32011
rect 25053 31977 25087 32011
rect 26617 31977 26651 32011
rect 28917 31977 28951 32011
rect 4721 31909 4755 31943
rect 6009 31909 6043 31943
rect 8493 31909 8527 31943
rect 9597 31909 9631 31943
rect 18337 31909 18371 31943
rect 19993 31909 20027 31943
rect 4261 31841 4295 31875
rect 5365 31841 5399 31875
rect 6101 31841 6135 31875
rect 8217 31841 8251 31875
rect 10241 31841 10275 31875
rect 18521 31841 18555 31875
rect 20085 31841 20119 31875
rect 24409 31841 24443 31875
rect 27077 31841 27111 31875
rect 27169 31841 27203 31875
rect 2513 31773 2547 31807
rect 4077 31773 4111 31807
rect 5457 31773 5491 31807
rect 6285 31773 6319 31807
rect 6377 31773 6411 31807
rect 7941 31773 7975 31807
rect 8309 31773 8343 31807
rect 8769 31773 8803 31807
rect 9137 31773 9171 31807
rect 9341 31773 9375 31807
rect 11989 31773 12023 31807
rect 12081 31773 12115 31807
rect 13277 31773 13311 31807
rect 14473 31773 14507 31807
rect 17141 31773 17175 31807
rect 17234 31773 17268 31807
rect 17417 31773 17451 31807
rect 17606 31773 17640 31807
rect 18613 31773 18647 31807
rect 18981 31773 19015 31807
rect 19257 31773 19291 31807
rect 19441 31773 19475 31807
rect 19717 31773 19751 31807
rect 19809 31773 19843 31807
rect 22017 31773 22051 31807
rect 27721 31773 27755 31807
rect 27905 31773 27939 31807
rect 28089 31773 28123 31807
rect 28365 31773 28399 31807
rect 28549 31773 28583 31807
rect 28733 31773 28767 31807
rect 4353 31705 4387 31739
rect 4997 31705 5031 31739
rect 5825 31705 5859 31739
rect 11713 31705 11747 31739
rect 12357 31705 12391 31739
rect 14289 31705 14323 31739
rect 17509 31705 17543 31739
rect 18889 31705 18923 31739
rect 22293 31705 22327 31739
rect 27997 31705 28031 31739
rect 28641 31705 28675 31739
rect 4553 31637 4587 31671
rect 4813 31637 4847 31671
rect 6101 31637 6135 31671
rect 7757 31637 7791 31671
rect 8677 31637 8711 31671
rect 9965 31637 9999 31671
rect 10149 31637 10183 31671
rect 19625 31637 19659 31671
rect 26985 31637 27019 31671
rect 28273 31637 28307 31671
rect 4537 31433 4571 31467
rect 5825 31433 5859 31467
rect 6469 31433 6503 31467
rect 8585 31433 8619 31467
rect 10149 31433 10183 31467
rect 10609 31433 10643 31467
rect 17141 31433 17175 31467
rect 19441 31433 19475 31467
rect 22569 31433 22603 31467
rect 22937 31433 22971 31467
rect 23397 31433 23431 31467
rect 27721 31433 27755 31467
rect 28457 31433 28491 31467
rect 6009 31365 6043 31399
rect 9781 31365 9815 31399
rect 15117 31365 15151 31399
rect 23305 31365 23339 31399
rect 2789 31297 2823 31331
rect 5733 31297 5767 31331
rect 7021 31297 7055 31331
rect 8125 31297 8159 31331
rect 9965 31297 9999 31331
rect 10425 31297 10459 31331
rect 14749 31297 14783 31331
rect 15393 31297 15427 31331
rect 17325 31297 17359 31331
rect 17601 31297 17635 31331
rect 17693 31297 17727 31331
rect 17877 31297 17911 31331
rect 19165 31297 19199 31331
rect 19257 31297 19291 31331
rect 20177 31297 20211 31331
rect 21189 31297 21223 31331
rect 21281 31297 21315 31331
rect 22753 31297 22787 31331
rect 24961 31297 24995 31331
rect 3065 31229 3099 31263
rect 9137 31229 9171 31263
rect 17509 31229 17543 31263
rect 19441 31229 19475 31263
rect 20453 31229 20487 31263
rect 20821 31229 20855 31263
rect 21005 31229 21039 31263
rect 21097 31229 21131 31263
rect 23489 31229 23523 31263
rect 27629 31229 27663 31263
rect 28365 31229 28399 31263
rect 29101 31229 29135 31263
rect 15301 31161 15335 31195
rect 20361 31161 20395 31195
rect 6009 31093 6043 31127
rect 7573 31093 7607 31127
rect 15117 31093 15151 31127
rect 15577 31093 15611 31127
rect 20269 31093 20303 31127
rect 24777 31093 24811 31127
rect 26985 31093 27019 31127
rect 3249 30889 3283 30923
rect 5444 30889 5478 30923
rect 6929 30889 6963 30923
rect 7284 30889 7318 30923
rect 12344 30889 12378 30923
rect 14105 30889 14139 30923
rect 14841 30889 14875 30923
rect 15025 30889 15059 30923
rect 17325 30889 17359 30923
rect 19349 30889 19383 30923
rect 20913 30889 20947 30923
rect 21465 30889 21499 30923
rect 24672 30889 24706 30923
rect 27997 30889 28031 30923
rect 17049 30821 17083 30855
rect 5181 30753 5215 30787
rect 7021 30753 7055 30787
rect 12081 30753 12115 30787
rect 15301 30753 15335 30787
rect 15577 30753 15611 30787
rect 24409 30753 24443 30787
rect 26249 30753 26283 30787
rect 28641 30753 28675 30787
rect 3433 30685 3467 30719
rect 9781 30685 9815 30719
rect 14289 30685 14323 30719
rect 14565 30685 14599 30719
rect 14749 30685 14783 30719
rect 17504 30685 17538 30719
rect 17693 30685 17727 30719
rect 17821 30685 17855 30719
rect 17969 30685 18003 30719
rect 19441 30685 19475 30719
rect 21097 30685 21131 30719
rect 21373 30685 21407 30719
rect 21557 30685 21591 30719
rect 9229 30617 9263 30651
rect 14993 30617 15027 30651
rect 15209 30617 15243 30651
rect 17601 30617 17635 30651
rect 21281 30617 21315 30651
rect 26525 30617 26559 30651
rect 8769 30549 8803 30583
rect 13829 30549 13863 30583
rect 26157 30549 26191 30583
rect 28089 30549 28123 30583
rect 14197 30345 14231 30379
rect 15209 30345 15243 30379
rect 25145 30345 25179 30379
rect 25605 30345 25639 30379
rect 26985 30345 27019 30379
rect 29745 30345 29779 30379
rect 6653 30277 6687 30311
rect 9413 30277 9447 30311
rect 9873 30277 9907 30311
rect 26157 30277 26191 30311
rect 8953 30209 8987 30243
rect 9505 30209 9539 30243
rect 13737 30209 13771 30243
rect 13829 30209 13863 30243
rect 13921 30209 13955 30243
rect 15577 30209 15611 30243
rect 15669 30209 15703 30243
rect 20269 30209 20303 30243
rect 21373 30209 21407 30243
rect 21557 30209 21591 30243
rect 24041 30209 24075 30243
rect 25513 30209 25547 30243
rect 25973 30209 26007 30243
rect 26249 30209 26283 30243
rect 26341 30209 26375 30243
rect 27997 30209 28031 30243
rect 6536 30141 6570 30175
rect 6745 30141 6779 30175
rect 7021 30141 7055 30175
rect 9137 30141 9171 30175
rect 14013 30141 14047 30175
rect 15393 30141 15427 30175
rect 15485 30141 15519 30175
rect 19993 30141 20027 30175
rect 20729 30141 20763 30175
rect 20913 30141 20947 30175
rect 21005 30141 21039 30175
rect 21097 30141 21131 30175
rect 21189 30141 21223 30175
rect 22109 30141 22143 30175
rect 22385 30141 22419 30175
rect 24317 30141 24351 30175
rect 25789 30141 25823 30175
rect 27537 30141 27571 30175
rect 28273 30141 28307 30175
rect 8769 30073 8803 30107
rect 21465 30073 21499 30107
rect 26525 30073 26559 30107
rect 6377 30005 6411 30039
rect 9321 30005 9355 30039
rect 9873 30005 9907 30039
rect 10057 30005 10091 30039
rect 20085 30005 20119 30039
rect 20177 30005 20211 30039
rect 23857 30005 23891 30039
rect 8769 29801 8803 29835
rect 9229 29801 9263 29835
rect 13921 29801 13955 29835
rect 18153 29801 18187 29835
rect 20821 29801 20855 29835
rect 22661 29801 22695 29835
rect 9413 29733 9447 29767
rect 23029 29733 23063 29767
rect 29377 29733 29411 29767
rect 3801 29665 3835 29699
rect 8401 29665 8435 29699
rect 8493 29665 8527 29699
rect 8585 29665 8619 29699
rect 9597 29665 9631 29699
rect 9781 29665 9815 29699
rect 9874 29665 9908 29699
rect 10057 29665 10091 29699
rect 11989 29665 12023 29699
rect 14197 29665 14231 29699
rect 15577 29665 15611 29699
rect 19901 29665 19935 29699
rect 23489 29665 23523 29699
rect 23673 29665 23707 29699
rect 26341 29665 26375 29699
rect 8309 29597 8343 29631
rect 9965 29597 9999 29631
rect 13001 29597 13035 29631
rect 13645 29597 13679 29631
rect 13737 29597 13771 29631
rect 15025 29597 15059 29631
rect 15117 29597 15151 29631
rect 17417 29597 17451 29631
rect 17601 29597 17635 29631
rect 17693 29597 17727 29631
rect 17785 29597 17819 29631
rect 17969 29597 18003 29631
rect 18705 29597 18739 29631
rect 18889 29597 18923 29631
rect 20085 29597 20119 29631
rect 20177 29597 20211 29631
rect 21189 29597 21223 29631
rect 22845 29597 22879 29631
rect 29193 29597 29227 29631
rect 29377 29597 29411 29631
rect 30113 29597 30147 29631
rect 30849 29597 30883 29631
rect 4077 29529 4111 29563
rect 9045 29529 9079 29563
rect 9245 29529 9279 29563
rect 11713 29529 11747 29563
rect 15853 29529 15887 29563
rect 19901 29529 19935 29563
rect 21005 29529 21039 29563
rect 26065 29529 26099 29563
rect 30297 29529 30331 29563
rect 5549 29461 5583 29495
rect 10241 29461 10275 29495
rect 12357 29461 12391 29495
rect 15301 29461 15335 29495
rect 17325 29461 17359 29495
rect 18797 29461 18831 29495
rect 23397 29461 23431 29495
rect 24593 29461 24627 29495
rect 29561 29461 29595 29495
rect 4077 29257 4111 29291
rect 6009 29257 6043 29291
rect 15485 29257 15519 29291
rect 17509 29257 17543 29291
rect 20453 29257 20487 29291
rect 25605 29257 25639 29291
rect 4537 29189 4571 29223
rect 7573 29189 7607 29223
rect 7757 29189 7791 29223
rect 8677 29189 8711 29223
rect 14105 29189 14139 29223
rect 15393 29189 15427 29223
rect 15669 29189 15703 29223
rect 17785 29189 17819 29223
rect 17877 29189 17911 29223
rect 18889 29189 18923 29223
rect 23121 29189 23155 29223
rect 25697 29189 25731 29223
rect 31125 29189 31159 29223
rect 3433 29121 3467 29155
rect 3617 29121 3651 29155
rect 3893 29121 3927 29155
rect 5181 29121 5215 29155
rect 5365 29121 5399 29155
rect 5733 29121 5767 29155
rect 7021 29121 7055 29155
rect 7113 29121 7147 29155
rect 7849 29121 7883 29155
rect 9045 29121 9079 29155
rect 9321 29121 9355 29155
rect 9505 29121 9539 29155
rect 9873 29121 9907 29155
rect 10609 29121 10643 29155
rect 11161 29121 11195 29155
rect 11345 29121 11379 29155
rect 11529 29121 11563 29155
rect 13830 29143 13864 29177
rect 14197 29121 14231 29155
rect 14381 29121 14415 29155
rect 16865 29121 16899 29155
rect 17049 29121 17083 29155
rect 17141 29121 17175 29155
rect 17688 29121 17722 29155
rect 18060 29121 18094 29155
rect 18153 29121 18187 29155
rect 18245 29121 18279 29155
rect 18429 29121 18463 29155
rect 18613 29121 18647 29155
rect 18705 29121 18739 29155
rect 19165 29121 19199 29155
rect 20637 29121 20671 29155
rect 22477 29121 22511 29155
rect 23029 29121 23063 29155
rect 24317 29121 24351 29155
rect 24501 29121 24535 29155
rect 24593 29121 24627 29155
rect 24685 29121 24719 29155
rect 26341 29121 26375 29155
rect 27169 29121 27203 29155
rect 29377 29121 29411 29155
rect 31401 29121 31435 29155
rect 5641 29053 5675 29087
rect 5850 29053 5884 29087
rect 10517 29053 10551 29087
rect 11805 29053 11839 29087
rect 13277 29053 13311 29087
rect 14105 29053 14139 29087
rect 14657 29053 14691 29087
rect 18889 29053 18923 29087
rect 19349 29053 19383 29087
rect 19533 29053 19567 29087
rect 19625 29053 19659 29087
rect 19717 29053 19751 29087
rect 19809 29053 19843 29087
rect 20729 29053 20763 29087
rect 20821 29053 20855 29087
rect 20913 29053 20947 29087
rect 23305 29053 23339 29087
rect 24961 29053 24995 29087
rect 27445 29053 27479 29087
rect 29009 29053 29043 29087
rect 29285 29053 29319 29087
rect 10793 28985 10827 29019
rect 16037 28985 16071 29019
rect 18521 28985 18555 29019
rect 19073 28985 19107 29019
rect 22661 28985 22695 29019
rect 24869 28985 24903 29019
rect 28917 28985 28951 29019
rect 7297 28917 7331 28951
rect 7389 28917 7423 28951
rect 8861 28917 8895 28951
rect 11345 28917 11379 28951
rect 13921 28917 13955 28951
rect 14197 28917 14231 28951
rect 15669 28917 15703 28951
rect 16681 28917 16715 28951
rect 22293 28917 22327 28951
rect 29653 28917 29687 28951
rect 3801 28713 3835 28747
rect 4629 28713 4663 28747
rect 5273 28713 5307 28747
rect 7297 28713 7331 28747
rect 10701 28713 10735 28747
rect 15853 28713 15887 28747
rect 16681 28713 16715 28747
rect 16865 28713 16899 28747
rect 18337 28713 18371 28747
rect 18797 28713 18831 28747
rect 19717 28713 19751 28747
rect 20821 28713 20855 28747
rect 21005 28713 21039 28747
rect 23489 28713 23523 28747
rect 29193 28713 29227 28747
rect 29377 28713 29411 28747
rect 30389 28713 30423 28747
rect 4813 28645 4847 28679
rect 6929 28645 6963 28679
rect 7481 28645 7515 28679
rect 19901 28645 19935 28679
rect 3617 28577 3651 28611
rect 4077 28577 4111 28611
rect 4169 28577 4203 28611
rect 5917 28577 5951 28611
rect 8953 28577 8987 28611
rect 12265 28577 12299 28611
rect 14105 28577 14139 28611
rect 18613 28577 18647 28611
rect 21741 28577 21775 28611
rect 28365 28577 28399 28611
rect 28549 28577 28583 28611
rect 28733 28577 28767 28611
rect 29653 28577 29687 28611
rect 2973 28509 3007 28543
rect 3157 28509 3191 28543
rect 3433 28509 3467 28543
rect 3985 28509 4019 28543
rect 4261 28509 4295 28543
rect 4905 28509 4939 28543
rect 5733 28509 5767 28543
rect 5825 28509 5859 28543
rect 6009 28509 6043 28543
rect 8769 28509 8803 28543
rect 18521 28509 18555 28543
rect 18797 28509 18831 28543
rect 19349 28509 19383 28543
rect 19809 28509 19843 28543
rect 19993 28509 20027 28543
rect 20453 28509 20487 28543
rect 20637 28509 20671 28543
rect 20913 28509 20947 28543
rect 21097 28509 21131 28543
rect 23581 28509 23615 28543
rect 23765 28509 23799 28543
rect 23949 28509 23983 28543
rect 25053 28509 25087 28543
rect 26525 28509 26559 28543
rect 26709 28509 26743 28543
rect 26801 28509 26835 28543
rect 28642 28509 28676 28543
rect 28825 28509 28859 28543
rect 30573 28509 30607 28543
rect 30665 28509 30699 28543
rect 4445 28441 4479 28475
rect 5273 28441 5307 28475
rect 7297 28441 7331 28475
rect 7665 28441 7699 28475
rect 8493 28441 8527 28475
rect 9229 28441 9263 28475
rect 14381 28441 14415 28475
rect 17049 28441 17083 28475
rect 19533 28441 19567 28475
rect 22017 28441 22051 28475
rect 23857 28441 23891 28475
rect 29009 28441 29043 28475
rect 30297 28441 30331 28475
rect 30389 28441 30423 28475
rect 3065 28373 3099 28407
rect 3249 28373 3283 28407
rect 4645 28373 4679 28407
rect 5457 28373 5491 28407
rect 5549 28373 5583 28407
rect 8585 28373 8619 28407
rect 12909 28373 12943 28407
rect 16849 28373 16883 28407
rect 24133 28373 24167 28407
rect 24409 28373 24443 28407
rect 26341 28373 26375 28407
rect 29209 28373 29243 28407
rect 3341 28169 3375 28203
rect 3801 28169 3835 28203
rect 7113 28169 7147 28203
rect 27721 28169 27755 28203
rect 1869 28101 1903 28135
rect 8585 28101 8619 28135
rect 12541 28101 12575 28135
rect 22569 28101 22603 28135
rect 3525 28033 3559 28067
rect 5549 28033 5583 28067
rect 8861 28033 8895 28067
rect 12265 28033 12299 28067
rect 12357 28033 12391 28067
rect 22477 28033 22511 28067
rect 22937 28033 22971 28067
rect 25605 28033 25639 28067
rect 26985 28033 27019 28067
rect 30113 28033 30147 28067
rect 30573 28033 30607 28067
rect 31125 28033 31159 28067
rect 34345 28033 34379 28067
rect 1593 27965 1627 27999
rect 3617 27965 3651 27999
rect 3801 27965 3835 27999
rect 22753 27965 22787 27999
rect 23489 27965 23523 27999
rect 25329 27965 25363 27999
rect 25697 27965 25731 27999
rect 26249 27965 26283 27999
rect 28273 27965 28307 27999
rect 30021 27965 30055 27999
rect 23857 27897 23891 27931
rect 30481 27897 30515 27931
rect 5365 27829 5399 27863
rect 12541 27829 12575 27863
rect 22109 27829 22143 27863
rect 27629 27829 27663 27863
rect 34161 27829 34195 27863
rect 5444 27625 5478 27659
rect 22293 27625 22327 27659
rect 23949 27625 23983 27659
rect 27641 27625 27675 27659
rect 30757 27625 30791 27659
rect 32241 27625 32275 27659
rect 34087 27625 34121 27659
rect 6929 27557 6963 27591
rect 16037 27557 16071 27591
rect 20545 27489 20579 27523
rect 23397 27489 23431 27523
rect 27905 27489 27939 27523
rect 32505 27489 32539 27523
rect 34345 27489 34379 27523
rect 5181 27421 5215 27455
rect 10333 27421 10367 27455
rect 11253 27421 11287 27455
rect 11529 27421 11563 27455
rect 13645 27421 13679 27455
rect 14473 27421 14507 27455
rect 15393 27421 15427 27455
rect 15853 27421 15887 27455
rect 16221 27421 16255 27455
rect 16313 27421 16347 27455
rect 17049 27421 17083 27455
rect 17601 27421 17635 27455
rect 17785 27421 17819 27455
rect 17969 27421 18003 27455
rect 18153 27421 18187 27455
rect 18797 27421 18831 27455
rect 19441 27421 19475 27455
rect 24685 27421 24719 27455
rect 28181 27421 28215 27455
rect 13369 27353 13403 27387
rect 16037 27353 16071 27387
rect 20821 27353 20855 27387
rect 25881 27353 25915 27387
rect 28917 27353 28951 27387
rect 10149 27285 10183 27319
rect 11069 27285 11103 27319
rect 11437 27285 11471 27319
rect 11897 27285 11931 27319
rect 14289 27285 14323 27319
rect 17877 27285 17911 27319
rect 19257 27285 19291 27319
rect 25329 27285 25363 27319
rect 32597 27285 32631 27319
rect 11345 27081 11379 27115
rect 11687 27081 11721 27115
rect 12725 27081 12759 27115
rect 13737 27081 13771 27115
rect 16681 27081 16715 27115
rect 18889 27081 18923 27115
rect 21833 27081 21867 27115
rect 23029 27081 23063 27115
rect 25513 27081 25547 27115
rect 26617 27081 26651 27115
rect 9873 27013 9907 27047
rect 11897 27013 11931 27047
rect 14105 27013 14139 27047
rect 17417 27013 17451 27047
rect 19349 27013 19383 27047
rect 24501 27013 24535 27047
rect 26157 27013 26191 27047
rect 12081 26945 12115 26979
rect 15945 26945 15979 26979
rect 16865 26945 16899 26979
rect 16957 26945 16991 26979
rect 21557 26945 21591 26979
rect 22017 26945 22051 26979
rect 24777 26945 24811 26979
rect 25237 26945 25271 26979
rect 25329 26945 25363 26979
rect 27169 26945 27203 26979
rect 27353 26945 27387 26979
rect 27629 26945 27663 26979
rect 27813 26945 27847 26979
rect 28273 26945 28307 26979
rect 7021 26877 7055 26911
rect 9597 26877 9631 26911
rect 13093 26877 13127 26911
rect 13829 26877 13863 26911
rect 16681 26877 16715 26911
rect 17141 26877 17175 26911
rect 19073 26877 19107 26911
rect 20821 26877 20855 26911
rect 24869 26877 24903 26911
rect 24961 26877 24995 26911
rect 28549 26877 28583 26911
rect 7297 26809 7331 26843
rect 26433 26809 26467 26843
rect 27905 26809 27939 26843
rect 7481 26741 7515 26775
rect 11529 26741 11563 26775
rect 11713 26741 11747 26775
rect 15577 26741 15611 26775
rect 16497 26741 16531 26775
rect 20913 26741 20947 26775
rect 30021 26741 30055 26775
rect 6469 26537 6503 26571
rect 10333 26537 10367 26571
rect 10517 26537 10551 26571
rect 12265 26537 12299 26571
rect 12633 26537 12667 26571
rect 14105 26537 14139 26571
rect 14289 26537 14323 26571
rect 16116 26537 16150 26571
rect 17601 26537 17635 26571
rect 19349 26537 19383 26571
rect 21189 26537 21223 26571
rect 26985 26537 27019 26571
rect 28825 26537 28859 26571
rect 10885 26469 10919 26503
rect 3801 26401 3835 26435
rect 6929 26401 6963 26435
rect 12173 26401 12207 26435
rect 15853 26401 15887 26435
rect 19993 26401 20027 26435
rect 21281 26401 21315 26435
rect 21557 26401 21591 26435
rect 23029 26401 23063 26435
rect 23765 26401 23799 26435
rect 27353 26401 27387 26435
rect 27997 26401 28031 26435
rect 30665 26401 30699 26435
rect 31861 26401 31895 26435
rect 33609 26401 33643 26435
rect 3433 26333 3467 26367
rect 5825 26333 5859 26367
rect 6009 26333 6043 26367
rect 6193 26333 6227 26367
rect 6285 26333 6319 26367
rect 12449 26333 12483 26367
rect 14657 26333 14691 26367
rect 14933 26333 14967 26367
rect 19717 26333 19751 26367
rect 21005 26333 21039 26367
rect 25053 26333 25087 26367
rect 25237 26333 25271 26367
rect 28181 26333 28215 26367
rect 28457 26333 28491 26367
rect 28549 26333 28583 26367
rect 29009 26333 29043 26367
rect 29193 26333 29227 26367
rect 29285 26333 29319 26367
rect 30573 26333 30607 26367
rect 31217 26333 31251 26367
rect 31493 26333 31527 26367
rect 31585 26333 31619 26367
rect 1409 26265 1443 26299
rect 1777 26265 1811 26299
rect 4077 26265 4111 26299
rect 7205 26265 7239 26299
rect 10517 26265 10551 26299
rect 14289 26265 14323 26299
rect 14749 26265 14783 26299
rect 15117 26265 15151 26299
rect 19809 26265 19843 26299
rect 24409 26265 24443 26299
rect 25513 26265 25547 26299
rect 28365 26265 28399 26299
rect 31401 26265 31435 26299
rect 33333 26265 33367 26299
rect 3617 26197 3651 26231
rect 5549 26197 5583 26231
rect 8677 26197 8711 26231
rect 23121 26197 23155 26231
rect 28733 26197 28767 26231
rect 30113 26197 30147 26231
rect 30481 26197 30515 26231
rect 31769 26197 31803 26231
rect 3801 25993 3835 26027
rect 3985 25993 4019 26027
rect 7389 25993 7423 26027
rect 21833 25993 21867 26027
rect 22201 25993 22235 26027
rect 25053 25993 25087 26027
rect 30389 25993 30423 26027
rect 32137 25993 32171 26027
rect 5365 25925 5399 25959
rect 7021 25925 7055 25959
rect 12357 25925 12391 25959
rect 23397 25925 23431 25959
rect 26341 25925 26375 25959
rect 4353 25857 4387 25891
rect 4997 25857 5031 25891
rect 5825 25857 5859 25891
rect 6561 25857 6595 25891
rect 7573 25857 7607 25891
rect 14381 25857 14415 25891
rect 23121 25857 23155 25891
rect 25329 25857 25363 25891
rect 25605 25857 25639 25891
rect 26433 25857 26467 25891
rect 26617 25857 26651 25891
rect 27077 25857 27111 25891
rect 27261 25857 27295 25891
rect 27445 25857 27479 25891
rect 30021 25857 30055 25891
rect 32321 25857 32355 25891
rect 32505 25857 32539 25891
rect 32597 25857 32631 25891
rect 4721 25789 4755 25823
rect 4813 25789 4847 25823
rect 4905 25789 4939 25823
rect 5641 25789 5675 25823
rect 6653 25789 6687 25823
rect 8769 25789 8803 25823
rect 14197 25789 14231 25823
rect 22293 25789 22327 25823
rect 22477 25789 22511 25823
rect 25053 25789 25087 25823
rect 26801 25789 26835 25823
rect 30113 25789 30147 25823
rect 6009 25721 6043 25755
rect 12173 25721 12207 25755
rect 12725 25721 12759 25755
rect 25237 25721 25271 25755
rect 27261 25721 27295 25755
rect 3985 25653 4019 25687
rect 4537 25653 4571 25687
rect 5825 25653 5859 25687
rect 6377 25653 6411 25687
rect 6929 25653 6963 25687
rect 9413 25653 9447 25687
rect 12357 25653 12391 25687
rect 14565 25653 14599 25687
rect 24869 25653 24903 25687
rect 27721 25653 27755 25687
rect 4629 25449 4663 25483
rect 4813 25449 4847 25483
rect 7205 25449 7239 25483
rect 7849 25449 7883 25483
rect 9045 25449 9079 25483
rect 15761 25449 15795 25483
rect 16037 25449 16071 25483
rect 21005 25449 21039 25483
rect 28825 25449 28859 25483
rect 29193 25449 29227 25483
rect 29837 25449 29871 25483
rect 30205 25449 30239 25483
rect 32781 25449 32815 25483
rect 9137 25381 9171 25415
rect 27169 25381 27203 25415
rect 4445 25313 4479 25347
rect 9229 25313 9263 25347
rect 9321 25313 9355 25347
rect 11069 25313 11103 25347
rect 17325 25313 17359 25347
rect 19257 25313 19291 25347
rect 32045 25313 32079 25347
rect 33425 25313 33459 25347
rect 3249 25245 3283 25279
rect 3433 25245 3467 25279
rect 3525 25245 3559 25279
rect 3801 25245 3835 25279
rect 6653 25245 6687 25279
rect 6929 25245 6963 25279
rect 7573 25245 7607 25279
rect 7941 25245 7975 25279
rect 8953 25245 8987 25279
rect 11713 25245 11747 25279
rect 11897 25245 11931 25279
rect 12081 25245 12115 25279
rect 13921 25245 13955 25279
rect 15577 25245 15611 25279
rect 16313 25245 16347 25279
rect 16497 25245 16531 25279
rect 26157 25245 26191 25279
rect 26249 25245 26283 25279
rect 26617 25245 26651 25279
rect 26985 25245 27019 25279
rect 28733 25245 28767 25279
rect 29561 25245 29595 25279
rect 30113 25245 30147 25279
rect 30297 25245 30331 25279
rect 30481 25245 30515 25279
rect 30665 25245 30699 25279
rect 32137 25245 32171 25279
rect 4997 25177 5031 25211
rect 7389 25177 7423 25211
rect 7849 25177 7883 25211
rect 9597 25177 9631 25211
rect 13645 25177 13679 25211
rect 15393 25177 15427 25211
rect 16221 25177 16255 25211
rect 16681 25177 16715 25211
rect 17601 25177 17635 25211
rect 19533 25177 19567 25211
rect 24685 25177 24719 25211
rect 25421 25177 25455 25211
rect 26433 25177 26467 25211
rect 27445 25177 27479 25211
rect 33241 25177 33275 25211
rect 3065 25109 3099 25143
rect 4797 25109 4831 25143
rect 6469 25109 6503 25143
rect 6837 25109 6871 25143
rect 7021 25109 7055 25143
rect 7189 25109 7223 25143
rect 7665 25109 7699 25143
rect 8585 25109 8619 25143
rect 11161 25109 11195 25143
rect 11989 25109 12023 25143
rect 12173 25109 12207 25143
rect 15853 25109 15887 25143
rect 16021 25109 16055 25143
rect 19073 25109 19107 25143
rect 27537 25109 27571 25143
rect 30021 25109 30055 25143
rect 30849 25109 30883 25143
rect 32505 25109 32539 25143
rect 33149 25109 33183 25143
rect 3617 24905 3651 24939
rect 3893 24905 3927 24939
rect 6561 24905 6595 24939
rect 7757 24905 7791 24939
rect 10241 24905 10275 24939
rect 12081 24905 12115 24939
rect 12373 24905 12407 24939
rect 12541 24905 12575 24939
rect 12909 24905 12943 24939
rect 16497 24905 16531 24939
rect 18061 24905 18095 24939
rect 18245 24905 18279 24939
rect 19533 24905 19567 24939
rect 21189 24905 21223 24939
rect 23673 24905 23707 24939
rect 24317 24905 24351 24939
rect 31861 24905 31895 24939
rect 4813 24837 4847 24871
rect 12173 24837 12207 24871
rect 22109 24837 22143 24871
rect 3801 24769 3835 24803
rect 4077 24769 4111 24803
rect 4997 24769 5031 24803
rect 5181 24769 5215 24803
rect 6929 24769 6963 24803
rect 9505 24769 9539 24803
rect 10425 24769 10459 24803
rect 10701 24769 10735 24803
rect 11161 24769 11195 24803
rect 11621 24769 11655 24803
rect 11713 24769 11747 24803
rect 12725 24769 12759 24803
rect 14749 24769 14783 24803
rect 16957 24769 16991 24803
rect 17509 24769 17543 24803
rect 18429 24769 18463 24803
rect 19349 24769 19383 24803
rect 21097 24769 21131 24803
rect 23857 24769 23891 24803
rect 26985 24769 27019 24803
rect 27169 24769 27203 24803
rect 27261 24769 27295 24803
rect 29469 24769 29503 24803
rect 30481 24769 30515 24803
rect 30665 24769 30699 24803
rect 30757 24769 30791 24803
rect 30941 24769 30975 24803
rect 31125 24769 31159 24803
rect 31309 24769 31343 24803
rect 31401 24769 31435 24803
rect 31493 24769 31527 24803
rect 31585 24769 31619 24803
rect 31769 24769 31803 24803
rect 31953 24769 31987 24803
rect 1869 24701 1903 24735
rect 2145 24701 2179 24735
rect 9229 24701 9263 24735
rect 10977 24701 11011 24735
rect 11805 24701 11839 24735
rect 11897 24701 11931 24735
rect 15025 24701 15059 24735
rect 21005 24701 21039 24735
rect 21833 24701 21867 24735
rect 24409 24701 24443 24735
rect 24593 24701 24627 24735
rect 27077 24701 27111 24735
rect 28089 24701 28123 24735
rect 28825 24701 28859 24735
rect 30205 24701 30239 24735
rect 4077 24633 4111 24667
rect 23949 24633 23983 24667
rect 29193 24633 29227 24667
rect 29285 24633 29319 24667
rect 6377 24565 6411 24599
rect 6561 24565 6595 24599
rect 10609 24565 10643 24599
rect 11345 24565 11379 24599
rect 12357 24565 12391 24599
rect 21557 24565 21591 24599
rect 23581 24565 23615 24599
rect 30481 24565 30515 24599
rect 4721 24361 4755 24395
rect 8033 24361 8067 24395
rect 11621 24361 11655 24395
rect 15485 24361 15519 24395
rect 17785 24361 17819 24395
rect 19257 24361 19291 24395
rect 21281 24361 21315 24395
rect 31401 24361 31435 24395
rect 31585 24361 31619 24395
rect 32597 24361 32631 24395
rect 11805 24293 11839 24327
rect 17233 24293 17267 24327
rect 26617 24293 26651 24327
rect 31769 24293 31803 24327
rect 4997 24225 5031 24259
rect 5825 24225 5859 24259
rect 6285 24225 6319 24259
rect 18797 24225 18831 24259
rect 24593 24225 24627 24259
rect 27261 24225 27295 24259
rect 4537 24157 4571 24191
rect 4813 24157 4847 24191
rect 4905 24157 4939 24191
rect 5089 24157 5123 24191
rect 11437 24157 11471 24191
rect 11713 24157 11747 24191
rect 12081 24157 12115 24191
rect 15669 24157 15703 24191
rect 17509 24157 17543 24191
rect 18705 24157 18739 24191
rect 19533 24157 19567 24191
rect 21097 24157 21131 24191
rect 26801 24157 26835 24191
rect 26985 24157 27019 24191
rect 27169 24157 27203 24191
rect 29561 24157 29595 24191
rect 31493 24157 31527 24191
rect 32045 24157 32079 24191
rect 34345 24157 34379 24191
rect 5273 24089 5307 24123
rect 6561 24089 6595 24123
rect 11805 24089 11839 24123
rect 17601 24089 17635 24123
rect 19625 24089 19659 24123
rect 19809 24089 19843 24123
rect 24869 24089 24903 24123
rect 26893 24089 26927 24123
rect 30297 24089 30331 24123
rect 34069 24089 34103 24123
rect 4353 24021 4387 24055
rect 11253 24021 11287 24055
rect 11989 24021 12023 24055
rect 17417 24021 17451 24055
rect 18337 24021 18371 24055
rect 19441 24021 19475 24055
rect 26341 24021 26375 24055
rect 27905 24021 27939 24055
rect 31033 24021 31067 24055
rect 5549 23817 5583 23851
rect 6561 23817 6595 23851
rect 12081 23817 12115 23851
rect 19349 23817 19383 23851
rect 19533 23817 19567 23851
rect 24777 23817 24811 23851
rect 27629 23817 27663 23851
rect 32689 23817 32723 23851
rect 33241 23817 33275 23851
rect 4077 23749 4111 23783
rect 13185 23749 13219 23783
rect 18981 23749 19015 23783
rect 25881 23749 25915 23783
rect 32321 23749 32355 23783
rect 3801 23681 3835 23715
rect 6745 23681 6779 23715
rect 8493 23681 8527 23715
rect 12633 23681 12667 23715
rect 12909 23681 12943 23715
rect 19165 23681 19199 23715
rect 19441 23681 19475 23715
rect 19625 23681 19659 23715
rect 22109 23681 22143 23715
rect 22385 23681 22419 23715
rect 25329 23681 25363 23715
rect 27445 23681 27479 23715
rect 27721 23681 27755 23715
rect 29745 23681 29779 23715
rect 29929 23681 29963 23715
rect 30021 23681 30055 23715
rect 30113 23681 30147 23715
rect 30297 23681 30331 23715
rect 32137 23681 32171 23715
rect 32413 23681 32447 23715
rect 32505 23681 32539 23715
rect 32781 23681 32815 23715
rect 32873 23681 32907 23715
rect 33057 23681 33091 23715
rect 8769 23613 8803 23647
rect 22661 23613 22695 23647
rect 24593 23613 24627 23647
rect 24685 23613 24719 23647
rect 27905 23613 27939 23647
rect 28549 23613 28583 23647
rect 22293 23545 22327 23579
rect 24133 23545 24167 23579
rect 10241 23477 10275 23511
rect 14657 23477 14691 23511
rect 25145 23477 25179 23511
rect 27261 23477 27295 23511
rect 29561 23477 29595 23511
rect 12357 23273 12391 23307
rect 21649 23273 21683 23307
rect 22477 23273 22511 23307
rect 24777 23273 24811 23307
rect 28365 23273 28399 23307
rect 19073 23205 19107 23239
rect 28273 23205 28307 23239
rect 10609 23137 10643 23171
rect 10885 23137 10919 23171
rect 18429 23137 18463 23171
rect 18797 23137 18831 23171
rect 23029 23137 23063 23171
rect 26525 23137 26559 23171
rect 26801 23137 26835 23171
rect 28917 23137 28951 23171
rect 30021 23137 30055 23171
rect 30389 23137 30423 23171
rect 30665 23137 30699 23171
rect 31217 23137 31251 23171
rect 5089 23069 5123 23103
rect 5273 23069 5307 23103
rect 5641 23069 5675 23103
rect 6009 23069 6043 23103
rect 10149 23069 10183 23103
rect 15945 23069 15979 23103
rect 16037 23069 16071 23103
rect 16405 23069 16439 23103
rect 19625 23069 19659 23103
rect 19901 23069 19935 23103
rect 22201 23069 22235 23103
rect 22845 23069 22879 23103
rect 24961 23069 24995 23103
rect 28825 23069 28859 23103
rect 29929 23069 29963 23103
rect 31125 23069 31159 23103
rect 31309 23069 31343 23103
rect 15669 23001 15703 23035
rect 17877 23001 17911 23035
rect 18914 23001 18948 23035
rect 20177 23001 20211 23035
rect 22293 23001 22327 23035
rect 28733 23001 28767 23035
rect 30874 23001 30908 23035
rect 5181 22933 5215 22967
rect 7435 22933 7469 22967
rect 9505 22933 9539 22967
rect 14197 22933 14231 22967
rect 18705 22933 18739 22967
rect 19809 22933 19843 22967
rect 22937 22933 22971 22967
rect 29561 22933 29595 22967
rect 30757 22933 30791 22967
rect 31033 22933 31067 22967
rect 16681 22729 16715 22763
rect 16865 22729 16899 22763
rect 17417 22729 17451 22763
rect 18797 22729 18831 22763
rect 19257 22729 19291 22763
rect 29377 22729 29411 22763
rect 30021 22729 30055 22763
rect 16957 22661 16991 22695
rect 19165 22661 19199 22695
rect 31217 22661 31251 22695
rect 7021 22593 7055 22627
rect 11989 22593 12023 22627
rect 16681 22593 16715 22627
rect 17049 22593 17083 22627
rect 18981 22593 19015 22627
rect 19441 22593 19475 22627
rect 19625 22593 19659 22627
rect 20821 22593 20855 22627
rect 28641 22593 28675 22627
rect 29285 22593 29319 22627
rect 29929 22593 29963 22627
rect 30113 22593 30147 22627
rect 7297 22525 7331 22559
rect 9045 22525 9079 22559
rect 12265 22525 12299 22559
rect 14013 22525 14047 22559
rect 18061 22525 18095 22559
rect 20913 22525 20947 22559
rect 24777 22525 24811 22559
rect 28733 22525 28767 22559
rect 33977 22525 34011 22559
rect 34253 22525 34287 22559
rect 21189 22457 21223 22491
rect 29009 22457 29043 22491
rect 31401 22457 31435 22491
rect 24133 22389 24167 22423
rect 32505 22389 32539 22423
rect 6193 22185 6227 22219
rect 12173 22185 12207 22219
rect 15595 22185 15629 22219
rect 32229 22185 32263 22219
rect 6561 22049 6595 22083
rect 8217 22049 8251 22083
rect 8677 22049 8711 22083
rect 9321 22049 9355 22083
rect 12725 22049 12759 22083
rect 23121 22049 23155 22083
rect 24869 22049 24903 22083
rect 28273 22049 28307 22083
rect 33333 22049 33367 22083
rect 33517 22049 33551 22083
rect 3801 21981 3835 22015
rect 6377 21981 6411 22015
rect 6653 21981 6687 22015
rect 7113 21981 7147 22015
rect 7757 21981 7791 22015
rect 8402 21981 8436 22015
rect 8553 21981 8587 22015
rect 8769 21981 8803 22015
rect 11989 21981 12023 22015
rect 12633 21981 12667 22015
rect 12909 21981 12943 22015
rect 13001 21981 13035 22015
rect 15853 21981 15887 22015
rect 18981 21981 19015 22015
rect 24041 21981 24075 22015
rect 24593 21981 24627 22015
rect 31309 21981 31343 22015
rect 31677 21981 31711 22015
rect 32413 21981 32447 22015
rect 32689 21981 32723 22015
rect 4077 21913 4111 21947
rect 5825 21913 5859 21947
rect 9597 21913 9631 21947
rect 11345 21913 11379 21947
rect 12265 21913 12299 21947
rect 12449 21913 12483 21947
rect 23397 21913 23431 21947
rect 25145 21913 25179 21947
rect 31493 21913 31527 21947
rect 31585 21913 31619 21947
rect 14105 21845 14139 21879
rect 18797 21845 18831 21879
rect 23305 21845 23339 21879
rect 23765 21845 23799 21879
rect 23857 21845 23891 21879
rect 24777 21845 24811 21879
rect 26617 21845 26651 21879
rect 28917 21845 28951 21879
rect 31861 21845 31895 21879
rect 32597 21845 32631 21879
rect 32873 21845 32907 21879
rect 33241 21845 33275 21879
rect 4813 21641 4847 21675
rect 7205 21641 7239 21675
rect 9597 21641 9631 21675
rect 10057 21641 10091 21675
rect 12909 21641 12943 21675
rect 20085 21641 20119 21675
rect 24869 21641 24903 21675
rect 25329 21641 25363 21675
rect 30389 21641 30423 21675
rect 31033 21641 31067 21675
rect 7941 21573 7975 21607
rect 9781 21573 9815 21607
rect 12357 21573 12391 21607
rect 12449 21573 12483 21607
rect 15301 21573 15335 21607
rect 17877 21573 17911 21607
rect 18613 21573 18647 21607
rect 21490 21573 21524 21607
rect 22017 21573 22051 21607
rect 25421 21573 25455 21607
rect 31401 21573 31435 21607
rect 4997 21505 5031 21539
rect 5089 21505 5123 21539
rect 5365 21505 5399 21539
rect 5549 21505 5583 21539
rect 5733 21505 5767 21539
rect 7389 21505 7423 21539
rect 7481 21505 7515 21539
rect 7757 21505 7791 21539
rect 7849 21505 7883 21539
rect 8033 21505 8067 21539
rect 9045 21505 9079 21539
rect 9321 21505 9355 21539
rect 9413 21505 9447 21539
rect 9689 21505 9723 21539
rect 9873 21505 9907 21539
rect 9965 21505 9999 21539
rect 10149 21505 10183 21539
rect 12173 21505 12207 21539
rect 12541 21505 12575 21539
rect 12817 21505 12851 21539
rect 13001 21505 13035 21539
rect 16313 21505 16347 21539
rect 17601 21505 17635 21539
rect 18337 21505 18371 21539
rect 20361 21505 20395 21539
rect 21373 21505 21407 21539
rect 21833 21505 21867 21539
rect 22201 21505 22235 21539
rect 26617 21505 26651 21539
rect 26985 21505 27019 21539
rect 29929 21505 29963 21539
rect 30481 21505 30515 21539
rect 31309 21505 31343 21539
rect 31677 21505 31711 21539
rect 32321 21505 32355 21539
rect 34345 21505 34379 21539
rect 5641 21437 5675 21471
rect 14841 21437 14875 21471
rect 17969 21437 18003 21471
rect 18086 21437 18120 21471
rect 20637 21437 20671 21471
rect 21005 21437 21039 21471
rect 21281 21437 21315 21471
rect 23121 21437 23155 21471
rect 23397 21437 23431 21471
rect 25605 21437 25639 21471
rect 27261 21437 27295 21471
rect 28733 21437 28767 21471
rect 29377 21437 29411 21471
rect 30757 21437 30791 21471
rect 31493 21437 31527 21471
rect 32229 21437 32263 21471
rect 32689 21437 32723 21471
rect 12725 21369 12759 21403
rect 15025 21369 15059 21403
rect 18245 21369 18279 21403
rect 24961 21369 24995 21403
rect 26801 21369 26835 21403
rect 5273 21301 5307 21335
rect 7665 21301 7699 21335
rect 9137 21301 9171 21335
rect 16129 21301 16163 21335
rect 20729 21301 20763 21335
rect 20913 21301 20947 21335
rect 21649 21301 21683 21335
rect 28825 21301 28859 21335
rect 30205 21301 30239 21335
rect 30573 21301 30607 21335
rect 34161 21301 34195 21335
rect 9873 21097 9907 21131
rect 13657 21097 13691 21131
rect 15840 21097 15874 21131
rect 17509 21097 17543 21131
rect 18981 21097 19015 21131
rect 20453 21097 20487 21131
rect 22109 21097 22143 21131
rect 26709 21097 26743 21131
rect 30205 21097 30239 21131
rect 30665 21097 30699 21131
rect 30849 21097 30883 21131
rect 31217 21097 31251 21131
rect 20269 21029 20303 21063
rect 22845 21029 22879 21063
rect 30573 21029 30607 21063
rect 11897 20961 11931 20995
rect 13921 20961 13955 20995
rect 15577 20961 15611 20995
rect 20821 20961 20855 20995
rect 21005 20961 21039 20995
rect 23305 20961 23339 20995
rect 27261 20961 27295 20995
rect 34069 20961 34103 20995
rect 34345 20961 34379 20995
rect 7297 20893 7331 20927
rect 11345 20893 11379 20927
rect 11529 20893 11563 20927
rect 17668 20893 17702 20927
rect 18153 20893 18187 20927
rect 18613 20893 18647 20927
rect 20177 20893 20211 20927
rect 20361 20893 20395 20927
rect 20453 20893 20487 20927
rect 20637 20893 20671 20927
rect 21189 20893 21223 20927
rect 21649 20893 21683 20927
rect 21741 20893 21775 20927
rect 22293 20893 22327 20927
rect 22661 20893 22695 20927
rect 22937 20893 22971 20927
rect 23121 20893 23155 20927
rect 23213 20893 23247 20927
rect 25053 20893 25087 20927
rect 25605 20893 25639 20927
rect 27077 20893 27111 20927
rect 28733 20893 28767 20927
rect 30113 20893 30147 20927
rect 31125 20893 31159 20927
rect 31309 20893 31343 20927
rect 4997 20825 5031 20859
rect 17877 20825 17911 20859
rect 18797 20825 18831 20859
rect 22477 20825 22511 20859
rect 22569 20825 22603 20859
rect 27169 20825 27203 20859
rect 30833 20825 30867 20859
rect 31033 20825 31067 20859
rect 4905 20757 4939 20791
rect 7113 20757 7147 20791
rect 17325 20757 17359 20791
rect 17785 20757 17819 20791
rect 23029 20757 23063 20791
rect 24409 20757 24443 20791
rect 25421 20757 25455 20791
rect 28181 20757 28215 20791
rect 32597 20757 32631 20791
rect 4997 20553 5031 20587
rect 6745 20553 6779 20587
rect 11621 20553 11655 20587
rect 17509 20553 17543 20587
rect 18153 20553 18187 20587
rect 22017 20553 22051 20587
rect 30481 20553 30515 20587
rect 32781 20553 32815 20587
rect 5365 20485 5399 20519
rect 9965 20485 9999 20519
rect 10793 20485 10827 20519
rect 17141 20485 17175 20519
rect 18305 20485 18339 20519
rect 18521 20485 18555 20519
rect 25329 20485 25363 20519
rect 4077 20417 4111 20451
rect 4537 20417 4571 20451
rect 5181 20417 5215 20451
rect 5549 20417 5583 20451
rect 5641 20417 5675 20451
rect 6377 20417 6411 20451
rect 6561 20417 6595 20451
rect 6653 20417 6687 20451
rect 6929 20417 6963 20451
rect 7021 20417 7055 20451
rect 7205 20417 7239 20451
rect 7297 20417 7331 20451
rect 7389 20417 7423 20451
rect 7481 20417 7515 20451
rect 8033 20417 8067 20451
rect 8953 20417 8987 20451
rect 9321 20417 9355 20451
rect 10149 20417 10183 20451
rect 10425 20417 10459 20451
rect 10701 20417 10735 20451
rect 10885 20417 10919 20451
rect 11713 20417 11747 20451
rect 12265 20417 12299 20451
rect 12461 20417 12495 20451
rect 16129 20417 16163 20451
rect 17325 20417 17359 20451
rect 21833 20417 21867 20451
rect 22201 20417 22235 20451
rect 22477 20417 22511 20451
rect 22569 20417 22603 20451
rect 22753 20417 22787 20451
rect 25053 20417 25087 20451
rect 27905 20417 27939 20451
rect 30010 20415 30044 20449
rect 33149 20417 33183 20451
rect 1961 20349 1995 20383
rect 2329 20349 2363 20383
rect 4629 20349 4663 20383
rect 4813 20349 4847 20383
rect 7941 20349 7975 20383
rect 9413 20349 9447 20383
rect 9781 20349 9815 20383
rect 10241 20349 10275 20383
rect 15853 20349 15887 20383
rect 33241 20349 33275 20383
rect 33425 20349 33459 20383
rect 8769 20281 8803 20315
rect 4169 20213 4203 20247
rect 5549 20213 5583 20247
rect 6469 20213 6503 20247
rect 7573 20213 7607 20247
rect 7757 20213 7791 20247
rect 10609 20213 10643 20247
rect 12449 20213 12483 20247
rect 14381 20213 14415 20247
rect 18337 20213 18371 20247
rect 22293 20213 22327 20247
rect 22661 20213 22695 20247
rect 26801 20213 26835 20247
rect 28168 20213 28202 20247
rect 29653 20213 29687 20247
rect 30297 20213 30331 20247
rect 2697 20009 2731 20043
rect 4353 20009 4387 20043
rect 4537 20009 4571 20043
rect 5089 20009 5123 20043
rect 7113 20009 7147 20043
rect 7297 20009 7331 20043
rect 13369 20009 13403 20043
rect 17141 20009 17175 20043
rect 17325 20009 17359 20043
rect 22569 20009 22603 20043
rect 25329 20009 25363 20043
rect 28089 20009 28123 20043
rect 30021 20009 30055 20043
rect 10057 19941 10091 19975
rect 27445 19941 27479 19975
rect 17417 19873 17451 19907
rect 20821 19873 20855 19907
rect 21097 19873 21131 19907
rect 23581 19873 23615 19907
rect 25973 19873 26007 19907
rect 28457 19873 28491 19907
rect 28549 19873 28583 19907
rect 1409 19805 1443 19839
rect 2881 19805 2915 19839
rect 3985 19805 4019 19839
rect 4353 19805 4387 19839
rect 4721 19805 4755 19839
rect 4905 19805 4939 19839
rect 5273 19805 5307 19839
rect 5549 19805 5583 19839
rect 5733 19805 5767 19839
rect 5917 19805 5951 19839
rect 7021 19805 7055 19839
rect 7205 19805 7239 19839
rect 7408 19805 7442 19839
rect 7573 19805 7607 19839
rect 8585 19805 8619 19839
rect 8769 19805 8803 19839
rect 9505 19805 9539 19839
rect 9873 19805 9907 19839
rect 10149 19805 10183 19839
rect 10333 19805 10367 19839
rect 10517 19805 10551 19839
rect 10977 19805 11011 19839
rect 13277 19805 13311 19839
rect 17785 19805 17819 19839
rect 22569 19805 22603 19839
rect 22753 19805 22787 19839
rect 23857 19805 23891 19839
rect 24593 19805 24627 19839
rect 24685 19805 24719 19839
rect 25697 19805 25731 19839
rect 26801 19805 26835 19839
rect 28273 19805 28307 19839
rect 28641 19805 28675 19839
rect 28825 19805 28859 19839
rect 29929 19805 29963 19839
rect 6009 19737 6043 19771
rect 9321 19737 9355 19771
rect 16957 19737 16991 19771
rect 17902 19737 17936 19771
rect 24777 19737 24811 19771
rect 25789 19737 25823 19771
rect 1593 19669 1627 19703
rect 4813 19669 4847 19703
rect 5457 19669 5491 19703
rect 8677 19669 8711 19703
rect 9137 19669 9171 19703
rect 10517 19669 10551 19703
rect 10885 19669 10919 19703
rect 17157 19669 17191 19703
rect 17693 19669 17727 19703
rect 18061 19669 18095 19703
rect 19349 19669 19383 19703
rect 23765 19669 23799 19703
rect 24225 19669 24259 19703
rect 24409 19669 24443 19703
rect 30389 19669 30423 19703
rect 3157 19465 3191 19499
rect 5181 19465 5215 19499
rect 15209 19465 15243 19499
rect 17417 19465 17451 19499
rect 31401 19465 31435 19499
rect 33149 19465 33183 19499
rect 1685 19397 1719 19431
rect 5365 19397 5399 19431
rect 9137 19397 9171 19431
rect 13737 19397 13771 19431
rect 17509 19397 17543 19431
rect 19717 19397 19751 19431
rect 1409 19329 1443 19363
rect 4261 19329 4295 19363
rect 4445 19329 4479 19363
rect 5457 19329 5491 19363
rect 7205 19329 7239 19363
rect 7389 19329 7423 19363
rect 11805 19329 11839 19363
rect 12449 19329 12483 19363
rect 12633 19329 12667 19363
rect 13093 19329 13127 19363
rect 13461 19329 13495 19363
rect 17049 19329 17083 19363
rect 17233 19329 17267 19363
rect 17693 19329 17727 19363
rect 17877 19329 17911 19363
rect 20545 19329 20579 19363
rect 20729 19329 20763 19363
rect 20821 19329 20855 19363
rect 21005 19329 21039 19363
rect 26525 19329 26559 19363
rect 26985 19329 27019 19363
rect 30021 19329 30055 19363
rect 31217 19329 31251 19363
rect 31493 19329 31527 19363
rect 31585 19329 31619 19363
rect 31769 19329 31803 19363
rect 32781 19329 32815 19363
rect 4629 19261 4663 19295
rect 4813 19261 4847 19295
rect 4997 19261 5031 19295
rect 5089 19261 5123 19295
rect 8493 19261 8527 19295
rect 12265 19261 12299 19295
rect 20361 19261 20395 19295
rect 23489 19261 23523 19295
rect 23765 19261 23799 19295
rect 25237 19261 25271 19295
rect 27261 19261 27295 19295
rect 28733 19261 28767 19295
rect 31033 19261 31067 19295
rect 31677 19261 31711 19295
rect 32689 19261 32723 19295
rect 26709 19193 26743 19227
rect 7573 19125 7607 19159
rect 18245 19125 18279 19159
rect 20821 19125 20855 19159
rect 30205 19125 30239 19159
rect 30481 19125 30515 19159
rect 18613 18921 18647 18955
rect 23213 18921 23247 18955
rect 26341 18921 26375 18955
rect 29929 18921 29963 18955
rect 31217 18921 31251 18955
rect 32781 18921 32815 18955
rect 8585 18853 8619 18887
rect 15577 18853 15611 18887
rect 21833 18853 21867 18887
rect 30941 18853 30975 18887
rect 32413 18853 32447 18887
rect 33701 18853 33735 18887
rect 1593 18785 1627 18819
rect 9045 18785 9079 18819
rect 12173 18785 12207 18819
rect 23121 18785 23155 18819
rect 23673 18785 23707 18819
rect 26801 18785 26835 18819
rect 26893 18785 26927 18819
rect 28457 18785 28491 18819
rect 6837 18717 6871 18751
rect 7389 18717 7423 18751
rect 7757 18717 7791 18751
rect 8401 18717 8435 18751
rect 9799 18717 9833 18751
rect 9965 18717 9999 18751
rect 10701 18717 10735 18751
rect 11069 18717 11103 18751
rect 12817 18717 12851 18751
rect 13369 18717 13403 18751
rect 13737 18717 13771 18751
rect 15761 18717 15795 18751
rect 16037 18717 16071 18751
rect 16313 18717 16347 18751
rect 16497 18717 16531 18751
rect 18429 18717 18463 18751
rect 18705 18717 18739 18751
rect 20545 18717 20579 18751
rect 22017 18717 22051 18751
rect 22109 18717 22143 18751
rect 22201 18717 22235 18751
rect 22569 18717 22603 18751
rect 22845 18717 22879 18751
rect 23581 18717 23615 18751
rect 24409 18717 24443 18751
rect 28641 18717 28675 18751
rect 30067 18717 30101 18751
rect 30297 18717 30331 18751
rect 30480 18717 30514 18751
rect 30573 18717 30607 18751
rect 30665 18717 30699 18751
rect 31401 18717 31435 18751
rect 31585 18717 31619 18751
rect 31677 18717 31711 18751
rect 31769 18717 31803 18751
rect 32413 18717 32447 18751
rect 32685 18695 32719 18729
rect 32965 18717 32999 18751
rect 33241 18717 33275 18751
rect 33333 18717 33367 18751
rect 1869 18649 1903 18683
rect 3617 18649 3651 18683
rect 8033 18649 8067 18683
rect 9321 18649 9355 18683
rect 12633 18649 12667 18683
rect 16681 18649 16715 18683
rect 19993 18649 20027 18683
rect 21833 18649 21867 18683
rect 22385 18649 22419 18683
rect 22477 18649 22511 18683
rect 26709 18649 26743 18683
rect 27813 18649 27847 18683
rect 30205 18649 30239 18683
rect 33517 18649 33551 18683
rect 7389 18581 7423 18615
rect 9229 18581 9263 18615
rect 9689 18581 9723 18615
rect 10149 18581 10183 18615
rect 18889 18581 18923 18615
rect 22753 18581 22787 18615
rect 23397 18581 23431 18615
rect 24593 18581 24627 18615
rect 29193 18581 29227 18615
rect 31125 18581 31159 18615
rect 31861 18581 31895 18615
rect 32597 18581 32631 18615
rect 33149 18581 33183 18615
rect 3433 18377 3467 18411
rect 5381 18377 5415 18411
rect 6101 18377 6135 18411
rect 9413 18377 9447 18411
rect 15485 18377 15519 18411
rect 17877 18377 17911 18411
rect 18245 18377 18279 18411
rect 32781 18377 32815 18411
rect 3801 18309 3835 18343
rect 5181 18309 5215 18343
rect 8125 18309 8159 18343
rect 8953 18309 8987 18343
rect 9597 18309 9631 18343
rect 11805 18309 11839 18343
rect 16129 18309 16163 18343
rect 17969 18309 18003 18343
rect 18797 18309 18831 18343
rect 24501 18309 24535 18343
rect 3617 18241 3651 18275
rect 3709 18241 3743 18275
rect 3985 18241 4019 18275
rect 5641 18241 5675 18275
rect 5917 18241 5951 18275
rect 6469 18241 6503 18275
rect 6837 18241 6871 18275
rect 7573 18241 7607 18275
rect 7849 18241 7883 18275
rect 9045 18241 9079 18275
rect 9137 18241 9171 18275
rect 9781 18241 9815 18275
rect 9873 18241 9907 18275
rect 11529 18241 11563 18275
rect 12541 18241 12575 18275
rect 12725 18241 12759 18275
rect 12817 18241 12851 18275
rect 12909 18241 12943 18275
rect 13277 18241 13311 18275
rect 13645 18241 13679 18275
rect 14197 18241 14231 18275
rect 14657 18241 14691 18275
rect 15117 18241 15151 18275
rect 15209 18241 15243 18275
rect 15945 18241 15979 18275
rect 17601 18241 17635 18275
rect 22385 18241 22419 18275
rect 22477 18241 22511 18275
rect 22753 18241 22787 18275
rect 22937 18241 22971 18275
rect 23305 18241 23339 18275
rect 23581 18241 23615 18275
rect 23673 18241 23707 18275
rect 23949 18241 23983 18275
rect 29745 18241 29779 18275
rect 29929 18241 29963 18275
rect 32689 18241 32723 18275
rect 32873 18241 32907 18275
rect 7941 18173 7975 18207
rect 11621 18173 11655 18207
rect 11805 18173 11839 18207
rect 14473 18173 14507 18207
rect 15025 18173 15059 18207
rect 15301 18173 15335 18207
rect 18086 18173 18120 18207
rect 18521 18173 18555 18207
rect 23397 18173 23431 18207
rect 24225 18173 24259 18207
rect 25973 18173 26007 18207
rect 27169 18173 27203 18207
rect 30205 18173 30239 18207
rect 5733 18105 5767 18139
rect 12817 18105 12851 18139
rect 14381 18105 14415 18139
rect 20269 18105 20303 18139
rect 5365 18037 5399 18071
rect 5549 18037 5583 18071
rect 9229 18037 9263 18071
rect 9597 18037 9631 18071
rect 14841 18037 14875 18071
rect 16313 18037 16347 18071
rect 21925 18037 21959 18071
rect 23857 18037 23891 18071
rect 27813 18037 27847 18071
rect 27997 18037 28031 18071
rect 29481 18037 29515 18071
rect 4537 17833 4571 17867
rect 10885 17833 10919 17867
rect 14841 17833 14875 17867
rect 16313 17833 16347 17867
rect 18337 17833 18371 17867
rect 20361 17833 20395 17867
rect 21373 17833 21407 17867
rect 22569 17833 22603 17867
rect 23305 17833 23339 17867
rect 24409 17833 24443 17867
rect 28733 17833 28767 17867
rect 31677 17833 31711 17867
rect 32597 17833 32631 17867
rect 33149 17833 33183 17867
rect 7389 17765 7423 17799
rect 18153 17765 18187 17799
rect 21557 17765 21591 17799
rect 3525 17697 3559 17731
rect 4997 17697 5031 17731
rect 7941 17697 7975 17731
rect 10977 17697 11011 17731
rect 13185 17697 13219 17731
rect 19993 17697 20027 17731
rect 24869 17697 24903 17731
rect 24961 17697 24995 17731
rect 26065 17697 26099 17731
rect 32689 17697 32723 17731
rect 3433 17629 3467 17663
rect 3617 17629 3651 17663
rect 3985 17629 4019 17663
rect 4169 17629 4203 17663
rect 4353 17629 4387 17663
rect 4445 17629 4479 17663
rect 4629 17629 4663 17663
rect 5273 17629 5307 17663
rect 6653 17629 6687 17663
rect 7297 17629 7331 17663
rect 7481 17629 7515 17663
rect 8769 17629 8803 17663
rect 8953 17629 8987 17663
rect 9229 17629 9263 17663
rect 9413 17629 9447 17663
rect 9505 17629 9539 17663
rect 9689 17629 9723 17663
rect 10701 17629 10735 17663
rect 10793 17629 10827 17663
rect 11069 17629 11103 17663
rect 11253 17629 11287 17663
rect 11437 17629 11471 17663
rect 11529 17629 11563 17663
rect 11621 17629 11655 17663
rect 13921 17629 13955 17663
rect 14565 17629 14599 17663
rect 14841 17629 14875 17663
rect 15853 17629 15887 17663
rect 16129 17629 16163 17663
rect 16497 17629 16531 17663
rect 16773 17629 16807 17663
rect 17325 17629 17359 17663
rect 18061 17629 18095 17663
rect 20177 17629 20211 17663
rect 20913 17629 20947 17663
rect 21005 17629 21039 17663
rect 21189 17629 21223 17663
rect 21465 17629 21499 17663
rect 21649 17629 21683 17663
rect 22753 17629 22787 17663
rect 23055 17629 23089 17663
rect 23213 17629 23247 17663
rect 23581 17629 23615 17663
rect 23857 17629 23891 17663
rect 24777 17629 24811 17663
rect 26893 17629 26927 17663
rect 27997 17629 28031 17663
rect 28181 17629 28215 17663
rect 28273 17629 28307 17663
rect 28365 17629 28399 17663
rect 28549 17629 28583 17663
rect 31953 17629 31987 17663
rect 32045 17629 32079 17663
rect 32137 17629 32171 17663
rect 32321 17629 32355 17663
rect 32597 17629 32631 17663
rect 33149 17629 33183 17663
rect 33241 17629 33275 17663
rect 4077 17561 4111 17595
rect 11897 17561 11931 17595
rect 17693 17561 17727 17595
rect 17877 17561 17911 17595
rect 18521 17561 18555 17595
rect 22845 17561 22879 17595
rect 22937 17561 22971 17595
rect 23305 17561 23339 17595
rect 23949 17561 23983 17595
rect 26157 17561 26191 17595
rect 26249 17561 26283 17595
rect 33057 17561 33091 17595
rect 3801 17493 3835 17527
rect 5917 17493 5951 17527
rect 9045 17493 9079 17527
rect 9597 17493 9631 17527
rect 14657 17493 14691 17527
rect 15945 17493 15979 17527
rect 17417 17493 17451 17527
rect 18321 17493 18355 17527
rect 23489 17493 23523 17527
rect 26617 17493 26651 17527
rect 26709 17493 26743 17527
rect 32413 17493 32447 17527
rect 33517 17493 33551 17527
rect 7849 17289 7883 17323
rect 12166 17289 12200 17323
rect 13553 17289 13587 17323
rect 17969 17289 18003 17323
rect 28273 17289 28307 17323
rect 31585 17289 31619 17323
rect 32873 17289 32907 17323
rect 12081 17221 12115 17255
rect 12909 17221 12943 17255
rect 17601 17221 17635 17255
rect 18429 17221 18463 17255
rect 33793 17221 33827 17255
rect 3433 17153 3467 17187
rect 3525 17153 3559 17187
rect 3617 17153 3651 17187
rect 3755 17153 3789 17187
rect 4997 17153 5031 17187
rect 5181 17153 5215 17187
rect 5273 17153 5307 17187
rect 7389 17153 7423 17187
rect 7573 17153 7607 17187
rect 7665 17153 7699 17187
rect 8033 17153 8067 17187
rect 9229 17153 9263 17187
rect 9505 17153 9539 17187
rect 9597 17153 9631 17187
rect 10885 17153 10919 17187
rect 11069 17153 11103 17187
rect 11161 17153 11195 17187
rect 11713 17153 11747 17187
rect 11897 17153 11931 17187
rect 11989 17153 12023 17187
rect 12265 17153 12299 17187
rect 12449 17153 12483 17187
rect 12633 17153 12667 17187
rect 12725 17153 12759 17187
rect 13093 17153 13127 17187
rect 13277 17153 13311 17187
rect 13645 17153 13679 17187
rect 13829 17153 13863 17187
rect 13921 17153 13955 17187
rect 14933 17153 14967 17187
rect 15577 17153 15611 17187
rect 17417 17153 17451 17187
rect 17693 17153 17727 17187
rect 18061 17153 18095 17187
rect 18613 17153 18647 17187
rect 21005 17153 21039 17187
rect 21189 17153 21223 17187
rect 28457 17153 28491 17187
rect 28549 17153 28583 17187
rect 28733 17153 28767 17187
rect 28825 17153 28859 17187
rect 29745 17153 29779 17187
rect 29929 17153 29963 17187
rect 30205 17153 30239 17187
rect 30389 17153 30423 17187
rect 31033 17153 31067 17187
rect 31125 17153 31159 17187
rect 31309 17153 31343 17187
rect 31401 17153 31435 17187
rect 32689 17153 32723 17187
rect 32965 17153 32999 17187
rect 33149 17153 33183 17187
rect 33701 17153 33735 17187
rect 33885 17153 33919 17187
rect 1409 17085 1443 17119
rect 1685 17085 1719 17119
rect 3249 17085 3283 17119
rect 3893 17085 3927 17119
rect 5089 17085 5123 17119
rect 7481 17085 7515 17119
rect 8125 17085 8159 17119
rect 13185 17085 13219 17119
rect 13369 17085 13403 17119
rect 15209 17085 15243 17119
rect 17233 17085 17267 17119
rect 18178 17085 18212 17119
rect 11345 17017 11379 17051
rect 12541 17017 12575 17051
rect 13645 17017 13679 17051
rect 30113 17017 30147 17051
rect 3157 16949 3191 16983
rect 5457 16949 5491 16983
rect 8217 16949 8251 16983
rect 8401 16949 8435 16983
rect 9321 16949 9355 16983
rect 9781 16949 9815 16983
rect 10885 16949 10919 16983
rect 11805 16949 11839 16983
rect 15301 16949 15335 16983
rect 15485 16949 15519 16983
rect 15669 16949 15703 16983
rect 18337 16949 18371 16983
rect 18797 16949 18831 16983
rect 21189 16949 21223 16983
rect 30297 16949 30331 16983
rect 5622 16745 5656 16779
rect 5917 16745 5951 16779
rect 6929 16745 6963 16779
rect 7481 16745 7515 16779
rect 13553 16745 13587 16779
rect 13921 16745 13955 16779
rect 15301 16745 15335 16779
rect 16129 16745 16163 16779
rect 21465 16745 21499 16779
rect 21833 16745 21867 16779
rect 22937 16745 22971 16779
rect 26144 16745 26178 16779
rect 27629 16745 27663 16779
rect 29285 16745 29319 16779
rect 30757 16745 30791 16779
rect 31125 16745 31159 16779
rect 31309 16745 31343 16779
rect 31677 16745 31711 16779
rect 32413 16745 32447 16779
rect 33793 16745 33827 16779
rect 5733 16677 5767 16711
rect 6745 16677 6779 16711
rect 7389 16677 7423 16711
rect 5825 16609 5859 16643
rect 8125 16609 8159 16643
rect 8585 16609 8619 16643
rect 12633 16609 12667 16643
rect 13829 16609 13863 16643
rect 15117 16609 15151 16643
rect 20361 16609 20395 16643
rect 21373 16609 21407 16643
rect 22569 16609 22603 16643
rect 24869 16609 24903 16643
rect 24961 16609 24995 16643
rect 25881 16609 25915 16643
rect 30573 16609 30607 16643
rect 32505 16609 32539 16643
rect 33517 16609 33551 16643
rect 33977 16609 34011 16643
rect 3341 16541 3375 16575
rect 5457 16541 5491 16575
rect 6285 16541 6319 16575
rect 6561 16541 6595 16575
rect 6745 16541 6779 16575
rect 6837 16541 6871 16575
rect 7113 16541 7147 16575
rect 7205 16541 7239 16575
rect 7665 16541 7699 16575
rect 7757 16541 7791 16575
rect 7849 16541 7883 16575
rect 7941 16541 7975 16575
rect 8309 16541 8343 16575
rect 8493 16541 8527 16575
rect 9505 16541 9539 16575
rect 9597 16541 9631 16575
rect 9781 16541 9815 16575
rect 13461 16541 13495 16575
rect 13737 16541 13771 16575
rect 15025 16541 15059 16575
rect 15393 16541 15427 16575
rect 15761 16541 15795 16575
rect 15945 16541 15979 16575
rect 16129 16541 16163 16575
rect 18061 16541 18095 16575
rect 19993 16541 20027 16575
rect 20131 16541 20165 16575
rect 20269 16541 20303 16575
rect 20453 16541 20487 16575
rect 21649 16541 21683 16575
rect 22753 16541 22787 16575
rect 28273 16541 28307 16575
rect 29193 16541 29227 16575
rect 30941 16541 30975 16575
rect 31033 16541 31067 16575
rect 31585 16541 31619 16575
rect 31769 16541 31803 16575
rect 32597 16541 32631 16575
rect 33425 16541 33459 16575
rect 33885 16541 33919 16575
rect 34069 16541 34103 16575
rect 3065 16473 3099 16507
rect 13369 16473 13403 16507
rect 15301 16473 15335 16507
rect 31277 16473 31311 16507
rect 31493 16473 31527 16507
rect 6377 16405 6411 16439
rect 9965 16405 9999 16439
rect 14841 16405 14875 16439
rect 18245 16405 18279 16439
rect 24409 16405 24443 16439
rect 24777 16405 24811 16439
rect 27721 16405 27755 16439
rect 32229 16405 32263 16439
rect 3249 16201 3283 16235
rect 4813 16201 4847 16235
rect 5457 16201 5491 16235
rect 8585 16201 8619 16235
rect 9505 16201 9539 16235
rect 13277 16201 13311 16235
rect 19993 16201 20027 16235
rect 22201 16201 22235 16235
rect 23489 16201 23523 16235
rect 26801 16201 26835 16235
rect 31493 16201 31527 16235
rect 5825 16133 5859 16167
rect 8401 16133 8435 16167
rect 18521 16133 18555 16167
rect 27445 16133 27479 16167
rect 29745 16133 29779 16167
rect 32321 16133 32355 16167
rect 32689 16133 32723 16167
rect 32873 16133 32907 16167
rect 2881 16065 2915 16099
rect 4169 16065 4203 16099
rect 4353 16065 4387 16099
rect 4721 16065 4755 16099
rect 4997 16065 5031 16099
rect 5273 16065 5307 16099
rect 8217 16065 8251 16099
rect 9413 16065 9447 16099
rect 9689 16065 9723 16099
rect 9873 16065 9907 16099
rect 10333 16065 10367 16099
rect 10517 16065 10551 16099
rect 10701 16065 10735 16099
rect 10885 16065 10919 16099
rect 13185 16065 13219 16099
rect 13369 16065 13403 16099
rect 15209 16065 15243 16099
rect 15393 16065 15427 16099
rect 15485 16065 15519 16099
rect 15669 16065 15703 16099
rect 22845 16065 22879 16099
rect 23029 16065 23063 16099
rect 23121 16065 23155 16099
rect 23213 16065 23247 16099
rect 23581 16065 23615 16099
rect 23765 16065 23799 16099
rect 23857 16065 23891 16099
rect 24133 16065 24167 16099
rect 27169 16065 27203 16099
rect 29648 16065 29682 16099
rect 29837 16065 29871 16099
rect 30020 16065 30054 16099
rect 30113 16065 30147 16099
rect 31309 16065 31343 16099
rect 31493 16065 31527 16099
rect 32505 16065 32539 16099
rect 32597 16065 32631 16099
rect 2973 15997 3007 16031
rect 5089 15997 5123 16031
rect 10609 15997 10643 16031
rect 15301 15997 15335 16031
rect 18245 15997 18279 16031
rect 22293 15997 22327 16031
rect 22477 15997 22511 16031
rect 23673 15997 23707 16031
rect 24409 15997 24443 16031
rect 25881 15997 25915 16031
rect 26157 15997 26191 16031
rect 21833 15929 21867 15963
rect 24041 15929 24075 15963
rect 32873 15929 32907 15963
rect 4537 15861 4571 15895
rect 5181 15861 5215 15895
rect 5733 15861 5767 15895
rect 11069 15861 11103 15895
rect 15669 15861 15703 15895
rect 28917 15861 28951 15895
rect 29469 15861 29503 15895
rect 32137 15861 32171 15895
rect 3267 15657 3301 15691
rect 7205 15657 7239 15691
rect 7389 15657 7423 15691
rect 8585 15657 8619 15691
rect 10333 15657 10367 15691
rect 10793 15657 10827 15691
rect 13277 15657 13311 15691
rect 14933 15657 14967 15691
rect 21465 15657 21499 15691
rect 22937 15657 22971 15691
rect 27721 15657 27755 15691
rect 29653 15657 29687 15691
rect 30205 15657 30239 15691
rect 30573 15657 30607 15691
rect 21097 15589 21131 15623
rect 23397 15589 23431 15623
rect 30021 15589 30055 15623
rect 3525 15521 3559 15555
rect 7573 15521 7607 15555
rect 10701 15521 10735 15555
rect 11897 15521 11931 15555
rect 16405 15521 16439 15555
rect 16497 15521 16531 15555
rect 16865 15521 16899 15555
rect 25789 15521 25823 15555
rect 28181 15521 28215 15555
rect 1501 15453 1535 15487
rect 6009 15453 6043 15487
rect 6101 15453 6135 15487
rect 7021 15453 7055 15487
rect 7205 15453 7239 15487
rect 7481 15453 7515 15487
rect 7665 15453 7699 15487
rect 7941 15453 7975 15487
rect 8034 15453 8068 15487
rect 8406 15453 8440 15487
rect 9229 15453 9263 15487
rect 9413 15453 9447 15487
rect 9505 15453 9539 15487
rect 9597 15453 9631 15487
rect 10609 15453 10643 15487
rect 10885 15453 10919 15487
rect 11069 15453 11103 15487
rect 11253 15453 11287 15487
rect 11437 15453 11471 15487
rect 11529 15453 11563 15487
rect 11621 15453 11655 15487
rect 12357 15453 12391 15487
rect 12633 15453 12667 15487
rect 12725 15453 12759 15487
rect 12909 15453 12943 15487
rect 13093 15453 13127 15487
rect 14749 15453 14783 15487
rect 14841 15453 14875 15487
rect 16589 15453 16623 15487
rect 16681 15453 16715 15487
rect 16957 15453 16991 15487
rect 17233 15453 17267 15487
rect 17417 15453 17451 15487
rect 17601 15453 17635 15487
rect 19533 15453 19567 15487
rect 19809 15453 19843 15487
rect 19993 15453 20027 15487
rect 21097 15453 21131 15487
rect 21189 15453 21223 15487
rect 21649 15453 21683 15487
rect 21741 15453 21775 15487
rect 22753 15453 22787 15487
rect 23489 15453 23523 15487
rect 23673 15453 23707 15487
rect 25513 15453 25547 15487
rect 27905 15453 27939 15487
rect 28089 15453 28123 15487
rect 28273 15453 28307 15487
rect 28457 15453 28491 15487
rect 29561 15453 29595 15487
rect 30113 15453 30147 15487
rect 6929 15385 6963 15419
rect 8217 15385 8251 15419
rect 8309 15385 8343 15419
rect 12173 15385 12207 15419
rect 13001 15385 13035 15419
rect 17877 15385 17911 15419
rect 22017 15385 22051 15419
rect 22109 15385 22143 15419
rect 22569 15385 22603 15419
rect 23029 15385 23063 15419
rect 23213 15385 23247 15419
rect 26065 15385 26099 15419
rect 9873 15317 9907 15351
rect 12541 15317 12575 15351
rect 15117 15317 15151 15351
rect 17049 15317 17083 15351
rect 19625 15317 19659 15351
rect 23581 15317 23615 15351
rect 25697 15317 25731 15351
rect 27537 15317 27571 15351
rect 3157 15113 3191 15147
rect 5733 15113 5767 15147
rect 6929 15113 6963 15147
rect 8309 15113 8343 15147
rect 9781 15113 9815 15147
rect 10885 15113 10919 15147
rect 17233 15113 17267 15147
rect 25789 15113 25823 15147
rect 26157 15113 26191 15147
rect 31401 15113 31435 15147
rect 5457 15045 5491 15079
rect 7205 15045 7239 15079
rect 7297 15045 7331 15079
rect 13829 15045 13863 15079
rect 16497 15045 16531 15079
rect 19625 15045 19659 15079
rect 26249 15045 26283 15079
rect 28273 15045 28307 15079
rect 30757 15045 30791 15079
rect 31953 15045 31987 15079
rect 33609 15045 33643 15079
rect 3341 14977 3375 15011
rect 3433 14977 3467 15011
rect 3617 14977 3651 15011
rect 4077 14977 4111 15011
rect 4261 14977 4295 15011
rect 4629 14977 4663 15011
rect 5181 14977 5215 15011
rect 7113 14977 7147 15011
rect 7389 14977 7423 15011
rect 7573 14977 7607 15011
rect 8861 14977 8895 15011
rect 9321 14977 9355 15011
rect 9597 14977 9631 15011
rect 10793 14977 10827 15011
rect 11069 14977 11103 15011
rect 12265 14977 12299 15011
rect 12449 14977 12483 15011
rect 13093 14977 13127 15011
rect 13185 14977 13219 15011
rect 13369 14977 13403 15011
rect 13461 14977 13495 15011
rect 13553 14977 13587 15011
rect 14013 14977 14047 15011
rect 14197 14977 14231 15011
rect 14289 14977 14323 15011
rect 15485 14977 15519 15011
rect 15669 14977 15703 15011
rect 16129 14977 16163 15011
rect 16313 14977 16347 15011
rect 16865 14977 16899 15011
rect 16957 14977 16991 15011
rect 17969 14977 18003 15011
rect 18337 14977 18371 15011
rect 19257 14977 19291 15011
rect 19441 14977 19475 15011
rect 19717 14977 19751 15011
rect 19809 14977 19843 15011
rect 20453 14977 20487 15011
rect 20729 14977 20763 15011
rect 21005 14977 21039 15011
rect 21097 14977 21131 15011
rect 23029 14977 23063 15011
rect 23489 14977 23523 15011
rect 23581 14977 23615 15011
rect 28457 14977 28491 15011
rect 31217 14977 31251 15011
rect 31677 14977 31711 15011
rect 33241 14977 33275 15011
rect 34345 14977 34379 15011
rect 8585 14909 8619 14943
rect 9413 14909 9447 14943
rect 16773 14909 16807 14943
rect 17049 14909 17083 14943
rect 17693 14909 17727 14943
rect 22661 14909 22695 14943
rect 23213 14909 23247 14943
rect 26341 14909 26375 14943
rect 31033 14909 31067 14943
rect 31861 14909 31895 14943
rect 3525 14841 3559 14875
rect 5181 14841 5215 14875
rect 14105 14841 14139 14875
rect 18429 14841 18463 14875
rect 20085 14841 20119 14875
rect 8493 14773 8527 14807
rect 11069 14773 11103 14807
rect 12449 14773 12483 14807
rect 13737 14773 13771 14807
rect 15577 14773 15611 14807
rect 28641 14773 28675 14807
rect 31217 14773 31251 14807
rect 31493 14773 31527 14807
rect 31861 14773 31895 14807
rect 34161 14773 34195 14807
rect 7021 14569 7055 14603
rect 13461 14569 13495 14603
rect 15209 14569 15243 14603
rect 16957 14569 16991 14603
rect 18521 14569 18555 14603
rect 19993 14569 20027 14603
rect 21005 14569 21039 14603
rect 29377 14569 29411 14603
rect 31217 14569 31251 14603
rect 34253 14569 34287 14603
rect 13553 14501 13587 14535
rect 16405 14501 16439 14535
rect 19441 14501 19475 14535
rect 19529 14501 19563 14535
rect 23397 14501 23431 14535
rect 32505 14501 32539 14535
rect 5917 14433 5951 14467
rect 7389 14433 7423 14467
rect 11345 14433 11379 14467
rect 11621 14433 11655 14467
rect 13001 14433 13035 14467
rect 17049 14433 17083 14467
rect 20637 14433 20671 14467
rect 21649 14433 21683 14467
rect 25973 14433 26007 14467
rect 26157 14433 26191 14467
rect 27629 14433 27663 14467
rect 4721 14365 4755 14399
rect 5181 14365 5215 14399
rect 6101 14365 6135 14399
rect 7205 14365 7239 14399
rect 7297 14365 7331 14399
rect 7481 14365 7515 14399
rect 7665 14365 7699 14399
rect 10977 14365 11011 14399
rect 11437 14365 11471 14399
rect 12725 14365 12759 14399
rect 12909 14365 12943 14399
rect 13093 14365 13127 14399
rect 13277 14365 13311 14399
rect 13553 14365 13587 14399
rect 13737 14365 13771 14399
rect 15393 14365 15427 14399
rect 15485 14365 15519 14399
rect 15669 14365 15703 14399
rect 15761 14365 15795 14399
rect 15853 14365 15887 14399
rect 15945 14365 15979 14399
rect 16129 14365 16163 14399
rect 16221 14365 16255 14399
rect 16957 14365 16991 14399
rect 18153 14365 18187 14399
rect 18337 14365 18371 14399
rect 19349 14365 19383 14399
rect 19625 14365 19659 14399
rect 20177 14365 20211 14399
rect 20361 14365 20395 14399
rect 20453 14365 20487 14399
rect 20821 14365 20855 14399
rect 21189 14365 21223 14399
rect 21465 14365 21499 14399
rect 21741 14365 21775 14399
rect 21925 14365 21959 14399
rect 22753 14365 22787 14399
rect 22937 14365 22971 14399
rect 23213 14365 23247 14399
rect 23305 14365 23339 14399
rect 23489 14365 23523 14399
rect 26893 14365 26927 14399
rect 31217 14365 31251 14399
rect 31493 14365 31527 14399
rect 31769 14365 31803 14399
rect 32137 14365 32171 14399
rect 32229 14365 32263 14399
rect 32505 14365 32539 14399
rect 34069 14365 34103 14399
rect 6285 14297 6319 14331
rect 18061 14297 18095 14331
rect 23121 14297 23155 14331
rect 27537 14297 27571 14331
rect 27905 14297 27939 14331
rect 31861 14297 31895 14331
rect 31953 14297 31987 14331
rect 4537 14229 4571 14263
rect 11069 14229 11103 14263
rect 11253 14229 11287 14263
rect 17325 14229 17359 14263
rect 19809 14229 19843 14263
rect 26249 14229 26283 14263
rect 26617 14229 26651 14263
rect 31401 14229 31435 14263
rect 31585 14229 31619 14263
rect 32321 14229 32355 14263
rect 4905 14025 4939 14059
rect 5457 14025 5491 14059
rect 6679 14025 6713 14059
rect 8217 14025 8251 14059
rect 10333 14025 10367 14059
rect 12909 14025 12943 14059
rect 15301 14025 15335 14059
rect 18889 14025 18923 14059
rect 25697 14025 25731 14059
rect 27905 14025 27939 14059
rect 30665 14025 30699 14059
rect 32137 14025 32171 14059
rect 4353 13957 4387 13991
rect 6469 13957 6503 13991
rect 10793 13957 10827 13991
rect 15669 13957 15703 13991
rect 16129 13957 16163 13991
rect 26709 13957 26743 13991
rect 31401 13957 31435 13991
rect 32321 13957 32355 13991
rect 3433 13889 3467 13923
rect 3985 13889 4019 13923
rect 4261 13889 4295 13923
rect 4537 13889 4571 13923
rect 4629 13889 4663 13923
rect 5089 13889 5123 13923
rect 5181 13889 5215 13923
rect 5549 13889 5583 13923
rect 6929 13889 6963 13923
rect 7113 13889 7147 13923
rect 8401 13889 8435 13923
rect 8585 13889 8619 13923
rect 8953 13889 8987 13923
rect 9689 13889 9723 13923
rect 9781 13889 9815 13923
rect 9965 13889 9999 13923
rect 10609 13889 10643 13923
rect 10701 13889 10735 13923
rect 11529 13889 11563 13923
rect 13093 13889 13127 13923
rect 13277 13889 13311 13923
rect 13737 13889 13771 13923
rect 13829 13889 13863 13923
rect 14013 13889 14047 13923
rect 14105 13889 14139 13923
rect 15485 13889 15519 13923
rect 15577 13889 15611 13923
rect 15853 13889 15887 13923
rect 15945 13889 15979 13923
rect 16037 13889 16071 13923
rect 18061 13889 18095 13923
rect 18245 13889 18279 13923
rect 18429 13889 18463 13923
rect 18613 13889 18647 13923
rect 19165 13889 19199 13923
rect 19257 13889 19291 13923
rect 20361 13889 20395 13923
rect 20545 13889 20579 13923
rect 20729 13889 20763 13923
rect 23673 13889 23707 13923
rect 23949 13889 23983 13923
rect 25881 13889 25915 13923
rect 26985 13889 27019 13923
rect 28089 13889 28123 13923
rect 28365 13889 28399 13923
rect 28457 13889 28491 13923
rect 28641 13889 28675 13923
rect 30205 13889 30239 13923
rect 31309 13889 31343 13923
rect 31493 13889 31527 13923
rect 32505 13889 32539 13923
rect 3709 13821 3743 13855
rect 4077 13821 4111 13855
rect 5641 13821 5675 13855
rect 7021 13821 7055 13855
rect 8677 13821 8711 13855
rect 8769 13821 8803 13855
rect 9045 13821 9079 13855
rect 9137 13821 9171 13855
rect 9229 13821 9263 13855
rect 10149 13821 10183 13855
rect 10333 13821 10367 13855
rect 11621 13821 11655 13855
rect 13185 13821 13219 13855
rect 13369 13821 13403 13855
rect 18153 13821 18187 13855
rect 18521 13821 18555 13855
rect 18705 13821 18739 13855
rect 18981 13821 19015 13855
rect 24225 13821 24259 13855
rect 28273 13821 28307 13855
rect 5917 13753 5951 13787
rect 9873 13753 9907 13787
rect 11897 13753 11931 13787
rect 19073 13753 19107 13787
rect 23857 13753 23891 13787
rect 4537 13685 4571 13719
rect 5273 13685 5307 13719
rect 5549 13685 5583 13719
rect 6653 13685 6687 13719
rect 6837 13685 6871 13719
rect 10517 13685 10551 13719
rect 11529 13685 11563 13719
rect 13553 13685 13587 13719
rect 27169 13685 27203 13719
rect 30297 13685 30331 13719
rect 4169 13481 4203 13515
rect 7757 13481 7791 13515
rect 9689 13481 9723 13515
rect 11621 13481 11655 13515
rect 12725 13481 12759 13515
rect 13461 13481 13495 13515
rect 15209 13481 15243 13515
rect 21741 13481 21775 13515
rect 22753 13481 22787 13515
rect 24409 13481 24443 13515
rect 25881 13481 25915 13515
rect 31309 13481 31343 13515
rect 31677 13481 31711 13515
rect 9321 13413 9355 13447
rect 9413 13413 9447 13447
rect 22109 13413 22143 13447
rect 22385 13413 22419 13447
rect 30481 13413 30515 13447
rect 31033 13413 31067 13447
rect 31217 13413 31251 13447
rect 15577 13345 15611 13379
rect 16129 13345 16163 13379
rect 19809 13345 19843 13379
rect 20453 13345 20487 13379
rect 21189 13345 21223 13379
rect 21833 13345 21867 13379
rect 24133 13345 24167 13379
rect 24961 13345 24995 13379
rect 27353 13345 27387 13379
rect 27629 13345 27663 13379
rect 30665 13345 30699 13379
rect 31585 13345 31619 13379
rect 1409 13277 1443 13311
rect 3801 13277 3835 13311
rect 4077 13277 4111 13311
rect 4261 13277 4295 13311
rect 5365 13277 5399 13311
rect 6469 13277 6503 13311
rect 6561 13277 6595 13311
rect 7665 13277 7699 13311
rect 7849 13277 7883 13311
rect 7941 13277 7975 13311
rect 8125 13277 8159 13311
rect 8953 13277 8987 13311
rect 9229 13277 9263 13311
rect 9781 13277 9815 13311
rect 9965 13277 9999 13311
rect 10333 13277 10367 13311
rect 11529 13277 11563 13311
rect 11805 13277 11839 13311
rect 12081 13277 12115 13311
rect 12174 13277 12208 13311
rect 12587 13277 12621 13311
rect 12817 13277 12851 13311
rect 13001 13277 13035 13311
rect 13093 13277 13127 13311
rect 13185 13277 13219 13311
rect 13553 13277 13587 13311
rect 13737 13277 13771 13311
rect 15393 13277 15427 13311
rect 15669 13277 15703 13311
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 16037 13277 16071 13311
rect 19717 13277 19751 13311
rect 20821 13277 20855 13311
rect 20913 13277 20947 13311
rect 21373 13277 21407 13311
rect 21649 13277 21683 13311
rect 21741 13277 21775 13311
rect 22201 13277 22235 13311
rect 22937 13277 22971 13311
rect 23213 13277 23247 13311
rect 23305 13277 23339 13311
rect 24777 13277 24811 13311
rect 28457 13277 28491 13311
rect 31677 13277 31711 13311
rect 5457 13209 5491 13243
rect 6193 13209 6227 13243
rect 8033 13209 8067 13243
rect 11989 13209 12023 13243
rect 12357 13209 12391 13243
rect 12449 13209 12483 13243
rect 20545 13209 20579 13243
rect 21557 13209 21591 13243
rect 24869 13209 24903 13243
rect 30205 13209 30239 13243
rect 30757 13209 30791 13243
rect 1593 13141 1627 13175
rect 3893 13141 3927 13175
rect 6377 13141 6411 13175
rect 6745 13141 6779 13175
rect 9045 13141 9079 13175
rect 9965 13141 9999 13175
rect 13553 13141 13587 13175
rect 20361 13141 20395 13175
rect 21097 13141 21131 13175
rect 23121 13141 23155 13175
rect 27905 13141 27939 13175
rect 9137 12937 9171 12971
rect 15577 12937 15611 12971
rect 31585 12937 31619 12971
rect 31953 12937 31987 12971
rect 33057 12937 33091 12971
rect 33517 12937 33551 12971
rect 16037 12869 16071 12903
rect 24593 12869 24627 12903
rect 28733 12869 28767 12903
rect 33609 12869 33643 12903
rect 9045 12801 9079 12835
rect 9229 12801 9263 12835
rect 15117 12801 15151 12835
rect 15669 12801 15703 12835
rect 15853 12801 15887 12835
rect 17141 12801 17175 12835
rect 17325 12801 17359 12835
rect 22845 12801 22879 12835
rect 22937 12801 22971 12835
rect 24869 12801 24903 12835
rect 27169 12801 27203 12835
rect 27353 12801 27387 12835
rect 27445 12801 27479 12835
rect 31493 12801 31527 12835
rect 31769 12801 31803 12835
rect 32689 12801 32723 12835
rect 33977 12801 34011 12835
rect 34161 12801 34195 12835
rect 22753 12733 22787 12767
rect 23029 12733 23063 12767
rect 23857 12733 23891 12767
rect 27997 12733 28031 12767
rect 32597 12733 32631 12767
rect 33701 12733 33735 12767
rect 34069 12733 34103 12767
rect 15393 12597 15427 12631
rect 17509 12597 17543 12631
rect 22569 12597 22603 12631
rect 24685 12597 24719 12631
rect 26985 12597 27019 12631
rect 33149 12597 33183 12631
rect 3617 12393 3651 12427
rect 4813 12393 4847 12427
rect 8953 12393 8987 12427
rect 11069 12393 11103 12427
rect 12541 12393 12575 12427
rect 18153 12393 18187 12427
rect 21925 12393 21959 12427
rect 23949 12393 23983 12427
rect 26157 12393 26191 12427
rect 31125 12393 31159 12427
rect 31861 12393 31895 12427
rect 33057 12393 33091 12427
rect 33793 12393 33827 12427
rect 4169 12325 4203 12359
rect 13461 12325 13495 12359
rect 17969 12325 18003 12359
rect 23765 12325 23799 12359
rect 30113 12325 30147 12359
rect 32045 12325 32079 12359
rect 33425 12325 33459 12359
rect 3525 12257 3559 12291
rect 7389 12257 7423 12291
rect 7941 12257 7975 12291
rect 13001 12257 13035 12291
rect 16773 12257 16807 12291
rect 17233 12257 17267 12291
rect 17718 12257 17752 12291
rect 22017 12257 22051 12291
rect 22385 12257 22419 12291
rect 23397 12257 23431 12291
rect 23489 12257 23523 12291
rect 23581 12257 23615 12291
rect 24409 12257 24443 12291
rect 26525 12257 26559 12291
rect 26801 12257 26835 12291
rect 28365 12257 28399 12291
rect 3617 12189 3651 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 4169 12189 4203 12223
rect 4445 12189 4479 12223
rect 4629 12189 4663 12223
rect 4997 12189 5031 12223
rect 5273 12189 5307 12223
rect 6101 12189 6135 12223
rect 6193 12189 6227 12223
rect 6377 12189 6411 12223
rect 6466 12189 6500 12223
rect 6745 12189 6779 12223
rect 6837 12189 6871 12223
rect 7021 12189 7055 12223
rect 7113 12189 7147 12223
rect 7573 12189 7607 12223
rect 9137 12189 9171 12223
rect 9229 12189 9263 12223
rect 9413 12189 9447 12223
rect 9515 12189 9549 12223
rect 11253 12189 11287 12223
rect 12725 12189 12759 12223
rect 12817 12189 12851 12223
rect 12909 12189 12943 12223
rect 13185 12189 13219 12223
rect 13461 12189 13495 12223
rect 17141 12189 17175 12223
rect 18613 12189 18647 12223
rect 20085 12189 20119 12223
rect 20269 12189 20303 12223
rect 21373 12189 21407 12223
rect 21557 12189 21591 12223
rect 21741 12189 21775 12223
rect 22201 12189 22235 12223
rect 22477 12189 22511 12223
rect 22661 12189 22695 12223
rect 22753 12189 22787 12223
rect 23305 12189 23339 12223
rect 24041 12189 24075 12223
rect 29561 12189 29595 12223
rect 29837 12189 29871 12223
rect 29929 12189 29963 12223
rect 30389 12189 30423 12223
rect 30665 12189 30699 12223
rect 31309 12189 31343 12223
rect 31401 12189 31435 12223
rect 31677 12189 31711 12223
rect 31769 12189 31803 12223
rect 32321 12189 32355 12223
rect 32965 12189 32999 12223
rect 33517 12189 33551 12223
rect 5457 12121 5491 12155
rect 7297 12121 7331 12155
rect 11437 12121 11471 12155
rect 16656 12121 16690 12155
rect 18337 12121 18371 12155
rect 21649 12121 21683 12155
rect 24685 12121 24719 12155
rect 29009 12121 29043 12155
rect 29745 12121 29779 12155
rect 31493 12121 31527 12155
rect 3249 12053 3283 12087
rect 5089 12053 5123 12087
rect 6653 12053 6687 12087
rect 7849 12053 7883 12087
rect 13277 12053 13311 12087
rect 16497 12053 16531 12087
rect 16865 12053 16899 12087
rect 17509 12053 17543 12087
rect 17601 12053 17635 12087
rect 17877 12053 17911 12087
rect 18137 12053 18171 12087
rect 18429 12053 18463 12087
rect 20177 12053 20211 12087
rect 28273 12053 28307 12087
rect 30205 12053 30239 12087
rect 30573 12053 30607 12087
rect 33977 12053 34011 12087
rect 3985 11849 4019 11883
rect 4537 11849 4571 11883
rect 6653 11849 6687 11883
rect 7389 11849 7423 11883
rect 7665 11849 7699 11883
rect 8861 11849 8895 11883
rect 12449 11849 12483 11883
rect 13369 11849 13403 11883
rect 17509 11849 17543 11883
rect 19717 11849 19751 11883
rect 21649 11849 21683 11883
rect 22477 11849 22511 11883
rect 24593 11849 24627 11883
rect 24961 11849 24995 11883
rect 3617 11781 3651 11815
rect 4905 11781 4939 11815
rect 8033 11781 8067 11815
rect 8401 11781 8435 11815
rect 9347 11781 9381 11815
rect 9597 11781 9631 11815
rect 17877 11781 17911 11815
rect 22109 11781 22143 11815
rect 22845 11781 22879 11815
rect 25053 11781 25087 11815
rect 30113 11781 30147 11815
rect 3249 11713 3283 11747
rect 3433 11713 3467 11747
rect 3525 11713 3559 11747
rect 3801 11713 3835 11747
rect 4169 11713 4203 11747
rect 4261 11713 4295 11747
rect 4721 11713 4755 11747
rect 5089 11713 5123 11747
rect 6469 11713 6503 11747
rect 6745 11713 6779 11747
rect 6837 11713 6871 11747
rect 7205 11713 7239 11747
rect 7297 11713 7331 11747
rect 7665 11713 7699 11747
rect 7849 11713 7883 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 9046 11713 9080 11747
rect 9137 11713 9171 11747
rect 9254 11713 9288 11747
rect 10426 11735 10460 11769
rect 10517 11713 10551 11747
rect 10793 11713 10827 11747
rect 10899 11713 10933 11747
rect 11069 11713 11103 11747
rect 11161 11713 11195 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 11897 11713 11931 11747
rect 12357 11713 12391 11747
rect 12633 11713 12667 11747
rect 12725 11713 12759 11747
rect 12909 11713 12943 11747
rect 13185 11713 13219 11747
rect 13461 11713 13495 11747
rect 13553 11713 13587 11747
rect 13737 11713 13771 11747
rect 13829 11713 13863 11747
rect 15577 11713 15611 11747
rect 16313 11713 16347 11747
rect 16773 11713 16807 11747
rect 17693 11713 17727 11747
rect 17969 11713 18003 11747
rect 20085 11713 20119 11747
rect 20361 11713 20395 11747
rect 20453 11713 20487 11747
rect 20545 11713 20579 11747
rect 21097 11713 21131 11747
rect 21465 11713 21499 11747
rect 21833 11713 21867 11747
rect 21926 11713 21960 11747
rect 22201 11713 22235 11747
rect 22339 11713 22373 11747
rect 22754 11735 22788 11769
rect 22937 11713 22971 11747
rect 23055 11713 23089 11747
rect 30389 11713 30423 11747
rect 31217 11713 31251 11747
rect 6377 11645 6411 11679
rect 9505 11645 9539 11679
rect 9744 11645 9778 11679
rect 9965 11645 9999 11679
rect 10701 11645 10735 11679
rect 12173 11645 12207 11679
rect 14013 11645 14047 11679
rect 16129 11645 16163 11679
rect 16497 11645 16531 11679
rect 17049 11645 17083 11679
rect 18245 11645 18279 11679
rect 20269 11645 20303 11679
rect 20729 11645 20763 11679
rect 21005 11645 21039 11679
rect 23213 11645 23247 11679
rect 25145 11645 25179 11679
rect 28641 11645 28675 11679
rect 13001 11577 13035 11611
rect 13093 11577 13127 11611
rect 3341 11509 3375 11543
rect 4353 11509 4387 11543
rect 7113 11509 7147 11543
rect 7573 11509 7607 11543
rect 8217 11509 8251 11543
rect 9873 11509 9907 11543
rect 10057 11509 10091 11543
rect 10609 11509 10643 11543
rect 11345 11509 11379 11543
rect 12633 11509 12667 11543
rect 15393 11509 15427 11543
rect 21465 11509 21499 11543
rect 22569 11509 22603 11543
rect 31309 11509 31343 11543
rect 31677 11509 31711 11543
rect 4261 11305 4295 11339
rect 6377 11305 6411 11339
rect 8677 11305 8711 11339
rect 9965 11305 9999 11339
rect 10425 11305 10459 11339
rect 12449 11305 12483 11339
rect 13553 11305 13587 11339
rect 16589 11305 16623 11339
rect 21005 11305 21039 11339
rect 22569 11305 22603 11339
rect 30573 11305 30607 11339
rect 30757 11305 30791 11339
rect 31677 11305 31711 11339
rect 6837 11237 6871 11271
rect 9689 11237 9723 11271
rect 23213 11237 23247 11271
rect 1409 11169 1443 11203
rect 1685 11169 1719 11203
rect 6469 11169 6503 11203
rect 12817 11169 12851 11203
rect 14841 11169 14875 11203
rect 15117 11169 15151 11203
rect 26985 11169 27019 11203
rect 30205 11169 30239 11203
rect 32045 11169 32079 11203
rect 6377 11101 6411 11135
rect 6653 11101 6687 11135
rect 8033 11101 8067 11135
rect 8126 11101 8160 11135
rect 8309 11101 8343 11135
rect 8498 11101 8532 11135
rect 9045 11101 9079 11135
rect 9229 11101 9263 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 9965 11101 9999 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 12633 11101 12667 11135
rect 12725 11101 12759 11135
rect 12909 11101 12943 11135
rect 13093 11101 13127 11135
rect 13369 11101 13403 11135
rect 20913 11101 20947 11135
rect 21097 11101 21131 11135
rect 22845 11101 22879 11135
rect 23121 11101 23155 11135
rect 23305 11101 23339 11135
rect 23673 11101 23707 11135
rect 26709 11101 26743 11135
rect 29561 11101 29595 11135
rect 30297 11101 30331 11135
rect 31217 11101 31251 11135
rect 31309 11101 31343 11135
rect 31493 11101 31527 11135
rect 31953 11101 31987 11135
rect 4077 11033 4111 11067
rect 4277 11033 4311 11067
rect 8401 11033 8435 11067
rect 13185 11033 13219 11067
rect 22569 11033 22603 11067
rect 23765 11033 23799 11067
rect 27261 11033 27295 11067
rect 3157 10965 3191 10999
rect 4445 10965 4479 10999
rect 22753 10965 22787 10999
rect 26893 10965 26927 10999
rect 28733 10965 28767 10999
rect 32321 10965 32355 10999
rect 5181 10761 5215 10795
rect 17693 10761 17727 10795
rect 18061 10761 18095 10795
rect 18337 10761 18371 10795
rect 20177 10761 20211 10795
rect 24685 10761 24719 10795
rect 26985 10761 27019 10795
rect 31953 10761 31987 10795
rect 32689 10761 32723 10795
rect 33057 10761 33091 10795
rect 5457 10693 5491 10727
rect 18705 10693 18739 10727
rect 25053 10693 25087 10727
rect 27445 10693 27479 10727
rect 30297 10693 30331 10727
rect 31677 10693 31711 10727
rect 3617 10625 3651 10659
rect 4905 10625 4939 10659
rect 4997 10625 5031 10659
rect 5273 10625 5307 10659
rect 5549 10625 5583 10659
rect 6561 10625 6595 10659
rect 6837 10625 6871 10659
rect 7021 10625 7055 10659
rect 17417 10625 17451 10659
rect 17785 10625 17819 10659
rect 18153 10625 18187 10659
rect 23121 10625 23155 10659
rect 24501 10625 24535 10659
rect 27353 10625 27387 10659
rect 28089 10625 28123 10659
rect 28733 10625 28767 10659
rect 31401 10625 31435 10659
rect 31585 10625 31619 10659
rect 31769 10625 31803 10659
rect 32321 10625 32355 10659
rect 32505 10625 32539 10659
rect 32597 10625 32631 10659
rect 4721 10557 4755 10591
rect 4813 10557 4847 10591
rect 6745 10557 6779 10591
rect 17902 10557 17936 10591
rect 18429 10557 18463 10591
rect 24777 10557 24811 10591
rect 27537 10557 27571 10591
rect 33149 10557 33183 10591
rect 33333 10557 33367 10591
rect 6653 10489 6687 10523
rect 30665 10489 30699 10523
rect 3065 10421 3099 10455
rect 5549 10421 5583 10455
rect 6377 10421 6411 10455
rect 22937 10421 22971 10455
rect 26525 10421 26559 10455
rect 30757 10421 30791 10455
rect 32137 10421 32171 10455
rect 6561 10217 6595 10251
rect 6929 10217 6963 10251
rect 7941 10217 7975 10251
rect 8953 10217 8987 10251
rect 11253 10217 11287 10251
rect 12909 10217 12943 10251
rect 17877 10217 17911 10251
rect 18153 10217 18187 10251
rect 22740 10217 22774 10251
rect 24961 10217 24995 10251
rect 31309 10217 31343 10251
rect 32854 10217 32888 10251
rect 34345 10217 34379 10251
rect 5641 10149 5675 10183
rect 6009 10149 6043 10183
rect 6101 10149 6135 10183
rect 8309 10149 8343 10183
rect 12357 10149 12391 10183
rect 17969 10149 18003 10183
rect 24225 10149 24259 10183
rect 27353 10149 27387 10183
rect 7481 10081 7515 10115
rect 10977 10081 11011 10115
rect 11069 10081 11103 10115
rect 11345 10081 11379 10115
rect 12817 10081 12851 10115
rect 22477 10081 22511 10115
rect 25421 10081 25455 10115
rect 25513 10081 25547 10115
rect 26617 10081 26651 10115
rect 26709 10081 26743 10115
rect 29561 10081 29595 10115
rect 32597 10081 32631 10115
rect 5368 10013 5402 10047
rect 5457 10013 5491 10047
rect 5917 10013 5951 10047
rect 6193 10013 6227 10047
rect 6469 10013 6503 10047
rect 6745 10013 6779 10047
rect 7573 10013 7607 10047
rect 8033 10013 8067 10047
rect 9137 10013 9171 10047
rect 9321 10013 9355 10047
rect 9413 10013 9447 10047
rect 10609 10013 10643 10047
rect 10701 10013 10735 10047
rect 11529 10013 11563 10047
rect 11621 10013 11655 10047
rect 12173 10013 12207 10047
rect 12357 10013 12391 10047
rect 12449 10013 12483 10047
rect 12633 10013 12667 10047
rect 13277 10013 13311 10047
rect 13553 10013 13587 10047
rect 17693 10013 17727 10047
rect 27997 10013 28031 10047
rect 28365 10013 28399 10047
rect 28457 10013 28491 10047
rect 28641 10013 28675 10047
rect 28733 10013 28767 10047
rect 28825 10013 28859 10047
rect 29009 10013 29043 10047
rect 5641 9945 5675 9979
rect 6377 9945 6411 9979
rect 7113 9945 7147 9979
rect 7297 9945 7331 9979
rect 7757 9945 7791 9979
rect 8125 9945 8159 9979
rect 8309 9945 8343 9979
rect 12725 9945 12759 9979
rect 13185 9945 13219 9979
rect 13737 9945 13771 9979
rect 17509 9945 17543 9979
rect 18121 9945 18155 9979
rect 18337 9945 18371 9979
rect 25329 9945 25363 9979
rect 25973 9945 26007 9979
rect 28181 9945 28215 9979
rect 29193 9945 29227 9979
rect 29837 9945 29871 9979
rect 10793 9877 10827 9911
rect 11345 9877 11379 9911
rect 12541 9877 12575 9911
rect 13093 9877 13127 9911
rect 13369 9877 13403 9911
rect 9137 9673 9171 9707
rect 10057 9673 10091 9707
rect 11529 9673 11563 9707
rect 13553 9673 13587 9707
rect 17877 9673 17911 9707
rect 22937 9673 22971 9707
rect 2973 9605 3007 9639
rect 8585 9605 8619 9639
rect 10701 9605 10735 9639
rect 12725 9605 12759 9639
rect 13461 9605 13495 9639
rect 14565 9605 14599 9639
rect 15761 9605 15795 9639
rect 17049 9605 17083 9639
rect 17417 9605 17451 9639
rect 17994 9605 18028 9639
rect 21005 9605 21039 9639
rect 21649 9605 21683 9639
rect 23397 9605 23431 9639
rect 27445 9605 27479 9639
rect 2697 9537 2731 9571
rect 8125 9537 8159 9571
rect 8217 9537 8251 9571
rect 8401 9537 8435 9571
rect 8953 9537 8987 9571
rect 9485 9537 9519 9571
rect 9597 9537 9631 9571
rect 9710 9537 9744 9571
rect 9873 9537 9907 9571
rect 9965 9537 9999 9571
rect 10425 9537 10459 9571
rect 10885 9537 10919 9571
rect 10977 9537 11011 9571
rect 11161 9537 11195 9571
rect 11345 9537 11379 9571
rect 11805 9537 11839 9571
rect 11897 9537 11931 9571
rect 11989 9537 12023 9571
rect 12149 9537 12183 9571
rect 12541 9537 12575 9571
rect 13186 9559 13220 9593
rect 13553 9537 13587 9571
rect 13737 9537 13771 9571
rect 14841 9537 14875 9571
rect 15117 9537 15151 9571
rect 16037 9537 16071 9571
rect 16129 9537 16163 9571
rect 17233 9537 17267 9571
rect 18429 9537 18463 9571
rect 20729 9537 20763 9571
rect 21087 9537 21121 9571
rect 21189 9537 21223 9571
rect 21373 9537 21407 9571
rect 21465 9537 21499 9571
rect 21833 9537 21867 9571
rect 22201 9537 22235 9571
rect 23305 9537 23339 9571
rect 23857 9537 23891 9571
rect 24409 9537 24443 9571
rect 26433 9537 26467 9571
rect 27353 9537 27387 9571
rect 29653 9537 29687 9571
rect 31125 9537 31159 9571
rect 8677 9469 8711 9503
rect 9229 9469 9263 9503
rect 10241 9469 10275 9503
rect 12265 9469 12299 9503
rect 13461 9469 13495 9503
rect 14749 9469 14783 9503
rect 15393 9469 15427 9503
rect 15761 9469 15795 9503
rect 17509 9469 17543 9503
rect 17785 9469 17819 9503
rect 18705 9469 18739 9503
rect 20177 9469 20211 9503
rect 21005 9469 21039 9503
rect 22017 9469 22051 9503
rect 23581 9469 23615 9503
rect 27537 9469 27571 9503
rect 29929 9469 29963 9503
rect 31401 9469 31435 9503
rect 11069 9401 11103 9435
rect 15025 9401 15059 9435
rect 21903 9401 21937 9435
rect 26985 9401 27019 9435
rect 30205 9401 30239 9435
rect 31677 9401 31711 9435
rect 4445 9333 4479 9367
rect 8769 9333 8803 9367
rect 12357 9333 12391 9367
rect 13277 9333 13311 9367
rect 14565 9333 14599 9367
rect 15209 9333 15243 9367
rect 15669 9333 15703 9367
rect 15945 9333 15979 9367
rect 16221 9333 16255 9367
rect 18153 9333 18187 9367
rect 20821 9333 20855 9367
rect 22109 9333 22143 9367
rect 26249 9333 26283 9367
rect 29837 9333 29871 9367
rect 31217 9333 31251 9367
rect 9045 9129 9079 9163
rect 9137 9129 9171 9163
rect 10241 9129 10275 9163
rect 11621 9129 11655 9163
rect 14657 9129 14691 9163
rect 15301 9129 15335 9163
rect 16405 9129 16439 9163
rect 17417 9129 17451 9163
rect 17601 9129 17635 9163
rect 18429 9129 18463 9163
rect 20913 9129 20947 9163
rect 21833 9129 21867 9163
rect 23581 9129 23615 9163
rect 27813 9129 27847 9163
rect 30849 9129 30883 9163
rect 31033 9129 31067 9163
rect 31769 9129 31803 9163
rect 32045 9129 32079 9163
rect 32689 9129 32723 9163
rect 11253 9061 11287 9095
rect 15209 9061 15243 9095
rect 15577 9061 15611 9095
rect 16497 9061 16531 9095
rect 32137 9061 32171 9095
rect 9229 8993 9263 9027
rect 11161 8993 11195 9027
rect 21833 8993 21867 9027
rect 21925 8993 21959 9027
rect 23765 8993 23799 9027
rect 24501 8993 24535 9027
rect 26341 8993 26375 9027
rect 28273 8993 28307 9027
rect 31953 8993 31987 9027
rect 33241 8993 33275 9027
rect 8953 8925 8987 8959
rect 10057 8925 10091 8959
rect 10241 8925 10275 8959
rect 11437 8925 11471 8959
rect 14841 8925 14875 8959
rect 15025 8925 15059 8959
rect 15485 8925 15519 8959
rect 15669 8925 15703 8959
rect 15761 8925 15795 8959
rect 15945 8925 15979 8959
rect 16037 8925 16071 8959
rect 16497 8925 16531 8959
rect 18245 8925 18279 8959
rect 21097 8925 21131 8959
rect 21281 8925 21315 8959
rect 21465 8925 21499 8959
rect 22017 8925 22051 8959
rect 23489 8925 23523 8959
rect 24409 8925 24443 8959
rect 24593 8925 24627 8959
rect 24961 8925 24995 8959
rect 25605 8925 25639 8959
rect 26065 8925 26099 8959
rect 27905 8925 27939 8959
rect 28181 8925 28215 8959
rect 28365 8925 28399 8959
rect 31309 8925 31343 8959
rect 31861 8925 31895 8959
rect 32229 8925 32263 8959
rect 14565 8857 14599 8891
rect 17785 8857 17819 8891
rect 21189 8857 21223 8891
rect 21649 8857 21683 8891
rect 28549 8857 28583 8891
rect 33149 8857 33183 8891
rect 16129 8789 16163 8823
rect 16221 8789 16255 8823
rect 17585 8789 17619 8823
rect 23765 8789 23799 8823
rect 28733 8789 28767 8823
rect 31401 8789 31435 8823
rect 33057 8789 33091 8823
rect 17509 8585 17543 8619
rect 21373 8585 21407 8619
rect 25237 8585 25271 8619
rect 29837 8585 29871 8619
rect 19717 8517 19751 8551
rect 19487 8483 19521 8517
rect 17693 8449 17727 8483
rect 21189 8449 21223 8483
rect 21373 8449 21407 8483
rect 23121 8449 23155 8483
rect 23213 8449 23247 8483
rect 23489 8449 23523 8483
rect 26985 8449 27019 8483
rect 31217 8449 31251 8483
rect 31401 8449 31435 8483
rect 32321 8449 32355 8483
rect 34345 8449 34379 8483
rect 17877 8381 17911 8415
rect 23765 8381 23799 8415
rect 25973 8381 26007 8415
rect 28089 8381 28123 8415
rect 28365 8381 28399 8415
rect 32229 8381 32263 8415
rect 32689 8381 32723 8415
rect 19349 8313 19383 8347
rect 23305 8313 23339 8347
rect 26617 8313 26651 8347
rect 19533 8245 19567 8279
rect 22937 8245 22971 8279
rect 27077 8245 27111 8279
rect 31309 8245 31343 8279
rect 34161 8245 34195 8279
rect 13921 8041 13955 8075
rect 15853 8041 15887 8075
rect 22845 8041 22879 8075
rect 27997 8041 28031 8075
rect 30849 8041 30883 8075
rect 17785 7973 17819 8007
rect 20177 7973 20211 8007
rect 32597 7973 32631 8007
rect 12173 7905 12207 7939
rect 17141 7905 17175 7939
rect 19533 7905 19567 7939
rect 22293 7905 22327 7939
rect 24869 7905 24903 7939
rect 25053 7905 25087 7939
rect 25237 7905 25271 7939
rect 25881 7905 25915 7939
rect 26433 7905 26467 7939
rect 26525 7905 26559 7939
rect 28365 7905 28399 7939
rect 28457 7905 28491 7939
rect 34069 7905 34103 7939
rect 15577 7837 15611 7871
rect 16129 7837 16163 7871
rect 17417 7837 17451 7871
rect 18245 7837 18279 7871
rect 20453 7837 20487 7871
rect 20729 7837 20763 7871
rect 23765 7837 23799 7871
rect 27253 7837 27287 7871
rect 28181 7837 28215 7871
rect 28549 7837 28583 7871
rect 28733 7837 28767 7871
rect 34345 7837 34379 7871
rect 12449 7769 12483 7803
rect 15853 7769 15887 7803
rect 17626 7769 17660 7803
rect 17877 7769 17911 7803
rect 18061 7769 18095 7803
rect 20018 7769 20052 7803
rect 20269 7769 20303 7803
rect 20637 7769 20671 7803
rect 22477 7769 22511 7803
rect 23121 7769 23155 7803
rect 26617 7769 26651 7803
rect 30665 7769 30699 7803
rect 15669 7701 15703 7735
rect 16037 7701 16071 7735
rect 17509 7701 17543 7735
rect 19809 7701 19843 7735
rect 19901 7701 19935 7735
rect 22385 7701 22419 7735
rect 24409 7701 24443 7735
rect 24777 7701 24811 7735
rect 26985 7701 27019 7735
rect 27077 7701 27111 7735
rect 30865 7701 30899 7735
rect 31033 7701 31067 7735
rect 11345 7497 11379 7531
rect 16313 7497 16347 7531
rect 16773 7497 16807 7531
rect 19809 7497 19843 7531
rect 21649 7497 21683 7531
rect 23673 7497 23707 7531
rect 26157 7497 26191 7531
rect 31861 7497 31895 7531
rect 8585 7429 8619 7463
rect 12633 7429 12667 7463
rect 20177 7429 20211 7463
rect 22201 7429 22235 7463
rect 30389 7429 30423 7463
rect 14565 7361 14599 7395
rect 16681 7361 16715 7395
rect 16865 7361 16899 7395
rect 17601 7361 17635 7395
rect 18797 7361 18831 7395
rect 18981 7361 19015 7395
rect 19625 7361 19659 7395
rect 24133 7361 24167 7395
rect 24409 7361 24443 7395
rect 29837 7361 29871 7395
rect 30941 7361 30975 7395
rect 31493 7361 31527 7395
rect 7941 7293 7975 7327
rect 10701 7293 10735 7327
rect 12357 7293 12391 7327
rect 14841 7293 14875 7327
rect 19901 7293 19935 7327
rect 21925 7293 21959 7327
rect 24685 7293 24719 7327
rect 30297 7293 30331 7327
rect 31401 7293 31435 7327
rect 31585 7293 31619 7327
rect 24317 7225 24351 7259
rect 30665 7225 30699 7259
rect 14105 7157 14139 7191
rect 17417 7157 17451 7191
rect 18889 7157 18923 7191
rect 29929 7157 29963 7191
rect 30849 7157 30883 7191
rect 31033 7157 31067 7191
rect 31493 7157 31527 7191
rect 16221 6953 16255 6987
rect 17312 6953 17346 6987
rect 18797 6953 18831 6987
rect 26328 6953 26362 6987
rect 27813 6953 27847 6987
rect 31033 6953 31067 6987
rect 19809 6885 19843 6919
rect 1409 6817 1443 6851
rect 3157 6817 3191 6851
rect 16129 6817 16163 6851
rect 17049 6817 17083 6851
rect 26065 6817 26099 6851
rect 31769 6817 31803 6851
rect 32413 6817 32447 6851
rect 32597 6817 32631 6851
rect 15945 6749 15979 6783
rect 19533 6749 19567 6783
rect 19625 6749 19659 6783
rect 23581 6749 23615 6783
rect 29561 6749 29595 6783
rect 30757 6749 30791 6783
rect 30849 6749 30883 6783
rect 31677 6749 31711 6783
rect 1685 6681 1719 6715
rect 16221 6681 16255 6715
rect 19441 6681 19475 6715
rect 31033 6681 31067 6715
rect 15761 6613 15795 6647
rect 19257 6613 19291 6647
rect 23397 6613 23431 6647
rect 29653 6613 29687 6647
rect 32045 6613 32079 6647
rect 32689 6613 32723 6647
rect 33057 6613 33091 6647
rect 1593 6409 1627 6443
rect 8953 6409 8987 6443
rect 15209 6409 15243 6443
rect 19257 6409 19291 6443
rect 22845 6409 22879 6443
rect 23305 6409 23339 6443
rect 24685 6409 24719 6443
rect 29561 6409 29595 6443
rect 29745 6409 29779 6443
rect 30481 6409 30515 6443
rect 30849 6409 30883 6443
rect 32597 6409 32631 6443
rect 11805 6341 11839 6375
rect 18889 6341 18923 6375
rect 19073 6341 19107 6375
rect 27997 6341 28031 6375
rect 1409 6273 1443 6307
rect 7205 6273 7239 6307
rect 13461 6273 13495 6307
rect 19349 6273 19383 6307
rect 20545 6273 20579 6307
rect 22385 6273 22419 6307
rect 22937 6273 22971 6307
rect 24317 6273 24351 6307
rect 27537 6273 27571 6307
rect 28549 6273 28583 6307
rect 29929 6273 29963 6307
rect 30021 6273 30055 6307
rect 30205 6273 30239 6307
rect 30297 6273 30331 6307
rect 30389 6273 30423 6307
rect 30665 6273 30699 6307
rect 34345 6273 34379 6307
rect 7481 6205 7515 6239
rect 11529 6205 11563 6239
rect 13737 6205 13771 6239
rect 22661 6205 22695 6239
rect 23489 6205 23523 6239
rect 24133 6205 24167 6239
rect 25881 6205 25915 6239
rect 27445 6205 27479 6239
rect 28457 6205 28491 6239
rect 29101 6205 29135 6239
rect 34069 6205 34103 6239
rect 28273 6137 28307 6171
rect 29009 6137 29043 6171
rect 29377 6137 29411 6171
rect 13277 6069 13311 6103
rect 19533 6069 19567 6103
rect 20361 6069 20395 6103
rect 21833 6069 21867 6103
rect 24685 6069 24719 6103
rect 24869 6069 24903 6103
rect 25329 6069 25363 6103
rect 27813 6069 27847 6103
rect 28641 6069 28675 6103
rect 14105 5865 14139 5899
rect 15945 5865 15979 5899
rect 21373 5865 21407 5899
rect 22740 5865 22774 5899
rect 26709 5865 26743 5899
rect 30021 5865 30055 5899
rect 32229 5865 32263 5899
rect 14657 5729 14691 5763
rect 17693 5729 17727 5763
rect 19257 5729 19291 5763
rect 19533 5729 19567 5763
rect 21925 5729 21959 5763
rect 22477 5729 22511 5763
rect 24961 5729 24995 5763
rect 25237 5729 25271 5763
rect 28089 5729 28123 5763
rect 21741 5661 21775 5695
rect 29561 5661 29595 5695
rect 29653 5661 29687 5695
rect 29837 5661 29871 5695
rect 31493 5661 31527 5695
rect 31769 5661 31803 5695
rect 31861 5661 31895 5695
rect 32413 5661 32447 5695
rect 32597 5661 32631 5695
rect 32689 5661 32723 5695
rect 17417 5593 17451 5627
rect 21281 5593 21315 5627
rect 27905 5593 27939 5627
rect 31677 5593 31711 5627
rect 21833 5525 21867 5559
rect 24225 5525 24259 5559
rect 27445 5525 27479 5559
rect 27813 5525 27847 5559
rect 32045 5525 32079 5559
rect 21649 5321 21683 5355
rect 23857 5321 23891 5355
rect 25421 5321 25455 5355
rect 26433 5321 26467 5355
rect 26985 5321 27019 5355
rect 28457 5321 28491 5355
rect 28825 5321 28859 5355
rect 30021 5321 30055 5355
rect 30849 5321 30883 5355
rect 20177 5253 20211 5287
rect 22293 5253 22327 5287
rect 25145 5253 25179 5287
rect 12909 5185 12943 5219
rect 16497 5185 16531 5219
rect 22201 5185 22235 5219
rect 23029 5185 23063 5219
rect 23673 5185 23707 5219
rect 24777 5185 24811 5219
rect 24870 5185 24904 5219
rect 25053 5185 25087 5219
rect 25242 5185 25276 5219
rect 26341 5185 26375 5219
rect 26617 5185 26651 5219
rect 27169 5185 27203 5219
rect 27261 5185 27295 5219
rect 27353 5185 27387 5219
rect 27537 5185 27571 5219
rect 28917 5185 28951 5219
rect 30389 5185 30423 5219
rect 30665 5185 30699 5219
rect 30849 5185 30883 5219
rect 13185 5117 13219 5151
rect 14657 5117 14691 5151
rect 14749 5117 14783 5151
rect 16221 5117 16255 5151
rect 19901 5117 19935 5151
rect 22477 5117 22511 5151
rect 24409 5117 24443 5151
rect 25513 5117 25547 5151
rect 26157 5117 26191 5151
rect 29009 5117 29043 5151
rect 30297 5117 30331 5151
rect 26801 5049 26835 5083
rect 21833 4981 21867 5015
rect 13277 4777 13311 4811
rect 15301 4777 15335 4811
rect 23673 4777 23707 4811
rect 29009 4777 29043 4811
rect 30021 4777 30055 4811
rect 30205 4777 30239 4811
rect 29377 4709 29411 4743
rect 29837 4709 29871 4743
rect 21925 4641 21959 4675
rect 25053 4641 25087 4675
rect 13829 4573 13863 4607
rect 14657 4573 14691 4607
rect 18153 4573 18187 4607
rect 21649 4573 21683 4607
rect 28917 4573 28951 4607
rect 29561 4573 29595 4607
rect 30113 4573 30147 4607
rect 22201 4505 22235 4539
rect 24869 4505 24903 4539
rect 18797 4437 18831 4471
rect 21833 4437 21867 4471
rect 24409 4437 24443 4471
rect 24777 4437 24811 4471
rect 14197 4233 14231 4267
rect 25973 4233 26007 4267
rect 28733 4233 28767 4267
rect 30205 4233 30239 4267
rect 27261 4165 27295 4199
rect 11897 4097 11931 4131
rect 19717 4097 19751 4131
rect 22109 4097 22143 4131
rect 22201 4097 22235 4131
rect 23949 4097 23983 4131
rect 24225 4097 24259 4131
rect 26985 4097 27019 4131
rect 31953 4097 31987 4131
rect 12173 4029 12207 4063
rect 13645 4029 13679 4063
rect 15669 4029 15703 4063
rect 15945 4029 15979 4063
rect 17969 4029 18003 4063
rect 19441 4029 19475 4063
rect 24501 4029 24535 4063
rect 31677 4029 31711 4063
rect 24133 3961 24167 3995
rect 16773 3689 16807 3723
rect 18521 3553 18555 3587
rect 18245 3417 18279 3451
rect 6101 2601 6135 2635
rect 12357 2601 12391 2635
rect 24593 2601 24627 2635
rect 31217 2601 31251 2635
rect 34161 2533 34195 2567
rect 1409 2397 1443 2431
rect 5917 2397 5951 2431
rect 12541 2397 12575 2431
rect 19349 2397 19383 2431
rect 24777 2397 24811 2431
rect 31033 2397 31067 2431
rect 34345 2397 34379 2431
rect 1593 2261 1627 2295
rect 19441 2261 19475 2295
<< metal1 >>
rect 1104 35386 34684 35408
rect 1104 35334 5147 35386
rect 5199 35334 5211 35386
rect 5263 35334 5275 35386
rect 5327 35334 5339 35386
rect 5391 35334 5403 35386
rect 5455 35334 13541 35386
rect 13593 35334 13605 35386
rect 13657 35334 13669 35386
rect 13721 35334 13733 35386
rect 13785 35334 13797 35386
rect 13849 35334 21935 35386
rect 21987 35334 21999 35386
rect 22051 35334 22063 35386
rect 22115 35334 22127 35386
rect 22179 35334 22191 35386
rect 22243 35334 30329 35386
rect 30381 35334 30393 35386
rect 30445 35334 30457 35386
rect 30509 35334 30521 35386
rect 30573 35334 30585 35386
rect 30637 35334 34684 35386
rect 1104 35312 34684 35334
rect 1302 35232 1308 35284
rect 1360 35272 1366 35284
rect 1489 35275 1547 35281
rect 1489 35272 1501 35275
rect 1360 35244 1501 35272
rect 1360 35232 1366 35244
rect 1489 35241 1501 35244
rect 1535 35241 1547 35275
rect 1489 35235 1547 35241
rect 26418 35232 26424 35284
rect 26476 35272 26482 35284
rect 27157 35275 27215 35281
rect 27157 35272 27169 35275
rect 26476 35244 27169 35272
rect 26476 35232 26482 35244
rect 27157 35241 27169 35244
rect 27203 35241 27215 35275
rect 27157 35235 27215 35241
rect 9214 35164 9220 35216
rect 9272 35204 9278 35216
rect 15746 35204 15752 35216
rect 9272 35176 15752 35204
rect 9272 35164 9278 35176
rect 15746 35164 15752 35176
rect 15804 35204 15810 35216
rect 15804 35176 16896 35204
rect 15804 35164 15810 35176
rect 13906 35096 13912 35148
rect 13964 35096 13970 35148
rect 16868 35145 16896 35176
rect 16853 35139 16911 35145
rect 16853 35105 16865 35139
rect 16899 35105 16911 35139
rect 16853 35099 16911 35105
rect 7742 35028 7748 35080
rect 7800 35028 7806 35080
rect 8110 35028 8116 35080
rect 8168 35028 8174 35080
rect 8205 35071 8263 35077
rect 8205 35037 8217 35071
rect 8251 35037 8263 35071
rect 8205 35031 8263 35037
rect 13817 35071 13875 35077
rect 13817 35037 13829 35071
rect 13863 35068 13875 35071
rect 13924 35068 13952 35096
rect 13863 35040 13952 35068
rect 16393 35071 16451 35077
rect 13863 35037 13875 35040
rect 13817 35031 13875 35037
rect 16393 35037 16405 35071
rect 16439 35068 16451 35071
rect 16574 35068 16580 35080
rect 16439 35040 16580 35068
rect 16439 35037 16451 35040
rect 16393 35031 16451 35037
rect 1762 34960 1768 35012
rect 1820 34960 1826 35012
rect 7760 35000 7788 35028
rect 8220 35000 8248 35031
rect 16574 35028 16580 35040
rect 16632 35028 16638 35080
rect 17126 35028 17132 35080
rect 17184 35028 17190 35080
rect 19978 35028 19984 35080
rect 20036 35068 20042 35080
rect 20073 35071 20131 35077
rect 20073 35068 20085 35071
rect 20036 35040 20085 35068
rect 20036 35028 20042 35040
rect 20073 35037 20085 35040
rect 20119 35037 20131 35071
rect 21913 35071 21971 35077
rect 21913 35068 21925 35071
rect 20073 35031 20131 35037
rect 20272 35040 21925 35068
rect 7760 34972 8248 35000
rect 12526 34960 12532 35012
rect 12584 35000 12590 35012
rect 12584 34972 13952 35000
rect 12584 34960 12590 34972
rect 13924 34944 13952 34972
rect 7926 34892 7932 34944
rect 7984 34892 7990 34944
rect 8389 34935 8447 34941
rect 8389 34901 8401 34935
rect 8435 34932 8447 34935
rect 9766 34932 9772 34944
rect 8435 34904 9772 34932
rect 8435 34901 8447 34904
rect 8389 34895 8447 34901
rect 9766 34892 9772 34904
rect 9824 34892 9830 34944
rect 13630 34892 13636 34944
rect 13688 34892 13694 34944
rect 13906 34892 13912 34944
rect 13964 34892 13970 34944
rect 15654 34892 15660 34944
rect 15712 34932 15718 34944
rect 15749 34935 15807 34941
rect 15749 34932 15761 34935
rect 15712 34904 15761 34932
rect 15712 34892 15718 34904
rect 15749 34901 15761 34904
rect 15795 34901 15807 34935
rect 17144 34932 17172 35028
rect 20272 34941 20300 35040
rect 21913 35037 21925 35040
rect 21959 35037 21971 35071
rect 21913 35031 21971 35037
rect 32858 35028 32864 35080
rect 32916 35068 32922 35080
rect 33137 35071 33195 35077
rect 33137 35068 33149 35071
rect 32916 35040 33149 35068
rect 32916 35028 32922 35040
rect 33137 35037 33149 35040
rect 33183 35037 33195 35071
rect 33137 35031 33195 35037
rect 22278 34960 22284 35012
rect 22336 35000 22342 35012
rect 22465 35003 22523 35009
rect 22465 35000 22477 35003
rect 22336 34972 22477 35000
rect 22336 34960 22342 34972
rect 22465 34969 22477 34972
rect 22511 35000 22523 35003
rect 24210 35000 24216 35012
rect 22511 34972 24216 35000
rect 22511 34969 22523 34972
rect 22465 34963 22523 34969
rect 24210 34960 24216 34972
rect 24268 34960 24274 35012
rect 27062 34960 27068 35012
rect 27120 34960 27126 35012
rect 20257 34935 20315 34941
rect 20257 34932 20269 34935
rect 17144 34904 20269 34932
rect 15749 34895 15807 34901
rect 20257 34901 20269 34904
rect 20303 34901 20315 34935
rect 20257 34895 20315 34901
rect 32674 34892 32680 34944
rect 32732 34932 32738 34944
rect 32953 34935 33011 34941
rect 32953 34932 32965 34935
rect 32732 34904 32965 34932
rect 32732 34892 32738 34904
rect 32953 34901 32965 34904
rect 32999 34901 33011 34935
rect 32953 34895 33011 34901
rect 1104 34842 34840 34864
rect 1104 34790 9344 34842
rect 9396 34790 9408 34842
rect 9460 34790 9472 34842
rect 9524 34790 9536 34842
rect 9588 34790 9600 34842
rect 9652 34790 17738 34842
rect 17790 34790 17802 34842
rect 17854 34790 17866 34842
rect 17918 34790 17930 34842
rect 17982 34790 17994 34842
rect 18046 34790 26132 34842
rect 26184 34790 26196 34842
rect 26248 34790 26260 34842
rect 26312 34790 26324 34842
rect 26376 34790 26388 34842
rect 26440 34790 34526 34842
rect 34578 34790 34590 34842
rect 34642 34790 34654 34842
rect 34706 34790 34718 34842
rect 34770 34790 34782 34842
rect 34834 34790 34840 34842
rect 1104 34768 34840 34790
rect 12526 34728 12532 34740
rect 12406 34700 12532 34728
rect 7926 34620 7932 34672
rect 7984 34620 7990 34672
rect 9214 34660 9220 34672
rect 9154 34632 9220 34660
rect 9214 34620 9220 34632
rect 9272 34660 9278 34672
rect 9582 34660 9588 34672
rect 9272 34632 9588 34660
rect 9272 34620 9278 34632
rect 9582 34620 9588 34632
rect 9640 34620 9646 34672
rect 9766 34620 9772 34672
rect 9824 34660 9830 34672
rect 9861 34663 9919 34669
rect 9861 34660 9873 34663
rect 9824 34632 9873 34660
rect 9824 34620 9830 34632
rect 9861 34629 9873 34632
rect 9907 34629 9919 34663
rect 12406 34660 12434 34700
rect 12526 34688 12532 34700
rect 12584 34688 12590 34740
rect 13630 34728 13636 34740
rect 12636 34700 13636 34728
rect 12636 34669 12664 34700
rect 13630 34688 13636 34700
rect 13688 34688 13694 34740
rect 19334 34728 19340 34740
rect 14844 34700 15608 34728
rect 11086 34646 12434 34660
rect 9861 34623 9919 34629
rect 11072 34632 12434 34646
rect 12621 34663 12679 34669
rect 5718 34592 5724 34604
rect 5014 34564 5724 34592
rect 5718 34552 5724 34564
rect 5776 34552 5782 34604
rect 3602 34484 3608 34536
rect 3660 34484 3666 34536
rect 5902 34484 5908 34536
rect 5960 34524 5966 34536
rect 6365 34527 6423 34533
rect 6365 34524 6377 34527
rect 5960 34496 6377 34524
rect 5960 34484 5966 34496
rect 6365 34493 6377 34496
rect 6411 34493 6423 34527
rect 6365 34487 6423 34493
rect 7653 34527 7711 34533
rect 7653 34493 7665 34527
rect 7699 34493 7711 34527
rect 9585 34527 9643 34533
rect 9585 34524 9597 34527
rect 7653 34487 7711 34493
rect 8956 34496 9597 34524
rect 7668 34400 7696 34487
rect 8956 34400 8984 34496
rect 9585 34493 9597 34496
rect 9631 34493 9643 34527
rect 9585 34487 9643 34493
rect 10594 34484 10600 34536
rect 10652 34524 10658 34536
rect 11072 34524 11100 34632
rect 12621 34629 12633 34663
rect 12667 34629 12679 34663
rect 13906 34660 13912 34672
rect 13846 34632 13912 34660
rect 12621 34623 12679 34629
rect 13906 34620 13912 34632
rect 13964 34660 13970 34672
rect 14844 34660 14872 34700
rect 13964 34632 14872 34660
rect 13964 34620 13970 34632
rect 14182 34552 14188 34604
rect 14240 34552 14246 34604
rect 10652 34496 11100 34524
rect 10652 34484 10658 34496
rect 11330 34484 11336 34536
rect 11388 34484 11394 34536
rect 12345 34527 12403 34533
rect 12345 34493 12357 34527
rect 12391 34524 12403 34527
rect 14200 34524 14228 34552
rect 12391 34496 14228 34524
rect 12391 34493 12403 34496
rect 12345 34487 12403 34493
rect 14458 34484 14464 34536
rect 14516 34484 14522 34536
rect 15580 34456 15608 34700
rect 17328 34700 19340 34728
rect 17328 34604 17356 34700
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 20548 34700 22140 34728
rect 20548 34660 20576 34700
rect 22112 34669 22140 34700
rect 22554 34688 22560 34740
rect 22612 34728 22618 34740
rect 24302 34728 24308 34740
rect 22612 34700 24308 34728
rect 22612 34688 22618 34700
rect 24302 34688 24308 34700
rect 24360 34688 24366 34740
rect 26053 34731 26111 34737
rect 26053 34697 26065 34731
rect 26099 34728 26111 34731
rect 27062 34728 27068 34740
rect 26099 34700 27068 34728
rect 26099 34697 26111 34700
rect 26053 34691 26111 34697
rect 27062 34688 27068 34700
rect 27120 34688 27126 34740
rect 22097 34663 22155 34669
rect 18814 34632 20654 34660
rect 22097 34629 22109 34663
rect 22143 34660 22155 34663
rect 23106 34660 23112 34672
rect 22143 34632 23112 34660
rect 22143 34629 22155 34632
rect 22097 34623 22155 34629
rect 23106 34620 23112 34632
rect 23164 34620 23170 34672
rect 32401 34663 32459 34669
rect 23952 34632 25070 34660
rect 15746 34552 15752 34604
rect 15804 34592 15810 34604
rect 16025 34595 16083 34601
rect 16025 34592 16037 34595
rect 15804 34564 16037 34592
rect 15804 34552 15810 34564
rect 16025 34561 16037 34564
rect 16071 34561 16083 34595
rect 16574 34592 16580 34604
rect 16025 34555 16083 34561
rect 16132 34564 16580 34592
rect 15933 34527 15991 34533
rect 15933 34493 15945 34527
rect 15979 34524 15991 34527
rect 16132 34524 16160 34564
rect 16574 34552 16580 34564
rect 16632 34592 16638 34604
rect 16632 34564 17080 34592
rect 16632 34552 16638 34564
rect 15979 34496 16160 34524
rect 16301 34527 16359 34533
rect 15979 34493 15991 34496
rect 15933 34487 15991 34493
rect 16301 34493 16313 34527
rect 16347 34524 16359 34527
rect 16482 34524 16488 34536
rect 16347 34496 16488 34524
rect 16347 34493 16359 34496
rect 16301 34487 16359 34493
rect 16316 34456 16344 34487
rect 16482 34484 16488 34496
rect 16540 34484 16546 34536
rect 16758 34484 16764 34536
rect 16816 34484 16822 34536
rect 17052 34465 17080 34564
rect 17310 34552 17316 34604
rect 17368 34552 17374 34604
rect 19610 34552 19616 34604
rect 19668 34552 19674 34604
rect 19889 34595 19947 34601
rect 19889 34592 19901 34595
rect 19720 34564 19901 34592
rect 17586 34484 17592 34536
rect 17644 34484 17650 34536
rect 19334 34484 19340 34536
rect 19392 34524 19398 34536
rect 19720 34524 19748 34564
rect 19889 34561 19901 34564
rect 19935 34561 19947 34595
rect 19889 34555 19947 34561
rect 21821 34595 21879 34601
rect 21821 34561 21833 34595
rect 21867 34592 21879 34595
rect 22278 34592 22284 34604
rect 21867 34564 22284 34592
rect 21867 34561 21879 34564
rect 21821 34555 21879 34561
rect 22278 34552 22284 34564
rect 22336 34552 22342 34604
rect 20165 34527 20223 34533
rect 20165 34524 20177 34527
rect 19392 34496 19748 34524
rect 19812 34496 20177 34524
rect 19392 34484 19398 34496
rect 19812 34465 19840 34496
rect 20165 34493 20177 34496
rect 20211 34493 20223 34527
rect 20165 34487 20223 34493
rect 22370 34484 22376 34536
rect 22428 34484 22434 34536
rect 22646 34484 22652 34536
rect 22704 34484 22710 34536
rect 23106 34484 23112 34536
rect 23164 34524 23170 34536
rect 23952 34524 23980 34632
rect 32401 34629 32413 34663
rect 32447 34660 32459 34663
rect 32674 34660 32680 34672
rect 32447 34632 32680 34660
rect 32447 34629 32459 34632
rect 32401 34623 32459 34629
rect 32674 34620 32680 34632
rect 32732 34620 32738 34672
rect 24302 34552 24308 34604
rect 24360 34552 24366 34604
rect 33428 34564 33534 34592
rect 24581 34527 24639 34533
rect 24581 34524 24593 34527
rect 23164 34496 23980 34524
rect 24412 34496 24593 34524
rect 23164 34484 23170 34496
rect 15580 34428 16344 34456
rect 17037 34459 17095 34465
rect 17037 34425 17049 34459
rect 17083 34425 17095 34459
rect 17037 34419 17095 34425
rect 19797 34459 19855 34465
rect 19797 34425 19809 34459
rect 19843 34425 19855 34459
rect 19797 34419 19855 34425
rect 21560 34428 21772 34456
rect 3868 34391 3926 34397
rect 3868 34357 3880 34391
rect 3914 34388 3926 34391
rect 4614 34388 4620 34400
rect 3914 34360 4620 34388
rect 3914 34357 3926 34360
rect 3868 34351 3926 34357
rect 4614 34348 4620 34360
rect 4672 34348 4678 34400
rect 5353 34391 5411 34397
rect 5353 34357 5365 34391
rect 5399 34388 5411 34391
rect 5626 34388 5632 34400
rect 5399 34360 5632 34388
rect 5399 34357 5411 34360
rect 5353 34351 5411 34357
rect 5626 34348 5632 34360
rect 5684 34348 5690 34400
rect 7006 34348 7012 34400
rect 7064 34348 7070 34400
rect 7650 34348 7656 34400
rect 7708 34388 7714 34400
rect 8938 34388 8944 34400
rect 7708 34360 8944 34388
rect 7708 34348 7714 34360
rect 8938 34348 8944 34360
rect 8996 34348 9002 34400
rect 9398 34348 9404 34400
rect 9456 34348 9462 34400
rect 14090 34348 14096 34400
rect 14148 34348 14154 34400
rect 17221 34391 17279 34397
rect 17221 34357 17233 34391
rect 17267 34388 17279 34391
rect 18782 34388 18788 34400
rect 17267 34360 18788 34388
rect 17267 34357 17279 34360
rect 17221 34351 17279 34357
rect 18782 34348 18788 34360
rect 18840 34348 18846 34400
rect 19061 34391 19119 34397
rect 19061 34357 19073 34391
rect 19107 34388 19119 34391
rect 19334 34388 19340 34400
rect 19107 34360 19340 34388
rect 19107 34357 19119 34360
rect 19061 34351 19119 34357
rect 19334 34348 19340 34360
rect 19392 34348 19398 34400
rect 19978 34348 19984 34400
rect 20036 34388 20042 34400
rect 21560 34388 21588 34428
rect 20036 34360 21588 34388
rect 20036 34348 20042 34360
rect 21634 34348 21640 34400
rect 21692 34348 21698 34400
rect 21744 34388 21772 34428
rect 21818 34416 21824 34468
rect 21876 34456 21882 34468
rect 22388 34456 22416 34484
rect 24412 34456 24440 34496
rect 24581 34493 24593 34496
rect 24627 34493 24639 34527
rect 24581 34487 24639 34493
rect 32125 34527 32183 34533
rect 32125 34493 32137 34527
rect 32171 34524 32183 34527
rect 32398 34524 32404 34536
rect 32171 34496 32404 34524
rect 32171 34493 32183 34496
rect 32125 34487 32183 34493
rect 32398 34484 32404 34496
rect 32456 34484 32462 34536
rect 21876 34428 22416 34456
rect 23676 34428 24440 34456
rect 21876 34416 21882 34428
rect 23676 34388 23704 34428
rect 21744 34360 23704 34388
rect 24118 34348 24124 34400
rect 24176 34348 24182 34400
rect 32950 34348 32956 34400
rect 33008 34388 33014 34400
rect 33428 34388 33456 34564
rect 33008 34360 33456 34388
rect 33008 34348 33014 34360
rect 33870 34348 33876 34400
rect 33928 34348 33934 34400
rect 1104 34298 34684 34320
rect 1104 34246 5147 34298
rect 5199 34246 5211 34298
rect 5263 34246 5275 34298
rect 5327 34246 5339 34298
rect 5391 34246 5403 34298
rect 5455 34246 13541 34298
rect 13593 34246 13605 34298
rect 13657 34246 13669 34298
rect 13721 34246 13733 34298
rect 13785 34246 13797 34298
rect 13849 34246 21935 34298
rect 21987 34246 21999 34298
rect 22051 34246 22063 34298
rect 22115 34246 22127 34298
rect 22179 34246 22191 34298
rect 22243 34246 30329 34298
rect 30381 34246 30393 34298
rect 30445 34246 30457 34298
rect 30509 34246 30521 34298
rect 30573 34246 30585 34298
rect 30637 34246 34684 34298
rect 1104 34224 34684 34246
rect 4341 34187 4399 34193
rect 4341 34153 4353 34187
rect 4387 34153 4399 34187
rect 4341 34147 4399 34153
rect 4154 34076 4160 34128
rect 4212 34116 4218 34128
rect 4356 34116 4384 34147
rect 4614 34144 4620 34196
rect 4672 34144 4678 34196
rect 7837 34187 7895 34193
rect 7837 34184 7849 34187
rect 4724 34156 7849 34184
rect 4724 34116 4752 34156
rect 7837 34153 7849 34156
rect 7883 34184 7895 34187
rect 7926 34184 7932 34196
rect 7883 34156 7932 34184
rect 7883 34153 7895 34156
rect 7837 34147 7895 34153
rect 7926 34144 7932 34156
rect 7984 34144 7990 34196
rect 8021 34187 8079 34193
rect 8021 34153 8033 34187
rect 8067 34184 8079 34187
rect 8110 34184 8116 34196
rect 8067 34156 8116 34184
rect 8067 34153 8079 34156
rect 8021 34147 8079 34153
rect 8110 34144 8116 34156
rect 8168 34144 8174 34196
rect 14458 34144 14464 34196
rect 14516 34184 14522 34196
rect 14921 34187 14979 34193
rect 14921 34184 14933 34187
rect 14516 34156 14933 34184
rect 14516 34144 14522 34156
rect 14921 34153 14933 34156
rect 14967 34153 14979 34187
rect 14921 34147 14979 34153
rect 16758 34144 16764 34196
rect 16816 34184 16822 34196
rect 17037 34187 17095 34193
rect 17037 34184 17049 34187
rect 16816 34156 17049 34184
rect 16816 34144 16822 34156
rect 17037 34153 17049 34156
rect 17083 34153 17095 34187
rect 17037 34147 17095 34153
rect 17586 34144 17592 34196
rect 17644 34184 17650 34196
rect 17865 34187 17923 34193
rect 17865 34184 17877 34187
rect 17644 34156 17877 34184
rect 17644 34144 17650 34156
rect 17865 34153 17877 34156
rect 17911 34153 17923 34187
rect 17865 34147 17923 34153
rect 19610 34144 19616 34196
rect 19668 34184 19674 34196
rect 19705 34187 19763 34193
rect 19705 34184 19717 34187
rect 19668 34156 19717 34184
rect 19668 34144 19674 34156
rect 19705 34153 19717 34156
rect 19751 34153 19763 34187
rect 19705 34147 19763 34153
rect 22646 34144 22652 34196
rect 22704 34184 22710 34196
rect 22925 34187 22983 34193
rect 22925 34184 22937 34187
rect 22704 34156 22937 34184
rect 22704 34144 22710 34156
rect 22925 34153 22937 34156
rect 22971 34153 22983 34187
rect 22925 34147 22983 34153
rect 9582 34116 9588 34128
rect 4212 34088 4752 34116
rect 7024 34088 9588 34116
rect 4212 34076 4218 34088
rect 7024 34048 7052 34088
rect 9582 34076 9588 34088
rect 9640 34076 9646 34128
rect 5736 34020 7052 34048
rect 7101 34051 7159 34057
rect 5736 33992 5764 34020
rect 7101 34017 7113 34051
rect 7147 34048 7159 34051
rect 7650 34048 7656 34060
rect 7147 34020 7656 34048
rect 7147 34017 7159 34020
rect 7101 34011 7159 34017
rect 7650 34008 7656 34020
rect 7708 34008 7714 34060
rect 14090 34008 14096 34060
rect 14148 34008 14154 34060
rect 14182 34008 14188 34060
rect 14240 34048 14246 34060
rect 15102 34048 15108 34060
rect 14240 34020 15108 34048
rect 14240 34008 14246 34020
rect 15102 34008 15108 34020
rect 15160 34048 15166 34060
rect 15289 34051 15347 34057
rect 15289 34048 15301 34051
rect 15160 34020 15301 34048
rect 15160 34008 15166 34020
rect 15289 34017 15301 34020
rect 15335 34048 15347 34051
rect 17310 34048 17316 34060
rect 15335 34020 17316 34048
rect 15335 34017 15347 34020
rect 15289 34011 15347 34017
rect 17310 34008 17316 34020
rect 17368 34008 17374 34060
rect 18782 34008 18788 34060
rect 18840 34048 18846 34060
rect 20257 34051 20315 34057
rect 20257 34048 20269 34051
rect 18840 34020 20269 34048
rect 18840 34008 18846 34020
rect 20257 34017 20269 34020
rect 20303 34017 20315 34051
rect 20257 34011 20315 34017
rect 23382 34008 23388 34060
rect 23440 34048 23446 34060
rect 23937 34051 23995 34057
rect 23440 34020 23520 34048
rect 23440 34008 23446 34020
rect 3970 33940 3976 33992
rect 4028 33940 4034 33992
rect 4801 33983 4859 33989
rect 4801 33980 4813 33983
rect 4540 33952 4813 33980
rect 4338 33804 4344 33856
rect 4396 33804 4402 33856
rect 4540 33853 4568 33952
rect 4801 33949 4813 33952
rect 4847 33949 4859 33983
rect 4801 33943 4859 33949
rect 5718 33940 5724 33992
rect 5776 33940 5782 33992
rect 7469 33983 7527 33989
rect 7469 33980 7481 33983
rect 7116 33952 7481 33980
rect 6822 33872 6828 33924
rect 6880 33872 6886 33924
rect 7116 33856 7144 33952
rect 7469 33949 7481 33952
rect 7515 33949 7527 33983
rect 8481 33983 8539 33989
rect 8481 33980 8493 33983
rect 7469 33943 7527 33949
rect 7852 33952 8493 33980
rect 7852 33921 7880 33952
rect 8481 33949 8493 33952
rect 8527 33949 8539 33983
rect 8481 33943 8539 33949
rect 9398 33940 9404 33992
rect 9456 33940 9462 33992
rect 14108 33980 14136 34008
rect 14277 33983 14335 33989
rect 14277 33980 14289 33983
rect 14108 33952 14289 33980
rect 14277 33949 14289 33952
rect 14323 33949 14335 33983
rect 18049 33983 18107 33989
rect 14277 33943 14335 33949
rect 7837 33915 7895 33921
rect 7837 33881 7849 33915
rect 7883 33881 7895 33915
rect 7837 33875 7895 33881
rect 8018 33872 8024 33924
rect 8076 33912 8082 33924
rect 8113 33915 8171 33921
rect 8113 33912 8125 33915
rect 8076 33884 8125 33912
rect 8076 33872 8082 33884
rect 8113 33881 8125 33884
rect 8159 33881 8171 33915
rect 8113 33875 8171 33881
rect 8294 33872 8300 33924
rect 8352 33912 8358 33924
rect 9416 33912 9444 33940
rect 8352 33884 9444 33912
rect 15565 33915 15623 33921
rect 8352 33872 8358 33884
rect 15565 33881 15577 33915
rect 15611 33912 15623 33915
rect 15654 33912 15660 33924
rect 15611 33884 15660 33912
rect 15611 33881 15623 33884
rect 15565 33875 15623 33881
rect 15654 33872 15660 33884
rect 15712 33872 15718 33924
rect 4525 33847 4583 33853
rect 4525 33813 4537 33847
rect 4571 33813 4583 33847
rect 4525 33807 4583 33813
rect 5353 33847 5411 33853
rect 5353 33813 5365 33847
rect 5399 33844 5411 33847
rect 5902 33844 5908 33856
rect 5399 33816 5908 33844
rect 5399 33813 5411 33816
rect 5353 33807 5411 33813
rect 5902 33804 5908 33816
rect 5960 33804 5966 33856
rect 7098 33804 7104 33856
rect 7156 33804 7162 33856
rect 16482 33804 16488 33856
rect 16540 33844 16546 33856
rect 16684 33844 16712 33966
rect 18049 33949 18061 33983
rect 18095 33980 18107 33983
rect 18095 33952 18276 33980
rect 18095 33949 18107 33952
rect 18049 33943 18107 33949
rect 18248 33853 18276 33952
rect 19334 33940 19340 33992
rect 19392 33980 19398 33992
rect 20533 33983 20591 33989
rect 20533 33980 20545 33983
rect 19392 33952 20545 33980
rect 19392 33940 19398 33952
rect 20533 33949 20545 33952
rect 20579 33949 20591 33983
rect 20533 33943 20591 33949
rect 23109 33983 23167 33989
rect 23109 33949 23121 33983
rect 23155 33980 23167 33983
rect 23492 33980 23520 34020
rect 23937 34017 23949 34051
rect 23983 34017 23995 34051
rect 23937 34011 23995 34017
rect 23952 33980 23980 34011
rect 24210 34008 24216 34060
rect 24268 34048 24274 34060
rect 33781 34051 33839 34057
rect 24268 34020 27844 34048
rect 24268 34008 24274 34020
rect 23155 33952 23428 33980
rect 23492 33952 23980 33980
rect 23155 33949 23167 33952
rect 23109 33943 23167 33949
rect 18693 33915 18751 33921
rect 18693 33881 18705 33915
rect 18739 33912 18751 33915
rect 20073 33915 20131 33921
rect 20073 33912 20085 33915
rect 18739 33884 20085 33912
rect 18739 33881 18751 33884
rect 18693 33875 18751 33881
rect 20073 33881 20085 33884
rect 20119 33912 20131 33915
rect 20119 33884 20760 33912
rect 20119 33881 20131 33884
rect 20073 33875 20131 33881
rect 20732 33856 20760 33884
rect 16540 33816 16712 33844
rect 18233 33847 18291 33853
rect 16540 33804 16546 33816
rect 18233 33813 18245 33847
rect 18279 33813 18291 33847
rect 18233 33807 18291 33813
rect 18601 33847 18659 33853
rect 18601 33813 18613 33847
rect 18647 33844 18659 33847
rect 19334 33844 19340 33856
rect 18647 33816 19340 33844
rect 18647 33813 18659 33816
rect 18601 33807 18659 33813
rect 19334 33804 19340 33816
rect 19392 33804 19398 33856
rect 20162 33804 20168 33856
rect 20220 33844 20226 33856
rect 20625 33847 20683 33853
rect 20625 33844 20637 33847
rect 20220 33816 20637 33844
rect 20220 33804 20226 33816
rect 20625 33813 20637 33816
rect 20671 33813 20683 33847
rect 20625 33807 20683 33813
rect 20714 33804 20720 33856
rect 20772 33804 20778 33856
rect 23400 33853 23428 33952
rect 24118 33940 24124 33992
rect 24176 33980 24182 33992
rect 24489 33983 24547 33989
rect 24489 33980 24501 33983
rect 24176 33952 24501 33980
rect 24176 33940 24182 33952
rect 24489 33949 24501 33952
rect 24535 33949 24547 33983
rect 24489 33943 24547 33949
rect 26786 33940 26792 33992
rect 26844 33940 26850 33992
rect 26082 33884 26464 33912
rect 23385 33847 23443 33853
rect 23385 33813 23397 33847
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 23750 33804 23756 33856
rect 23808 33804 23814 33856
rect 23845 33847 23903 33853
rect 23845 33813 23857 33847
rect 23891 33844 23903 33847
rect 23934 33844 23940 33856
rect 23891 33816 23940 33844
rect 23891 33813 23903 33816
rect 23845 33807 23903 33813
rect 23934 33804 23940 33816
rect 23992 33844 23998 33856
rect 24581 33847 24639 33853
rect 24581 33844 24593 33847
rect 23992 33816 24593 33844
rect 23992 33804 23998 33816
rect 24581 33813 24593 33816
rect 24627 33813 24639 33847
rect 24581 33807 24639 33813
rect 25038 33804 25044 33856
rect 25096 33804 25102 33856
rect 26436 33844 26464 33884
rect 26510 33872 26516 33924
rect 26568 33872 26574 33924
rect 27816 33921 27844 34020
rect 33781 34017 33793 34051
rect 33827 34048 33839 34051
rect 33870 34048 33876 34060
rect 33827 34020 33876 34048
rect 33827 34017 33839 34020
rect 33781 34011 33839 34017
rect 33870 34008 33876 34020
rect 33928 34008 33934 34060
rect 26973 33915 27031 33921
rect 26973 33881 26985 33915
rect 27019 33881 27031 33915
rect 26973 33875 27031 33881
rect 27801 33915 27859 33921
rect 27801 33881 27813 33915
rect 27847 33912 27859 33915
rect 32950 33912 32956 33924
rect 27847 33884 32956 33912
rect 27847 33881 27859 33884
rect 27801 33875 27859 33881
rect 26988 33844 27016 33875
rect 32950 33872 32956 33884
rect 33008 33872 33014 33924
rect 27154 33844 27160 33856
rect 26436 33816 27160 33844
rect 27154 33804 27160 33816
rect 27212 33804 27218 33856
rect 34330 33804 34336 33856
rect 34388 33804 34394 33856
rect 1104 33754 34840 33776
rect 1104 33702 9344 33754
rect 9396 33702 9408 33754
rect 9460 33702 9472 33754
rect 9524 33702 9536 33754
rect 9588 33702 9600 33754
rect 9652 33702 17738 33754
rect 17790 33702 17802 33754
rect 17854 33702 17866 33754
rect 17918 33702 17930 33754
rect 17982 33702 17994 33754
rect 18046 33702 26132 33754
rect 26184 33702 26196 33754
rect 26248 33702 26260 33754
rect 26312 33702 26324 33754
rect 26376 33702 26388 33754
rect 26440 33702 34526 33754
rect 34578 33702 34590 33754
rect 34642 33702 34654 33754
rect 34706 33702 34718 33754
rect 34770 33702 34782 33754
rect 34834 33702 34840 33754
rect 1104 33680 34840 33702
rect 4338 33600 4344 33652
rect 4396 33640 4402 33652
rect 5629 33643 5687 33649
rect 5629 33640 5641 33643
rect 4396 33612 5641 33640
rect 4396 33600 4402 33612
rect 5629 33609 5641 33612
rect 5675 33609 5687 33643
rect 5902 33640 5908 33652
rect 5629 33603 5687 33609
rect 5736 33612 5908 33640
rect 5337 33575 5395 33581
rect 5337 33541 5349 33575
rect 5383 33572 5395 33575
rect 5537 33575 5595 33581
rect 5383 33544 5488 33572
rect 5383 33541 5395 33544
rect 5337 33535 5395 33541
rect 5460 33504 5488 33544
rect 5537 33541 5549 33575
rect 5583 33572 5595 33575
rect 5736 33572 5764 33612
rect 5902 33600 5908 33612
rect 5960 33600 5966 33652
rect 6365 33643 6423 33649
rect 6365 33609 6377 33643
rect 6411 33640 6423 33643
rect 6822 33640 6828 33652
rect 6411 33612 6828 33640
rect 6411 33609 6423 33612
rect 6365 33603 6423 33609
rect 6822 33600 6828 33612
rect 6880 33600 6886 33652
rect 17494 33640 17500 33652
rect 17420 33612 17500 33640
rect 5583 33544 5764 33572
rect 5583 33541 5595 33544
rect 5537 33535 5595 33541
rect 5810 33532 5816 33584
rect 5868 33572 5874 33584
rect 17420 33581 17448 33612
rect 17494 33600 17500 33612
rect 17552 33640 17558 33652
rect 18325 33643 18383 33649
rect 18325 33640 18337 33643
rect 17552 33612 18337 33640
rect 17552 33600 17558 33612
rect 18325 33609 18337 33612
rect 18371 33609 18383 33643
rect 19978 33640 19984 33652
rect 18325 33603 18383 33609
rect 18616 33612 19984 33640
rect 17405 33575 17463 33581
rect 5868 33544 7328 33572
rect 5868 33532 5874 33544
rect 5460 33476 6500 33504
rect 5810 33396 5816 33448
rect 5868 33396 5874 33448
rect 5902 33396 5908 33448
rect 5960 33396 5966 33448
rect 5994 33396 6000 33448
rect 6052 33396 6058 33448
rect 6089 33439 6147 33445
rect 6089 33405 6101 33439
rect 6135 33405 6147 33439
rect 6472 33436 6500 33476
rect 6546 33464 6552 33516
rect 6604 33464 6610 33516
rect 6825 33507 6883 33513
rect 6825 33473 6837 33507
rect 6871 33473 6883 33507
rect 6825 33467 6883 33473
rect 6840 33436 6868 33467
rect 7006 33464 7012 33516
rect 7064 33464 7070 33516
rect 7300 33513 7328 33544
rect 17405 33541 17417 33575
rect 17451 33541 17463 33575
rect 17405 33535 17463 33541
rect 17865 33575 17923 33581
rect 17865 33541 17877 33575
rect 17911 33572 17923 33575
rect 18616 33572 18644 33612
rect 19978 33600 19984 33612
rect 20036 33600 20042 33652
rect 20162 33600 20168 33652
rect 20220 33600 20226 33652
rect 20533 33643 20591 33649
rect 20533 33609 20545 33643
rect 20579 33640 20591 33643
rect 21082 33640 21088 33652
rect 20579 33612 21088 33640
rect 20579 33609 20591 33612
rect 20533 33603 20591 33609
rect 21082 33600 21088 33612
rect 21140 33600 21146 33652
rect 21634 33600 21640 33652
rect 21692 33600 21698 33652
rect 23750 33600 23756 33652
rect 23808 33640 23814 33652
rect 24762 33640 24768 33652
rect 23808 33612 24768 33640
rect 23808 33600 23814 33612
rect 24762 33600 24768 33612
rect 24820 33640 24826 33652
rect 24949 33643 25007 33649
rect 24949 33640 24961 33643
rect 24820 33612 24961 33640
rect 24820 33600 24826 33612
rect 24949 33609 24961 33612
rect 24995 33609 25007 33643
rect 24949 33603 25007 33609
rect 25038 33600 25044 33652
rect 25096 33600 25102 33652
rect 26510 33600 26516 33652
rect 26568 33640 26574 33652
rect 26605 33643 26663 33649
rect 26605 33640 26617 33643
rect 26568 33612 26617 33640
rect 26568 33600 26574 33612
rect 26605 33609 26617 33612
rect 26651 33609 26663 33643
rect 26605 33603 26663 33609
rect 17911 33544 18644 33572
rect 18693 33575 18751 33581
rect 17911 33541 17923 33544
rect 17865 33535 17923 33541
rect 18693 33541 18705 33575
rect 18739 33572 18751 33575
rect 19702 33572 19708 33584
rect 18739 33544 19708 33572
rect 18739 33541 18751 33544
rect 18693 33535 18751 33541
rect 19702 33532 19708 33544
rect 19760 33532 19766 33584
rect 20180 33572 20208 33600
rect 20180 33544 20852 33572
rect 7285 33507 7343 33513
rect 7285 33473 7297 33507
rect 7331 33473 7343 33507
rect 7285 33467 7343 33473
rect 7469 33507 7527 33513
rect 7469 33473 7481 33507
rect 7515 33504 7527 33507
rect 8294 33504 8300 33516
rect 7515 33476 8300 33504
rect 7515 33473 7527 33476
rect 7469 33467 7527 33473
rect 7098 33436 7104 33448
rect 6472 33408 7104 33436
rect 6089 33399 6147 33405
rect 6104 33368 6132 33399
rect 7098 33396 7104 33408
rect 7156 33396 7162 33448
rect 5644 33340 6132 33368
rect 5644 33312 5672 33340
rect 6178 33328 6184 33380
rect 6236 33368 6242 33380
rect 7484 33368 7512 33467
rect 8294 33464 8300 33476
rect 8352 33464 8358 33516
rect 8846 33464 8852 33516
rect 8904 33464 8910 33516
rect 16666 33464 16672 33516
rect 16724 33504 16730 33516
rect 17497 33507 17555 33513
rect 17497 33504 17509 33507
rect 16724 33476 17509 33504
rect 16724 33464 16730 33476
rect 17497 33473 17509 33476
rect 17543 33473 17555 33507
rect 17497 33467 17555 33473
rect 18785 33507 18843 33513
rect 18785 33473 18797 33507
rect 18831 33504 18843 33507
rect 19153 33507 19211 33513
rect 19153 33504 19165 33507
rect 18831 33476 19165 33504
rect 18831 33473 18843 33476
rect 18785 33467 18843 33473
rect 19153 33473 19165 33476
rect 19199 33473 19211 33507
rect 19153 33467 19211 33473
rect 19242 33464 19248 33516
rect 19300 33504 19306 33516
rect 19337 33507 19395 33513
rect 19337 33504 19349 33507
rect 19300 33476 19349 33504
rect 19300 33464 19306 33476
rect 19337 33473 19349 33476
rect 19383 33504 19395 33507
rect 20073 33507 20131 33513
rect 19383 33476 20024 33504
rect 19383 33473 19395 33476
rect 19337 33467 19395 33473
rect 17218 33396 17224 33448
rect 17276 33396 17282 33448
rect 17773 33439 17831 33445
rect 17773 33405 17785 33439
rect 17819 33405 17831 33439
rect 17773 33399 17831 33405
rect 18969 33439 19027 33445
rect 18969 33405 18981 33439
rect 19015 33436 19027 33439
rect 19613 33439 19671 33445
rect 19613 33436 19625 33439
rect 19015 33408 19288 33436
rect 19015 33405 19027 33408
rect 18969 33399 19027 33405
rect 6236 33340 7512 33368
rect 6236 33328 6242 33340
rect 13446 33328 13452 33380
rect 13504 33368 13510 33380
rect 17788 33368 17816 33399
rect 13504 33340 17816 33368
rect 13504 33328 13510 33340
rect 3970 33260 3976 33312
rect 4028 33300 4034 33312
rect 5169 33303 5227 33309
rect 5169 33300 5181 33303
rect 4028 33272 5181 33300
rect 4028 33260 4034 33272
rect 5169 33269 5181 33272
rect 5215 33269 5227 33303
rect 5169 33263 5227 33269
rect 5353 33303 5411 33309
rect 5353 33269 5365 33303
rect 5399 33300 5411 33303
rect 5626 33300 5632 33312
rect 5399 33272 5632 33300
rect 5399 33269 5411 33272
rect 5353 33263 5411 33269
rect 5626 33260 5632 33272
rect 5684 33260 5690 33312
rect 5902 33260 5908 33312
rect 5960 33300 5966 33312
rect 6362 33300 6368 33312
rect 5960 33272 6368 33300
rect 5960 33260 5966 33272
rect 6362 33260 6368 33272
rect 6420 33260 6426 33312
rect 9033 33303 9091 33309
rect 9033 33269 9045 33303
rect 9079 33300 9091 33303
rect 9122 33300 9128 33312
rect 9079 33272 9128 33300
rect 9079 33269 9091 33272
rect 9033 33263 9091 33269
rect 9122 33260 9128 33272
rect 9180 33260 9186 33312
rect 17034 33260 17040 33312
rect 17092 33300 17098 33312
rect 17681 33303 17739 33309
rect 17681 33300 17693 33303
rect 17092 33272 17693 33300
rect 17092 33260 17098 33272
rect 17681 33269 17693 33272
rect 17727 33269 17739 33303
rect 19260 33300 19288 33408
rect 19352 33408 19625 33436
rect 19352 33380 19380 33408
rect 19613 33405 19625 33408
rect 19659 33405 19671 33439
rect 19996 33436 20024 33476
rect 20073 33473 20085 33507
rect 20119 33504 20131 33507
rect 20180 33504 20208 33544
rect 20119 33476 20208 33504
rect 20257 33507 20315 33513
rect 20119 33473 20131 33476
rect 20073 33467 20131 33473
rect 20257 33473 20269 33507
rect 20303 33504 20315 33507
rect 20530 33504 20536 33516
rect 20303 33476 20536 33504
rect 20303 33473 20315 33476
rect 20257 33467 20315 33473
rect 20530 33464 20536 33476
rect 20588 33464 20594 33516
rect 20824 33513 20852 33544
rect 20809 33507 20867 33513
rect 20809 33473 20821 33507
rect 20855 33473 20867 33507
rect 20809 33467 20867 33473
rect 20993 33507 21051 33513
rect 20993 33473 21005 33507
rect 21039 33504 21051 33507
rect 21652 33504 21680 33600
rect 23106 33532 23112 33584
rect 23164 33532 23170 33584
rect 21039 33476 21680 33504
rect 25056 33504 25084 33600
rect 25501 33507 25559 33513
rect 25501 33504 25513 33507
rect 25056 33476 25513 33504
rect 21039 33473 21051 33476
rect 20993 33467 21051 33473
rect 25501 33473 25513 33476
rect 25547 33473 25559 33507
rect 25501 33467 25559 33473
rect 20625 33439 20683 33445
rect 20625 33436 20637 33439
rect 19996 33408 20637 33436
rect 19613 33399 19671 33405
rect 20625 33405 20637 33408
rect 20671 33436 20683 33439
rect 20714 33436 20720 33448
rect 20671 33408 20720 33436
rect 20671 33405 20683 33408
rect 20625 33399 20683 33405
rect 20714 33396 20720 33408
rect 20772 33436 20778 33448
rect 21008 33436 21036 33467
rect 20772 33408 21036 33436
rect 20772 33396 20778 33408
rect 21818 33396 21824 33448
rect 21876 33396 21882 33448
rect 22097 33439 22155 33445
rect 22097 33405 22109 33439
rect 22143 33436 22155 33439
rect 22186 33436 22192 33448
rect 22143 33408 22192 33436
rect 22143 33405 22155 33408
rect 22097 33399 22155 33405
rect 22186 33396 22192 33408
rect 22244 33396 22250 33448
rect 25958 33396 25964 33448
rect 26016 33396 26022 33448
rect 19334 33328 19340 33380
rect 19392 33328 19398 33380
rect 19444 33340 20576 33368
rect 19444 33300 19472 33340
rect 20548 33312 20576 33340
rect 19260 33272 19472 33300
rect 17681 33263 17739 33269
rect 19518 33260 19524 33312
rect 19576 33260 19582 33312
rect 20530 33260 20536 33312
rect 20588 33260 20594 33312
rect 20990 33260 20996 33312
rect 21048 33300 21054 33312
rect 21177 33303 21235 33309
rect 21177 33300 21189 33303
rect 21048 33272 21189 33300
rect 21048 33260 21054 33272
rect 21177 33269 21189 33272
rect 21223 33269 21235 33303
rect 21177 33263 21235 33269
rect 23566 33260 23572 33312
rect 23624 33260 23630 33312
rect 1104 33210 34684 33232
rect 1104 33158 5147 33210
rect 5199 33158 5211 33210
rect 5263 33158 5275 33210
rect 5327 33158 5339 33210
rect 5391 33158 5403 33210
rect 5455 33158 13541 33210
rect 13593 33158 13605 33210
rect 13657 33158 13669 33210
rect 13721 33158 13733 33210
rect 13785 33158 13797 33210
rect 13849 33158 21935 33210
rect 21987 33158 21999 33210
rect 22051 33158 22063 33210
rect 22115 33158 22127 33210
rect 22179 33158 22191 33210
rect 22243 33158 30329 33210
rect 30381 33158 30393 33210
rect 30445 33158 30457 33210
rect 30509 33158 30521 33210
rect 30573 33158 30585 33210
rect 30637 33158 34684 33210
rect 1104 33136 34684 33158
rect 6546 33056 6552 33108
rect 6604 33096 6610 33108
rect 6641 33099 6699 33105
rect 6641 33096 6653 33099
rect 6604 33068 6653 33096
rect 6604 33056 6610 33068
rect 6641 33065 6653 33068
rect 6687 33065 6699 33099
rect 6641 33059 6699 33065
rect 7926 33056 7932 33108
rect 7984 33096 7990 33108
rect 8294 33096 8300 33108
rect 7984 33068 8300 33096
rect 7984 33056 7990 33068
rect 8294 33056 8300 33068
rect 8352 33096 8358 33108
rect 8481 33099 8539 33105
rect 8481 33096 8493 33099
rect 8352 33068 8493 33096
rect 8352 33056 8358 33068
rect 8481 33065 8493 33068
rect 8527 33065 8539 33099
rect 8481 33059 8539 33065
rect 8665 33099 8723 33105
rect 8665 33065 8677 33099
rect 8711 33096 8723 33099
rect 8846 33096 8852 33108
rect 8711 33068 8852 33096
rect 8711 33065 8723 33068
rect 8665 33059 8723 33065
rect 8846 33056 8852 33068
rect 8904 33056 8910 33108
rect 9048 33068 13032 33096
rect 6178 32988 6184 33040
rect 6236 33028 6242 33040
rect 9048 33028 9076 33068
rect 6236 33000 9076 33028
rect 6236 32988 6242 33000
rect 1673 32963 1731 32969
rect 1673 32929 1685 32963
rect 1719 32960 1731 32963
rect 1719 32932 12848 32960
rect 1719 32929 1731 32932
rect 1673 32923 1731 32929
rect 12820 32904 12848 32932
rect 934 32852 940 32904
rect 992 32892 998 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 992 32864 1409 32892
rect 992 32852 998 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 3970 32852 3976 32904
rect 4028 32892 4034 32904
rect 4249 32895 4307 32901
rect 4249 32892 4261 32895
rect 4028 32864 4261 32892
rect 4028 32852 4034 32864
rect 4249 32861 4261 32864
rect 4295 32861 4307 32895
rect 4249 32855 4307 32861
rect 5810 32852 5816 32904
rect 5868 32852 5874 32904
rect 6178 32852 6184 32904
rect 6236 32852 6242 32904
rect 6270 32852 6276 32904
rect 6328 32852 6334 32904
rect 6362 32852 6368 32904
rect 6420 32852 6426 32904
rect 6457 32895 6515 32901
rect 6457 32861 6469 32895
rect 6503 32892 6515 32895
rect 8018 32892 8024 32904
rect 6503 32864 8024 32892
rect 6503 32861 6515 32864
rect 6457 32855 6515 32861
rect 4065 32827 4123 32833
rect 4065 32824 4077 32827
rect 3528 32796 4077 32824
rect 3528 32768 3556 32796
rect 4065 32793 4077 32796
rect 4111 32793 4123 32827
rect 5828 32824 5856 32852
rect 6472 32824 6500 32855
rect 8018 32852 8024 32864
rect 8076 32892 8082 32904
rect 8113 32895 8171 32901
rect 8113 32892 8125 32895
rect 8076 32864 8125 32892
rect 8076 32852 8082 32864
rect 8113 32861 8125 32864
rect 8159 32861 8171 32895
rect 8113 32855 8171 32861
rect 8938 32852 8944 32904
rect 8996 32852 9002 32904
rect 12802 32852 12808 32904
rect 12860 32852 12866 32904
rect 13004 32901 13032 33068
rect 14936 33068 16712 33096
rect 13446 32920 13452 32972
rect 13504 32920 13510 32972
rect 12989 32895 13047 32901
rect 12989 32861 13001 32895
rect 13035 32892 13047 32895
rect 13464 32892 13492 32920
rect 13035 32864 13492 32892
rect 13035 32861 13047 32864
rect 12989 32855 13047 32861
rect 14734 32852 14740 32904
rect 14792 32852 14798 32904
rect 14829 32895 14887 32901
rect 14829 32861 14841 32895
rect 14875 32892 14887 32895
rect 14936 32892 14964 33068
rect 16684 33040 16712 33068
rect 19702 33056 19708 33108
rect 19760 33096 19766 33108
rect 19797 33099 19855 33105
rect 19797 33096 19809 33099
rect 19760 33068 19809 33096
rect 19760 33056 19766 33068
rect 19797 33065 19809 33068
rect 19843 33065 19855 33099
rect 19797 33059 19855 33065
rect 22005 33099 22063 33105
rect 22005 33065 22017 33099
rect 22051 33096 22063 33099
rect 22278 33096 22284 33108
rect 22051 33068 22284 33096
rect 22051 33065 22063 33068
rect 22005 33059 22063 33065
rect 22278 33056 22284 33068
rect 22336 33056 22342 33108
rect 23014 33056 23020 33108
rect 23072 33096 23078 33108
rect 24578 33096 24584 33108
rect 23072 33068 24584 33096
rect 23072 33056 23078 33068
rect 24578 33056 24584 33068
rect 24636 33056 24642 33108
rect 25317 33099 25375 33105
rect 25317 33065 25329 33099
rect 25363 33096 25375 33099
rect 25958 33096 25964 33108
rect 25363 33068 25964 33096
rect 25363 33065 25375 33068
rect 25317 33059 25375 33065
rect 25958 33056 25964 33068
rect 26016 33056 26022 33108
rect 15013 33031 15071 33037
rect 15013 32997 15025 33031
rect 15059 33028 15071 33031
rect 15059 33000 15240 33028
rect 15059 32997 15071 33000
rect 15013 32991 15071 32997
rect 15102 32920 15108 32972
rect 15160 32920 15166 32972
rect 15212 32960 15240 33000
rect 16666 32988 16672 33040
rect 16724 32988 16730 33040
rect 15381 32963 15439 32969
rect 15381 32960 15393 32963
rect 15212 32932 15393 32960
rect 15381 32929 15393 32932
rect 15427 32929 15439 32963
rect 15381 32923 15439 32929
rect 16574 32920 16580 32972
rect 16632 32920 16638 32972
rect 16853 32963 16911 32969
rect 16853 32929 16865 32963
rect 16899 32960 16911 32963
rect 17218 32960 17224 32972
rect 16899 32932 17224 32960
rect 16899 32929 16911 32932
rect 16853 32923 16911 32929
rect 17218 32920 17224 32932
rect 17276 32920 17282 32972
rect 23109 32963 23167 32969
rect 22066 32932 22968 32960
rect 16592 32892 16620 32920
rect 14875 32864 14964 32892
rect 16514 32864 16620 32892
rect 14875 32861 14887 32864
rect 14829 32855 14887 32861
rect 19242 32852 19248 32904
rect 19300 32852 19306 32904
rect 19705 32895 19763 32901
rect 19705 32892 19717 32895
rect 19536 32864 19717 32892
rect 5828 32796 6500 32824
rect 8404 32796 9076 32824
rect 4065 32787 4123 32793
rect 3510 32716 3516 32768
rect 3568 32716 3574 32768
rect 3878 32716 3884 32768
rect 3936 32716 3942 32768
rect 4890 32716 4896 32768
rect 4948 32756 4954 32768
rect 8404 32756 8432 32796
rect 4948 32728 8432 32756
rect 4948 32716 4954 32728
rect 8478 32716 8484 32768
rect 8536 32716 8542 32768
rect 9048 32756 9076 32796
rect 9122 32784 9128 32836
rect 9180 32824 9186 32836
rect 9217 32827 9275 32833
rect 9217 32824 9229 32827
rect 9180 32796 9229 32824
rect 9180 32784 9186 32796
rect 9217 32793 9229 32796
rect 9263 32793 9275 32827
rect 9217 32787 9275 32793
rect 9674 32784 9680 32836
rect 9732 32784 9738 32836
rect 15013 32827 15071 32833
rect 15013 32793 15025 32827
rect 15059 32824 15071 32827
rect 15378 32824 15384 32836
rect 15059 32796 15384 32824
rect 15059 32793 15071 32796
rect 15013 32787 15071 32793
rect 15378 32784 15384 32796
rect 15436 32784 15442 32836
rect 19334 32784 19340 32836
rect 19392 32824 19398 32836
rect 19429 32827 19487 32833
rect 19429 32824 19441 32827
rect 19392 32796 19441 32824
rect 19392 32784 19398 32796
rect 19429 32793 19441 32796
rect 19475 32793 19487 32827
rect 19429 32787 19487 32793
rect 19536 32824 19564 32864
rect 19705 32861 19717 32864
rect 19751 32861 19763 32895
rect 19705 32855 19763 32861
rect 19889 32895 19947 32901
rect 19889 32861 19901 32895
rect 19935 32892 19947 32895
rect 20990 32892 20996 32904
rect 19935 32864 20996 32892
rect 19935 32861 19947 32864
rect 19889 32855 19947 32861
rect 20990 32852 20996 32864
rect 21048 32852 21054 32904
rect 22066 32824 22094 32932
rect 22940 32901 22968 32932
rect 23109 32929 23121 32963
rect 23155 32960 23167 32963
rect 23382 32960 23388 32972
rect 23155 32932 23388 32960
rect 23155 32929 23167 32932
rect 23109 32923 23167 32929
rect 23382 32920 23388 32932
rect 23440 32920 23446 32972
rect 23566 32920 23572 32972
rect 23624 32920 23630 32972
rect 24302 32920 24308 32972
rect 24360 32960 24366 32972
rect 24360 32932 26372 32960
rect 24360 32920 24366 32932
rect 22189 32895 22247 32901
rect 22189 32861 22201 32895
rect 22235 32892 22247 32895
rect 22925 32895 22983 32901
rect 22235 32864 22508 32892
rect 22235 32861 22247 32864
rect 22189 32855 22247 32861
rect 19536 32796 22094 32824
rect 19536 32768 19564 32796
rect 9858 32756 9864 32768
rect 9048 32728 9864 32756
rect 9858 32716 9864 32728
rect 9916 32716 9922 32768
rect 10686 32716 10692 32768
rect 10744 32716 10750 32768
rect 17586 32716 17592 32768
rect 17644 32756 17650 32768
rect 17865 32759 17923 32765
rect 17865 32756 17877 32759
rect 17644 32728 17877 32756
rect 17644 32716 17650 32728
rect 17865 32725 17877 32728
rect 17911 32725 17923 32759
rect 17865 32719 17923 32725
rect 19518 32716 19524 32768
rect 19576 32716 19582 32768
rect 19610 32716 19616 32768
rect 19668 32716 19674 32768
rect 22480 32765 22508 32864
rect 22925 32861 22937 32895
rect 22971 32892 22983 32895
rect 23584 32892 23612 32920
rect 22971 32864 23612 32892
rect 22971 32861 22983 32864
rect 22925 32855 22983 32861
rect 24762 32852 24768 32904
rect 24820 32852 24826 32904
rect 25133 32895 25191 32901
rect 25133 32892 25145 32895
rect 24872 32864 25145 32892
rect 24394 32784 24400 32836
rect 24452 32824 24458 32836
rect 24872 32824 24900 32864
rect 25133 32861 25145 32864
rect 25179 32861 25191 32895
rect 25133 32855 25191 32861
rect 24452 32796 24900 32824
rect 24452 32784 24458 32796
rect 24946 32784 24952 32836
rect 25004 32784 25010 32836
rect 25038 32784 25044 32836
rect 25096 32784 25102 32836
rect 22465 32759 22523 32765
rect 22465 32725 22477 32759
rect 22511 32725 22523 32759
rect 22465 32719 22523 32725
rect 22833 32759 22891 32765
rect 22833 32725 22845 32759
rect 22879 32756 22891 32759
rect 25056 32756 25084 32784
rect 26344 32765 26372 32932
rect 32398 32920 32404 32972
rect 32456 32960 32462 32972
rect 34333 32963 34391 32969
rect 34333 32960 34345 32963
rect 32456 32932 34345 32960
rect 32456 32920 32462 32932
rect 34333 32929 34345 32932
rect 34379 32929 34391 32963
rect 34333 32923 34391 32929
rect 26970 32852 26976 32904
rect 27028 32852 27034 32904
rect 32950 32852 32956 32904
rect 33008 32852 33014 32904
rect 34057 32827 34115 32833
rect 34057 32793 34069 32827
rect 34103 32824 34115 32827
rect 34330 32824 34336 32836
rect 34103 32796 34336 32824
rect 34103 32793 34115 32796
rect 34057 32787 34115 32793
rect 34330 32784 34336 32796
rect 34388 32784 34394 32836
rect 22879 32728 25084 32756
rect 26329 32759 26387 32765
rect 22879 32725 22891 32728
rect 22833 32719 22891 32725
rect 26329 32725 26341 32759
rect 26375 32756 26387 32759
rect 28350 32756 28356 32768
rect 26375 32728 28356 32756
rect 26375 32725 26387 32728
rect 26329 32719 26387 32725
rect 28350 32716 28356 32728
rect 28408 32716 28414 32768
rect 32582 32716 32588 32768
rect 32640 32716 32646 32768
rect 1104 32666 34840 32688
rect 1104 32614 9344 32666
rect 9396 32614 9408 32666
rect 9460 32614 9472 32666
rect 9524 32614 9536 32666
rect 9588 32614 9600 32666
rect 9652 32614 17738 32666
rect 17790 32614 17802 32666
rect 17854 32614 17866 32666
rect 17918 32614 17930 32666
rect 17982 32614 17994 32666
rect 18046 32614 26132 32666
rect 26184 32614 26196 32666
rect 26248 32614 26260 32666
rect 26312 32614 26324 32666
rect 26376 32614 26388 32666
rect 26440 32614 34526 32666
rect 34578 32614 34590 32666
rect 34642 32614 34654 32666
rect 34706 32614 34718 32666
rect 34770 32614 34782 32666
rect 34834 32614 34840 32666
rect 1104 32592 34840 32614
rect 3878 32512 3884 32564
rect 3936 32512 3942 32564
rect 8018 32512 8024 32564
rect 8076 32512 8082 32564
rect 8478 32512 8484 32564
rect 8536 32552 8542 32564
rect 8941 32555 8999 32561
rect 8941 32552 8953 32555
rect 8536 32524 8953 32552
rect 8536 32512 8542 32524
rect 8941 32521 8953 32524
rect 8987 32521 8999 32555
rect 8941 32515 8999 32521
rect 9674 32512 9680 32564
rect 9732 32552 9738 32564
rect 10318 32552 10324 32564
rect 9732 32524 10324 32552
rect 9732 32512 9738 32524
rect 10318 32512 10324 32524
rect 10376 32512 10382 32564
rect 10686 32512 10692 32564
rect 10744 32512 10750 32564
rect 15102 32552 15108 32564
rect 12360 32524 15108 32552
rect 4338 32484 4344 32496
rect 3358 32456 4344 32484
rect 4338 32444 4344 32456
rect 4396 32444 4402 32496
rect 6270 32444 6276 32496
rect 6328 32484 6334 32496
rect 8202 32493 8208 32496
rect 6708 32487 6766 32493
rect 6708 32484 6720 32487
rect 6328 32456 6720 32484
rect 6328 32444 6334 32456
rect 6708 32453 6720 32456
rect 6754 32453 6766 32487
rect 6708 32447 6766 32453
rect 8189 32487 8208 32493
rect 8189 32453 8201 32487
rect 8189 32447 8208 32453
rect 8202 32444 8208 32447
rect 8260 32444 8266 32496
rect 8389 32487 8447 32493
rect 8389 32453 8401 32487
rect 8435 32484 8447 32487
rect 9030 32484 9036 32496
rect 8435 32456 9036 32484
rect 8435 32453 8447 32456
rect 8389 32447 8447 32453
rect 9030 32444 9036 32456
rect 9088 32444 9094 32496
rect 4433 32419 4491 32425
rect 4433 32416 4445 32419
rect 4264 32388 4445 32416
rect 1857 32351 1915 32357
rect 1857 32317 1869 32351
rect 1903 32317 1915 32351
rect 1857 32311 1915 32317
rect 1872 32212 1900 32311
rect 2130 32308 2136 32360
rect 2188 32308 2194 32360
rect 3602 32348 3608 32360
rect 3160 32320 3608 32348
rect 2774 32212 2780 32224
rect 1872 32184 2780 32212
rect 2774 32172 2780 32184
rect 2832 32212 2838 32224
rect 3160 32212 3188 32320
rect 3602 32308 3608 32320
rect 3660 32308 3666 32360
rect 4264 32357 4292 32388
rect 4433 32385 4445 32388
rect 4479 32385 4491 32419
rect 4433 32379 4491 32385
rect 4614 32376 4620 32428
rect 4672 32376 4678 32428
rect 6825 32419 6883 32425
rect 6825 32385 6837 32419
rect 6871 32416 6883 32419
rect 9401 32419 9459 32425
rect 9401 32416 9413 32419
rect 6871 32388 9413 32416
rect 6871 32385 6883 32388
rect 6825 32379 6883 32385
rect 4249 32351 4307 32357
rect 4249 32317 4261 32351
rect 4295 32317 4307 32351
rect 4249 32311 4307 32317
rect 4264 32224 4292 32311
rect 6914 32308 6920 32360
rect 6972 32308 6978 32360
rect 7193 32351 7251 32357
rect 7193 32317 7205 32351
rect 7239 32317 7251 32351
rect 7193 32311 7251 32317
rect 6362 32240 6368 32292
rect 6420 32280 6426 32292
rect 7208 32280 7236 32311
rect 6420 32252 7236 32280
rect 6420 32240 6426 32252
rect 2832 32184 3188 32212
rect 2832 32172 2838 32184
rect 3602 32172 3608 32224
rect 3660 32172 3666 32224
rect 3694 32172 3700 32224
rect 3752 32172 3758 32224
rect 3881 32215 3939 32221
rect 3881 32181 3893 32215
rect 3927 32212 3939 32215
rect 4154 32212 4160 32224
rect 3927 32184 4160 32212
rect 3927 32181 3939 32184
rect 3881 32175 3939 32181
rect 4154 32172 4160 32184
rect 4212 32172 4218 32224
rect 4246 32172 4252 32224
rect 4304 32172 4310 32224
rect 4801 32215 4859 32221
rect 4801 32181 4813 32215
rect 4847 32212 4859 32215
rect 4982 32212 4988 32224
rect 4847 32184 4988 32212
rect 4847 32181 4859 32184
rect 4801 32175 4859 32181
rect 4982 32172 4988 32184
rect 5040 32172 5046 32224
rect 6546 32172 6552 32224
rect 6604 32172 6610 32224
rect 8220 32221 8248 32388
rect 9401 32385 9413 32388
rect 9447 32416 9459 32419
rect 10704 32416 10732 32512
rect 12360 32428 12388 32524
rect 15102 32512 15108 32524
rect 15160 32512 15166 32564
rect 15378 32512 15384 32564
rect 15436 32512 15442 32564
rect 16666 32512 16672 32564
rect 16724 32512 16730 32564
rect 17034 32512 17040 32564
rect 17092 32512 17098 32564
rect 17586 32512 17592 32564
rect 17644 32512 17650 32564
rect 19610 32552 19616 32564
rect 19444 32524 19616 32552
rect 14090 32444 14096 32496
rect 14148 32484 14154 32496
rect 14461 32487 14519 32493
rect 14461 32484 14473 32487
rect 14148 32456 14473 32484
rect 14148 32444 14154 32456
rect 14461 32453 14473 32456
rect 14507 32453 14519 32487
rect 14461 32447 14519 32453
rect 14734 32444 14740 32496
rect 14792 32484 14798 32496
rect 14921 32487 14979 32493
rect 14921 32484 14933 32487
rect 14792 32456 14933 32484
rect 14792 32444 14798 32456
rect 9447 32388 10732 32416
rect 9447 32385 9459 32388
rect 9401 32379 9459 32385
rect 12342 32376 12348 32428
rect 12400 32416 12406 32428
rect 12437 32419 12495 32425
rect 12437 32416 12449 32419
rect 12400 32388 12449 32416
rect 12400 32376 12406 32388
rect 12437 32385 12449 32388
rect 12483 32385 12495 32419
rect 12437 32379 12495 32385
rect 13814 32376 13820 32428
rect 13872 32376 13878 32428
rect 14844 32425 14872 32456
rect 14921 32453 14933 32456
rect 14967 32484 14979 32487
rect 14967 32456 15608 32484
rect 14967 32453 14979 32456
rect 14921 32447 14979 32453
rect 14829 32419 14887 32425
rect 14829 32385 14841 32419
rect 14875 32416 14887 32419
rect 14875 32388 14909 32416
rect 14875 32385 14887 32388
rect 14829 32379 14887 32385
rect 15010 32376 15016 32428
rect 15068 32416 15074 32428
rect 15580 32425 15608 32456
rect 15105 32419 15163 32425
rect 15105 32416 15117 32419
rect 15068 32388 15117 32416
rect 15068 32376 15074 32388
rect 15105 32385 15117 32388
rect 15151 32385 15163 32419
rect 15565 32419 15623 32425
rect 15105 32379 15163 32385
rect 15304 32388 15516 32416
rect 9122 32308 9128 32360
rect 9180 32308 9186 32360
rect 9217 32351 9275 32357
rect 9217 32317 9229 32351
rect 9263 32317 9275 32351
rect 9217 32311 9275 32317
rect 9309 32351 9367 32357
rect 9309 32317 9321 32351
rect 9355 32348 9367 32351
rect 9674 32348 9680 32360
rect 9355 32320 9680 32348
rect 9355 32317 9367 32320
rect 9309 32311 9367 32317
rect 9232 32280 9260 32311
rect 9674 32308 9680 32320
rect 9732 32308 9738 32360
rect 12710 32308 12716 32360
rect 12768 32308 12774 32360
rect 15304 32357 15332 32388
rect 15289 32351 15347 32357
rect 15289 32348 15301 32351
rect 13924 32320 15301 32348
rect 9140 32252 9260 32280
rect 9140 32224 9168 32252
rect 8205 32215 8263 32221
rect 8205 32181 8217 32215
rect 8251 32181 8263 32215
rect 8205 32175 8263 32181
rect 9122 32172 9128 32224
rect 9180 32172 9186 32224
rect 13924 32212 13952 32320
rect 15289 32317 15301 32320
rect 15335 32317 15347 32351
rect 15289 32311 15347 32317
rect 15381 32351 15439 32357
rect 15381 32317 15393 32351
rect 15427 32317 15439 32351
rect 15488 32348 15516 32388
rect 15565 32385 15577 32419
rect 15611 32385 15623 32419
rect 15565 32379 15623 32385
rect 15657 32419 15715 32425
rect 15657 32385 15669 32419
rect 15703 32416 15715 32419
rect 16684 32416 16712 32512
rect 17604 32484 17632 32512
rect 19444 32493 19472 32524
rect 19610 32512 19616 32524
rect 19668 32512 19674 32564
rect 24213 32555 24271 32561
rect 24213 32552 24225 32555
rect 23584 32524 24225 32552
rect 17512 32456 17632 32484
rect 19429 32487 19487 32493
rect 17512 32425 17540 32456
rect 19429 32453 19441 32487
rect 19475 32453 19487 32487
rect 19429 32447 19487 32453
rect 20364 32456 21680 32484
rect 20364 32428 20392 32456
rect 17221 32419 17279 32425
rect 17221 32416 17233 32419
rect 15703 32388 16712 32416
rect 16776 32388 17233 32416
rect 15703 32385 15715 32388
rect 15657 32379 15715 32385
rect 16776 32348 16804 32388
rect 17221 32385 17233 32388
rect 17267 32385 17279 32419
rect 17221 32379 17279 32385
rect 17497 32419 17555 32425
rect 17497 32385 17509 32419
rect 17543 32385 17555 32419
rect 17497 32379 17555 32385
rect 17586 32376 17592 32428
rect 17644 32376 17650 32428
rect 17770 32376 17776 32428
rect 17828 32376 17834 32428
rect 20346 32376 20352 32428
rect 20404 32376 20410 32428
rect 20530 32376 20536 32428
rect 20588 32416 20594 32428
rect 20714 32416 20720 32428
rect 20588 32388 20720 32416
rect 20588 32376 20594 32388
rect 20714 32376 20720 32388
rect 20772 32376 20778 32428
rect 21652 32425 21680 32456
rect 23584 32425 23612 32524
rect 24213 32521 24225 32524
rect 24259 32552 24271 32555
rect 25038 32552 25044 32564
rect 24259 32524 25044 32552
rect 24259 32521 24271 32524
rect 24213 32515 24271 32521
rect 25038 32512 25044 32524
rect 25096 32512 25102 32564
rect 26697 32555 26755 32561
rect 26697 32521 26709 32555
rect 26743 32552 26755 32555
rect 26743 32524 28488 32552
rect 26743 32521 26755 32524
rect 26697 32515 26755 32521
rect 23842 32444 23848 32496
rect 23900 32484 23906 32496
rect 24302 32484 24308 32496
rect 23900 32456 24308 32484
rect 23900 32444 23906 32456
rect 24302 32444 24308 32456
rect 24360 32444 24366 32496
rect 26970 32444 26976 32496
rect 27028 32444 27034 32496
rect 27154 32444 27160 32496
rect 27212 32484 27218 32496
rect 28460 32493 28488 32524
rect 28736 32524 30604 32552
rect 28445 32487 28503 32493
rect 27212 32456 27278 32484
rect 27212 32444 27218 32456
rect 28445 32453 28457 32487
rect 28491 32453 28503 32487
rect 28445 32447 28503 32453
rect 28534 32444 28540 32496
rect 28592 32484 28598 32496
rect 28736 32484 28764 32524
rect 28592 32456 28764 32484
rect 28592 32444 28598 32456
rect 20901 32419 20959 32425
rect 20901 32385 20913 32419
rect 20947 32416 20959 32419
rect 21269 32419 21327 32425
rect 21269 32416 21281 32419
rect 20947 32388 21281 32416
rect 20947 32385 20959 32388
rect 20901 32379 20959 32385
rect 21269 32385 21281 32388
rect 21315 32385 21327 32419
rect 21269 32379 21327 32385
rect 21453 32419 21511 32425
rect 21453 32385 21465 32419
rect 21499 32385 21511 32419
rect 21453 32379 21511 32385
rect 21637 32419 21695 32425
rect 21637 32385 21649 32419
rect 21683 32385 21695 32419
rect 21637 32379 21695 32385
rect 23569 32419 23627 32425
rect 23569 32385 23581 32419
rect 23615 32385 23627 32419
rect 23569 32379 23627 32385
rect 15488 32320 16804 32348
rect 15381 32311 15439 32317
rect 13998 32240 14004 32292
rect 14056 32280 14062 32292
rect 14056 32252 14504 32280
rect 14056 32240 14062 32252
rect 14182 32212 14188 32224
rect 13924 32184 14188 32212
rect 14182 32172 14188 32184
rect 14240 32172 14246 32224
rect 14274 32172 14280 32224
rect 14332 32172 14338 32224
rect 14476 32221 14504 32252
rect 14461 32215 14519 32221
rect 14461 32181 14473 32215
rect 14507 32212 14519 32215
rect 15396 32212 15424 32311
rect 17402 32308 17408 32360
rect 17460 32308 17466 32360
rect 20441 32351 20499 32357
rect 20441 32317 20453 32351
rect 20487 32348 20499 32351
rect 20809 32351 20867 32357
rect 20809 32348 20821 32351
rect 20487 32320 20821 32348
rect 20487 32317 20499 32320
rect 20441 32311 20499 32317
rect 20809 32317 20821 32320
rect 20855 32317 20867 32351
rect 20809 32311 20867 32317
rect 20990 32308 20996 32360
rect 21048 32308 21054 32360
rect 21082 32308 21088 32360
rect 21140 32308 21146 32360
rect 17586 32240 17592 32292
rect 17644 32280 17650 32292
rect 19978 32280 19984 32292
rect 17644 32252 19984 32280
rect 17644 32240 17650 32252
rect 19978 32240 19984 32252
rect 20036 32240 20042 32292
rect 20714 32240 20720 32292
rect 20772 32280 20778 32292
rect 21468 32280 21496 32379
rect 21652 32348 21680 32379
rect 23750 32376 23756 32428
rect 23808 32376 23814 32428
rect 23937 32419 23995 32425
rect 23937 32385 23949 32419
rect 23983 32416 23995 32419
rect 24394 32416 24400 32428
rect 23983 32388 24400 32416
rect 23983 32385 23995 32388
rect 23937 32379 23995 32385
rect 24394 32376 24400 32388
rect 24452 32376 24458 32428
rect 24578 32376 24584 32428
rect 24636 32376 24642 32428
rect 26510 32376 26516 32428
rect 26568 32376 26574 32428
rect 26786 32376 26792 32428
rect 26844 32376 26850 32428
rect 24596 32348 24624 32376
rect 25130 32348 25136 32360
rect 21652 32320 24440 32348
rect 24596 32320 25136 32348
rect 20772 32252 21496 32280
rect 20772 32240 20778 32252
rect 14507 32184 15424 32212
rect 19337 32215 19395 32221
rect 14507 32181 14519 32184
rect 14461 32175 14519 32181
rect 19337 32181 19349 32215
rect 19383 32212 19395 32215
rect 20162 32212 20168 32224
rect 19383 32184 20168 32212
rect 19383 32181 19395 32184
rect 19337 32175 19395 32181
rect 20162 32172 20168 32184
rect 20220 32172 20226 32224
rect 20622 32172 20628 32224
rect 20680 32172 20686 32224
rect 21468 32212 21496 32252
rect 23934 32212 23940 32224
rect 21468 32184 23940 32212
rect 23934 32172 23940 32184
rect 23992 32172 23998 32224
rect 24118 32172 24124 32224
rect 24176 32172 24182 32224
rect 24412 32212 24440 32320
rect 25130 32308 25136 32320
rect 25188 32308 25194 32360
rect 25682 32308 25688 32360
rect 25740 32308 25746 32360
rect 25961 32351 26019 32357
rect 25961 32317 25973 32351
rect 26007 32348 26019 32351
rect 26804 32348 26832 32376
rect 26007 32320 26832 32348
rect 26988 32348 27016 32444
rect 28736 32425 28764 32456
rect 28810 32444 28816 32496
rect 28868 32484 28874 32496
rect 28868 32456 29118 32484
rect 28868 32444 28874 32456
rect 30576 32425 30604 32524
rect 28721 32419 28779 32425
rect 28721 32385 28733 32419
rect 28767 32385 28779 32419
rect 28721 32379 28779 32385
rect 30561 32419 30619 32425
rect 30561 32385 30573 32419
rect 30607 32416 30619 32419
rect 32398 32416 32404 32428
rect 30607 32388 32404 32416
rect 30607 32385 30619 32388
rect 30561 32379 30619 32385
rect 32398 32376 32404 32388
rect 32456 32376 32462 32428
rect 28813 32351 28871 32357
rect 28813 32348 28825 32351
rect 26988 32320 28825 32348
rect 26007 32317 26019 32320
rect 25961 32311 26019 32317
rect 28813 32317 28825 32320
rect 28859 32317 28871 32351
rect 28813 32311 28871 32317
rect 28902 32308 28908 32360
rect 28960 32348 28966 32360
rect 30285 32351 30343 32357
rect 30285 32348 30297 32351
rect 28960 32320 30297 32348
rect 28960 32308 28966 32320
rect 30285 32317 30297 32320
rect 30331 32317 30343 32351
rect 30285 32311 30343 32317
rect 26970 32212 26976 32224
rect 24412 32184 26976 32212
rect 26970 32172 26976 32184
rect 27028 32172 27034 32224
rect 27154 32172 27160 32224
rect 27212 32212 27218 32224
rect 27982 32212 27988 32224
rect 27212 32184 27988 32212
rect 27212 32172 27218 32184
rect 27982 32172 27988 32184
rect 28040 32212 28046 32224
rect 28810 32212 28816 32224
rect 28040 32184 28816 32212
rect 28040 32172 28046 32184
rect 28810 32172 28816 32184
rect 28868 32172 28874 32224
rect 1104 32122 34684 32144
rect 1104 32070 5147 32122
rect 5199 32070 5211 32122
rect 5263 32070 5275 32122
rect 5327 32070 5339 32122
rect 5391 32070 5403 32122
rect 5455 32070 13541 32122
rect 13593 32070 13605 32122
rect 13657 32070 13669 32122
rect 13721 32070 13733 32122
rect 13785 32070 13797 32122
rect 13849 32070 21935 32122
rect 21987 32070 21999 32122
rect 22051 32070 22063 32122
rect 22115 32070 22127 32122
rect 22179 32070 22191 32122
rect 22243 32070 30329 32122
rect 30381 32070 30393 32122
rect 30445 32070 30457 32122
rect 30509 32070 30521 32122
rect 30573 32070 30585 32122
rect 30637 32070 34684 32122
rect 1104 32048 34684 32070
rect 2130 31968 2136 32020
rect 2188 32008 2194 32020
rect 2317 32011 2375 32017
rect 2317 32008 2329 32011
rect 2188 31980 2329 32008
rect 2188 31968 2194 31980
rect 2317 31977 2329 31980
rect 2363 31977 2375 32011
rect 3694 32008 3700 32020
rect 2317 31971 2375 31977
rect 2746 31980 3700 32008
rect 2501 31807 2559 31813
rect 2501 31773 2513 31807
rect 2547 31804 2559 31807
rect 2746 31804 2774 31980
rect 3694 31968 3700 31980
rect 3752 31968 3758 32020
rect 3881 32011 3939 32017
rect 3881 31977 3893 32011
rect 3927 32008 3939 32011
rect 4246 32008 4252 32020
rect 3927 31980 4252 32008
rect 3927 31977 3939 31980
rect 3881 31971 3939 31977
rect 4246 31968 4252 31980
rect 4304 31968 4310 32020
rect 4525 32011 4583 32017
rect 4525 31977 4537 32011
rect 4571 32008 4583 32011
rect 4571 31980 4844 32008
rect 4571 31977 4583 31980
rect 4525 31971 4583 31977
rect 3602 31832 3608 31884
rect 3660 31872 3666 31884
rect 4249 31875 4307 31881
rect 4249 31872 4261 31875
rect 3660 31844 4261 31872
rect 3660 31832 3666 31844
rect 4249 31841 4261 31844
rect 4295 31872 4307 31875
rect 4540 31872 4568 31971
rect 4709 31943 4767 31949
rect 4709 31909 4721 31943
rect 4755 31909 4767 31943
rect 4709 31903 4767 31909
rect 4295 31844 4568 31872
rect 4295 31841 4307 31844
rect 4249 31835 4307 31841
rect 2547 31776 2774 31804
rect 2547 31773 2559 31776
rect 2501 31767 2559 31773
rect 3970 31764 3976 31816
rect 4028 31804 4034 31816
rect 4065 31807 4123 31813
rect 4065 31804 4077 31807
rect 4028 31776 4077 31804
rect 4028 31764 4034 31776
rect 4065 31773 4077 31776
rect 4111 31804 4123 31807
rect 4724 31804 4752 31903
rect 4816 31872 4844 31980
rect 4890 31968 4896 32020
rect 4948 32008 4954 32020
rect 4985 32011 5043 32017
rect 4985 32008 4997 32011
rect 4948 31980 4997 32008
rect 4948 31968 4954 31980
rect 4985 31977 4997 31980
rect 5031 31977 5043 32011
rect 4985 31971 5043 31977
rect 5813 32011 5871 32017
rect 5813 31977 5825 32011
rect 5859 31977 5871 32011
rect 5813 31971 5871 31977
rect 8113 32011 8171 32017
rect 8113 31977 8125 32011
rect 8159 32008 8171 32011
rect 8202 32008 8208 32020
rect 8159 31980 8208 32008
rect 8159 31977 8171 31980
rect 8113 31971 8171 31977
rect 5828 31940 5856 31971
rect 8202 31968 8208 31980
rect 8260 32008 8266 32020
rect 9493 32011 9551 32017
rect 9493 32008 9505 32011
rect 8260 31980 9505 32008
rect 8260 31968 8266 31980
rect 5092 31912 5856 31940
rect 5997 31943 6055 31949
rect 5092 31872 5120 31912
rect 5997 31909 6009 31943
rect 6043 31940 6055 31943
rect 6270 31940 6276 31952
rect 6043 31912 6276 31940
rect 6043 31909 6055 31912
rect 5997 31903 6055 31909
rect 6270 31900 6276 31912
rect 6328 31900 6334 31952
rect 8481 31943 8539 31949
rect 8481 31940 8493 31943
rect 7944 31912 8493 31940
rect 4816 31844 5120 31872
rect 5353 31875 5411 31881
rect 5353 31841 5365 31875
rect 5399 31872 5411 31875
rect 5399 31844 5580 31872
rect 5399 31841 5411 31844
rect 5353 31835 5411 31841
rect 5368 31804 5396 31835
rect 5552 31816 5580 31844
rect 5810 31832 5816 31884
rect 5868 31872 5874 31884
rect 6089 31875 6147 31881
rect 6089 31872 6101 31875
rect 5868 31844 6101 31872
rect 5868 31832 5874 31844
rect 6089 31841 6101 31844
rect 6135 31872 6147 31875
rect 6135 31844 6500 31872
rect 6135 31841 6147 31844
rect 6089 31835 6147 31841
rect 4111 31776 4292 31804
rect 4724 31776 5396 31804
rect 5445 31807 5503 31813
rect 4111 31773 4123 31776
rect 4065 31767 4123 31773
rect 4264 31668 4292 31776
rect 5445 31773 5457 31807
rect 5491 31773 5503 31807
rect 5445 31767 5503 31773
rect 4341 31739 4399 31745
rect 4341 31705 4353 31739
rect 4387 31736 4399 31739
rect 4430 31736 4436 31748
rect 4387 31708 4436 31736
rect 4387 31705 4399 31708
rect 4341 31699 4399 31705
rect 4430 31696 4436 31708
rect 4488 31736 4494 31748
rect 4488 31708 4936 31736
rect 4488 31696 4494 31708
rect 4541 31671 4599 31677
rect 4541 31668 4553 31671
rect 4264 31640 4553 31668
rect 4541 31637 4553 31640
rect 4587 31637 4599 31671
rect 4541 31631 4599 31637
rect 4798 31628 4804 31680
rect 4856 31628 4862 31680
rect 4908 31668 4936 31708
rect 4982 31696 4988 31748
rect 5040 31696 5046 31748
rect 5460 31668 5488 31767
rect 5534 31764 5540 31816
rect 5592 31804 5598 31816
rect 6273 31807 6331 31813
rect 6273 31804 6285 31807
rect 5592 31776 6285 31804
rect 5592 31764 5598 31776
rect 6273 31773 6285 31776
rect 6319 31773 6331 31807
rect 6273 31767 6331 31773
rect 6362 31764 6368 31816
rect 6420 31764 6426 31816
rect 5626 31696 5632 31748
rect 5684 31736 5690 31748
rect 5813 31739 5871 31745
rect 5813 31736 5825 31739
rect 5684 31708 5825 31736
rect 5684 31696 5690 31708
rect 5813 31705 5825 31708
rect 5859 31705 5871 31739
rect 6472 31736 6500 31844
rect 7944 31813 7972 31912
rect 8481 31909 8493 31912
rect 8527 31909 8539 31943
rect 8481 31903 8539 31909
rect 8205 31875 8263 31881
rect 8205 31841 8217 31875
rect 8251 31872 8263 31875
rect 8570 31872 8576 31884
rect 8251 31844 8576 31872
rect 8251 31841 8263 31844
rect 8205 31835 8263 31841
rect 8570 31832 8576 31844
rect 8628 31832 8634 31884
rect 7929 31807 7987 31813
rect 7929 31773 7941 31807
rect 7975 31773 7987 31807
rect 7929 31767 7987 31773
rect 8294 31764 8300 31816
rect 8352 31764 8358 31816
rect 8772 31813 8800 31980
rect 9493 31977 9505 31980
rect 9539 31977 9551 32011
rect 9493 31971 9551 31977
rect 9214 31900 9220 31952
rect 9272 31900 9278 31952
rect 9508 31940 9536 31971
rect 9858 31968 9864 32020
rect 9916 32008 9922 32020
rect 9953 32011 10011 32017
rect 9953 32008 9965 32011
rect 9916 31980 9965 32008
rect 9916 31968 9922 31980
rect 9953 31977 9965 31980
rect 9999 32008 10011 32011
rect 9999 31980 12434 32008
rect 9999 31977 10011 31980
rect 9953 31971 10011 31977
rect 9585 31943 9643 31949
rect 9585 31940 9597 31943
rect 9508 31912 9597 31940
rect 9585 31909 9597 31912
rect 9631 31909 9643 31943
rect 12406 31940 12434 31980
rect 12710 31968 12716 32020
rect 12768 32008 12774 32020
rect 13081 32011 13139 32017
rect 13081 32008 13093 32011
rect 12768 31980 13093 32008
rect 12768 31968 12774 31980
rect 13081 31977 13093 31980
rect 13127 31977 13139 32011
rect 13081 31971 13139 31977
rect 14090 31968 14096 32020
rect 14148 31968 14154 32020
rect 14274 31968 14280 32020
rect 14332 31968 14338 32020
rect 17402 31968 17408 32020
rect 17460 31968 17466 32020
rect 17770 31968 17776 32020
rect 17828 31968 17834 32020
rect 19518 32008 19524 32020
rect 18432 31980 19524 32008
rect 13998 31940 14004 31952
rect 12406 31912 14004 31940
rect 9585 31903 9643 31909
rect 9232 31872 9260 31900
rect 10229 31875 10287 31881
rect 9232 31844 9352 31872
rect 9324 31813 9352 31844
rect 10229 31841 10241 31875
rect 10275 31841 10287 31875
rect 12342 31872 12348 31884
rect 10229 31835 10287 31841
rect 11992 31844 12348 31872
rect 8757 31807 8815 31813
rect 8757 31773 8769 31807
rect 8803 31773 8815 31807
rect 8757 31767 8815 31773
rect 9125 31807 9183 31813
rect 9125 31773 9137 31807
rect 9171 31773 9183 31807
rect 9324 31807 9387 31813
rect 9324 31776 9341 31807
rect 9125 31767 9183 31773
rect 9329 31773 9341 31776
rect 9375 31773 9387 31807
rect 9674 31804 9680 31816
rect 9329 31767 9387 31773
rect 9416 31776 9680 31804
rect 8312 31736 8340 31764
rect 6472 31708 8340 31736
rect 9140 31736 9168 31767
rect 9416 31736 9444 31776
rect 9674 31764 9680 31776
rect 9732 31804 9738 31816
rect 10244 31804 10272 31835
rect 9732 31776 10272 31804
rect 9732 31764 9738 31776
rect 10594 31764 10600 31816
rect 10652 31764 10658 31816
rect 11992 31813 12020 31844
rect 12342 31832 12348 31844
rect 12400 31832 12406 31884
rect 11977 31807 12035 31813
rect 11977 31773 11989 31807
rect 12023 31773 12035 31807
rect 11977 31767 12035 31773
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31773 12127 31807
rect 12452 31804 12480 31912
rect 13998 31900 14004 31912
rect 14056 31900 14062 31952
rect 14292 31872 14320 31968
rect 17420 31940 17448 31968
rect 18325 31943 18383 31949
rect 18325 31940 18337 31943
rect 17420 31912 18337 31940
rect 13280 31844 14320 31872
rect 14384 31844 17264 31872
rect 13280 31813 13308 31844
rect 12069 31767 12127 31773
rect 12360 31776 12480 31804
rect 13265 31807 13323 31813
rect 9140 31708 9444 31736
rect 5813 31699 5871 31705
rect 11698 31696 11704 31748
rect 11756 31696 11762 31748
rect 4908 31640 5488 31668
rect 5718 31628 5724 31680
rect 5776 31668 5782 31680
rect 5902 31668 5908 31680
rect 5776 31640 5908 31668
rect 5776 31628 5782 31640
rect 5902 31628 5908 31640
rect 5960 31628 5966 31680
rect 6086 31628 6092 31680
rect 6144 31628 6150 31680
rect 7745 31671 7803 31677
rect 7745 31637 7757 31671
rect 7791 31668 7803 31671
rect 8110 31668 8116 31680
rect 7791 31640 8116 31668
rect 7791 31637 7803 31640
rect 7745 31631 7803 31637
rect 8110 31628 8116 31640
rect 8168 31628 8174 31680
rect 8665 31671 8723 31677
rect 8665 31637 8677 31671
rect 8711 31668 8723 31671
rect 9122 31668 9128 31680
rect 8711 31640 9128 31668
rect 8711 31637 8723 31640
rect 8665 31631 8723 31637
rect 9122 31628 9128 31640
rect 9180 31628 9186 31680
rect 9950 31628 9956 31680
rect 10008 31628 10014 31680
rect 10137 31671 10195 31677
rect 10137 31637 10149 31671
rect 10183 31668 10195 31671
rect 10410 31668 10416 31680
rect 10183 31640 10416 31668
rect 10183 31637 10195 31640
rect 10137 31631 10195 31637
rect 10410 31628 10416 31640
rect 10468 31628 10474 31680
rect 12084 31668 12112 31767
rect 12360 31745 12388 31776
rect 13265 31773 13277 31807
rect 13311 31773 13323 31807
rect 13265 31767 13323 31773
rect 14182 31764 14188 31816
rect 14240 31804 14246 31816
rect 14384 31804 14412 31844
rect 14240 31776 14412 31804
rect 14240 31764 14246 31776
rect 12345 31739 12403 31745
rect 12345 31705 12357 31739
rect 12391 31736 12403 31739
rect 14277 31739 14335 31745
rect 12391 31708 12425 31736
rect 12391 31705 12403 31708
rect 12345 31699 12403 31705
rect 14277 31705 14289 31739
rect 14323 31736 14335 31739
rect 14384 31736 14412 31776
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31804 14519 31807
rect 15010 31804 15016 31816
rect 14507 31776 15016 31804
rect 14507 31773 14519 31776
rect 14461 31767 14519 31773
rect 15010 31764 15016 31776
rect 15068 31764 15074 31816
rect 17126 31764 17132 31816
rect 17184 31764 17190 31816
rect 17236 31813 17264 31844
rect 17420 31813 17448 31912
rect 18325 31909 18337 31912
rect 18371 31909 18383 31943
rect 18325 31903 18383 31909
rect 18432 31872 18460 31980
rect 19518 31968 19524 31980
rect 19576 31968 19582 32020
rect 19889 32011 19947 32017
rect 19889 32008 19901 32011
rect 19628 31980 19901 32008
rect 18509 31875 18567 31881
rect 18509 31872 18521 31875
rect 18432 31844 18521 31872
rect 18509 31841 18521 31844
rect 18555 31841 18567 31875
rect 19628 31872 19656 31980
rect 19889 31977 19901 31980
rect 19935 32008 19947 32011
rect 19935 31980 20208 32008
rect 19935 31977 19947 31980
rect 19889 31971 19947 31977
rect 20180 31952 20208 31980
rect 20622 31968 20628 32020
rect 20680 31968 20686 32020
rect 23382 32008 23388 32020
rect 20732 31980 23388 32008
rect 19978 31900 19984 31952
rect 20036 31900 20042 31952
rect 20162 31900 20168 31952
rect 20220 31900 20226 31952
rect 18509 31835 18567 31841
rect 18616 31844 19656 31872
rect 20073 31875 20131 31881
rect 17222 31807 17280 31813
rect 17222 31773 17234 31807
rect 17268 31773 17280 31807
rect 17222 31767 17280 31773
rect 17405 31807 17463 31813
rect 17405 31773 17417 31807
rect 17451 31773 17463 31807
rect 17405 31767 17463 31773
rect 17586 31764 17592 31816
rect 17644 31813 17650 31816
rect 18616 31813 18644 31844
rect 20073 31841 20085 31875
rect 20119 31872 20131 31875
rect 20640 31872 20668 31968
rect 20119 31844 20668 31872
rect 20119 31841 20131 31844
rect 20073 31835 20131 31841
rect 17644 31804 17652 31813
rect 18601 31807 18659 31813
rect 17644 31776 17689 31804
rect 17644 31767 17652 31776
rect 18601 31773 18613 31807
rect 18647 31773 18659 31807
rect 18601 31767 18659 31773
rect 18969 31807 19027 31813
rect 18969 31773 18981 31807
rect 19015 31804 19027 31807
rect 19245 31807 19303 31813
rect 19245 31804 19257 31807
rect 19015 31776 19257 31804
rect 19015 31773 19027 31776
rect 18969 31767 19027 31773
rect 19245 31773 19257 31776
rect 19291 31773 19303 31807
rect 19245 31767 19303 31773
rect 17644 31764 17650 31767
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 19702 31804 19708 31816
rect 19663 31776 19708 31804
rect 19702 31764 19708 31776
rect 19760 31804 19766 31816
rect 19797 31807 19855 31813
rect 19797 31804 19809 31807
rect 19760 31776 19809 31804
rect 19760 31764 19766 31776
rect 19797 31773 19809 31776
rect 19843 31773 19855 31807
rect 20732 31804 20760 31980
rect 23382 31968 23388 31980
rect 23440 32008 23446 32020
rect 23753 32011 23811 32017
rect 23753 32008 23765 32011
rect 23440 31980 23765 32008
rect 23440 31968 23446 31980
rect 23753 31977 23765 31980
rect 23799 31977 23811 32011
rect 23753 31971 23811 31977
rect 25041 32011 25099 32017
rect 25041 31977 25053 32011
rect 25087 32008 25099 32011
rect 25682 32008 25688 32020
rect 25087 31980 25688 32008
rect 25087 31977 25099 31980
rect 25041 31971 25099 31977
rect 25682 31968 25688 31980
rect 25740 31968 25746 32020
rect 26510 31968 26516 32020
rect 26568 32008 26574 32020
rect 26605 32011 26663 32017
rect 26605 32008 26617 32011
rect 26568 31980 26617 32008
rect 26568 31968 26574 31980
rect 26605 31977 26617 31980
rect 26651 31977 26663 32011
rect 26605 31971 26663 31977
rect 28074 31968 28080 32020
rect 28132 32008 28138 32020
rect 28132 31980 28764 32008
rect 28132 31968 28138 31980
rect 24118 31832 24124 31884
rect 24176 31872 24182 31884
rect 24397 31875 24455 31881
rect 24397 31872 24409 31875
rect 24176 31844 24409 31872
rect 24176 31832 24182 31844
rect 24397 31841 24409 31844
rect 24443 31841 24455 31875
rect 24397 31835 24455 31841
rect 26970 31832 26976 31884
rect 27028 31872 27034 31884
rect 27065 31875 27123 31881
rect 27065 31872 27077 31875
rect 27028 31844 27077 31872
rect 27028 31832 27034 31844
rect 27065 31841 27077 31844
rect 27111 31841 27123 31875
rect 27065 31835 27123 31841
rect 27154 31832 27160 31884
rect 27212 31832 27218 31884
rect 27632 31844 28580 31872
rect 19797 31767 19855 31773
rect 20180 31776 20760 31804
rect 14323 31708 14412 31736
rect 14323 31705 14335 31708
rect 14277 31699 14335 31705
rect 17494 31696 17500 31748
rect 17552 31696 17558 31748
rect 18874 31696 18880 31748
rect 18932 31696 18938 31748
rect 19812 31736 19840 31767
rect 20180 31736 20208 31776
rect 21818 31764 21824 31816
rect 21876 31804 21882 31816
rect 22005 31807 22063 31813
rect 22005 31804 22017 31807
rect 21876 31776 22017 31804
rect 21876 31764 21882 31776
rect 22005 31773 22017 31776
rect 22051 31773 22063 31807
rect 27632 31804 27660 31844
rect 27908 31813 27936 31844
rect 22005 31767 22063 31773
rect 25792 31776 27660 31804
rect 27709 31807 27767 31813
rect 19812 31708 20208 31736
rect 20530 31696 20536 31748
rect 20588 31696 20594 31748
rect 22278 31696 22284 31748
rect 22336 31696 22342 31748
rect 23014 31696 23020 31748
rect 23072 31696 23078 31748
rect 12802 31668 12808 31680
rect 12084 31640 12808 31668
rect 12802 31628 12808 31640
rect 12860 31628 12866 31680
rect 19610 31628 19616 31680
rect 19668 31668 19674 31680
rect 20548 31668 20576 31696
rect 19668 31640 20576 31668
rect 19668 31628 19674 31640
rect 23750 31628 23756 31680
rect 23808 31668 23814 31680
rect 24854 31668 24860 31680
rect 23808 31640 24860 31668
rect 23808 31628 23814 31640
rect 24854 31628 24860 31640
rect 24912 31668 24918 31680
rect 25792 31668 25820 31776
rect 27709 31773 27721 31807
rect 27755 31773 27767 31807
rect 27709 31767 27767 31773
rect 27893 31807 27951 31813
rect 27893 31773 27905 31807
rect 27939 31773 27951 31807
rect 27893 31767 27951 31773
rect 24912 31640 25820 31668
rect 24912 31628 24918 31640
rect 26970 31628 26976 31680
rect 27028 31628 27034 31680
rect 27724 31668 27752 31767
rect 28074 31764 28080 31816
rect 28132 31764 28138 31816
rect 28350 31764 28356 31816
rect 28408 31764 28414 31816
rect 28552 31813 28580 31844
rect 28736 31813 28764 31980
rect 28902 31968 28908 32020
rect 28960 31968 28966 32020
rect 28537 31807 28595 31813
rect 28537 31773 28549 31807
rect 28583 31773 28595 31807
rect 28537 31767 28595 31773
rect 28721 31807 28779 31813
rect 28721 31773 28733 31807
rect 28767 31773 28779 31807
rect 28721 31767 28779 31773
rect 27798 31696 27804 31748
rect 27856 31736 27862 31748
rect 27985 31739 28043 31745
rect 27985 31736 27997 31739
rect 27856 31708 27997 31736
rect 27856 31696 27862 31708
rect 27985 31705 27997 31708
rect 28031 31705 28043 31739
rect 28442 31736 28448 31748
rect 27985 31699 28043 31705
rect 28184 31708 28448 31736
rect 28184 31668 28212 31708
rect 28442 31696 28448 31708
rect 28500 31736 28506 31748
rect 28629 31739 28687 31745
rect 28629 31736 28641 31739
rect 28500 31708 28641 31736
rect 28500 31696 28506 31708
rect 28629 31705 28641 31708
rect 28675 31705 28687 31739
rect 28629 31699 28687 31705
rect 27724 31640 28212 31668
rect 28261 31671 28319 31677
rect 28261 31637 28273 31671
rect 28307 31668 28319 31671
rect 28350 31668 28356 31680
rect 28307 31640 28356 31668
rect 28307 31637 28319 31640
rect 28261 31631 28319 31637
rect 28350 31628 28356 31640
rect 28408 31628 28414 31680
rect 1104 31578 34840 31600
rect 1104 31526 9344 31578
rect 9396 31526 9408 31578
rect 9460 31526 9472 31578
rect 9524 31526 9536 31578
rect 9588 31526 9600 31578
rect 9652 31526 17738 31578
rect 17790 31526 17802 31578
rect 17854 31526 17866 31578
rect 17918 31526 17930 31578
rect 17982 31526 17994 31578
rect 18046 31526 26132 31578
rect 26184 31526 26196 31578
rect 26248 31526 26260 31578
rect 26312 31526 26324 31578
rect 26376 31526 26388 31578
rect 26440 31526 34526 31578
rect 34578 31526 34590 31578
rect 34642 31526 34654 31578
rect 34706 31526 34718 31578
rect 34770 31526 34782 31578
rect 34834 31526 34840 31578
rect 1104 31504 34840 31526
rect 4430 31424 4436 31476
rect 4488 31464 4494 31476
rect 4525 31467 4583 31473
rect 4525 31464 4537 31467
rect 4488 31436 4537 31464
rect 4488 31424 4494 31436
rect 4525 31433 4537 31436
rect 4571 31433 4583 31467
rect 4525 31427 4583 31433
rect 5813 31467 5871 31473
rect 5813 31433 5825 31467
rect 5859 31464 5871 31467
rect 6362 31464 6368 31476
rect 5859 31436 6368 31464
rect 5859 31433 5871 31436
rect 5813 31427 5871 31433
rect 6362 31424 6368 31436
rect 6420 31464 6426 31476
rect 6457 31467 6515 31473
rect 6457 31464 6469 31467
rect 6420 31436 6469 31464
rect 6420 31424 6426 31436
rect 6457 31433 6469 31436
rect 6503 31433 6515 31467
rect 6457 31427 6515 31433
rect 8570 31424 8576 31476
rect 8628 31424 8634 31476
rect 9950 31424 9956 31476
rect 10008 31464 10014 31476
rect 10137 31467 10195 31473
rect 10137 31464 10149 31467
rect 10008 31436 10149 31464
rect 10008 31424 10014 31436
rect 10137 31433 10149 31436
rect 10183 31433 10195 31467
rect 10137 31427 10195 31433
rect 10597 31467 10655 31473
rect 10597 31433 10609 31467
rect 10643 31464 10655 31467
rect 11698 31464 11704 31476
rect 10643 31436 11704 31464
rect 10643 31433 10655 31436
rect 10597 31427 10655 31433
rect 11698 31424 11704 31436
rect 11756 31424 11762 31476
rect 17126 31424 17132 31476
rect 17184 31424 17190 31476
rect 19426 31424 19432 31476
rect 19484 31424 19490 31476
rect 20346 31424 20352 31476
rect 20404 31424 20410 31476
rect 22278 31424 22284 31476
rect 22336 31464 22342 31476
rect 22557 31467 22615 31473
rect 22557 31464 22569 31467
rect 22336 31436 22569 31464
rect 22336 31424 22342 31436
rect 22557 31433 22569 31436
rect 22603 31433 22615 31467
rect 22557 31427 22615 31433
rect 22925 31467 22983 31473
rect 22925 31433 22937 31467
rect 22971 31433 22983 31467
rect 22925 31427 22983 31433
rect 4338 31396 4344 31408
rect 4278 31368 4344 31396
rect 4338 31356 4344 31368
rect 4396 31396 4402 31408
rect 5902 31396 5908 31408
rect 4396 31368 5908 31396
rect 4396 31356 4402 31368
rect 5902 31356 5908 31368
rect 5960 31356 5966 31408
rect 5997 31399 6055 31405
rect 5997 31365 6009 31399
rect 6043 31396 6055 31399
rect 6086 31396 6092 31408
rect 6043 31368 6092 31396
rect 6043 31365 6055 31368
rect 5997 31359 6055 31365
rect 6086 31356 6092 31368
rect 6144 31356 6150 31408
rect 9214 31356 9220 31408
rect 9272 31396 9278 31408
rect 9769 31399 9827 31405
rect 9769 31396 9781 31399
rect 9272 31368 9781 31396
rect 9272 31356 9278 31368
rect 9769 31365 9781 31368
rect 9815 31365 9827 31399
rect 9769 31359 9827 31365
rect 15105 31399 15163 31405
rect 15105 31365 15117 31399
rect 15151 31396 15163 31399
rect 15194 31396 15200 31408
rect 15151 31368 15200 31396
rect 15151 31365 15163 31368
rect 15105 31359 15163 31365
rect 15194 31356 15200 31368
rect 15252 31356 15258 31408
rect 17494 31356 17500 31408
rect 17552 31356 17558 31408
rect 19610 31396 19616 31408
rect 19168 31368 19616 31396
rect 2774 31288 2780 31340
rect 2832 31288 2838 31340
rect 5718 31288 5724 31340
rect 5776 31288 5782 31340
rect 6914 31288 6920 31340
rect 6972 31328 6978 31340
rect 7009 31331 7067 31337
rect 7009 31328 7021 31331
rect 6972 31300 7021 31328
rect 6972 31288 6978 31300
rect 7009 31297 7021 31300
rect 7055 31297 7067 31331
rect 7009 31291 7067 31297
rect 8110 31288 8116 31340
rect 8168 31288 8174 31340
rect 9674 31288 9680 31340
rect 9732 31328 9738 31340
rect 9953 31331 10011 31337
rect 9953 31328 9965 31331
rect 9732 31300 9965 31328
rect 9732 31288 9738 31300
rect 9953 31297 9965 31300
rect 9999 31297 10011 31331
rect 9953 31291 10011 31297
rect 10410 31288 10416 31340
rect 10468 31288 10474 31340
rect 14737 31331 14795 31337
rect 14737 31297 14749 31331
rect 14783 31328 14795 31331
rect 14826 31328 14832 31340
rect 14783 31300 14832 31328
rect 14783 31297 14795 31300
rect 14737 31291 14795 31297
rect 14826 31288 14832 31300
rect 14884 31328 14890 31340
rect 15010 31328 15016 31340
rect 14884 31300 15016 31328
rect 14884 31288 14890 31300
rect 15010 31288 15016 31300
rect 15068 31288 15074 31340
rect 15381 31331 15439 31337
rect 15381 31328 15393 31331
rect 15304 31300 15393 31328
rect 3050 31220 3056 31272
rect 3108 31220 3114 31272
rect 8754 31220 8760 31272
rect 8812 31260 8818 31272
rect 9122 31260 9128 31272
rect 8812 31232 9128 31260
rect 8812 31220 8818 31232
rect 9122 31220 9128 31232
rect 9180 31220 9186 31272
rect 15304 31201 15332 31300
rect 15381 31297 15393 31300
rect 15427 31297 15439 31331
rect 15381 31291 15439 31297
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31297 17371 31331
rect 17512 31328 17540 31356
rect 17589 31331 17647 31337
rect 17589 31328 17601 31331
rect 17512 31300 17601 31328
rect 17313 31291 17371 31297
rect 17589 31297 17601 31300
rect 17635 31297 17647 31331
rect 17589 31291 17647 31297
rect 15289 31195 15347 31201
rect 15289 31161 15301 31195
rect 15335 31161 15347 31195
rect 15289 31155 15347 31161
rect 5994 31084 6000 31136
rect 6052 31084 6058 31136
rect 7374 31084 7380 31136
rect 7432 31124 7438 31136
rect 7561 31127 7619 31133
rect 7561 31124 7573 31127
rect 7432 31096 7573 31124
rect 7432 31084 7438 31096
rect 7561 31093 7573 31096
rect 7607 31093 7619 31127
rect 7561 31087 7619 31093
rect 13998 31084 14004 31136
rect 14056 31124 14062 31136
rect 14366 31124 14372 31136
rect 14056 31096 14372 31124
rect 14056 31084 14062 31096
rect 14366 31084 14372 31096
rect 14424 31124 14430 31136
rect 15105 31127 15163 31133
rect 15105 31124 15117 31127
rect 14424 31096 15117 31124
rect 14424 31084 14430 31096
rect 15105 31093 15117 31096
rect 15151 31093 15163 31127
rect 15105 31087 15163 31093
rect 15562 31084 15568 31136
rect 15620 31084 15626 31136
rect 17328 31124 17356 31291
rect 17678 31288 17684 31340
rect 17736 31288 17742 31340
rect 17862 31288 17868 31340
rect 17920 31288 17926 31340
rect 19168 31337 19196 31368
rect 19610 31356 19616 31368
rect 19668 31356 19674 31408
rect 20364 31396 20392 31424
rect 20180 31368 20392 31396
rect 19153 31331 19211 31337
rect 19153 31297 19165 31331
rect 19199 31297 19211 31331
rect 19153 31291 19211 31297
rect 19245 31331 19303 31337
rect 19245 31297 19257 31331
rect 19291 31328 19303 31331
rect 19702 31328 19708 31340
rect 19291 31300 19708 31328
rect 19291 31297 19303 31300
rect 19245 31291 19303 31297
rect 19702 31288 19708 31300
rect 19760 31288 19766 31340
rect 20180 31337 20208 31368
rect 20990 31356 20996 31408
rect 21048 31356 21054 31408
rect 21082 31356 21088 31408
rect 21140 31396 21146 31408
rect 21140 31368 21312 31396
rect 21140 31356 21146 31368
rect 20165 31331 20223 31337
rect 20165 31297 20177 31331
rect 20211 31297 20223 31331
rect 21008 31328 21036 31356
rect 21284 31337 21312 31368
rect 21177 31331 21235 31337
rect 21177 31328 21189 31331
rect 20165 31291 20223 31297
rect 20364 31300 21189 31328
rect 17497 31263 17555 31269
rect 17497 31229 17509 31263
rect 17543 31229 17555 31263
rect 17497 31223 17555 31229
rect 19429 31263 19487 31269
rect 19429 31229 19441 31263
rect 19475 31260 19487 31263
rect 20364 31260 20392 31300
rect 21177 31297 21189 31300
rect 21223 31297 21235 31331
rect 21177 31291 21235 31297
rect 21269 31331 21327 31337
rect 21269 31297 21281 31331
rect 21315 31297 21327 31331
rect 21269 31291 21327 31297
rect 22741 31331 22799 31337
rect 22741 31297 22753 31331
rect 22787 31328 22799 31331
rect 22940 31328 22968 31427
rect 23382 31424 23388 31476
rect 23440 31424 23446 31476
rect 23842 31424 23848 31476
rect 23900 31424 23906 31476
rect 26970 31424 26976 31476
rect 27028 31464 27034 31476
rect 27709 31467 27767 31473
rect 27709 31464 27721 31467
rect 27028 31436 27721 31464
rect 27028 31424 27034 31436
rect 27709 31433 27721 31436
rect 27755 31433 27767 31467
rect 27709 31427 27767 31433
rect 28442 31424 28448 31476
rect 28500 31424 28506 31476
rect 23293 31399 23351 31405
rect 23293 31365 23305 31399
rect 23339 31396 23351 31399
rect 23860 31396 23888 31424
rect 23339 31368 23888 31396
rect 23339 31365 23351 31368
rect 23293 31359 23351 31365
rect 22787 31300 22968 31328
rect 22787 31297 22799 31300
rect 22741 31291 22799 31297
rect 24946 31288 24952 31340
rect 25004 31288 25010 31340
rect 19475 31232 20392 31260
rect 20441 31263 20499 31269
rect 19475 31229 19487 31232
rect 19429 31223 19487 31229
rect 20441 31229 20453 31263
rect 20487 31260 20499 31263
rect 20809 31263 20867 31269
rect 20809 31260 20821 31263
rect 20487 31232 20821 31260
rect 20487 31229 20499 31232
rect 20441 31223 20499 31229
rect 20809 31229 20821 31232
rect 20855 31229 20867 31263
rect 20809 31223 20867 31229
rect 20993 31263 21051 31269
rect 20993 31229 21005 31263
rect 21039 31229 21051 31263
rect 20993 31223 21051 31229
rect 17512 31192 17540 31223
rect 17678 31192 17684 31204
rect 17512 31164 17684 31192
rect 17678 31152 17684 31164
rect 17736 31192 17742 31204
rect 20349 31195 20407 31201
rect 20349 31192 20361 31195
rect 17736 31164 20361 31192
rect 17736 31152 17742 31164
rect 20349 31161 20361 31164
rect 20395 31161 20407 31195
rect 21008 31192 21036 31223
rect 21082 31220 21088 31272
rect 21140 31220 21146 31272
rect 23382 31220 23388 31272
rect 23440 31260 23446 31272
rect 23477 31263 23535 31269
rect 23477 31260 23489 31263
rect 23440 31232 23489 31260
rect 23440 31220 23446 31232
rect 23477 31229 23489 31232
rect 23523 31229 23535 31263
rect 23477 31223 23535 31229
rect 27614 31220 27620 31272
rect 27672 31220 27678 31272
rect 28353 31263 28411 31269
rect 28353 31229 28365 31263
rect 28399 31260 28411 31263
rect 29089 31263 29147 31269
rect 29089 31260 29101 31263
rect 28399 31232 29101 31260
rect 28399 31229 28411 31232
rect 28353 31223 28411 31229
rect 29089 31229 29101 31232
rect 29135 31260 29147 31263
rect 29730 31260 29736 31272
rect 29135 31232 29736 31260
rect 29135 31229 29147 31232
rect 29089 31223 29147 31229
rect 29730 31220 29736 31232
rect 29788 31220 29794 31272
rect 21358 31192 21364 31204
rect 21008 31164 21364 31192
rect 20349 31155 20407 31161
rect 21358 31152 21364 31164
rect 21416 31152 21422 31204
rect 17770 31124 17776 31136
rect 17328 31096 17776 31124
rect 17770 31084 17776 31096
rect 17828 31084 17834 31136
rect 20162 31084 20168 31136
rect 20220 31124 20226 31136
rect 20257 31127 20315 31133
rect 20257 31124 20269 31127
rect 20220 31096 20269 31124
rect 20220 31084 20226 31096
rect 20257 31093 20269 31096
rect 20303 31093 20315 31127
rect 20257 31087 20315 31093
rect 24762 31084 24768 31136
rect 24820 31084 24826 31136
rect 25866 31084 25872 31136
rect 25924 31124 25930 31136
rect 26973 31127 27031 31133
rect 26973 31124 26985 31127
rect 25924 31096 26985 31124
rect 25924 31084 25930 31096
rect 26973 31093 26985 31096
rect 27019 31093 27031 31127
rect 26973 31087 27031 31093
rect 1104 31034 34684 31056
rect 1104 30982 5147 31034
rect 5199 30982 5211 31034
rect 5263 30982 5275 31034
rect 5327 30982 5339 31034
rect 5391 30982 5403 31034
rect 5455 30982 13541 31034
rect 13593 30982 13605 31034
rect 13657 30982 13669 31034
rect 13721 30982 13733 31034
rect 13785 30982 13797 31034
rect 13849 30982 21935 31034
rect 21987 30982 21999 31034
rect 22051 30982 22063 31034
rect 22115 30982 22127 31034
rect 22179 30982 22191 31034
rect 22243 30982 30329 31034
rect 30381 30982 30393 31034
rect 30445 30982 30457 31034
rect 30509 30982 30521 31034
rect 30573 30982 30585 31034
rect 30637 30982 34684 31034
rect 1104 30960 34684 30982
rect 3050 30880 3056 30932
rect 3108 30920 3114 30932
rect 3237 30923 3295 30929
rect 3237 30920 3249 30923
rect 3108 30892 3249 30920
rect 3108 30880 3114 30892
rect 3237 30889 3249 30892
rect 3283 30889 3295 30923
rect 3237 30883 3295 30889
rect 5432 30923 5490 30929
rect 5432 30889 5444 30923
rect 5478 30920 5490 30923
rect 5994 30920 6000 30932
rect 5478 30892 6000 30920
rect 5478 30889 5490 30892
rect 5432 30883 5490 30889
rect 5994 30880 6000 30892
rect 6052 30880 6058 30932
rect 6914 30880 6920 30932
rect 6972 30880 6978 30932
rect 7272 30923 7330 30929
rect 7272 30889 7284 30923
rect 7318 30920 7330 30923
rect 7374 30920 7380 30932
rect 7318 30892 7380 30920
rect 7318 30889 7330 30892
rect 7272 30883 7330 30889
rect 7374 30880 7380 30892
rect 7432 30880 7438 30932
rect 12332 30923 12390 30929
rect 12332 30889 12344 30923
rect 12378 30920 12390 30923
rect 14093 30923 14151 30929
rect 14093 30920 14105 30923
rect 12378 30892 14105 30920
rect 12378 30889 12390 30892
rect 12332 30883 12390 30889
rect 14093 30889 14105 30892
rect 14139 30889 14151 30923
rect 14093 30883 14151 30889
rect 14826 30880 14832 30932
rect 14884 30880 14890 30932
rect 15013 30923 15071 30929
rect 15013 30889 15025 30923
rect 15059 30920 15071 30923
rect 17313 30923 17371 30929
rect 15059 30892 15148 30920
rect 15059 30889 15071 30892
rect 15013 30883 15071 30889
rect 5169 30787 5227 30793
rect 5169 30784 5181 30787
rect 2792 30756 5181 30784
rect 2792 30728 2820 30756
rect 5169 30753 5181 30756
rect 5215 30784 5227 30787
rect 7009 30787 7067 30793
rect 7009 30784 7021 30787
rect 5215 30756 7021 30784
rect 5215 30753 5227 30756
rect 5169 30747 5227 30753
rect 7009 30753 7021 30756
rect 7055 30784 7067 30787
rect 8938 30784 8944 30796
rect 7055 30756 8944 30784
rect 7055 30753 7067 30756
rect 7009 30747 7067 30753
rect 8938 30744 8944 30756
rect 8996 30744 9002 30796
rect 12069 30787 12127 30793
rect 12069 30753 12081 30787
rect 12115 30784 12127 30787
rect 12342 30784 12348 30796
rect 12115 30756 12348 30784
rect 12115 30753 12127 30756
rect 12069 30747 12127 30753
rect 12342 30744 12348 30756
rect 12400 30744 12406 30796
rect 2774 30676 2780 30728
rect 2832 30676 2838 30728
rect 3421 30719 3479 30725
rect 3421 30685 3433 30719
rect 3467 30716 3479 30719
rect 4798 30716 4804 30728
rect 3467 30688 4804 30716
rect 3467 30685 3479 30688
rect 3421 30679 3479 30685
rect 4798 30676 4804 30688
rect 4856 30676 4862 30728
rect 9769 30719 9827 30725
rect 9769 30685 9781 30719
rect 9815 30716 9827 30719
rect 10318 30716 10324 30728
rect 9815 30688 10324 30716
rect 9815 30685 9827 30688
rect 9769 30679 9827 30685
rect 10318 30676 10324 30688
rect 10376 30676 10382 30728
rect 13906 30716 13912 30728
rect 13478 30702 13912 30716
rect 13464 30688 13912 30702
rect 5902 30608 5908 30660
rect 5960 30608 5966 30660
rect 9217 30651 9275 30657
rect 9217 30648 9229 30651
rect 8510 30620 9229 30648
rect 9217 30617 9229 30620
rect 9263 30617 9275 30651
rect 9217 30611 9275 30617
rect 8754 30540 8760 30592
rect 8812 30540 8818 30592
rect 9232 30580 9260 30611
rect 9766 30580 9772 30592
rect 9232 30552 9772 30580
rect 9766 30540 9772 30552
rect 9824 30540 9830 30592
rect 10594 30540 10600 30592
rect 10652 30580 10658 30592
rect 13464 30580 13492 30688
rect 13906 30676 13912 30688
rect 13964 30676 13970 30728
rect 14274 30676 14280 30728
rect 14332 30676 14338 30728
rect 14550 30676 14556 30728
rect 14608 30718 14614 30728
rect 14737 30719 14795 30725
rect 14608 30690 14688 30718
rect 14608 30676 14614 30690
rect 14660 30648 14688 30690
rect 14737 30685 14749 30719
rect 14783 30716 14795 30719
rect 15120 30716 15148 30892
rect 17313 30889 17325 30923
rect 17359 30920 17371 30923
rect 17862 30920 17868 30932
rect 17359 30892 17868 30920
rect 17359 30889 17371 30892
rect 17313 30883 17371 30889
rect 17862 30880 17868 30892
rect 17920 30880 17926 30932
rect 18874 30880 18880 30932
rect 18932 30920 18938 30932
rect 19337 30923 19395 30929
rect 19337 30920 19349 30923
rect 18932 30892 19349 30920
rect 18932 30880 18938 30892
rect 19337 30889 19349 30892
rect 19383 30889 19395 30923
rect 19337 30883 19395 30889
rect 20901 30923 20959 30929
rect 20901 30889 20913 30923
rect 20947 30920 20959 30923
rect 21082 30920 21088 30932
rect 20947 30892 21088 30920
rect 20947 30889 20959 30892
rect 20901 30883 20959 30889
rect 21082 30880 21088 30892
rect 21140 30880 21146 30932
rect 21358 30880 21364 30932
rect 21416 30920 21422 30932
rect 21453 30923 21511 30929
rect 21453 30920 21465 30923
rect 21416 30892 21465 30920
rect 21416 30880 21422 30892
rect 21453 30889 21465 30892
rect 21499 30889 21511 30923
rect 21453 30883 21511 30889
rect 24660 30923 24718 30929
rect 24660 30889 24672 30923
rect 24706 30920 24718 30923
rect 24762 30920 24768 30932
rect 24706 30892 24768 30920
rect 24706 30889 24718 30892
rect 24660 30883 24718 30889
rect 24762 30880 24768 30892
rect 24820 30880 24826 30932
rect 27614 30880 27620 30932
rect 27672 30920 27678 30932
rect 27985 30923 28043 30929
rect 27985 30920 27997 30923
rect 27672 30892 27997 30920
rect 27672 30880 27678 30892
rect 27985 30889 27997 30892
rect 28031 30889 28043 30923
rect 27985 30883 28043 30889
rect 17034 30812 17040 30864
rect 17092 30852 17098 30864
rect 17494 30852 17500 30864
rect 17092 30824 17500 30852
rect 17092 30812 17098 30824
rect 17494 30812 17500 30824
rect 17552 30812 17558 30864
rect 17678 30812 17684 30864
rect 17736 30812 17742 30864
rect 17770 30812 17776 30864
rect 17828 30812 17834 30864
rect 21174 30852 21180 30864
rect 19444 30824 21180 30852
rect 15286 30744 15292 30796
rect 15344 30744 15350 30796
rect 15562 30744 15568 30796
rect 15620 30744 15626 30796
rect 17586 30744 17592 30796
rect 17644 30744 17650 30796
rect 14783 30688 15148 30716
rect 14783 30685 14795 30688
rect 14737 30679 14795 30685
rect 14981 30651 15039 30657
rect 14981 30648 14993 30651
rect 14660 30620 14993 30648
rect 14981 30617 14993 30620
rect 15027 30617 15039 30651
rect 14981 30611 15039 30617
rect 10652 30552 13492 30580
rect 10652 30540 10658 30552
rect 13814 30540 13820 30592
rect 13872 30580 13878 30592
rect 15120 30580 15148 30688
rect 16666 30676 16672 30728
rect 16724 30676 16730 30728
rect 17492 30719 17550 30725
rect 17492 30685 17504 30719
rect 17538 30716 17550 30719
rect 17604 30716 17632 30744
rect 17696 30725 17724 30812
rect 17788 30725 17816 30812
rect 17538 30688 17632 30716
rect 17681 30719 17739 30725
rect 17538 30685 17550 30688
rect 17492 30679 17550 30685
rect 17681 30685 17693 30719
rect 17727 30685 17739 30719
rect 17681 30679 17739 30685
rect 17788 30719 17867 30725
rect 17788 30685 17821 30719
rect 17855 30685 17867 30719
rect 17788 30679 17867 30685
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30716 18015 30719
rect 18138 30716 18144 30728
rect 18003 30688 18144 30716
rect 18003 30685 18015 30688
rect 17957 30679 18015 30685
rect 15197 30651 15255 30657
rect 15197 30617 15209 30651
rect 15243 30648 15255 30651
rect 15654 30648 15660 30660
rect 15243 30620 15660 30648
rect 15243 30617 15255 30620
rect 15197 30611 15255 30617
rect 15654 30608 15660 30620
rect 15712 30608 15718 30660
rect 17402 30608 17408 30660
rect 17460 30648 17466 30660
rect 17589 30651 17647 30657
rect 17589 30648 17601 30651
rect 17460 30620 17601 30648
rect 17460 30608 17466 30620
rect 17589 30617 17601 30620
rect 17635 30617 17647 30651
rect 17589 30611 17647 30617
rect 15562 30580 15568 30592
rect 13872 30552 15568 30580
rect 13872 30540 13878 30552
rect 15562 30540 15568 30552
rect 15620 30580 15626 30592
rect 17788 30580 17816 30679
rect 18138 30676 18144 30688
rect 18196 30676 18202 30728
rect 19444 30725 19472 30824
rect 21174 30812 21180 30824
rect 21232 30812 21238 30864
rect 20530 30744 20536 30796
rect 20588 30744 20594 30796
rect 21818 30744 21824 30796
rect 21876 30784 21882 30796
rect 24397 30787 24455 30793
rect 24397 30784 24409 30787
rect 21876 30756 24409 30784
rect 21876 30744 21882 30756
rect 24397 30753 24409 30756
rect 24443 30784 24455 30787
rect 26237 30787 26295 30793
rect 26237 30784 26249 30787
rect 24443 30756 26249 30784
rect 24443 30753 24455 30756
rect 24397 30747 24455 30753
rect 26237 30753 26249 30756
rect 26283 30753 26295 30787
rect 28000 30784 28028 30883
rect 28629 30787 28687 30793
rect 28629 30784 28641 30787
rect 28000 30756 28641 30784
rect 26237 30747 26295 30753
rect 28629 30753 28641 30756
rect 28675 30753 28687 30787
rect 28629 30747 28687 30753
rect 19429 30719 19487 30725
rect 19429 30685 19441 30719
rect 19475 30685 19487 30719
rect 20548 30716 20576 30744
rect 21085 30719 21143 30725
rect 21085 30716 21097 30719
rect 20548 30688 21097 30716
rect 19429 30679 19487 30685
rect 21085 30685 21097 30688
rect 21131 30716 21143 30719
rect 21358 30716 21364 30728
rect 21131 30688 21364 30716
rect 21131 30685 21143 30688
rect 21085 30679 21143 30685
rect 21358 30676 21364 30688
rect 21416 30676 21422 30728
rect 21545 30719 21603 30725
rect 21545 30685 21557 30719
rect 21591 30685 21603 30719
rect 21545 30679 21603 30685
rect 21266 30608 21272 30660
rect 21324 30648 21330 30660
rect 21560 30648 21588 30679
rect 21324 30620 22094 30648
rect 21324 30608 21330 30620
rect 15620 30552 17816 30580
rect 22066 30580 22094 30620
rect 25130 30608 25136 30660
rect 25188 30608 25194 30660
rect 26510 30608 26516 30660
rect 26568 30608 26574 30660
rect 27982 30648 27988 30660
rect 27738 30620 27988 30648
rect 27982 30608 27988 30620
rect 28040 30648 28046 30660
rect 28902 30648 28908 30660
rect 28040 30620 28908 30648
rect 28040 30608 28046 30620
rect 28902 30608 28908 30620
rect 28960 30608 28966 30660
rect 25590 30580 25596 30592
rect 22066 30552 25596 30580
rect 15620 30540 15626 30552
rect 25590 30540 25596 30552
rect 25648 30580 25654 30592
rect 26145 30583 26203 30589
rect 26145 30580 26157 30583
rect 25648 30552 26157 30580
rect 25648 30540 25654 30552
rect 26145 30549 26157 30552
rect 26191 30549 26203 30583
rect 26145 30543 26203 30549
rect 27798 30540 27804 30592
rect 27856 30580 27862 30592
rect 28074 30580 28080 30592
rect 27856 30552 28080 30580
rect 27856 30540 27862 30552
rect 28074 30540 28080 30552
rect 28132 30540 28138 30592
rect 1104 30490 34840 30512
rect 1104 30438 9344 30490
rect 9396 30438 9408 30490
rect 9460 30438 9472 30490
rect 9524 30438 9536 30490
rect 9588 30438 9600 30490
rect 9652 30438 17738 30490
rect 17790 30438 17802 30490
rect 17854 30438 17866 30490
rect 17918 30438 17930 30490
rect 17982 30438 17994 30490
rect 18046 30438 26132 30490
rect 26184 30438 26196 30490
rect 26248 30438 26260 30490
rect 26312 30438 26324 30490
rect 26376 30438 26388 30490
rect 26440 30438 34526 30490
rect 34578 30438 34590 30490
rect 34642 30438 34654 30490
rect 34706 30438 34718 30490
rect 34770 30438 34782 30490
rect 34834 30438 34840 30490
rect 1104 30416 34840 30438
rect 14185 30379 14243 30385
rect 14185 30345 14197 30379
rect 14231 30376 14243 30379
rect 14274 30376 14280 30388
rect 14231 30348 14280 30376
rect 14231 30345 14243 30348
rect 14185 30339 14243 30345
rect 14274 30336 14280 30348
rect 14332 30336 14338 30388
rect 15194 30336 15200 30388
rect 15252 30336 15258 30388
rect 15562 30336 15568 30388
rect 15620 30336 15626 30388
rect 15654 30336 15660 30388
rect 15712 30376 15718 30388
rect 17034 30376 17040 30388
rect 15712 30348 17040 30376
rect 15712 30336 15718 30348
rect 17034 30336 17040 30348
rect 17092 30336 17098 30388
rect 21358 30336 21364 30388
rect 21416 30336 21422 30388
rect 24946 30336 24952 30388
rect 25004 30376 25010 30388
rect 25133 30379 25191 30385
rect 25133 30376 25145 30379
rect 25004 30348 25145 30376
rect 25004 30336 25010 30348
rect 25133 30345 25145 30348
rect 25179 30345 25191 30379
rect 25133 30339 25191 30345
rect 25590 30336 25596 30388
rect 25648 30336 25654 30388
rect 25976 30348 26280 30376
rect 6546 30268 6552 30320
rect 6604 30308 6610 30320
rect 6641 30311 6699 30317
rect 6641 30308 6653 30311
rect 6604 30280 6653 30308
rect 6604 30268 6610 30280
rect 6641 30277 6653 30280
rect 6687 30277 6699 30311
rect 6641 30271 6699 30277
rect 8754 30268 8760 30320
rect 8812 30308 8818 30320
rect 9401 30311 9459 30317
rect 9401 30308 9413 30311
rect 8812 30280 9413 30308
rect 8812 30268 8818 30280
rect 9401 30277 9413 30280
rect 9447 30277 9459 30311
rect 9401 30271 9459 30277
rect 9861 30311 9919 30317
rect 9861 30277 9873 30311
rect 9907 30277 9919 30311
rect 9861 30271 9919 30277
rect 8941 30243 8999 30249
rect 8941 30209 8953 30243
rect 8987 30209 8999 30243
rect 8941 30203 8999 30209
rect 6270 30132 6276 30184
rect 6328 30172 6334 30184
rect 6524 30175 6582 30181
rect 6524 30172 6536 30175
rect 6328 30144 6536 30172
rect 6328 30132 6334 30144
rect 6524 30141 6536 30144
rect 6570 30141 6582 30175
rect 6524 30135 6582 30141
rect 6730 30132 6736 30184
rect 6788 30132 6794 30184
rect 7009 30175 7067 30181
rect 7009 30141 7021 30175
rect 7055 30141 7067 30175
rect 7009 30135 7067 30141
rect 7024 30104 7052 30135
rect 8757 30107 8815 30113
rect 8757 30104 8769 30107
rect 7024 30076 8769 30104
rect 8757 30073 8769 30076
rect 8803 30073 8815 30107
rect 8757 30067 8815 30073
rect 6365 30039 6423 30045
rect 6365 30005 6377 30039
rect 6411 30036 6423 30039
rect 6914 30036 6920 30048
rect 6411 30008 6920 30036
rect 6411 30005 6423 30008
rect 6365 29999 6423 30005
rect 6914 29996 6920 30008
rect 6972 29996 6978 30048
rect 8956 30036 8984 30203
rect 9214 30200 9220 30252
rect 9272 30240 9278 30252
rect 9493 30243 9551 30249
rect 9493 30240 9505 30243
rect 9272 30212 9505 30240
rect 9272 30200 9278 30212
rect 9493 30209 9505 30212
rect 9539 30209 9551 30243
rect 9493 30203 9551 30209
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30172 9183 30175
rect 9674 30172 9680 30184
rect 9171 30144 9680 30172
rect 9171 30141 9183 30144
rect 9125 30135 9183 30141
rect 9674 30132 9680 30144
rect 9732 30132 9738 30184
rect 9030 30064 9036 30116
rect 9088 30104 9094 30116
rect 9876 30104 9904 30271
rect 13446 30200 13452 30252
rect 13504 30240 13510 30252
rect 13725 30243 13783 30249
rect 13725 30240 13737 30243
rect 13504 30212 13737 30240
rect 13504 30200 13510 30212
rect 13725 30209 13737 30212
rect 13771 30209 13783 30243
rect 13725 30203 13783 30209
rect 13814 30200 13820 30252
rect 13872 30200 13878 30252
rect 13906 30200 13912 30252
rect 13964 30240 13970 30252
rect 15580 30249 15608 30336
rect 15672 30249 15700 30336
rect 15565 30243 15623 30249
rect 13964 30212 15516 30240
rect 13964 30200 13970 30212
rect 13998 30132 14004 30184
rect 14056 30172 14062 30184
rect 15488 30181 15516 30212
rect 15565 30209 15577 30243
rect 15611 30209 15623 30243
rect 15565 30203 15623 30209
rect 15657 30243 15715 30249
rect 15657 30209 15669 30243
rect 15703 30209 15715 30243
rect 20257 30243 20315 30249
rect 15657 30203 15715 30209
rect 15764 30212 17448 30240
rect 15764 30184 15792 30212
rect 17420 30184 17448 30212
rect 20257 30209 20269 30243
rect 20303 30240 20315 30243
rect 21266 30240 21272 30252
rect 20303 30212 21272 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 21266 30200 21272 30212
rect 21324 30200 21330 30252
rect 21376 30249 21404 30336
rect 23106 30268 23112 30320
rect 23164 30268 23170 30320
rect 24670 30268 24676 30320
rect 24728 30308 24734 30320
rect 25976 30308 26004 30348
rect 24728 30280 26004 30308
rect 24728 30268 24734 30280
rect 26050 30268 26056 30320
rect 26108 30308 26114 30320
rect 26145 30311 26203 30317
rect 26145 30308 26157 30311
rect 26108 30280 26157 30308
rect 26108 30268 26114 30280
rect 26145 30277 26157 30280
rect 26191 30277 26203 30311
rect 26252 30308 26280 30348
rect 26510 30336 26516 30388
rect 26568 30376 26574 30388
rect 26973 30379 27031 30385
rect 26973 30376 26985 30379
rect 26568 30348 26985 30376
rect 26568 30336 26574 30348
rect 26973 30345 26985 30348
rect 27019 30345 27031 30379
rect 28166 30376 28172 30388
rect 26973 30339 27031 30345
rect 27908 30348 28172 30376
rect 27908 30308 27936 30348
rect 28166 30336 28172 30348
rect 28224 30336 28230 30388
rect 29730 30336 29736 30388
rect 29788 30336 29794 30388
rect 28258 30308 28264 30320
rect 26252 30280 27936 30308
rect 28000 30280 28264 30308
rect 26145 30271 26203 30277
rect 21361 30243 21419 30249
rect 21361 30209 21373 30243
rect 21407 30209 21419 30243
rect 21361 30203 21419 30209
rect 21545 30243 21603 30249
rect 21545 30209 21557 30243
rect 21591 30209 21603 30243
rect 21545 30203 21603 30209
rect 24029 30243 24087 30249
rect 24029 30209 24041 30243
rect 24075 30240 24087 30243
rect 24210 30240 24216 30252
rect 24075 30212 24216 30240
rect 24075 30209 24087 30212
rect 24029 30203 24087 30209
rect 15381 30175 15439 30181
rect 15381 30172 15393 30175
rect 14056 30144 15393 30172
rect 14056 30132 14062 30144
rect 15381 30141 15393 30144
rect 15427 30141 15439 30175
rect 15381 30135 15439 30141
rect 15473 30175 15531 30181
rect 15473 30141 15485 30175
rect 15519 30172 15531 30175
rect 15746 30172 15752 30184
rect 15519 30144 15752 30172
rect 15519 30141 15531 30144
rect 15473 30135 15531 30141
rect 9088 30076 9904 30104
rect 15396 30104 15424 30135
rect 15746 30132 15752 30144
rect 15804 30132 15810 30184
rect 16574 30132 16580 30184
rect 16632 30132 16638 30184
rect 17402 30132 17408 30184
rect 17460 30132 17466 30184
rect 19981 30175 20039 30181
rect 19981 30141 19993 30175
rect 20027 30172 20039 30175
rect 20717 30175 20775 30181
rect 20717 30172 20729 30175
rect 20027 30144 20729 30172
rect 20027 30141 20039 30144
rect 19981 30135 20039 30141
rect 20717 30141 20729 30144
rect 20763 30141 20775 30175
rect 20717 30135 20775 30141
rect 20901 30175 20959 30181
rect 20901 30141 20913 30175
rect 20947 30141 20959 30175
rect 20901 30135 20959 30141
rect 16592 30104 16620 30132
rect 15396 30076 16620 30104
rect 20916 30104 20944 30135
rect 20990 30132 20996 30184
rect 21048 30132 21054 30184
rect 21082 30132 21088 30184
rect 21140 30132 21146 30184
rect 21174 30132 21180 30184
rect 21232 30132 21238 30184
rect 21453 30107 21511 30113
rect 21453 30104 21465 30107
rect 20916 30076 21465 30104
rect 9088 30064 9094 30076
rect 21453 30073 21465 30076
rect 21499 30073 21511 30107
rect 21453 30067 21511 30073
rect 9122 30036 9128 30048
rect 8956 30008 9128 30036
rect 9122 29996 9128 30008
rect 9180 29996 9186 30048
rect 9309 30039 9367 30045
rect 9309 30005 9321 30039
rect 9355 30036 9367 30039
rect 9674 30036 9680 30048
rect 9355 30008 9680 30036
rect 9355 30005 9367 30008
rect 9309 29999 9367 30005
rect 9674 29996 9680 30008
rect 9732 29996 9738 30048
rect 9858 29996 9864 30048
rect 9916 29996 9922 30048
rect 10042 29996 10048 30048
rect 10100 29996 10106 30048
rect 17586 29996 17592 30048
rect 17644 30036 17650 30048
rect 20073 30039 20131 30045
rect 20073 30036 20085 30039
rect 17644 30008 20085 30036
rect 17644 29996 17650 30008
rect 20073 30005 20085 30008
rect 20119 30005 20131 30039
rect 20073 29999 20131 30005
rect 20162 29996 20168 30048
rect 20220 29996 20226 30048
rect 21560 30036 21588 30203
rect 24210 30200 24216 30212
rect 24268 30240 24274 30252
rect 24762 30240 24768 30252
rect 24268 30212 24768 30240
rect 24268 30200 24274 30212
rect 24762 30200 24768 30212
rect 24820 30200 24826 30252
rect 25501 30243 25559 30249
rect 25501 30209 25513 30243
rect 25547 30240 25559 30243
rect 25866 30240 25872 30252
rect 25547 30212 25872 30240
rect 25547 30209 25559 30212
rect 25501 30203 25559 30209
rect 25866 30200 25872 30212
rect 25924 30200 25930 30252
rect 25961 30243 26019 30249
rect 25961 30209 25973 30243
rect 26007 30240 26019 30243
rect 26007 30212 26188 30240
rect 26007 30209 26019 30212
rect 25961 30203 26019 30209
rect 21818 30132 21824 30184
rect 21876 30172 21882 30184
rect 22097 30175 22155 30181
rect 22097 30172 22109 30175
rect 21876 30144 22109 30172
rect 21876 30132 21882 30144
rect 22097 30141 22109 30144
rect 22143 30141 22155 30175
rect 22097 30135 22155 30141
rect 22370 30132 22376 30184
rect 22428 30132 22434 30184
rect 23106 30132 23112 30184
rect 23164 30172 23170 30184
rect 24305 30175 24363 30181
rect 24305 30172 24317 30175
rect 23164 30144 24317 30172
rect 23164 30132 23170 30144
rect 24305 30141 24317 30144
rect 24351 30141 24363 30175
rect 24305 30135 24363 30141
rect 25777 30175 25835 30181
rect 25777 30141 25789 30175
rect 25823 30141 25835 30175
rect 25777 30135 25835 30141
rect 25792 30104 25820 30135
rect 25792 30076 25912 30104
rect 25884 30048 25912 30076
rect 23842 30036 23848 30048
rect 21560 30008 23848 30036
rect 23842 29996 23848 30008
rect 23900 29996 23906 30048
rect 25866 29996 25872 30048
rect 25924 29996 25930 30048
rect 26160 30036 26188 30212
rect 26234 30200 26240 30252
rect 26292 30200 26298 30252
rect 26344 30249 26372 30280
rect 28000 30249 28028 30280
rect 28258 30268 28264 30280
rect 28316 30308 28322 30320
rect 28534 30308 28540 30320
rect 28316 30280 28540 30308
rect 28316 30268 28322 30280
rect 28534 30268 28540 30280
rect 28592 30268 28598 30320
rect 26329 30243 26387 30249
rect 26329 30209 26341 30243
rect 26375 30209 26387 30243
rect 26329 30203 26387 30209
rect 27985 30243 28043 30249
rect 27985 30209 27997 30243
rect 28031 30209 28043 30243
rect 27985 30203 28043 30209
rect 29270 30200 29276 30252
rect 29328 30240 29334 30252
rect 29328 30212 29394 30240
rect 29328 30200 29334 30212
rect 27525 30175 27583 30181
rect 27525 30172 27537 30175
rect 26528 30144 27537 30172
rect 26528 30113 26556 30144
rect 27525 30141 27537 30144
rect 27571 30141 27583 30175
rect 27525 30135 27583 30141
rect 28261 30175 28319 30181
rect 28261 30141 28273 30175
rect 28307 30172 28319 30175
rect 28350 30172 28356 30184
rect 28307 30144 28356 30172
rect 28307 30141 28319 30144
rect 28261 30135 28319 30141
rect 28350 30132 28356 30144
rect 28408 30132 28414 30184
rect 26513 30107 26571 30113
rect 26513 30073 26525 30107
rect 26559 30073 26571 30107
rect 26513 30067 26571 30073
rect 28074 30036 28080 30048
rect 26160 30008 28080 30036
rect 28074 29996 28080 30008
rect 28132 29996 28138 30048
rect 1104 29946 34684 29968
rect 1104 29894 5147 29946
rect 5199 29894 5211 29946
rect 5263 29894 5275 29946
rect 5327 29894 5339 29946
rect 5391 29894 5403 29946
rect 5455 29894 13541 29946
rect 13593 29894 13605 29946
rect 13657 29894 13669 29946
rect 13721 29894 13733 29946
rect 13785 29894 13797 29946
rect 13849 29894 21935 29946
rect 21987 29894 21999 29946
rect 22051 29894 22063 29946
rect 22115 29894 22127 29946
rect 22179 29894 22191 29946
rect 22243 29894 30329 29946
rect 30381 29894 30393 29946
rect 30445 29894 30457 29946
rect 30509 29894 30521 29946
rect 30573 29894 30585 29946
rect 30637 29894 34684 29946
rect 1104 29872 34684 29894
rect 8757 29835 8815 29841
rect 8757 29801 8769 29835
rect 8803 29832 8815 29835
rect 9030 29832 9036 29844
rect 8803 29804 9036 29832
rect 8803 29801 8815 29804
rect 8757 29795 8815 29801
rect 9030 29792 9036 29804
rect 9088 29792 9094 29844
rect 9217 29835 9275 29841
rect 9217 29801 9229 29835
rect 9263 29832 9275 29835
rect 9674 29832 9680 29844
rect 9263 29804 9680 29832
rect 9263 29801 9275 29804
rect 9217 29795 9275 29801
rect 9232 29764 9260 29795
rect 9674 29792 9680 29804
rect 9732 29832 9738 29844
rect 13909 29835 13967 29841
rect 9732 29804 10732 29832
rect 9732 29792 9738 29804
rect 8220 29736 8432 29764
rect 2774 29656 2780 29708
rect 2832 29696 2838 29708
rect 3789 29699 3847 29705
rect 3789 29696 3801 29699
rect 2832 29668 3801 29696
rect 2832 29656 2838 29668
rect 3789 29665 3801 29668
rect 3835 29665 3847 29699
rect 3789 29659 3847 29665
rect 4062 29520 4068 29572
rect 4120 29520 4126 29572
rect 4982 29452 4988 29504
rect 5040 29492 5046 29504
rect 5184 29492 5212 29614
rect 5040 29464 5212 29492
rect 5040 29452 5046 29464
rect 5534 29452 5540 29504
rect 5592 29452 5598 29504
rect 7650 29452 7656 29504
rect 7708 29492 7714 29504
rect 8220 29492 8248 29736
rect 8404 29705 8432 29736
rect 8496 29736 9260 29764
rect 8496 29705 8524 29736
rect 9306 29724 9312 29776
rect 9364 29764 9370 29776
rect 9401 29767 9459 29773
rect 9401 29764 9413 29767
rect 9364 29736 9413 29764
rect 9364 29724 9370 29736
rect 9401 29733 9413 29736
rect 9447 29733 9459 29767
rect 9401 29727 9459 29733
rect 9508 29736 9812 29764
rect 8389 29699 8447 29705
rect 8389 29665 8401 29699
rect 8435 29665 8447 29699
rect 8389 29659 8447 29665
rect 8481 29699 8539 29705
rect 8481 29665 8493 29699
rect 8527 29665 8539 29699
rect 8481 29659 8539 29665
rect 8570 29656 8576 29708
rect 8628 29696 8634 29708
rect 9508 29696 9536 29736
rect 8628 29668 9536 29696
rect 8628 29656 8634 29668
rect 9582 29656 9588 29708
rect 9640 29656 9646 29708
rect 9784 29705 9812 29736
rect 9769 29699 9827 29705
rect 9769 29665 9781 29699
rect 9815 29665 9827 29699
rect 9769 29659 9827 29665
rect 9862 29699 9920 29705
rect 9862 29665 9874 29699
rect 9908 29696 9920 29699
rect 9968 29696 9996 29804
rect 10704 29776 10732 29804
rect 13909 29801 13921 29835
rect 13955 29832 13967 29835
rect 14550 29832 14556 29844
rect 13955 29804 14556 29832
rect 13955 29801 13967 29804
rect 13909 29795 13967 29801
rect 14550 29792 14556 29804
rect 14608 29792 14614 29844
rect 18138 29792 18144 29844
rect 18196 29792 18202 29844
rect 20809 29835 20867 29841
rect 20809 29801 20821 29835
rect 20855 29832 20867 29835
rect 20990 29832 20996 29844
rect 20855 29804 20996 29832
rect 20855 29801 20867 29804
rect 20809 29795 20867 29801
rect 20990 29792 20996 29804
rect 21048 29792 21054 29844
rect 22370 29792 22376 29844
rect 22428 29832 22434 29844
rect 22649 29835 22707 29841
rect 22649 29832 22661 29835
rect 22428 29804 22661 29832
rect 22428 29792 22434 29804
rect 22649 29801 22661 29804
rect 22695 29801 22707 29835
rect 23842 29832 23848 29844
rect 22649 29795 22707 29801
rect 23492 29804 23848 29832
rect 10686 29724 10692 29776
rect 10744 29724 10750 29776
rect 23017 29767 23075 29773
rect 23017 29733 23029 29767
rect 23063 29733 23075 29767
rect 23017 29727 23075 29733
rect 9908 29668 9996 29696
rect 10045 29699 10103 29705
rect 9908 29665 9920 29668
rect 9862 29659 9920 29665
rect 10045 29665 10057 29699
rect 10091 29696 10103 29699
rect 11238 29696 11244 29708
rect 10091 29668 11244 29696
rect 10091 29665 10103 29668
rect 10045 29659 10103 29665
rect 11238 29656 11244 29668
rect 11296 29656 11302 29708
rect 11698 29656 11704 29708
rect 11756 29696 11762 29708
rect 11977 29699 12035 29705
rect 11977 29696 11989 29699
rect 11756 29668 11989 29696
rect 11756 29656 11762 29668
rect 11977 29665 11989 29668
rect 12023 29696 12035 29699
rect 12342 29696 12348 29708
rect 12023 29668 12348 29696
rect 12023 29665 12035 29668
rect 11977 29659 12035 29665
rect 12342 29656 12348 29668
rect 12400 29696 12406 29708
rect 14090 29696 14096 29708
rect 12400 29668 14096 29696
rect 12400 29656 12406 29668
rect 14090 29656 14096 29668
rect 14148 29696 14154 29708
rect 14185 29699 14243 29705
rect 14185 29696 14197 29699
rect 14148 29668 14197 29696
rect 14148 29656 14154 29668
rect 14185 29665 14197 29668
rect 14231 29696 14243 29699
rect 15565 29699 15623 29705
rect 15565 29696 15577 29699
rect 14231 29668 15577 29696
rect 14231 29665 14243 29668
rect 14185 29659 14243 29665
rect 15565 29665 15577 29668
rect 15611 29665 15623 29699
rect 19242 29696 19248 29708
rect 15565 29659 15623 29665
rect 17328 29668 18000 29696
rect 8297 29631 8355 29637
rect 8297 29597 8309 29631
rect 8343 29597 8355 29631
rect 9953 29631 10011 29637
rect 9692 29628 9812 29630
rect 9953 29628 9965 29631
rect 8297 29591 8355 29597
rect 9344 29602 9965 29628
rect 9344 29600 9720 29602
rect 9784 29600 9965 29602
rect 8312 29560 8340 29591
rect 9033 29563 9091 29569
rect 9033 29560 9045 29563
rect 8312 29532 9045 29560
rect 9033 29529 9045 29532
rect 9079 29560 9091 29563
rect 9122 29560 9128 29572
rect 9079 29532 9128 29560
rect 9079 29529 9091 29532
rect 9033 29523 9091 29529
rect 9122 29520 9128 29532
rect 9180 29520 9186 29572
rect 9214 29520 9220 29572
rect 9272 29569 9278 29572
rect 9272 29563 9291 29569
rect 9279 29529 9291 29563
rect 9272 29523 9291 29529
rect 9272 29520 9278 29523
rect 9344 29492 9372 29600
rect 9953 29597 9965 29600
rect 9999 29597 10011 29631
rect 9953 29591 10011 29597
rect 10594 29588 10600 29640
rect 10652 29588 10658 29640
rect 12989 29631 13047 29637
rect 12989 29597 13001 29631
rect 13035 29597 13047 29631
rect 12989 29591 13047 29597
rect 13633 29631 13691 29637
rect 13633 29597 13645 29631
rect 13679 29597 13691 29631
rect 13633 29591 13691 29597
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29628 13783 29631
rect 13998 29628 14004 29640
rect 13771 29600 14004 29628
rect 13771 29597 13783 29600
rect 13725 29591 13783 29597
rect 11422 29520 11428 29572
rect 11480 29560 11486 29572
rect 11701 29563 11759 29569
rect 11701 29560 11713 29563
rect 11480 29532 11713 29560
rect 11480 29520 11486 29532
rect 11701 29529 11713 29532
rect 11747 29529 11759 29563
rect 11701 29523 11759 29529
rect 13004 29504 13032 29591
rect 13648 29560 13676 29591
rect 13998 29588 14004 29600
rect 14056 29588 14062 29640
rect 15013 29631 15071 29637
rect 15013 29597 15025 29631
rect 15059 29597 15071 29631
rect 15013 29591 15071 29597
rect 15105 29631 15163 29637
rect 15105 29597 15117 29631
rect 15151 29628 15163 29631
rect 15470 29628 15476 29640
rect 15151 29600 15476 29628
rect 15151 29597 15163 29600
rect 15105 29591 15163 29597
rect 13906 29560 13912 29572
rect 13648 29532 13912 29560
rect 13906 29520 13912 29532
rect 13964 29520 13970 29572
rect 15028 29504 15056 29591
rect 15470 29588 15476 29600
rect 15528 29588 15534 29640
rect 15841 29563 15899 29569
rect 15841 29560 15853 29563
rect 15304 29532 15853 29560
rect 7708 29464 9372 29492
rect 7708 29452 7714 29464
rect 10226 29452 10232 29504
rect 10284 29452 10290 29504
rect 11514 29452 11520 29504
rect 11572 29492 11578 29504
rect 12250 29492 12256 29504
rect 11572 29464 12256 29492
rect 11572 29452 11578 29464
rect 12250 29452 12256 29464
rect 12308 29492 12314 29504
rect 12345 29495 12403 29501
rect 12345 29492 12357 29495
rect 12308 29464 12357 29492
rect 12308 29452 12314 29464
rect 12345 29461 12357 29464
rect 12391 29461 12403 29495
rect 12345 29455 12403 29461
rect 12986 29452 12992 29504
rect 13044 29452 13050 29504
rect 15010 29452 15016 29504
rect 15068 29452 15074 29504
rect 15304 29501 15332 29532
rect 15841 29529 15853 29532
rect 15887 29529 15899 29563
rect 15841 29523 15899 29529
rect 15289 29495 15347 29501
rect 15289 29461 15301 29495
rect 15335 29461 15347 29495
rect 15289 29455 15347 29461
rect 16666 29452 16672 29504
rect 16724 29492 16730 29504
rect 16960 29492 16988 29614
rect 16724 29464 16988 29492
rect 16724 29452 16730 29464
rect 17126 29452 17132 29504
rect 17184 29492 17190 29504
rect 17328 29501 17356 29668
rect 17402 29588 17408 29640
rect 17460 29588 17466 29640
rect 17494 29588 17500 29640
rect 17552 29588 17558 29640
rect 17586 29588 17592 29640
rect 17644 29588 17650 29640
rect 17972 29637 18000 29668
rect 18708 29668 19248 29696
rect 18708 29637 18736 29668
rect 19242 29656 19248 29668
rect 19300 29656 19306 29708
rect 19886 29656 19892 29708
rect 19944 29656 19950 29708
rect 17681 29631 17739 29637
rect 17681 29597 17693 29631
rect 17727 29597 17739 29631
rect 17681 29591 17739 29597
rect 17773 29631 17831 29637
rect 17773 29597 17785 29631
rect 17819 29597 17831 29631
rect 17773 29591 17831 29597
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29597 18015 29631
rect 17957 29591 18015 29597
rect 18693 29631 18751 29637
rect 18693 29597 18705 29631
rect 18739 29597 18751 29631
rect 18693 29591 18751 29597
rect 18877 29631 18935 29637
rect 18877 29597 18889 29631
rect 18923 29628 18935 29631
rect 19334 29628 19340 29640
rect 18923 29600 19340 29628
rect 18923 29597 18935 29600
rect 18877 29591 18935 29597
rect 17512 29560 17540 29588
rect 17696 29560 17724 29591
rect 17512 29532 17724 29560
rect 17788 29560 17816 29591
rect 19334 29588 19340 29600
rect 19392 29588 19398 29640
rect 20070 29588 20076 29640
rect 20128 29588 20134 29640
rect 20165 29631 20223 29637
rect 20165 29597 20177 29631
rect 20211 29628 20223 29631
rect 21177 29631 21235 29637
rect 21177 29628 21189 29631
rect 20211 29600 21189 29628
rect 20211 29597 20223 29600
rect 20165 29591 20223 29597
rect 21177 29597 21189 29600
rect 21223 29628 21235 29631
rect 22833 29631 22891 29637
rect 21223 29600 22094 29628
rect 21223 29597 21235 29600
rect 21177 29591 21235 29597
rect 18138 29560 18144 29572
rect 17788 29532 18144 29560
rect 18138 29520 18144 29532
rect 18196 29560 18202 29572
rect 19889 29563 19947 29569
rect 19889 29560 19901 29563
rect 18196 29532 19901 29560
rect 18196 29520 18202 29532
rect 19889 29529 19901 29532
rect 19935 29529 19947 29563
rect 19889 29523 19947 29529
rect 20806 29520 20812 29572
rect 20864 29560 20870 29572
rect 20993 29563 21051 29569
rect 20993 29560 21005 29563
rect 20864 29532 21005 29560
rect 20864 29520 20870 29532
rect 20993 29529 21005 29532
rect 21039 29560 21051 29563
rect 21358 29560 21364 29572
rect 21039 29532 21364 29560
rect 21039 29529 21051 29532
rect 20993 29523 21051 29529
rect 21358 29520 21364 29532
rect 21416 29520 21422 29572
rect 22066 29560 22094 29600
rect 22833 29597 22845 29631
rect 22879 29628 22891 29631
rect 23032 29628 23060 29727
rect 23492 29705 23520 29804
rect 23842 29792 23848 29804
rect 23900 29792 23906 29844
rect 25866 29832 25872 29844
rect 24596 29804 25872 29832
rect 23477 29699 23535 29705
rect 23477 29665 23489 29699
rect 23523 29665 23535 29699
rect 23477 29659 23535 29665
rect 22879 29600 23060 29628
rect 22879 29597 22891 29600
rect 22833 29591 22891 29597
rect 23492 29560 23520 29659
rect 23566 29656 23572 29708
rect 23624 29696 23630 29708
rect 23661 29699 23719 29705
rect 23661 29696 23673 29699
rect 23624 29668 23673 29696
rect 23624 29656 23630 29668
rect 23661 29665 23673 29668
rect 23707 29696 23719 29699
rect 24596 29696 24624 29804
rect 25866 29792 25872 29804
rect 25924 29832 25930 29844
rect 27338 29832 27344 29844
rect 25924 29804 27344 29832
rect 25924 29792 25930 29804
rect 27338 29792 27344 29804
rect 27396 29792 27402 29844
rect 29365 29767 29423 29773
rect 29365 29733 29377 29767
rect 29411 29764 29423 29767
rect 31110 29764 31116 29776
rect 29411 29736 31116 29764
rect 29411 29733 29423 29736
rect 29365 29727 29423 29733
rect 31110 29724 31116 29736
rect 31168 29724 31174 29776
rect 23707 29668 24624 29696
rect 23707 29665 23719 29668
rect 23661 29659 23719 29665
rect 24854 29656 24860 29708
rect 24912 29696 24918 29708
rect 26050 29696 26056 29708
rect 24912 29668 26056 29696
rect 24912 29656 24918 29668
rect 26050 29656 26056 29668
rect 26108 29656 26114 29708
rect 26329 29699 26387 29705
rect 26329 29665 26341 29699
rect 26375 29696 26387 29699
rect 26786 29696 26792 29708
rect 26375 29668 26792 29696
rect 26375 29665 26387 29668
rect 26329 29659 26387 29665
rect 26786 29656 26792 29668
rect 26844 29656 26850 29708
rect 24486 29588 24492 29640
rect 24544 29628 24550 29640
rect 24872 29628 24900 29656
rect 25038 29628 25044 29640
rect 24544 29600 24900 29628
rect 24978 29600 25044 29628
rect 24544 29588 24550 29600
rect 25038 29588 25044 29600
rect 25096 29588 25102 29640
rect 29181 29631 29239 29637
rect 29181 29597 29193 29631
rect 29227 29597 29239 29631
rect 29181 29591 29239 29597
rect 29365 29631 29423 29637
rect 29365 29597 29377 29631
rect 29411 29597 29423 29631
rect 29365 29591 29423 29597
rect 22066 29532 23520 29560
rect 26050 29520 26056 29572
rect 26108 29520 26114 29572
rect 26510 29520 26516 29572
rect 26568 29520 26574 29572
rect 17313 29495 17371 29501
rect 17313 29492 17325 29495
rect 17184 29464 17325 29492
rect 17184 29452 17190 29464
rect 17313 29461 17325 29464
rect 17359 29461 17371 29495
rect 17313 29455 17371 29461
rect 18598 29452 18604 29504
rect 18656 29492 18662 29504
rect 18785 29495 18843 29501
rect 18785 29492 18797 29495
rect 18656 29464 18797 29492
rect 18656 29452 18662 29464
rect 18785 29461 18797 29464
rect 18831 29461 18843 29495
rect 18785 29455 18843 29461
rect 20346 29452 20352 29504
rect 20404 29492 20410 29504
rect 21174 29492 21180 29504
rect 20404 29464 21180 29492
rect 20404 29452 20410 29464
rect 21174 29452 21180 29464
rect 21232 29452 21238 29504
rect 23385 29495 23443 29501
rect 23385 29461 23397 29495
rect 23431 29492 23443 29495
rect 24581 29495 24639 29501
rect 24581 29492 24593 29495
rect 23431 29464 24593 29492
rect 23431 29461 23443 29464
rect 23385 29455 23443 29461
rect 24581 29461 24593 29464
rect 24627 29492 24639 29495
rect 26528 29492 26556 29520
rect 24627 29464 26556 29492
rect 29196 29492 29224 29591
rect 29380 29560 29408 29591
rect 29454 29588 29460 29640
rect 29512 29628 29518 29640
rect 30101 29631 30159 29637
rect 30101 29628 30113 29631
rect 29512 29600 30113 29628
rect 29512 29588 29518 29600
rect 30101 29597 30113 29600
rect 30147 29597 30159 29631
rect 30101 29591 30159 29597
rect 30834 29588 30840 29640
rect 30892 29588 30898 29640
rect 30285 29563 30343 29569
rect 30285 29560 30297 29563
rect 29380 29532 30297 29560
rect 30285 29529 30297 29532
rect 30331 29529 30343 29563
rect 30285 29523 30343 29529
rect 29362 29492 29368 29504
rect 29196 29464 29368 29492
rect 24627 29461 24639 29464
rect 24581 29455 24639 29461
rect 29362 29452 29368 29464
rect 29420 29452 29426 29504
rect 29546 29452 29552 29504
rect 29604 29452 29610 29504
rect 1104 29402 34840 29424
rect 1104 29350 9344 29402
rect 9396 29350 9408 29402
rect 9460 29350 9472 29402
rect 9524 29350 9536 29402
rect 9588 29350 9600 29402
rect 9652 29350 17738 29402
rect 17790 29350 17802 29402
rect 17854 29350 17866 29402
rect 17918 29350 17930 29402
rect 17982 29350 17994 29402
rect 18046 29350 26132 29402
rect 26184 29350 26196 29402
rect 26248 29350 26260 29402
rect 26312 29350 26324 29402
rect 26376 29350 26388 29402
rect 26440 29350 34526 29402
rect 34578 29350 34590 29402
rect 34642 29350 34654 29402
rect 34706 29350 34718 29402
rect 34770 29350 34782 29402
rect 34834 29350 34840 29402
rect 1104 29328 34840 29350
rect 4062 29248 4068 29300
rect 4120 29248 4126 29300
rect 5997 29291 6055 29297
rect 5997 29257 6009 29291
rect 6043 29288 6055 29291
rect 6730 29288 6736 29300
rect 6043 29260 6736 29288
rect 6043 29257 6055 29260
rect 5997 29251 6055 29257
rect 6730 29248 6736 29260
rect 6788 29248 6794 29300
rect 15010 29288 15016 29300
rect 8588 29260 15016 29288
rect 4525 29223 4583 29229
rect 4525 29220 4537 29223
rect 3436 29192 4537 29220
rect 3234 29112 3240 29164
rect 3292 29112 3298 29164
rect 3436 29161 3464 29192
rect 4525 29189 4537 29192
rect 4571 29189 4583 29223
rect 7561 29223 7619 29229
rect 7561 29220 7573 29223
rect 4525 29183 4583 29189
rect 7024 29192 7573 29220
rect 7024 29164 7052 29192
rect 7561 29189 7573 29192
rect 7607 29220 7619 29223
rect 7650 29220 7656 29232
rect 7607 29192 7656 29220
rect 7607 29189 7619 29192
rect 7561 29183 7619 29189
rect 7650 29180 7656 29192
rect 7708 29180 7714 29232
rect 7745 29223 7803 29229
rect 7745 29189 7757 29223
rect 7791 29220 7803 29223
rect 8478 29220 8484 29232
rect 7791 29192 8484 29220
rect 7791 29189 7803 29192
rect 7745 29183 7803 29189
rect 3421 29155 3479 29161
rect 3421 29121 3433 29155
rect 3467 29121 3479 29155
rect 3421 29115 3479 29121
rect 3605 29155 3663 29161
rect 3605 29121 3617 29155
rect 3651 29121 3663 29155
rect 3605 29115 3663 29121
rect 3252 29084 3280 29112
rect 3620 29084 3648 29115
rect 3878 29112 3884 29164
rect 3936 29112 3942 29164
rect 4430 29112 4436 29164
rect 4488 29152 4494 29164
rect 5169 29155 5227 29161
rect 5169 29152 5181 29155
rect 4488 29124 5181 29152
rect 4488 29112 4494 29124
rect 5169 29121 5181 29124
rect 5215 29152 5227 29155
rect 5353 29155 5411 29161
rect 5353 29152 5365 29155
rect 5215 29124 5365 29152
rect 5215 29121 5227 29124
rect 5169 29115 5227 29121
rect 5353 29121 5365 29124
rect 5399 29152 5411 29155
rect 5534 29152 5540 29164
rect 5399 29124 5540 29152
rect 5399 29121 5411 29124
rect 5353 29115 5411 29121
rect 5534 29112 5540 29124
rect 5592 29112 5598 29164
rect 5721 29155 5779 29161
rect 5721 29121 5733 29155
rect 5767 29152 5779 29155
rect 7006 29152 7012 29164
rect 5767 29124 7012 29152
rect 5767 29121 5779 29124
rect 5721 29115 5779 29121
rect 7006 29112 7012 29124
rect 7064 29112 7070 29164
rect 7101 29155 7159 29161
rect 7101 29121 7113 29155
rect 7147 29152 7159 29155
rect 7760 29152 7788 29183
rect 8478 29180 8484 29192
rect 8536 29180 8542 29232
rect 7147 29124 7788 29152
rect 7837 29155 7895 29161
rect 7147 29121 7159 29124
rect 7101 29115 7159 29121
rect 7837 29121 7849 29155
rect 7883 29152 7895 29155
rect 8588 29152 8616 29260
rect 15010 29248 15016 29260
rect 15068 29288 15074 29300
rect 15068 29260 15424 29288
rect 15068 29248 15074 29260
rect 8665 29223 8723 29229
rect 8665 29189 8677 29223
rect 8711 29220 8723 29223
rect 8938 29220 8944 29232
rect 8711 29192 8944 29220
rect 8711 29189 8723 29192
rect 8665 29183 8723 29189
rect 8938 29180 8944 29192
rect 8996 29180 9002 29232
rect 9674 29220 9680 29232
rect 9048 29192 9680 29220
rect 8846 29152 8852 29164
rect 7883 29124 8852 29152
rect 7883 29121 7895 29124
rect 7837 29115 7895 29121
rect 3252 29056 3648 29084
rect 5626 29044 5632 29096
rect 5684 29044 5690 29096
rect 5838 29087 5896 29093
rect 5838 29053 5850 29087
rect 5884 29084 5896 29087
rect 5994 29084 6000 29096
rect 5884 29056 6000 29084
rect 5884 29053 5896 29056
rect 5838 29047 5896 29053
rect 5994 29044 6000 29056
rect 6052 29044 6058 29096
rect 4890 28976 4896 29028
rect 4948 29016 4954 29028
rect 7116 29016 7144 29115
rect 8846 29112 8852 29124
rect 8904 29112 8910 29164
rect 9048 29161 9076 29192
rect 9674 29180 9680 29192
rect 9732 29180 9738 29232
rect 10042 29180 10048 29232
rect 10100 29180 10106 29232
rect 11422 29220 11428 29232
rect 10796 29192 11428 29220
rect 9033 29155 9091 29161
rect 9033 29121 9045 29155
rect 9079 29121 9091 29155
rect 9033 29115 9091 29121
rect 9214 29112 9220 29164
rect 9272 29152 9278 29164
rect 9309 29155 9367 29161
rect 9309 29152 9321 29155
rect 9272 29124 9321 29152
rect 9272 29112 9278 29124
rect 9309 29121 9321 29124
rect 9355 29121 9367 29155
rect 9309 29115 9367 29121
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29152 9551 29155
rect 9861 29155 9919 29161
rect 9861 29152 9873 29155
rect 9539 29124 9873 29152
rect 9539 29121 9551 29124
rect 9493 29115 9551 29121
rect 9861 29121 9873 29124
rect 9907 29121 9919 29155
rect 10060 29152 10088 29180
rect 10597 29155 10655 29161
rect 10597 29152 10609 29155
rect 10060 29124 10609 29152
rect 9861 29115 9919 29121
rect 10597 29121 10609 29124
rect 10643 29121 10655 29155
rect 10597 29115 10655 29121
rect 9324 29084 9352 29115
rect 4948 28988 7144 29016
rect 7300 29056 9352 29084
rect 10505 29087 10563 29093
rect 4948 28976 4954 28988
rect 4154 28908 4160 28960
rect 4212 28948 4218 28960
rect 5718 28948 5724 28960
rect 4212 28920 5724 28948
rect 4212 28908 4218 28920
rect 5718 28908 5724 28920
rect 5776 28908 5782 28960
rect 7190 28908 7196 28960
rect 7248 28948 7254 28960
rect 7300 28957 7328 29056
rect 10505 29053 10517 29087
rect 10551 29084 10563 29087
rect 10686 29084 10692 29096
rect 10551 29056 10692 29084
rect 10551 29053 10563 29056
rect 10505 29047 10563 29053
rect 10686 29044 10692 29056
rect 10744 29044 10750 29096
rect 10796 29025 10824 29192
rect 11422 29180 11428 29192
rect 11480 29180 11486 29232
rect 11698 29220 11704 29232
rect 11532 29192 11704 29220
rect 11149 29155 11207 29161
rect 11149 29121 11161 29155
rect 11195 29152 11207 29155
rect 11238 29152 11244 29164
rect 11195 29124 11244 29152
rect 11195 29121 11207 29124
rect 11149 29115 11207 29121
rect 11238 29112 11244 29124
rect 11296 29112 11302 29164
rect 11532 29161 11560 29192
rect 11698 29180 11704 29192
rect 11756 29180 11762 29232
rect 13814 29180 13820 29232
rect 13872 29180 13878 29232
rect 15396 29229 15424 29260
rect 15470 29248 15476 29300
rect 15528 29248 15534 29300
rect 17402 29248 17408 29300
rect 17460 29288 17466 29300
rect 17497 29291 17555 29297
rect 17497 29288 17509 29291
rect 17460 29260 17509 29288
rect 17460 29248 17466 29260
rect 17497 29257 17509 29260
rect 17543 29257 17555 29291
rect 17497 29251 17555 29257
rect 18138 29248 18144 29300
rect 18196 29248 18202 29300
rect 19886 29248 19892 29300
rect 19944 29288 19950 29300
rect 20441 29291 20499 29297
rect 20441 29288 20453 29291
rect 19944 29260 20453 29288
rect 19944 29248 19950 29260
rect 20441 29257 20453 29260
rect 20487 29257 20499 29291
rect 20441 29251 20499 29257
rect 25593 29291 25651 29297
rect 25593 29257 25605 29291
rect 25639 29288 25651 29291
rect 26050 29288 26056 29300
rect 25639 29260 26056 29288
rect 25639 29257 25651 29260
rect 25593 29251 25651 29257
rect 26050 29248 26056 29260
rect 26108 29248 26114 29300
rect 26510 29248 26516 29300
rect 26568 29248 26574 29300
rect 28258 29248 28264 29300
rect 28316 29288 28322 29300
rect 28316 29260 31432 29288
rect 28316 29248 28322 29260
rect 14093 29223 14151 29229
rect 14093 29189 14105 29223
rect 14139 29189 14151 29223
rect 14093 29183 14151 29189
rect 15381 29223 15439 29229
rect 15381 29189 15393 29223
rect 15427 29189 15439 29223
rect 15381 29183 15439 29189
rect 15657 29223 15715 29229
rect 15657 29189 15669 29223
rect 15703 29189 15715 29223
rect 17773 29223 17831 29229
rect 17773 29220 17785 29223
rect 15657 29183 15715 29189
rect 17512 29192 17785 29220
rect 13818 29177 13876 29180
rect 11333 29155 11391 29161
rect 11333 29121 11345 29155
rect 11379 29121 11391 29155
rect 11333 29115 11391 29121
rect 11517 29155 11575 29161
rect 11517 29121 11529 29155
rect 11563 29121 11575 29155
rect 11517 29115 11575 29121
rect 10781 29019 10839 29025
rect 10781 28985 10793 29019
rect 10827 28985 10839 29019
rect 11348 29016 11376 29115
rect 12894 29112 12900 29164
rect 12952 29112 12958 29164
rect 13818 29143 13830 29177
rect 13864 29143 13876 29177
rect 13818 29137 13876 29143
rect 13998 29112 14004 29164
rect 14056 29112 14062 29164
rect 14108 29152 14136 29183
rect 14185 29155 14243 29161
rect 14185 29152 14197 29155
rect 14108 29124 14197 29152
rect 14185 29121 14197 29124
rect 14231 29121 14243 29155
rect 14185 29115 14243 29121
rect 14369 29155 14427 29161
rect 14369 29121 14381 29155
rect 14415 29152 14427 29155
rect 14415 29124 14596 29152
rect 14415 29121 14427 29124
rect 14369 29115 14427 29121
rect 11793 29087 11851 29093
rect 11793 29084 11805 29087
rect 11624 29056 11805 29084
rect 11514 29016 11520 29028
rect 11348 28988 11520 29016
rect 10781 28979 10839 28985
rect 11514 28976 11520 28988
rect 11572 28976 11578 29028
rect 7285 28951 7343 28957
rect 7285 28948 7297 28951
rect 7248 28920 7297 28948
rect 7248 28908 7254 28920
rect 7285 28917 7297 28920
rect 7331 28917 7343 28951
rect 7285 28911 7343 28917
rect 7374 28908 7380 28960
rect 7432 28908 7438 28960
rect 8849 28951 8907 28957
rect 8849 28917 8861 28951
rect 8895 28948 8907 28951
rect 9122 28948 9128 28960
rect 8895 28920 9128 28948
rect 8895 28917 8907 28920
rect 8849 28911 8907 28917
rect 9122 28908 9128 28920
rect 9180 28908 9186 28960
rect 11333 28951 11391 28957
rect 11333 28917 11345 28951
rect 11379 28948 11391 28951
rect 11624 28948 11652 29056
rect 11793 29053 11805 29056
rect 11839 29053 11851 29087
rect 11793 29047 11851 29053
rect 12342 29044 12348 29096
rect 12400 29084 12406 29096
rect 12986 29084 12992 29096
rect 12400 29056 12992 29084
rect 12400 29044 12406 29056
rect 12986 29044 12992 29056
rect 13044 29084 13050 29096
rect 13265 29087 13323 29093
rect 13265 29084 13277 29087
rect 13044 29056 13277 29084
rect 13044 29044 13050 29056
rect 13265 29053 13277 29056
rect 13311 29053 13323 29087
rect 13265 29047 13323 29053
rect 11379 28920 11652 28948
rect 13909 28951 13967 28957
rect 11379 28917 11391 28920
rect 11333 28911 11391 28917
rect 13909 28917 13921 28951
rect 13955 28948 13967 28951
rect 14016 28948 14044 29112
rect 14568 29096 14596 29124
rect 14093 29087 14151 29093
rect 14093 29053 14105 29087
rect 14139 29084 14151 29087
rect 14139 29056 14320 29084
rect 14139 29053 14151 29056
rect 14093 29047 14151 29053
rect 14292 29016 14320 29056
rect 14550 29044 14556 29096
rect 14608 29044 14614 29096
rect 14642 29044 14648 29096
rect 14700 29044 14706 29096
rect 14366 29016 14372 29028
rect 14292 28988 14372 29016
rect 14366 28976 14372 28988
rect 14424 29016 14430 29028
rect 15672 29016 15700 29183
rect 16853 29155 16911 29161
rect 16853 29121 16865 29155
rect 16899 29121 16911 29155
rect 16853 29115 16911 29121
rect 16868 29084 16896 29115
rect 16942 29112 16948 29164
rect 17000 29152 17006 29164
rect 17037 29155 17095 29161
rect 17037 29152 17049 29155
rect 17000 29124 17049 29152
rect 17000 29112 17006 29124
rect 17037 29121 17049 29124
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 17129 29155 17187 29161
rect 17129 29121 17141 29155
rect 17175 29152 17187 29155
rect 17512 29152 17540 29192
rect 17773 29189 17785 29192
rect 17819 29189 17831 29223
rect 17773 29183 17831 29189
rect 17865 29223 17923 29229
rect 17865 29189 17877 29223
rect 17911 29220 17923 29223
rect 18156 29220 18184 29248
rect 17911 29192 18184 29220
rect 18877 29223 18935 29229
rect 17911 29189 17923 29192
rect 17865 29183 17923 29189
rect 18877 29189 18889 29223
rect 18923 29189 18935 29223
rect 18877 29183 18935 29189
rect 17175 29124 17540 29152
rect 17175 29121 17187 29124
rect 17129 29115 17187 29121
rect 17512 29096 17540 29124
rect 17676 29155 17734 29161
rect 17676 29121 17688 29155
rect 17722 29152 17734 29155
rect 18048 29155 18106 29161
rect 17722 29124 17816 29152
rect 17722 29121 17734 29124
rect 17676 29115 17734 29121
rect 17788 29096 17816 29124
rect 18048 29121 18060 29155
rect 18094 29121 18106 29155
rect 18048 29115 18106 29121
rect 18141 29155 18199 29161
rect 18141 29121 18153 29155
rect 18187 29152 18199 29155
rect 18233 29155 18291 29161
rect 18233 29152 18245 29155
rect 18187 29124 18245 29152
rect 18187 29121 18199 29124
rect 18141 29115 18199 29121
rect 18233 29121 18245 29124
rect 18279 29121 18291 29155
rect 18233 29115 18291 29121
rect 18417 29155 18475 29161
rect 18417 29121 18429 29155
rect 18463 29152 18475 29155
rect 18506 29152 18512 29164
rect 18463 29124 18512 29152
rect 18463 29121 18475 29124
rect 18417 29115 18475 29121
rect 16868 29056 17080 29084
rect 17052 29028 17080 29056
rect 17494 29044 17500 29096
rect 17552 29044 17558 29096
rect 17770 29044 17776 29096
rect 17828 29044 17834 29096
rect 14424 28988 15700 29016
rect 16025 29019 16083 29025
rect 14424 28976 14430 28988
rect 16025 28985 16037 29019
rect 16071 29016 16083 29019
rect 16574 29016 16580 29028
rect 16071 28988 16580 29016
rect 16071 28985 16083 28988
rect 16025 28979 16083 28985
rect 16574 28976 16580 28988
rect 16632 28976 16638 29028
rect 17034 28976 17040 29028
rect 17092 29016 17098 29028
rect 18064 29016 18092 29115
rect 18506 29112 18512 29124
rect 18564 29112 18570 29164
rect 18598 29112 18604 29164
rect 18656 29112 18662 29164
rect 18693 29155 18751 29161
rect 18693 29121 18705 29155
rect 18739 29152 18751 29155
rect 18782 29152 18788 29164
rect 18739 29124 18788 29152
rect 18739 29121 18751 29124
rect 18693 29115 18751 29121
rect 18782 29112 18788 29124
rect 18840 29152 18846 29164
rect 18892 29152 18920 29183
rect 19702 29180 19708 29232
rect 19760 29220 19766 29232
rect 23106 29220 23112 29232
rect 19760 29192 20576 29220
rect 19760 29180 19766 29192
rect 18840 29124 18920 29152
rect 19153 29155 19211 29161
rect 18840 29112 18846 29124
rect 19153 29121 19165 29155
rect 19199 29152 19211 29155
rect 20438 29152 20444 29164
rect 19199 29124 20444 29152
rect 19199 29121 19211 29124
rect 19153 29115 19211 29121
rect 20438 29112 20444 29124
rect 20496 29112 20502 29164
rect 18877 29087 18935 29093
rect 18877 29053 18889 29087
rect 18923 29084 18935 29087
rect 19337 29087 19395 29093
rect 19337 29084 19349 29087
rect 18923 29056 19349 29084
rect 18923 29053 18935 29056
rect 18877 29047 18935 29053
rect 19337 29053 19349 29056
rect 19383 29053 19395 29087
rect 19337 29047 19395 29053
rect 19518 29044 19524 29096
rect 19576 29044 19582 29096
rect 19610 29044 19616 29096
rect 19668 29044 19674 29096
rect 19702 29044 19708 29096
rect 19760 29044 19766 29096
rect 19797 29087 19855 29093
rect 19797 29053 19809 29087
rect 19843 29084 19855 29087
rect 20346 29084 20352 29096
rect 19843 29056 20352 29084
rect 19843 29053 19855 29056
rect 19797 29047 19855 29053
rect 20346 29044 20352 29056
rect 20404 29044 20410 29096
rect 17092 28988 18092 29016
rect 18509 29019 18567 29025
rect 17092 28976 17098 28988
rect 18509 28985 18521 29019
rect 18555 29016 18567 29019
rect 19061 29019 19119 29025
rect 18555 28988 18920 29016
rect 18555 28985 18567 28988
rect 18509 28979 18567 28985
rect 18892 28960 18920 28988
rect 19061 28985 19073 29019
rect 19107 29016 19119 29019
rect 20070 29016 20076 29028
rect 19107 28988 20076 29016
rect 19107 28985 19119 28988
rect 19061 28979 19119 28985
rect 20070 28976 20076 28988
rect 20128 28976 20134 29028
rect 13955 28920 14044 28948
rect 14185 28951 14243 28957
rect 13955 28917 13967 28920
rect 13909 28911 13967 28917
rect 14185 28917 14197 28951
rect 14231 28948 14243 28951
rect 14274 28948 14280 28960
rect 14231 28920 14280 28948
rect 14231 28917 14243 28920
rect 14185 28911 14243 28917
rect 14274 28908 14280 28920
rect 14332 28908 14338 28960
rect 15657 28951 15715 28957
rect 15657 28917 15669 28951
rect 15703 28948 15715 28951
rect 16669 28951 16727 28957
rect 16669 28948 16681 28951
rect 15703 28920 16681 28948
rect 15703 28917 15715 28920
rect 15657 28911 15715 28917
rect 16669 28917 16681 28920
rect 16715 28917 16727 28951
rect 16669 28911 16727 28917
rect 18874 28908 18880 28960
rect 18932 28908 18938 28960
rect 20456 28948 20484 29112
rect 20548 29016 20576 29192
rect 22066 29192 23112 29220
rect 20625 29155 20683 29161
rect 20625 29121 20637 29155
rect 20671 29152 20683 29155
rect 20990 29152 20996 29164
rect 20671 29124 20996 29152
rect 20671 29121 20683 29124
rect 20625 29115 20683 29121
rect 20990 29112 20996 29124
rect 21048 29112 21054 29164
rect 21174 29112 21180 29164
rect 21232 29112 21238 29164
rect 20714 29044 20720 29096
rect 20772 29044 20778 29096
rect 20809 29087 20867 29093
rect 20809 29053 20821 29087
rect 20855 29053 20867 29087
rect 20809 29047 20867 29053
rect 20901 29087 20959 29093
rect 20901 29053 20913 29087
rect 20947 29084 20959 29087
rect 21192 29084 21220 29112
rect 20947 29056 21220 29084
rect 20947 29053 20959 29056
rect 20901 29047 20959 29053
rect 20824 29016 20852 29047
rect 21082 29016 21088 29028
rect 20548 28988 21088 29016
rect 21082 28976 21088 28988
rect 21140 28976 21146 29028
rect 22066 28948 22094 29192
rect 23106 29180 23112 29192
rect 23164 29180 23170 29232
rect 25685 29223 25743 29229
rect 25685 29220 25697 29223
rect 24320 29192 25697 29220
rect 22465 29155 22523 29161
rect 22465 29121 22477 29155
rect 22511 29152 22523 29155
rect 23017 29155 23075 29161
rect 22511 29124 22692 29152
rect 22511 29121 22523 29124
rect 22465 29115 22523 29121
rect 22664 29025 22692 29124
rect 23017 29121 23029 29155
rect 23063 29152 23075 29155
rect 23566 29152 23572 29164
rect 23063 29124 23572 29152
rect 23063 29121 23075 29124
rect 23017 29115 23075 29121
rect 23566 29112 23572 29124
rect 23624 29152 23630 29164
rect 24320 29161 24348 29192
rect 25685 29189 25697 29192
rect 25731 29189 25743 29223
rect 25685 29183 25743 29189
rect 24305 29155 24363 29161
rect 23624 29124 23796 29152
rect 23624 29112 23630 29124
rect 23293 29087 23351 29093
rect 23293 29053 23305 29087
rect 23339 29084 23351 29087
rect 23382 29084 23388 29096
rect 23339 29056 23388 29084
rect 23339 29053 23351 29056
rect 23293 29047 23351 29053
rect 23382 29044 23388 29056
rect 23440 29044 23446 29096
rect 23768 29084 23796 29124
rect 24305 29121 24317 29155
rect 24351 29121 24363 29155
rect 24305 29115 24363 29121
rect 24486 29112 24492 29164
rect 24544 29112 24550 29164
rect 24581 29155 24639 29161
rect 24581 29121 24593 29155
rect 24627 29121 24639 29155
rect 24581 29115 24639 29121
rect 24596 29084 24624 29115
rect 24670 29112 24676 29164
rect 24728 29112 24734 29164
rect 24762 29112 24768 29164
rect 24820 29152 24826 29164
rect 26329 29155 26387 29161
rect 24820 29124 25084 29152
rect 24820 29112 24826 29124
rect 24949 29087 25007 29093
rect 24949 29084 24961 29087
rect 23768 29056 24624 29084
rect 24872 29056 24961 29084
rect 24872 29025 24900 29056
rect 24949 29053 24961 29056
rect 24995 29053 25007 29087
rect 25056 29084 25084 29124
rect 26329 29121 26341 29155
rect 26375 29152 26387 29155
rect 26528 29152 26556 29248
rect 29178 29220 29184 29232
rect 28658 29192 29184 29220
rect 29178 29180 29184 29192
rect 29236 29180 29242 29232
rect 29454 29220 29460 29232
rect 29288 29192 29460 29220
rect 26375 29124 26556 29152
rect 26375 29121 26387 29124
rect 26329 29115 26387 29121
rect 26786 29112 26792 29164
rect 26844 29152 26850 29164
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 26844 29124 27169 29152
rect 26844 29112 26850 29124
rect 27157 29121 27169 29124
rect 27203 29121 27215 29155
rect 29288 29152 29316 29192
rect 29454 29180 29460 29192
rect 29512 29180 29518 29232
rect 31110 29180 31116 29232
rect 31168 29180 31174 29232
rect 27157 29115 27215 29121
rect 29196 29124 29316 29152
rect 29365 29155 29423 29161
rect 27433 29087 27491 29093
rect 25056 29056 27200 29084
rect 24949 29047 25007 29053
rect 27172 29028 27200 29056
rect 27433 29053 27445 29087
rect 27479 29084 27491 29087
rect 28997 29087 29055 29093
rect 28997 29084 29009 29087
rect 27479 29056 29009 29084
rect 27479 29053 27491 29056
rect 27433 29047 27491 29053
rect 28997 29053 29009 29056
rect 29043 29053 29055 29087
rect 28997 29047 29055 29053
rect 22649 29019 22707 29025
rect 22649 28985 22661 29019
rect 22695 28985 22707 29019
rect 22649 28979 22707 28985
rect 24857 29019 24915 29025
rect 24857 28985 24869 29019
rect 24903 28985 24915 29019
rect 24857 28979 24915 28985
rect 27154 28976 27160 29028
rect 27212 28976 27218 29028
rect 28905 29019 28963 29025
rect 28905 28985 28917 29019
rect 28951 29016 28963 29019
rect 29196 29016 29224 29124
rect 29365 29121 29377 29155
rect 29411 29152 29423 29155
rect 29546 29152 29552 29164
rect 29411 29124 29552 29152
rect 29411 29121 29423 29124
rect 29365 29115 29423 29121
rect 29546 29112 29552 29124
rect 29604 29112 29610 29164
rect 31404 29161 31432 29260
rect 31389 29155 31447 29161
rect 29273 29087 29331 29093
rect 29273 29053 29285 29087
rect 29319 29053 29331 29087
rect 30024 29084 30052 29138
rect 31389 29121 31401 29155
rect 31435 29121 31447 29155
rect 31389 29115 31447 29121
rect 29273 29047 29331 29053
rect 29472 29056 30052 29084
rect 28951 28988 29224 29016
rect 29288 29016 29316 29047
rect 29362 29016 29368 29028
rect 29288 28988 29368 29016
rect 28951 28985 28963 28988
rect 28905 28979 28963 28985
rect 29362 28976 29368 28988
rect 29420 28976 29426 29028
rect 20456 28920 22094 28948
rect 22278 28908 22284 28960
rect 22336 28908 22342 28960
rect 29178 28908 29184 28960
rect 29236 28948 29242 28960
rect 29472 28948 29500 29056
rect 29236 28920 29500 28948
rect 29236 28908 29242 28920
rect 29638 28908 29644 28960
rect 29696 28908 29702 28960
rect 1104 28858 34684 28880
rect 1104 28806 5147 28858
rect 5199 28806 5211 28858
rect 5263 28806 5275 28858
rect 5327 28806 5339 28858
rect 5391 28806 5403 28858
rect 5455 28806 13541 28858
rect 13593 28806 13605 28858
rect 13657 28806 13669 28858
rect 13721 28806 13733 28858
rect 13785 28806 13797 28858
rect 13849 28806 21935 28858
rect 21987 28806 21999 28858
rect 22051 28806 22063 28858
rect 22115 28806 22127 28858
rect 22179 28806 22191 28858
rect 22243 28806 30329 28858
rect 30381 28806 30393 28858
rect 30445 28806 30457 28858
rect 30509 28806 30521 28858
rect 30573 28806 30585 28858
rect 30637 28806 34684 28858
rect 1104 28784 34684 28806
rect 3789 28747 3847 28753
rect 3789 28713 3801 28747
rect 3835 28744 3847 28747
rect 3878 28744 3884 28756
rect 3835 28716 3884 28744
rect 3835 28713 3847 28716
rect 3789 28707 3847 28713
rect 3878 28704 3884 28716
rect 3936 28704 3942 28756
rect 4617 28747 4675 28753
rect 4617 28713 4629 28747
rect 4663 28713 4675 28747
rect 4617 28707 4675 28713
rect 5261 28747 5319 28753
rect 5261 28713 5273 28747
rect 5307 28744 5319 28747
rect 5810 28744 5816 28756
rect 5307 28716 5816 28744
rect 5307 28713 5319 28716
rect 5261 28707 5319 28713
rect 4080 28648 4568 28676
rect 3602 28568 3608 28620
rect 3660 28608 3666 28620
rect 4080 28617 4108 28648
rect 4065 28611 4123 28617
rect 4065 28608 4077 28611
rect 3660 28580 4077 28608
rect 3660 28568 3666 28580
rect 4065 28577 4077 28580
rect 4111 28577 4123 28611
rect 4065 28571 4123 28577
rect 4157 28611 4215 28617
rect 4157 28577 4169 28611
rect 4203 28608 4215 28611
rect 4203 28580 4476 28608
rect 4203 28577 4215 28580
rect 4157 28571 4215 28577
rect 2961 28543 3019 28549
rect 2961 28509 2973 28543
rect 3007 28509 3019 28543
rect 2961 28503 3019 28509
rect 3145 28543 3203 28549
rect 3145 28509 3157 28543
rect 3191 28540 3203 28543
rect 3234 28540 3240 28552
rect 3191 28512 3240 28540
rect 3191 28509 3203 28512
rect 3145 28503 3203 28509
rect 2976 28472 3004 28503
rect 3234 28500 3240 28512
rect 3292 28500 3298 28552
rect 3421 28543 3479 28549
rect 3421 28509 3433 28543
rect 3467 28540 3479 28543
rect 3970 28540 3976 28552
rect 3467 28512 3976 28540
rect 3467 28509 3479 28512
rect 3421 28503 3479 28509
rect 3970 28500 3976 28512
rect 4028 28500 4034 28552
rect 4249 28543 4307 28549
rect 4249 28509 4261 28543
rect 4295 28540 4307 28543
rect 4338 28540 4344 28552
rect 4295 28512 4344 28540
rect 4295 28509 4307 28512
rect 4249 28503 4307 28509
rect 4338 28500 4344 28512
rect 4396 28500 4402 28552
rect 4448 28484 4476 28580
rect 3694 28472 3700 28484
rect 2976 28444 3700 28472
rect 3694 28432 3700 28444
rect 3752 28432 3758 28484
rect 4430 28432 4436 28484
rect 4488 28432 4494 28484
rect 4540 28472 4568 28648
rect 4632 28608 4660 28707
rect 5810 28704 5816 28716
rect 5868 28744 5874 28756
rect 7282 28744 7288 28756
rect 5868 28716 7288 28744
rect 5868 28704 5874 28716
rect 7282 28704 7288 28716
rect 7340 28704 7346 28756
rect 10686 28704 10692 28756
rect 10744 28704 10750 28756
rect 15746 28704 15752 28756
rect 15804 28744 15810 28756
rect 15841 28747 15899 28753
rect 15841 28744 15853 28747
rect 15804 28716 15853 28744
rect 15804 28704 15810 28716
rect 15841 28713 15853 28716
rect 15887 28713 15899 28747
rect 15841 28707 15899 28713
rect 16574 28704 16580 28756
rect 16632 28744 16638 28756
rect 16669 28747 16727 28753
rect 16669 28744 16681 28747
rect 16632 28716 16681 28744
rect 16632 28704 16638 28716
rect 16669 28713 16681 28716
rect 16715 28713 16727 28747
rect 16669 28707 16727 28713
rect 16853 28747 16911 28753
rect 16853 28713 16865 28747
rect 16899 28713 16911 28747
rect 16853 28707 16911 28713
rect 4801 28679 4859 28685
rect 4801 28645 4813 28679
rect 4847 28676 4859 28679
rect 4890 28676 4896 28688
rect 4847 28648 4896 28676
rect 4847 28645 4859 28648
rect 4801 28639 4859 28645
rect 4890 28636 4896 28648
rect 4948 28636 4954 28688
rect 6917 28679 6975 28685
rect 5368 28648 6040 28676
rect 5368 28608 5396 28648
rect 4632 28580 5396 28608
rect 5534 28568 5540 28620
rect 5592 28608 5598 28620
rect 5905 28611 5963 28617
rect 5905 28608 5917 28611
rect 5592 28580 5917 28608
rect 5592 28568 5598 28580
rect 5905 28577 5917 28580
rect 5951 28577 5963 28611
rect 5905 28571 5963 28577
rect 6012 28552 6040 28648
rect 6917 28645 6929 28679
rect 6963 28676 6975 28679
rect 7190 28676 7196 28688
rect 6963 28648 7196 28676
rect 6963 28645 6975 28648
rect 6917 28639 6975 28645
rect 7190 28636 7196 28648
rect 7248 28636 7254 28688
rect 7469 28679 7527 28685
rect 7469 28645 7481 28679
rect 7515 28645 7527 28679
rect 16868 28676 16896 28707
rect 17954 28704 17960 28756
rect 18012 28744 18018 28756
rect 18325 28747 18383 28753
rect 18325 28744 18337 28747
rect 18012 28716 18337 28744
rect 18012 28704 18018 28716
rect 18325 28713 18337 28716
rect 18371 28713 18383 28747
rect 18325 28707 18383 28713
rect 18785 28747 18843 28753
rect 18785 28713 18797 28747
rect 18831 28744 18843 28747
rect 18874 28744 18880 28756
rect 18831 28716 18880 28744
rect 18831 28713 18843 28716
rect 18785 28707 18843 28713
rect 18874 28704 18880 28716
rect 18932 28704 18938 28756
rect 19518 28704 19524 28756
rect 19576 28704 19582 28756
rect 19610 28704 19616 28756
rect 19668 28744 19674 28756
rect 19705 28747 19763 28753
rect 19705 28744 19717 28747
rect 19668 28716 19717 28744
rect 19668 28704 19674 28716
rect 19705 28713 19717 28716
rect 19751 28713 19763 28747
rect 19705 28707 19763 28713
rect 20714 28704 20720 28756
rect 20772 28744 20778 28756
rect 20809 28747 20867 28753
rect 20809 28744 20821 28747
rect 20772 28716 20821 28744
rect 20772 28704 20778 28716
rect 20809 28713 20821 28716
rect 20855 28713 20867 28747
rect 20809 28707 20867 28713
rect 20990 28704 20996 28756
rect 21048 28704 21054 28756
rect 21818 28704 21824 28756
rect 21876 28704 21882 28756
rect 23106 28704 23112 28756
rect 23164 28744 23170 28756
rect 23477 28747 23535 28753
rect 23477 28744 23489 28747
rect 23164 28716 23489 28744
rect 23164 28704 23170 28716
rect 23477 28713 23489 28716
rect 23523 28713 23535 28747
rect 23477 28707 23535 28713
rect 28442 28704 28448 28756
rect 28500 28704 28506 28756
rect 28534 28704 28540 28756
rect 28592 28744 28598 28756
rect 29181 28747 29239 28753
rect 28592 28716 28764 28744
rect 28592 28704 28598 28716
rect 16942 28676 16948 28688
rect 16868 28648 16948 28676
rect 7469 28639 7527 28645
rect 4890 28500 4896 28552
rect 4948 28500 4954 28552
rect 5626 28540 5632 28552
rect 5000 28512 5632 28540
rect 5000 28472 5028 28512
rect 5626 28500 5632 28512
rect 5684 28500 5690 28552
rect 5718 28500 5724 28552
rect 5776 28500 5782 28552
rect 5813 28543 5871 28549
rect 5813 28509 5825 28543
rect 5859 28509 5871 28543
rect 5813 28503 5871 28509
rect 4540 28444 5028 28472
rect 5261 28475 5319 28481
rect 5261 28441 5273 28475
rect 5307 28472 5319 28475
rect 5644 28472 5672 28500
rect 5828 28472 5856 28503
rect 5994 28500 6000 28552
rect 6052 28540 6058 28552
rect 6454 28540 6460 28552
rect 6052 28512 6460 28540
rect 6052 28500 6058 28512
rect 6454 28500 6460 28512
rect 6512 28500 6518 28552
rect 7484 28540 7512 28639
rect 16942 28636 16948 28648
rect 17000 28676 17006 28688
rect 19536 28676 19564 28704
rect 19889 28679 19947 28685
rect 19889 28676 19901 28679
rect 17000 28648 18552 28676
rect 19536 28648 19901 28676
rect 17000 28636 17006 28648
rect 8938 28568 8944 28620
rect 8996 28568 9002 28620
rect 11330 28568 11336 28620
rect 11388 28608 11394 28620
rect 12253 28611 12311 28617
rect 12253 28608 12265 28611
rect 11388 28580 12265 28608
rect 11388 28568 11394 28580
rect 12253 28577 12265 28580
rect 12299 28577 12311 28611
rect 12253 28571 12311 28577
rect 14090 28568 14096 28620
rect 14148 28568 14154 28620
rect 18524 28552 18552 28648
rect 19889 28645 19901 28648
rect 19935 28645 19947 28679
rect 19889 28639 19947 28645
rect 18598 28568 18604 28620
rect 18656 28568 18662 28620
rect 21729 28611 21787 28617
rect 19812 28580 20208 28608
rect 8757 28543 8815 28549
rect 8757 28540 8769 28543
rect 7484 28512 8769 28540
rect 8757 28509 8769 28512
rect 8803 28509 8815 28543
rect 8757 28503 8815 28509
rect 18506 28500 18512 28552
rect 18564 28500 18570 28552
rect 18782 28500 18788 28552
rect 18840 28500 18846 28552
rect 18874 28500 18880 28552
rect 18932 28500 18938 28552
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 19812 28549 19840 28580
rect 19797 28543 19855 28549
rect 19392 28512 19748 28540
rect 19392 28500 19398 28512
rect 5307 28444 5580 28472
rect 5644 28444 5856 28472
rect 7285 28475 7343 28481
rect 5307 28441 5319 28444
rect 5261 28435 5319 28441
rect 2498 28364 2504 28416
rect 2556 28404 2562 28416
rect 3053 28407 3111 28413
rect 3053 28404 3065 28407
rect 2556 28376 3065 28404
rect 2556 28364 2562 28376
rect 3053 28373 3065 28376
rect 3099 28373 3111 28407
rect 3053 28367 3111 28373
rect 3234 28364 3240 28416
rect 3292 28404 3298 28416
rect 4633 28407 4691 28413
rect 4633 28404 4645 28407
rect 3292 28376 4645 28404
rect 3292 28364 3298 28376
rect 4633 28373 4645 28376
rect 4679 28373 4691 28407
rect 4633 28367 4691 28373
rect 5442 28364 5448 28416
rect 5500 28364 5506 28416
rect 5552 28413 5580 28444
rect 7285 28441 7297 28475
rect 7331 28472 7343 28475
rect 7374 28472 7380 28484
rect 7331 28444 7380 28472
rect 7331 28441 7343 28444
rect 7285 28435 7343 28441
rect 7374 28432 7380 28444
rect 7432 28432 7438 28484
rect 7650 28432 7656 28484
rect 7708 28432 7714 28484
rect 8481 28475 8539 28481
rect 8481 28441 8493 28475
rect 8527 28472 8539 28475
rect 8846 28472 8852 28484
rect 8527 28444 8852 28472
rect 8527 28441 8539 28444
rect 8481 28435 8539 28441
rect 8846 28432 8852 28444
rect 8904 28432 8910 28484
rect 9122 28432 9128 28484
rect 9180 28472 9186 28484
rect 9217 28475 9275 28481
rect 9217 28472 9229 28475
rect 9180 28444 9229 28472
rect 9180 28432 9186 28444
rect 9217 28441 9229 28444
rect 9263 28441 9275 28475
rect 9217 28435 9275 28441
rect 9766 28432 9772 28484
rect 9824 28432 9830 28484
rect 14274 28432 14280 28484
rect 14332 28472 14338 28484
rect 14369 28475 14427 28481
rect 14369 28472 14381 28475
rect 14332 28444 14381 28472
rect 14332 28432 14338 28444
rect 14369 28441 14381 28444
rect 14415 28441 14427 28475
rect 16574 28472 16580 28484
rect 15594 28444 16580 28472
rect 14369 28435 14427 28441
rect 16574 28432 16580 28444
rect 16632 28432 16638 28484
rect 17034 28432 17040 28484
rect 17092 28432 17098 28484
rect 18524 28472 18552 28500
rect 18892 28472 18920 28500
rect 18524 28444 18920 28472
rect 19521 28475 19579 28481
rect 19521 28441 19533 28475
rect 19567 28441 19579 28475
rect 19720 28472 19748 28512
rect 19797 28509 19809 28543
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 19981 28543 20039 28549
rect 19981 28509 19993 28543
rect 20027 28540 20039 28543
rect 20027 28512 20116 28540
rect 20027 28509 20039 28512
rect 19981 28503 20039 28509
rect 20088 28484 20116 28512
rect 20070 28472 20076 28484
rect 19720 28444 20076 28472
rect 19521 28435 19579 28441
rect 5537 28407 5595 28413
rect 5537 28373 5549 28407
rect 5583 28373 5595 28407
rect 5537 28367 5595 28373
rect 8570 28364 8576 28416
rect 8628 28364 8634 28416
rect 12897 28407 12955 28413
rect 12897 28373 12909 28407
rect 12943 28404 12955 28407
rect 13170 28404 13176 28416
rect 12943 28376 13176 28404
rect 12943 28373 12955 28376
rect 12897 28367 12955 28373
rect 13170 28364 13176 28376
rect 13228 28364 13234 28416
rect 16837 28407 16895 28413
rect 16837 28373 16849 28407
rect 16883 28404 16895 28407
rect 17494 28404 17500 28416
rect 16883 28376 17500 28404
rect 16883 28373 16895 28376
rect 16837 28367 16895 28373
rect 17494 28364 17500 28376
rect 17552 28364 17558 28416
rect 19536 28404 19564 28435
rect 20070 28432 20076 28444
rect 20128 28432 20134 28484
rect 20180 28404 20208 28580
rect 20456 28580 21128 28608
rect 20456 28552 20484 28580
rect 20438 28500 20444 28552
rect 20496 28500 20502 28552
rect 20625 28543 20683 28549
rect 20625 28509 20637 28543
rect 20671 28540 20683 28543
rect 20806 28540 20812 28552
rect 20671 28512 20812 28540
rect 20671 28509 20683 28512
rect 20625 28503 20683 28509
rect 20640 28404 20668 28503
rect 20806 28500 20812 28512
rect 20864 28540 20870 28552
rect 21100 28549 21128 28580
rect 21729 28577 21741 28611
rect 21775 28608 21787 28611
rect 21836 28608 21864 28704
rect 24486 28608 24492 28620
rect 21775 28580 21864 28608
rect 23768 28580 24492 28608
rect 21775 28577 21787 28580
rect 21729 28571 21787 28577
rect 20901 28543 20959 28549
rect 20901 28540 20913 28543
rect 20864 28512 20913 28540
rect 20864 28500 20870 28512
rect 20901 28509 20913 28512
rect 20947 28509 20959 28543
rect 20901 28503 20959 28509
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28509 21143 28543
rect 21085 28503 21143 28509
rect 23566 28500 23572 28552
rect 23624 28500 23630 28552
rect 23768 28549 23796 28580
rect 24486 28568 24492 28580
rect 24544 28568 24550 28620
rect 28353 28611 28411 28617
rect 28353 28608 28365 28611
rect 26528 28580 28365 28608
rect 23753 28543 23811 28549
rect 23753 28509 23765 28543
rect 23799 28509 23811 28543
rect 23753 28503 23811 28509
rect 23937 28543 23995 28549
rect 23937 28509 23949 28543
rect 23983 28540 23995 28543
rect 24670 28540 24676 28552
rect 23983 28512 24676 28540
rect 23983 28509 23995 28512
rect 23937 28503 23995 28509
rect 24670 28500 24676 28512
rect 24728 28500 24734 28552
rect 25041 28543 25099 28549
rect 25041 28509 25053 28543
rect 25087 28540 25099 28543
rect 25130 28540 25136 28552
rect 25087 28512 25136 28540
rect 25087 28509 25099 28512
rect 25041 28503 25099 28509
rect 25130 28500 25136 28512
rect 25188 28500 25194 28552
rect 26528 28549 26556 28580
rect 28353 28577 28365 28580
rect 28399 28577 28411 28611
rect 28460 28608 28488 28704
rect 28736 28617 28764 28716
rect 29181 28713 29193 28747
rect 29227 28713 29239 28747
rect 29181 28707 29239 28713
rect 28810 28636 28816 28688
rect 28868 28676 28874 28688
rect 29196 28676 29224 28707
rect 29362 28704 29368 28756
rect 29420 28704 29426 28756
rect 30377 28747 30435 28753
rect 30377 28713 30389 28747
rect 30423 28744 30435 28747
rect 30834 28744 30840 28756
rect 30423 28716 30840 28744
rect 30423 28713 30435 28716
rect 30377 28707 30435 28713
rect 30834 28704 30840 28716
rect 30892 28704 30898 28756
rect 28868 28648 29684 28676
rect 28868 28636 28874 28648
rect 29656 28620 29684 28648
rect 28537 28611 28595 28617
rect 28537 28608 28549 28611
rect 28460 28580 28549 28608
rect 28353 28571 28411 28577
rect 28537 28577 28549 28580
rect 28583 28577 28595 28611
rect 28537 28571 28595 28577
rect 28721 28611 28779 28617
rect 28721 28577 28733 28611
rect 28767 28577 28779 28611
rect 28721 28571 28779 28577
rect 28948 28568 28954 28620
rect 29006 28608 29012 28620
rect 29546 28608 29552 28620
rect 29006 28580 29552 28608
rect 29006 28568 29012 28580
rect 29546 28568 29552 28580
rect 29604 28568 29610 28620
rect 29638 28568 29644 28620
rect 29696 28568 29702 28620
rect 26513 28543 26571 28549
rect 26513 28509 26525 28543
rect 26559 28509 26571 28543
rect 26513 28503 26571 28509
rect 26694 28500 26700 28552
rect 26752 28500 26758 28552
rect 26789 28543 26847 28549
rect 26789 28509 26801 28543
rect 26835 28540 26847 28543
rect 27706 28540 27712 28552
rect 26835 28512 27712 28540
rect 26835 28509 26847 28512
rect 26789 28503 26847 28509
rect 27706 28500 27712 28512
rect 27764 28500 27770 28552
rect 28626 28500 28632 28552
rect 28684 28500 28690 28552
rect 28813 28543 28871 28549
rect 28813 28509 28825 28543
rect 28859 28509 28871 28543
rect 30558 28540 30564 28552
rect 28813 28503 28871 28509
rect 29012 28512 30564 28540
rect 22005 28475 22063 28481
rect 22005 28441 22017 28475
rect 22051 28472 22063 28475
rect 22278 28472 22284 28484
rect 22051 28444 22284 28472
rect 22051 28441 22063 28444
rect 22005 28435 22063 28441
rect 22278 28432 22284 28444
rect 22336 28432 22342 28484
rect 23290 28472 23296 28484
rect 23230 28444 23296 28472
rect 23290 28432 23296 28444
rect 23348 28432 23354 28484
rect 23842 28432 23848 28484
rect 23900 28432 23906 28484
rect 25774 28472 25780 28484
rect 24136 28444 25780 28472
rect 24136 28413 24164 28444
rect 25774 28432 25780 28444
rect 25832 28432 25838 28484
rect 19536 28376 20668 28404
rect 24121 28407 24179 28413
rect 24121 28373 24133 28407
rect 24167 28373 24179 28407
rect 24121 28367 24179 28373
rect 24302 28364 24308 28416
rect 24360 28404 24366 28416
rect 24397 28407 24455 28413
rect 24397 28404 24409 28407
rect 24360 28376 24409 28404
rect 24360 28364 24366 28376
rect 24397 28373 24409 28376
rect 24443 28373 24455 28407
rect 24397 28367 24455 28373
rect 26329 28407 26387 28413
rect 26329 28373 26341 28407
rect 26375 28404 26387 28407
rect 26970 28404 26976 28416
rect 26375 28376 26976 28404
rect 26375 28373 26387 28376
rect 26329 28367 26387 28373
rect 26970 28364 26976 28376
rect 27028 28364 27034 28416
rect 28350 28364 28356 28416
rect 28408 28404 28414 28416
rect 28828 28404 28856 28503
rect 29012 28484 29040 28512
rect 30558 28500 30564 28512
rect 30616 28500 30622 28552
rect 30653 28543 30711 28549
rect 30653 28509 30665 28543
rect 30699 28509 30711 28543
rect 30653 28503 30711 28509
rect 28948 28472 28954 28484
rect 28907 28444 28954 28472
rect 28948 28432 28954 28444
rect 29006 28481 29040 28484
rect 29006 28475 29055 28481
rect 29006 28441 29009 28475
rect 29043 28441 29055 28475
rect 29006 28435 29055 28441
rect 30285 28475 30343 28481
rect 30285 28441 30297 28475
rect 30331 28472 30343 28475
rect 30377 28475 30435 28481
rect 30377 28472 30389 28475
rect 30331 28444 30389 28472
rect 30331 28441 30343 28444
rect 30285 28435 30343 28441
rect 30377 28441 30389 28444
rect 30423 28441 30435 28475
rect 30377 28435 30435 28441
rect 29006 28432 29012 28435
rect 30668 28416 30696 28503
rect 28408 28376 28856 28404
rect 28408 28364 28414 28376
rect 29086 28364 29092 28416
rect 29144 28404 29150 28416
rect 29197 28407 29255 28413
rect 29197 28404 29209 28407
rect 29144 28376 29209 28404
rect 29144 28364 29150 28376
rect 29197 28373 29209 28376
rect 29243 28373 29255 28407
rect 29197 28367 29255 28373
rect 30650 28364 30656 28416
rect 30708 28364 30714 28416
rect 1104 28314 34840 28336
rect 1104 28262 9344 28314
rect 9396 28262 9408 28314
rect 9460 28262 9472 28314
rect 9524 28262 9536 28314
rect 9588 28262 9600 28314
rect 9652 28262 17738 28314
rect 17790 28262 17802 28314
rect 17854 28262 17866 28314
rect 17918 28262 17930 28314
rect 17982 28262 17994 28314
rect 18046 28262 26132 28314
rect 26184 28262 26196 28314
rect 26248 28262 26260 28314
rect 26312 28262 26324 28314
rect 26376 28262 26388 28314
rect 26440 28262 34526 28314
rect 34578 28262 34590 28314
rect 34642 28262 34654 28314
rect 34706 28262 34718 28314
rect 34770 28262 34782 28314
rect 34834 28262 34840 28314
rect 1104 28240 34840 28262
rect 2498 28200 2504 28212
rect 1872 28172 2504 28200
rect 1872 28141 1900 28172
rect 2498 28160 2504 28172
rect 2556 28160 2562 28212
rect 3329 28203 3387 28209
rect 3329 28169 3341 28203
rect 3375 28200 3387 28203
rect 3602 28200 3608 28212
rect 3375 28172 3608 28200
rect 3375 28169 3387 28172
rect 3329 28163 3387 28169
rect 1857 28135 1915 28141
rect 1857 28101 1869 28135
rect 1903 28101 1915 28135
rect 1857 28095 1915 28101
rect 3528 28073 3556 28172
rect 3602 28160 3608 28172
rect 3660 28160 3666 28212
rect 3694 28160 3700 28212
rect 3752 28200 3758 28212
rect 3789 28203 3847 28209
rect 3789 28200 3801 28203
rect 3752 28172 3801 28200
rect 3752 28160 3758 28172
rect 3789 28169 3801 28172
rect 3835 28169 3847 28203
rect 3789 28163 3847 28169
rect 5442 28160 5448 28212
rect 5500 28160 5506 28212
rect 7006 28160 7012 28212
rect 7064 28200 7070 28212
rect 7101 28203 7159 28209
rect 7101 28200 7113 28203
rect 7064 28172 7113 28200
rect 7064 28160 7070 28172
rect 7101 28169 7113 28172
rect 7147 28169 7159 28203
rect 7101 28163 7159 28169
rect 7650 28160 7656 28212
rect 7708 28200 7714 28212
rect 7708 28172 8892 28200
rect 7708 28160 7714 28172
rect 3513 28067 3571 28073
rect 1581 27999 1639 28005
rect 1581 27965 1593 27999
rect 1627 27965 1639 27999
rect 1581 27959 1639 27965
rect 1596 27860 1624 27959
rect 2976 27928 3004 28050
rect 3513 28033 3525 28067
rect 3559 28033 3571 28067
rect 4154 28064 4160 28076
rect 3513 28027 3571 28033
rect 3712 28036 4160 28064
rect 3605 27999 3663 28005
rect 3605 27965 3617 27999
rect 3651 27996 3663 27999
rect 3712 27996 3740 28036
rect 4154 28024 4160 28036
rect 4212 28024 4218 28076
rect 5460 28064 5488 28160
rect 8570 28092 8576 28144
rect 8628 28092 8634 28144
rect 5537 28067 5595 28073
rect 5537 28064 5549 28067
rect 5460 28036 5549 28064
rect 5537 28033 5549 28036
rect 5583 28033 5595 28067
rect 5537 28027 5595 28033
rect 5810 28024 5816 28076
rect 5868 28024 5874 28076
rect 5902 28024 5908 28076
rect 5960 28064 5966 28076
rect 8864 28073 8892 28172
rect 12342 28160 12348 28212
rect 12400 28160 12406 28212
rect 21818 28160 21824 28212
rect 21876 28200 21882 28212
rect 21876 28172 25636 28200
rect 21876 28160 21882 28172
rect 9766 28092 9772 28144
rect 9824 28092 9830 28144
rect 12360 28132 12388 28160
rect 12268 28104 12388 28132
rect 12529 28135 12587 28141
rect 8849 28067 8907 28073
rect 5960 28050 7498 28064
rect 5960 28036 7512 28050
rect 5960 28024 5966 28036
rect 3651 27968 3740 27996
rect 3789 27999 3847 28005
rect 3651 27965 3663 27968
rect 3605 27959 3663 27965
rect 3789 27965 3801 27999
rect 3835 27996 3847 27999
rect 3970 27996 3976 28008
rect 3835 27968 3976 27996
rect 3835 27965 3847 27968
rect 3789 27959 3847 27965
rect 3970 27956 3976 27968
rect 4028 27996 4034 28008
rect 5828 27996 5856 28024
rect 4028 27968 5856 27996
rect 4028 27956 4034 27968
rect 6178 27956 6184 28008
rect 6236 27956 6242 28008
rect 7484 27996 7512 28036
rect 8849 28033 8861 28067
rect 8895 28033 8907 28067
rect 8849 28027 8907 28033
rect 9784 27996 9812 28092
rect 11974 28024 11980 28076
rect 12032 28064 12038 28076
rect 12268 28073 12296 28104
rect 12529 28101 12541 28135
rect 12575 28132 12587 28135
rect 13446 28132 13452 28144
rect 12575 28104 13452 28132
rect 12575 28101 12587 28104
rect 12529 28095 12587 28101
rect 12253 28067 12311 28073
rect 12253 28064 12265 28067
rect 12032 28036 12265 28064
rect 12032 28024 12038 28036
rect 12253 28033 12265 28036
rect 12299 28033 12311 28067
rect 12253 28027 12311 28033
rect 12342 28024 12348 28076
rect 12400 28024 12406 28076
rect 7484 27968 9812 27996
rect 11238 27956 11244 28008
rect 11296 27996 11302 28008
rect 12158 27996 12164 28008
rect 11296 27968 12164 27996
rect 11296 27956 11302 27968
rect 12158 27956 12164 27968
rect 12216 27996 12222 28008
rect 12544 27996 12572 28095
rect 13446 28092 13452 28104
rect 13504 28132 13510 28144
rect 17034 28132 17040 28144
rect 13504 28104 17040 28132
rect 13504 28092 13510 28104
rect 17034 28092 17040 28104
rect 17092 28092 17098 28144
rect 20070 28092 20076 28144
rect 20128 28132 20134 28144
rect 22370 28132 22376 28144
rect 20128 28104 22376 28132
rect 20128 28092 20134 28104
rect 22370 28092 22376 28104
rect 22428 28132 22434 28144
rect 22557 28135 22615 28141
rect 22557 28132 22569 28135
rect 22428 28104 22569 28132
rect 22428 28092 22434 28104
rect 22557 28101 22569 28104
rect 22603 28101 22615 28135
rect 23382 28132 23388 28144
rect 22557 28095 22615 28101
rect 23124 28104 23388 28132
rect 22465 28067 22523 28073
rect 22465 28033 22477 28067
rect 22511 28064 22523 28067
rect 22925 28067 22983 28073
rect 22925 28064 22937 28067
rect 22511 28036 22937 28064
rect 22511 28033 22523 28036
rect 22465 28027 22523 28033
rect 22925 28033 22937 28036
rect 22971 28033 22983 28067
rect 22925 28027 22983 28033
rect 12216 27968 12572 27996
rect 22741 27999 22799 28005
rect 12216 27956 12222 27968
rect 22741 27965 22753 27999
rect 22787 27996 22799 27999
rect 23124 27996 23152 28104
rect 23382 28092 23388 28104
rect 23440 28092 23446 28144
rect 25608 28076 25636 28172
rect 26970 28160 26976 28212
rect 27028 28160 27034 28212
rect 27706 28160 27712 28212
rect 27764 28160 27770 28212
rect 30558 28160 30564 28212
rect 30616 28160 30622 28212
rect 32582 28200 32588 28212
rect 31726 28172 32588 28200
rect 22787 27968 23152 27996
rect 23216 28050 24242 28064
rect 23216 28036 24256 28050
rect 22787 27965 22799 27968
rect 22741 27959 22799 27965
rect 2976 27900 4292 27928
rect 3234 27860 3240 27872
rect 1596 27832 3240 27860
rect 3234 27820 3240 27832
rect 3292 27820 3298 27872
rect 4264 27860 4292 27900
rect 4338 27888 4344 27940
rect 4396 27928 4402 27940
rect 6196 27928 6224 27956
rect 4396 27900 6224 27928
rect 4396 27888 4402 27900
rect 18966 27888 18972 27940
rect 19024 27928 19030 27940
rect 23216 27928 23244 28036
rect 23474 27956 23480 28008
rect 23532 27956 23538 28008
rect 24228 27996 24256 28036
rect 25590 28024 25596 28076
rect 25648 28064 25654 28076
rect 26786 28064 26792 28076
rect 25648 28036 26792 28064
rect 25648 28024 25654 28036
rect 26786 28024 26792 28036
rect 26844 28024 26850 28076
rect 26988 28073 27016 28160
rect 30576 28132 30604 28160
rect 30742 28132 30748 28144
rect 30576 28104 30748 28132
rect 30742 28092 30748 28104
rect 30800 28132 30806 28144
rect 30800 28104 31156 28132
rect 30800 28092 30806 28104
rect 31128 28073 31156 28104
rect 26973 28067 27031 28073
rect 26973 28033 26985 28067
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 30101 28067 30159 28073
rect 30101 28033 30113 28067
rect 30147 28064 30159 28067
rect 30561 28067 30619 28073
rect 30561 28064 30573 28067
rect 30147 28036 30573 28064
rect 30147 28033 30159 28036
rect 30101 28027 30159 28033
rect 30561 28033 30573 28036
rect 30607 28033 30619 28067
rect 30561 28027 30619 28033
rect 31113 28067 31171 28073
rect 31113 28033 31125 28067
rect 31159 28033 31171 28067
rect 31113 28027 31171 28033
rect 24946 27996 24952 28008
rect 24228 27968 24952 27996
rect 24946 27956 24952 27968
rect 25004 27956 25010 28008
rect 25317 27999 25375 28005
rect 25317 27965 25329 27999
rect 25363 27996 25375 27999
rect 25685 27999 25743 28005
rect 25685 27996 25697 27999
rect 25363 27968 25697 27996
rect 25363 27965 25375 27968
rect 25317 27959 25375 27965
rect 25685 27965 25697 27968
rect 25731 27965 25743 27999
rect 25685 27959 25743 27965
rect 25774 27956 25780 28008
rect 25832 27996 25838 28008
rect 26237 27999 26295 28005
rect 26237 27996 26249 27999
rect 25832 27968 26249 27996
rect 25832 27956 25838 27968
rect 26237 27965 26249 27968
rect 26283 27965 26295 27999
rect 26237 27959 26295 27965
rect 27890 27956 27896 28008
rect 27948 27996 27954 28008
rect 28261 27999 28319 28005
rect 28261 27996 28273 27999
rect 27948 27968 28273 27996
rect 27948 27956 27954 27968
rect 28261 27965 28273 27968
rect 28307 27965 28319 27999
rect 28261 27959 28319 27965
rect 28350 27956 28356 28008
rect 28408 27996 28414 28008
rect 30009 27999 30067 28005
rect 30009 27996 30021 27999
rect 28408 27968 30021 27996
rect 28408 27956 28414 27968
rect 30009 27965 30021 27968
rect 30055 27965 30067 27999
rect 31726 27996 31754 28172
rect 32582 28160 32588 28172
rect 32640 28160 32646 28212
rect 34333 28067 34391 28073
rect 34333 28033 34345 28067
rect 34379 28033 34391 28067
rect 34333 28027 34391 28033
rect 30009 27959 30067 27965
rect 30392 27968 31754 27996
rect 34348 27996 34376 28027
rect 34790 27996 34796 28008
rect 34348 27968 34796 27996
rect 19024 27900 23244 27928
rect 19024 27888 19030 27900
rect 23566 27888 23572 27940
rect 23624 27928 23630 27940
rect 23845 27931 23903 27937
rect 23845 27928 23857 27931
rect 23624 27900 23857 27928
rect 23624 27888 23630 27900
rect 23845 27897 23857 27900
rect 23891 27897 23903 27931
rect 30392 27928 30420 27968
rect 34790 27956 34796 27968
rect 34848 27956 34854 28008
rect 23845 27891 23903 27897
rect 27540 27900 30420 27928
rect 30469 27931 30527 27937
rect 4982 27860 4988 27872
rect 4264 27832 4988 27860
rect 4982 27820 4988 27832
rect 5040 27820 5046 27872
rect 5353 27863 5411 27869
rect 5353 27829 5365 27863
rect 5399 27860 5411 27863
rect 5534 27860 5540 27872
rect 5399 27832 5540 27860
rect 5399 27829 5411 27832
rect 5353 27823 5411 27829
rect 5534 27820 5540 27832
rect 5592 27820 5598 27872
rect 12526 27820 12532 27872
rect 12584 27820 12590 27872
rect 22097 27863 22155 27869
rect 22097 27829 22109 27863
rect 22143 27860 22155 27863
rect 22278 27860 22284 27872
rect 22143 27832 22284 27860
rect 22143 27829 22155 27832
rect 22097 27823 22155 27829
rect 22278 27820 22284 27832
rect 22336 27820 22342 27872
rect 25130 27820 25136 27872
rect 25188 27860 25194 27872
rect 27540 27860 27568 27900
rect 30469 27897 30481 27931
rect 30515 27928 30527 27931
rect 30926 27928 30932 27940
rect 30515 27900 30932 27928
rect 30515 27897 30527 27900
rect 30469 27891 30527 27897
rect 30926 27888 30932 27900
rect 30984 27888 30990 27940
rect 25188 27832 27568 27860
rect 25188 27820 25194 27832
rect 27614 27820 27620 27872
rect 27672 27820 27678 27872
rect 34149 27863 34207 27869
rect 34149 27829 34161 27863
rect 34195 27860 34207 27863
rect 34195 27832 34744 27860
rect 34195 27829 34207 27832
rect 34149 27823 34207 27829
rect 1104 27770 34684 27792
rect 1104 27718 5147 27770
rect 5199 27718 5211 27770
rect 5263 27718 5275 27770
rect 5327 27718 5339 27770
rect 5391 27718 5403 27770
rect 5455 27718 13541 27770
rect 13593 27718 13605 27770
rect 13657 27718 13669 27770
rect 13721 27718 13733 27770
rect 13785 27718 13797 27770
rect 13849 27718 21935 27770
rect 21987 27718 21999 27770
rect 22051 27718 22063 27770
rect 22115 27718 22127 27770
rect 22179 27718 22191 27770
rect 22243 27718 30329 27770
rect 30381 27718 30393 27770
rect 30445 27718 30457 27770
rect 30509 27718 30521 27770
rect 30573 27718 30585 27770
rect 30637 27718 34684 27770
rect 1104 27696 34684 27718
rect 5432 27659 5490 27665
rect 5432 27625 5444 27659
rect 5478 27656 5490 27659
rect 5534 27656 5540 27668
rect 5478 27628 5540 27656
rect 5478 27625 5490 27628
rect 5432 27619 5490 27625
rect 5534 27616 5540 27628
rect 5592 27616 5598 27668
rect 22281 27659 22339 27665
rect 22281 27625 22293 27659
rect 22327 27656 22339 27659
rect 22370 27656 22376 27668
rect 22327 27628 22376 27656
rect 22327 27625 22339 27628
rect 22281 27619 22339 27625
rect 22370 27616 22376 27628
rect 22428 27616 22434 27668
rect 23842 27616 23848 27668
rect 23900 27656 23906 27668
rect 23937 27659 23995 27665
rect 23937 27656 23949 27659
rect 23900 27628 23949 27656
rect 23900 27616 23906 27628
rect 23937 27625 23949 27628
rect 23983 27625 23995 27659
rect 23937 27619 23995 27625
rect 27614 27616 27620 27668
rect 27672 27665 27678 27668
rect 27672 27659 27687 27665
rect 27675 27625 27687 27659
rect 27672 27619 27687 27625
rect 27672 27616 27678 27619
rect 30742 27616 30748 27668
rect 30800 27616 30806 27668
rect 30926 27616 30932 27668
rect 30984 27656 30990 27668
rect 32229 27659 32287 27665
rect 32229 27656 32241 27659
rect 30984 27628 32241 27656
rect 30984 27616 30990 27628
rect 32229 27625 32241 27628
rect 32275 27625 32287 27659
rect 32229 27619 32287 27625
rect 34075 27659 34133 27665
rect 34075 27625 34087 27659
rect 34121 27656 34133 27659
rect 34716 27656 34744 27832
rect 34121 27628 34744 27656
rect 34121 27625 34133 27628
rect 34075 27619 34133 27625
rect 6454 27548 6460 27600
rect 6512 27588 6518 27600
rect 6917 27591 6975 27597
rect 6917 27588 6929 27591
rect 6512 27560 6929 27588
rect 6512 27548 6518 27560
rect 6917 27557 6929 27560
rect 6963 27557 6975 27591
rect 6917 27551 6975 27557
rect 16022 27548 16028 27600
rect 16080 27548 16086 27600
rect 28902 27588 28908 27600
rect 28184 27560 28908 27588
rect 14642 27520 14648 27532
rect 13924 27492 14648 27520
rect 13924 27464 13952 27492
rect 14642 27480 14648 27492
rect 14700 27480 14706 27532
rect 20533 27523 20591 27529
rect 20533 27520 20545 27523
rect 16224 27492 18000 27520
rect 3234 27412 3240 27464
rect 3292 27452 3298 27464
rect 5169 27455 5227 27461
rect 5169 27452 5181 27455
rect 3292 27424 5181 27452
rect 3292 27412 3298 27424
rect 5169 27421 5181 27424
rect 5215 27421 5227 27455
rect 5169 27415 5227 27421
rect 10318 27412 10324 27464
rect 10376 27412 10382 27464
rect 11238 27412 11244 27464
rect 11296 27412 11302 27464
rect 11517 27455 11575 27461
rect 11517 27421 11529 27455
rect 11563 27452 11575 27455
rect 11974 27452 11980 27464
rect 11563 27424 11980 27452
rect 11563 27421 11575 27424
rect 11517 27415 11575 27421
rect 11974 27412 11980 27424
rect 12032 27412 12038 27464
rect 13633 27455 13691 27461
rect 13633 27421 13645 27455
rect 13679 27452 13691 27455
rect 13906 27452 13912 27464
rect 13679 27424 13912 27452
rect 13679 27421 13691 27424
rect 13633 27415 13691 27421
rect 13906 27412 13912 27424
rect 13964 27412 13970 27464
rect 14090 27412 14096 27464
rect 14148 27452 14154 27464
rect 14461 27455 14519 27461
rect 14461 27452 14473 27455
rect 14148 27424 14473 27452
rect 14148 27412 14154 27424
rect 14461 27421 14473 27424
rect 14507 27421 14519 27455
rect 14461 27415 14519 27421
rect 15378 27412 15384 27464
rect 15436 27412 15442 27464
rect 15838 27412 15844 27464
rect 15896 27412 15902 27464
rect 16224 27461 16252 27492
rect 16209 27455 16267 27461
rect 16209 27421 16221 27455
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 16301 27455 16359 27461
rect 16301 27421 16313 27455
rect 16347 27452 16359 27455
rect 16850 27452 16856 27464
rect 16347 27424 16856 27452
rect 16347 27421 16359 27424
rect 16301 27415 16359 27421
rect 16850 27412 16856 27424
rect 16908 27452 16914 27464
rect 17037 27455 17095 27461
rect 17037 27452 17049 27455
rect 16908 27424 17049 27452
rect 16908 27412 16914 27424
rect 17037 27421 17049 27424
rect 17083 27421 17095 27455
rect 17037 27415 17095 27421
rect 17494 27412 17500 27464
rect 17552 27452 17558 27464
rect 17972 27461 18000 27492
rect 19076 27492 20545 27520
rect 19076 27464 19104 27492
rect 20533 27489 20545 27492
rect 20579 27489 20591 27523
rect 20533 27483 20591 27489
rect 23385 27523 23443 27529
rect 23385 27489 23397 27523
rect 23431 27520 23443 27523
rect 23474 27520 23480 27532
rect 23431 27492 23480 27520
rect 23431 27489 23443 27492
rect 23385 27483 23443 27489
rect 23474 27480 23480 27492
rect 23532 27480 23538 27532
rect 26878 27480 26884 27532
rect 26936 27520 26942 27532
rect 27893 27523 27951 27529
rect 27893 27520 27905 27523
rect 26936 27492 27905 27520
rect 26936 27480 26942 27492
rect 27893 27489 27905 27492
rect 27939 27489 27951 27523
rect 27893 27483 27951 27489
rect 28074 27480 28080 27532
rect 28132 27480 28138 27532
rect 17589 27455 17647 27461
rect 17589 27452 17601 27455
rect 17552 27424 17601 27452
rect 17552 27412 17558 27424
rect 17589 27421 17601 27424
rect 17635 27421 17647 27455
rect 17589 27415 17647 27421
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27421 17831 27455
rect 17773 27415 17831 27421
rect 17957 27455 18015 27461
rect 17957 27421 17969 27455
rect 18003 27452 18015 27455
rect 18141 27455 18199 27461
rect 18141 27452 18153 27455
rect 18003 27424 18153 27452
rect 18003 27421 18015 27424
rect 17957 27415 18015 27421
rect 18141 27421 18153 27424
rect 18187 27421 18199 27455
rect 18141 27415 18199 27421
rect 18785 27455 18843 27461
rect 18785 27421 18797 27455
rect 18831 27452 18843 27455
rect 18874 27452 18880 27464
rect 18831 27424 18880 27452
rect 18831 27421 18843 27424
rect 18785 27415 18843 27421
rect 4982 27344 4988 27396
rect 5040 27384 5046 27396
rect 5902 27384 5908 27396
rect 5040 27356 5908 27384
rect 5040 27344 5046 27356
rect 5902 27344 5908 27356
rect 5960 27344 5966 27396
rect 12894 27344 12900 27396
rect 12952 27344 12958 27396
rect 13354 27344 13360 27396
rect 13412 27344 13418 27396
rect 16025 27387 16083 27393
rect 16025 27353 16037 27387
rect 16071 27384 16083 27387
rect 16666 27384 16672 27396
rect 16071 27356 16672 27384
rect 16071 27353 16083 27356
rect 16025 27347 16083 27353
rect 16666 27344 16672 27356
rect 16724 27344 16730 27396
rect 17788 27384 17816 27415
rect 18874 27412 18880 27424
rect 18932 27412 18938 27464
rect 19058 27412 19064 27464
rect 19116 27412 19122 27464
rect 19426 27412 19432 27464
rect 19484 27412 19490 27464
rect 22922 27412 22928 27464
rect 22980 27452 22986 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 22980 27424 24685 27452
rect 22980 27412 22986 27424
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 17052 27356 17816 27384
rect 17052 27328 17080 27356
rect 20806 27344 20812 27396
rect 20864 27344 20870 27396
rect 23290 27384 23296 27396
rect 22034 27356 23296 27384
rect 23290 27344 23296 27356
rect 23348 27344 23354 27396
rect 25866 27344 25872 27396
rect 25924 27344 25930 27396
rect 27154 27344 27160 27396
rect 27212 27384 27218 27396
rect 27522 27384 27528 27396
rect 27212 27356 27528 27384
rect 27212 27344 27218 27356
rect 27522 27344 27528 27356
rect 27580 27344 27586 27396
rect 27706 27344 27712 27396
rect 27764 27384 27770 27396
rect 28092 27384 28120 27480
rect 28184 27464 28212 27560
rect 28902 27548 28908 27560
rect 28960 27548 28966 27600
rect 28258 27480 28264 27532
rect 28316 27520 28322 27532
rect 32493 27523 32551 27529
rect 32493 27520 32505 27523
rect 28316 27492 32505 27520
rect 28316 27480 28322 27492
rect 32493 27489 32505 27492
rect 32539 27520 32551 27523
rect 33594 27520 33600 27532
rect 32539 27492 33600 27520
rect 32539 27489 32551 27492
rect 32493 27483 32551 27489
rect 33594 27480 33600 27492
rect 33652 27520 33658 27532
rect 34333 27523 34391 27529
rect 34333 27520 34345 27523
rect 33652 27492 34345 27520
rect 33652 27480 33658 27492
rect 34333 27489 34345 27492
rect 34379 27489 34391 27523
rect 34333 27483 34391 27489
rect 28166 27412 28172 27464
rect 28224 27412 28230 27464
rect 32950 27412 32956 27464
rect 33008 27412 33014 27464
rect 28905 27387 28963 27393
rect 28905 27384 28917 27387
rect 27764 27356 28917 27384
rect 27764 27344 27770 27356
rect 28905 27353 28917 27356
rect 28951 27384 28963 27387
rect 29086 27384 29092 27396
rect 28951 27356 29092 27384
rect 28951 27353 28963 27356
rect 28905 27347 28963 27353
rect 29086 27344 29092 27356
rect 29144 27384 29150 27396
rect 30650 27384 30656 27396
rect 29144 27356 30656 27384
rect 29144 27344 29150 27356
rect 30650 27344 30656 27356
rect 30708 27344 30714 27396
rect 31754 27344 31760 27396
rect 31812 27384 31818 27396
rect 32766 27384 32772 27396
rect 31812 27356 32772 27384
rect 31812 27344 31818 27356
rect 32766 27344 32772 27356
rect 32824 27344 32830 27396
rect 10134 27276 10140 27328
rect 10192 27276 10198 27328
rect 11054 27276 11060 27328
rect 11112 27276 11118 27328
rect 11425 27319 11483 27325
rect 11425 27285 11437 27319
rect 11471 27316 11483 27319
rect 11882 27316 11888 27328
rect 11471 27288 11888 27316
rect 11471 27285 11483 27288
rect 11425 27279 11483 27285
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 14274 27276 14280 27328
rect 14332 27276 14338 27328
rect 17034 27276 17040 27328
rect 17092 27276 17098 27328
rect 17586 27276 17592 27328
rect 17644 27316 17650 27328
rect 17865 27319 17923 27325
rect 17865 27316 17877 27319
rect 17644 27288 17877 27316
rect 17644 27276 17650 27288
rect 17865 27285 17877 27288
rect 17911 27285 17923 27319
rect 17865 27279 17923 27285
rect 19242 27276 19248 27328
rect 19300 27276 19306 27328
rect 25317 27319 25375 27325
rect 25317 27285 25329 27319
rect 25363 27316 25375 27319
rect 28442 27316 28448 27328
rect 25363 27288 28448 27316
rect 25363 27285 25375 27288
rect 25317 27279 25375 27285
rect 28442 27276 28448 27288
rect 28500 27276 28506 27328
rect 32582 27276 32588 27328
rect 32640 27276 32646 27328
rect 1104 27226 34840 27248
rect 1104 27174 9344 27226
rect 9396 27174 9408 27226
rect 9460 27174 9472 27226
rect 9524 27174 9536 27226
rect 9588 27174 9600 27226
rect 9652 27174 17738 27226
rect 17790 27174 17802 27226
rect 17854 27174 17866 27226
rect 17918 27174 17930 27226
rect 17982 27174 17994 27226
rect 18046 27174 26132 27226
rect 26184 27174 26196 27226
rect 26248 27174 26260 27226
rect 26312 27174 26324 27226
rect 26376 27174 26388 27226
rect 26440 27174 34526 27226
rect 34578 27174 34590 27226
rect 34642 27174 34654 27226
rect 34706 27174 34718 27226
rect 34770 27174 34782 27226
rect 34834 27174 34840 27226
rect 1104 27152 34840 27174
rect 10134 27112 10140 27124
rect 9876 27084 10140 27112
rect 9876 27053 9904 27084
rect 10134 27072 10140 27084
rect 10192 27072 10198 27124
rect 11238 27072 11244 27124
rect 11296 27112 11302 27124
rect 11333 27115 11391 27121
rect 11333 27112 11345 27115
rect 11296 27084 11345 27112
rect 11296 27072 11302 27084
rect 11333 27081 11345 27084
rect 11379 27112 11391 27115
rect 11675 27115 11733 27121
rect 11675 27112 11687 27115
rect 11379 27084 11687 27112
rect 11379 27081 11391 27084
rect 11333 27075 11391 27081
rect 11675 27081 11687 27084
rect 11721 27081 11733 27115
rect 11675 27075 11733 27081
rect 12342 27072 12348 27124
rect 12400 27112 12406 27124
rect 12713 27115 12771 27121
rect 12713 27112 12725 27115
rect 12400 27084 12725 27112
rect 12400 27072 12406 27084
rect 12713 27081 12725 27084
rect 12759 27081 12771 27115
rect 12713 27075 12771 27081
rect 13354 27072 13360 27124
rect 13412 27112 13418 27124
rect 13725 27115 13783 27121
rect 13725 27112 13737 27115
rect 13412 27084 13737 27112
rect 13412 27072 13418 27084
rect 13725 27081 13737 27084
rect 13771 27081 13783 27115
rect 14274 27112 14280 27124
rect 13725 27075 13783 27081
rect 14108 27084 14280 27112
rect 9861 27047 9919 27053
rect 9861 27013 9873 27047
rect 9907 27013 9919 27047
rect 9861 27007 9919 27013
rect 11882 27004 11888 27056
rect 11940 27044 11946 27056
rect 14108 27053 14136 27084
rect 14274 27072 14280 27084
rect 14332 27072 14338 27124
rect 16022 27072 16028 27124
rect 16080 27072 16086 27124
rect 16666 27072 16672 27124
rect 16724 27072 16730 27124
rect 16850 27072 16856 27124
rect 16908 27072 16914 27124
rect 16942 27072 16948 27124
rect 17000 27072 17006 27124
rect 17586 27112 17592 27124
rect 17420 27084 17592 27112
rect 14093 27047 14151 27053
rect 11940 27016 12112 27044
rect 11940 27004 11946 27016
rect 12084 26985 12112 27016
rect 14093 27013 14105 27047
rect 14139 27013 14151 27047
rect 15378 27044 15384 27056
rect 15318 27016 15384 27044
rect 14093 27007 14151 27013
rect 15378 27004 15384 27016
rect 15436 27004 15442 27056
rect 12069 26979 12127 26985
rect 7006 26868 7012 26920
rect 7064 26868 7070 26920
rect 7650 26868 7656 26920
rect 7708 26908 7714 26920
rect 9214 26908 9220 26920
rect 7708 26880 9220 26908
rect 7708 26868 7714 26880
rect 9214 26868 9220 26880
rect 9272 26908 9278 26920
rect 9585 26911 9643 26917
rect 9585 26908 9597 26911
rect 9272 26880 9597 26908
rect 9272 26868 9278 26880
rect 9585 26877 9597 26880
rect 9631 26877 9643 26911
rect 9585 26871 9643 26877
rect 10870 26868 10876 26920
rect 10928 26908 10934 26920
rect 10980 26908 11008 26962
rect 12069 26945 12081 26979
rect 12115 26945 12127 26979
rect 12069 26939 12127 26945
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26976 15991 26979
rect 16040 26976 16068 27072
rect 16868 26985 16896 27072
rect 16960 26985 16988 27072
rect 17420 27053 17448 27084
rect 17586 27072 17592 27084
rect 17644 27072 17650 27124
rect 18874 27072 18880 27124
rect 18932 27072 18938 27124
rect 19242 27072 19248 27124
rect 19300 27112 19306 27124
rect 19300 27084 19380 27112
rect 19300 27072 19306 27084
rect 17405 27047 17463 27053
rect 17405 27013 17417 27047
rect 17451 27013 17463 27047
rect 18966 27044 18972 27056
rect 18630 27016 18972 27044
rect 17405 27007 17463 27013
rect 18966 27004 18972 27016
rect 19024 27004 19030 27056
rect 19352 27053 19380 27084
rect 20806 27072 20812 27124
rect 20864 27112 20870 27124
rect 21821 27115 21879 27121
rect 21821 27112 21833 27115
rect 20864 27084 21833 27112
rect 20864 27072 20870 27084
rect 21821 27081 21833 27084
rect 21867 27081 21879 27115
rect 22922 27112 22928 27124
rect 21821 27075 21879 27081
rect 22066 27084 22928 27112
rect 19337 27047 19395 27053
rect 19337 27013 19349 27047
rect 19383 27013 19395 27047
rect 19337 27007 19395 27013
rect 20070 27004 20076 27056
rect 20128 27004 20134 27056
rect 22066 27044 22094 27084
rect 22922 27072 22928 27084
rect 22980 27072 22986 27124
rect 23017 27115 23075 27121
rect 23017 27081 23029 27115
rect 23063 27112 23075 27115
rect 23474 27112 23480 27124
rect 23063 27084 23480 27112
rect 23063 27081 23075 27084
rect 23017 27075 23075 27081
rect 23474 27072 23480 27084
rect 23532 27072 23538 27124
rect 25501 27115 25559 27121
rect 25501 27112 25513 27115
rect 24504 27084 25513 27112
rect 24504 27053 24532 27084
rect 25501 27081 25513 27084
rect 25547 27081 25559 27115
rect 25501 27075 25559 27081
rect 25866 27072 25872 27124
rect 25924 27072 25930 27124
rect 26605 27115 26663 27121
rect 26605 27081 26617 27115
rect 26651 27112 26663 27115
rect 26694 27112 26700 27124
rect 26651 27084 26700 27112
rect 26651 27081 26663 27084
rect 26605 27075 26663 27081
rect 26694 27072 26700 27084
rect 26752 27072 26758 27124
rect 29178 27112 29184 27124
rect 28920 27084 29184 27112
rect 21560 27016 22094 27044
rect 24489 27047 24547 27053
rect 21560 26985 21588 27016
rect 24489 27013 24501 27047
rect 24535 27013 24547 27047
rect 25884 27044 25912 27072
rect 26145 27047 26203 27053
rect 26145 27044 26157 27047
rect 24489 27007 24547 27013
rect 24780 27016 25636 27044
rect 25884 27016 26157 27044
rect 15979 26948 16068 26976
rect 16853 26979 16911 26985
rect 15979 26945 15991 26948
rect 15933 26939 15991 26945
rect 16853 26945 16865 26979
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 16945 26979 17003 26985
rect 16945 26945 16957 26979
rect 16991 26945 17003 26979
rect 21545 26979 21603 26985
rect 21545 26976 21557 26979
rect 16945 26939 17003 26945
rect 20824 26948 21557 26976
rect 12894 26908 12900 26920
rect 10928 26880 12900 26908
rect 10928 26868 10934 26880
rect 12894 26868 12900 26880
rect 12952 26868 12958 26920
rect 13078 26868 13084 26920
rect 13136 26868 13142 26920
rect 13817 26911 13875 26917
rect 13817 26877 13829 26911
rect 13863 26908 13875 26911
rect 13863 26880 13952 26908
rect 13863 26877 13875 26880
rect 13817 26871 13875 26877
rect 7282 26800 7288 26852
rect 7340 26800 7346 26852
rect 13924 26784 13952 26880
rect 14458 26868 14464 26920
rect 14516 26908 14522 26920
rect 16206 26908 16212 26920
rect 14516 26880 16212 26908
rect 14516 26868 14522 26880
rect 16206 26868 16212 26880
rect 16264 26908 16270 26920
rect 16669 26911 16727 26917
rect 16669 26908 16681 26911
rect 16264 26880 16681 26908
rect 16264 26868 16270 26880
rect 16669 26877 16681 26880
rect 16715 26877 16727 26911
rect 16669 26871 16727 26877
rect 16758 26868 16764 26920
rect 16816 26908 16822 26920
rect 17129 26911 17187 26917
rect 17129 26908 17141 26911
rect 16816 26880 17141 26908
rect 16816 26868 16822 26880
rect 17129 26877 17141 26880
rect 17175 26908 17187 26911
rect 19058 26908 19064 26920
rect 17175 26880 19064 26908
rect 17175 26877 17187 26880
rect 17129 26871 17187 26877
rect 19058 26868 19064 26880
rect 19116 26868 19122 26920
rect 20824 26917 20852 26948
rect 21545 26945 21557 26948
rect 21591 26945 21603 26979
rect 21545 26939 21603 26945
rect 22005 26979 22063 26985
rect 22005 26945 22017 26979
rect 22051 26976 22063 26979
rect 22278 26976 22284 26988
rect 22051 26948 22284 26976
rect 22051 26945 22063 26948
rect 22005 26939 22063 26945
rect 22278 26936 22284 26948
rect 22336 26936 22342 26988
rect 24780 26985 24808 27016
rect 25608 26988 25636 27016
rect 26145 27013 26157 27016
rect 26191 27013 26203 27047
rect 27890 27044 27896 27056
rect 26145 27007 26203 27013
rect 27172 27016 27896 27044
rect 24765 26979 24823 26985
rect 23308 26948 23414 26976
rect 20809 26911 20867 26917
rect 20809 26877 20821 26911
rect 20855 26877 20867 26911
rect 20809 26871 20867 26877
rect 23308 26784 23336 26948
rect 24765 26945 24777 26979
rect 24811 26945 24823 26979
rect 24765 26939 24823 26945
rect 25222 26936 25228 26988
rect 25280 26936 25286 26988
rect 25314 26936 25320 26988
rect 25372 26936 25378 26988
rect 25590 26936 25596 26988
rect 25648 26936 25654 26988
rect 23842 26868 23848 26920
rect 23900 26908 23906 26920
rect 23900 26880 24808 26908
rect 23900 26868 23906 26880
rect 24780 26840 24808 26880
rect 24854 26868 24860 26920
rect 24912 26868 24918 26920
rect 24949 26911 25007 26917
rect 24949 26877 24961 26911
rect 24995 26877 25007 26911
rect 26160 26908 26188 27007
rect 27172 26985 27200 27016
rect 27157 26979 27215 26985
rect 27157 26945 27169 26979
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27338 26936 27344 26988
rect 27396 26936 27402 26988
rect 27816 26985 27844 27016
rect 27890 27004 27896 27016
rect 27948 27004 27954 27056
rect 28920 27044 28948 27084
rect 29178 27072 29184 27084
rect 29236 27112 29242 27124
rect 29236 27084 31754 27112
rect 29236 27072 29242 27084
rect 31726 27056 31754 27084
rect 28000 27016 29026 27044
rect 31726 27016 31760 27056
rect 28000 26988 28028 27016
rect 31754 27004 31760 27016
rect 31812 27004 31818 27056
rect 27617 26979 27675 26985
rect 27617 26945 27629 26979
rect 27663 26945 27675 26979
rect 27617 26939 27675 26945
rect 27801 26979 27859 26985
rect 27801 26945 27813 26979
rect 27847 26945 27859 26979
rect 27801 26939 27859 26945
rect 26510 26908 26516 26920
rect 26160 26880 26516 26908
rect 24949 26871 25007 26877
rect 24964 26840 24992 26871
rect 26510 26868 26516 26880
rect 26568 26908 26574 26920
rect 27246 26908 27252 26920
rect 26568 26880 27252 26908
rect 26568 26868 26574 26880
rect 27246 26868 27252 26880
rect 27304 26908 27310 26920
rect 27632 26908 27660 26939
rect 27982 26936 27988 26988
rect 28040 26936 28046 26988
rect 28258 26936 28264 26988
rect 28316 26936 28322 26988
rect 30650 26936 30656 26988
rect 30708 26976 30714 26988
rect 32490 26976 32496 26988
rect 30708 26948 32496 26976
rect 30708 26936 30714 26948
rect 32490 26936 32496 26948
rect 32548 26936 32554 26988
rect 27304 26880 27660 26908
rect 27304 26868 27310 26880
rect 28534 26868 28540 26920
rect 28592 26868 28598 26920
rect 28626 26868 28632 26920
rect 28684 26908 28690 26920
rect 28684 26880 31616 26908
rect 28684 26868 28690 26880
rect 24780 26812 24992 26840
rect 25682 26800 25688 26852
rect 25740 26840 25746 26852
rect 26421 26843 26479 26849
rect 26421 26840 26433 26843
rect 25740 26812 26433 26840
rect 25740 26800 25746 26812
rect 26421 26809 26433 26812
rect 26467 26809 26479 26843
rect 26421 26803 26479 26809
rect 27154 26800 27160 26852
rect 27212 26840 27218 26852
rect 27893 26843 27951 26849
rect 27893 26840 27905 26843
rect 27212 26812 27905 26840
rect 27212 26800 27218 26812
rect 27893 26809 27905 26812
rect 27939 26809 27951 26843
rect 27893 26803 27951 26809
rect 31588 26784 31616 26880
rect 7466 26732 7472 26784
rect 7524 26732 7530 26784
rect 11514 26732 11520 26784
rect 11572 26732 11578 26784
rect 11701 26775 11759 26781
rect 11701 26741 11713 26775
rect 11747 26772 11759 26775
rect 11974 26772 11980 26784
rect 11747 26744 11980 26772
rect 11747 26741 11759 26744
rect 11701 26735 11759 26741
rect 11974 26732 11980 26744
rect 12032 26732 12038 26784
rect 13906 26732 13912 26784
rect 13964 26732 13970 26784
rect 14826 26732 14832 26784
rect 14884 26772 14890 26784
rect 15565 26775 15623 26781
rect 15565 26772 15577 26775
rect 14884 26744 15577 26772
rect 14884 26732 14890 26744
rect 15565 26741 15577 26744
rect 15611 26741 15623 26775
rect 15565 26735 15623 26741
rect 16482 26732 16488 26784
rect 16540 26732 16546 26784
rect 20898 26732 20904 26784
rect 20956 26732 20962 26784
rect 23290 26732 23296 26784
rect 23348 26732 23354 26784
rect 28074 26732 28080 26784
rect 28132 26772 28138 26784
rect 29914 26772 29920 26784
rect 28132 26744 29920 26772
rect 28132 26732 28138 26744
rect 29914 26732 29920 26744
rect 29972 26772 29978 26784
rect 30009 26775 30067 26781
rect 30009 26772 30021 26775
rect 29972 26744 30021 26772
rect 29972 26732 29978 26744
rect 30009 26741 30021 26744
rect 30055 26741 30067 26775
rect 30009 26735 30067 26741
rect 31570 26732 31576 26784
rect 31628 26732 31634 26784
rect 1104 26682 34684 26704
rect 1104 26630 5147 26682
rect 5199 26630 5211 26682
rect 5263 26630 5275 26682
rect 5327 26630 5339 26682
rect 5391 26630 5403 26682
rect 5455 26630 13541 26682
rect 13593 26630 13605 26682
rect 13657 26630 13669 26682
rect 13721 26630 13733 26682
rect 13785 26630 13797 26682
rect 13849 26630 21935 26682
rect 21987 26630 21999 26682
rect 22051 26630 22063 26682
rect 22115 26630 22127 26682
rect 22179 26630 22191 26682
rect 22243 26630 30329 26682
rect 30381 26630 30393 26682
rect 30445 26630 30457 26682
rect 30509 26630 30521 26682
rect 30573 26630 30585 26682
rect 30637 26630 34684 26682
rect 1104 26608 34684 26630
rect 6457 26571 6515 26577
rect 6457 26537 6469 26571
rect 6503 26568 6515 26571
rect 7282 26568 7288 26580
rect 6503 26540 7288 26568
rect 6503 26537 6515 26540
rect 6457 26531 6515 26537
rect 7282 26528 7288 26540
rect 7340 26528 7346 26580
rect 9950 26528 9956 26580
rect 10008 26528 10014 26580
rect 10318 26528 10324 26580
rect 10376 26528 10382 26580
rect 10505 26571 10563 26577
rect 10505 26537 10517 26571
rect 10551 26537 10563 26571
rect 10505 26531 10563 26537
rect 9968 26500 9996 26528
rect 10520 26500 10548 26531
rect 12250 26528 12256 26580
rect 12308 26528 12314 26580
rect 12621 26571 12679 26577
rect 12621 26537 12633 26571
rect 12667 26568 12679 26571
rect 13078 26568 13084 26580
rect 12667 26540 13084 26568
rect 12667 26537 12679 26540
rect 12621 26531 12679 26537
rect 13078 26528 13084 26540
rect 13136 26528 13142 26580
rect 14090 26528 14096 26580
rect 14148 26528 14154 26580
rect 14277 26571 14335 26577
rect 14277 26537 14289 26571
rect 14323 26568 14335 26571
rect 14366 26568 14372 26580
rect 14323 26540 14372 26568
rect 14323 26537 14335 26540
rect 14277 26531 14335 26537
rect 14366 26528 14372 26540
rect 14424 26528 14430 26580
rect 16104 26571 16162 26577
rect 16104 26537 16116 26571
rect 16150 26568 16162 26571
rect 16482 26568 16488 26580
rect 16150 26540 16488 26568
rect 16150 26537 16162 26540
rect 16104 26531 16162 26537
rect 16482 26528 16488 26540
rect 16540 26528 16546 26580
rect 17494 26528 17500 26580
rect 17552 26568 17558 26580
rect 17589 26571 17647 26577
rect 17589 26568 17601 26571
rect 17552 26540 17601 26568
rect 17552 26528 17558 26540
rect 17589 26537 17601 26540
rect 17635 26537 17647 26571
rect 17589 26531 17647 26537
rect 19337 26571 19395 26577
rect 19337 26537 19349 26571
rect 19383 26568 19395 26571
rect 19426 26568 19432 26580
rect 19383 26540 19432 26568
rect 19383 26537 19395 26540
rect 19337 26531 19395 26537
rect 19426 26528 19432 26540
rect 19484 26528 19490 26580
rect 21177 26571 21235 26577
rect 21177 26537 21189 26571
rect 21223 26568 21235 26571
rect 21223 26540 21404 26568
rect 21223 26537 21235 26540
rect 21177 26531 21235 26537
rect 9968 26472 10548 26500
rect 10873 26503 10931 26509
rect 10873 26469 10885 26503
rect 10919 26500 10931 26503
rect 11514 26500 11520 26512
rect 10919 26472 11520 26500
rect 10919 26469 10931 26472
rect 10873 26463 10931 26469
rect 11514 26460 11520 26472
rect 11572 26460 11578 26512
rect 19076 26472 21312 26500
rect 19076 26444 19104 26472
rect 3234 26392 3240 26444
rect 3292 26432 3298 26444
rect 3789 26435 3847 26441
rect 3789 26432 3801 26435
rect 3292 26404 3801 26432
rect 3292 26392 3298 26404
rect 3789 26401 3801 26404
rect 3835 26432 3847 26435
rect 6917 26435 6975 26441
rect 6917 26432 6929 26435
rect 3835 26404 6929 26432
rect 3835 26401 3847 26404
rect 3789 26395 3847 26401
rect 6917 26401 6929 26404
rect 6963 26432 6975 26435
rect 7650 26432 7656 26444
rect 6963 26404 7656 26432
rect 6963 26401 6975 26404
rect 6917 26395 6975 26401
rect 7650 26392 7656 26404
rect 7708 26392 7714 26444
rect 11054 26392 11060 26444
rect 11112 26392 11118 26444
rect 12161 26435 12219 26441
rect 12161 26401 12173 26435
rect 12207 26432 12219 26435
rect 12342 26432 12348 26444
rect 12207 26404 12348 26432
rect 12207 26401 12219 26404
rect 12161 26395 12219 26401
rect 12342 26392 12348 26404
rect 12400 26392 12406 26444
rect 15841 26435 15899 26441
rect 15841 26432 15853 26435
rect 13924 26404 15853 26432
rect 3418 26324 3424 26376
rect 3476 26324 3482 26376
rect 5074 26324 5080 26376
rect 5132 26364 5138 26376
rect 5132 26336 5198 26364
rect 5132 26324 5138 26336
rect 5626 26324 5632 26376
rect 5684 26364 5690 26376
rect 5813 26367 5871 26373
rect 5813 26364 5825 26367
rect 5684 26336 5825 26364
rect 5684 26324 5690 26336
rect 5813 26333 5825 26336
rect 5859 26333 5871 26367
rect 5997 26367 6055 26373
rect 5997 26364 6009 26367
rect 5813 26327 5871 26333
rect 5920 26336 6009 26364
rect 1394 26256 1400 26308
rect 1452 26256 1458 26308
rect 1765 26299 1823 26305
rect 1765 26265 1777 26299
rect 1811 26296 1823 26299
rect 1854 26296 1860 26308
rect 1811 26268 1860 26296
rect 1811 26265 1823 26268
rect 1765 26259 1823 26265
rect 1854 26256 1860 26268
rect 1912 26256 1918 26308
rect 4065 26299 4123 26305
rect 4065 26296 4077 26299
rect 3620 26268 4077 26296
rect 3620 26237 3648 26268
rect 4065 26265 4077 26268
rect 4111 26265 4123 26299
rect 4065 26259 4123 26265
rect 5920 26240 5948 26336
rect 5997 26333 6009 26336
rect 6043 26333 6055 26367
rect 5997 26327 6055 26333
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26364 6239 26367
rect 6273 26367 6331 26373
rect 6273 26364 6285 26367
rect 6227 26336 6285 26364
rect 6227 26333 6239 26336
rect 6181 26327 6239 26333
rect 6273 26333 6285 26336
rect 6319 26333 6331 26367
rect 9766 26364 9772 26376
rect 8326 26336 9772 26364
rect 6273 26327 6331 26333
rect 9766 26324 9772 26336
rect 9824 26324 9830 26376
rect 7190 26256 7196 26308
rect 7248 26256 7254 26308
rect 10505 26299 10563 26305
rect 10505 26265 10517 26299
rect 10551 26296 10563 26299
rect 11072 26296 11100 26392
rect 13924 26376 13952 26404
rect 15841 26401 15853 26404
rect 15887 26432 15899 26435
rect 16758 26432 16764 26444
rect 15887 26404 16764 26432
rect 15887 26401 15899 26404
rect 15841 26395 15899 26401
rect 16758 26392 16764 26404
rect 16816 26392 16822 26444
rect 19058 26392 19064 26444
rect 19116 26392 19122 26444
rect 19978 26392 19984 26444
rect 20036 26392 20042 26444
rect 20898 26392 20904 26444
rect 20956 26392 20962 26444
rect 21284 26441 21312 26472
rect 21269 26435 21327 26441
rect 21269 26401 21281 26435
rect 21315 26401 21327 26435
rect 21376 26432 21404 26540
rect 25222 26528 25228 26580
rect 25280 26568 25286 26580
rect 26973 26571 27031 26577
rect 25280 26540 26924 26568
rect 25280 26528 25286 26540
rect 26896 26500 26924 26540
rect 26973 26537 26985 26571
rect 27019 26568 27031 26571
rect 27890 26568 27896 26580
rect 27019 26540 27896 26568
rect 27019 26537 27031 26540
rect 26973 26531 27031 26537
rect 27890 26528 27896 26540
rect 27948 26528 27954 26580
rect 28534 26528 28540 26580
rect 28592 26568 28598 26580
rect 28813 26571 28871 26577
rect 28813 26568 28825 26571
rect 28592 26540 28825 26568
rect 28592 26528 28598 26540
rect 28813 26537 28825 26540
rect 28859 26537 28871 26571
rect 28813 26531 28871 26537
rect 30024 26540 30236 26568
rect 28902 26500 28908 26512
rect 26896 26472 28908 26500
rect 28902 26460 28908 26472
rect 28960 26500 28966 26512
rect 30024 26500 30052 26540
rect 28960 26472 30052 26500
rect 28960 26460 28966 26472
rect 21545 26435 21603 26441
rect 21545 26432 21557 26435
rect 21376 26404 21557 26432
rect 21269 26395 21327 26401
rect 21545 26401 21557 26404
rect 21591 26401 21603 26435
rect 21545 26395 21603 26401
rect 23017 26435 23075 26441
rect 23017 26401 23029 26435
rect 23063 26432 23075 26435
rect 23753 26435 23811 26441
rect 23753 26432 23765 26435
rect 23063 26404 23765 26432
rect 23063 26401 23075 26404
rect 23017 26395 23075 26401
rect 23753 26401 23765 26404
rect 23799 26432 23811 26435
rect 27341 26435 27399 26441
rect 27341 26432 27353 26435
rect 23799 26404 27353 26432
rect 23799 26401 23811 26404
rect 23753 26395 23811 26401
rect 27341 26401 27353 26404
rect 27387 26401 27399 26435
rect 27341 26395 27399 26401
rect 27985 26435 28043 26441
rect 27985 26401 27997 26435
rect 28031 26432 28043 26435
rect 30208 26432 30236 26540
rect 33594 26528 33600 26580
rect 33652 26528 33658 26580
rect 33612 26441 33640 26528
rect 30653 26435 30711 26441
rect 30653 26432 30665 26435
rect 28031 26404 29776 26432
rect 30208 26404 30665 26432
rect 28031 26401 28043 26404
rect 27985 26395 28043 26401
rect 12437 26367 12495 26373
rect 12437 26333 12449 26367
rect 12483 26364 12495 26367
rect 12526 26364 12532 26376
rect 12483 26336 12532 26364
rect 12483 26333 12495 26336
rect 12437 26327 12495 26333
rect 12526 26324 12532 26336
rect 12584 26324 12590 26376
rect 13906 26324 13912 26376
rect 13964 26324 13970 26376
rect 14550 26324 14556 26376
rect 14608 26364 14614 26376
rect 14645 26367 14703 26373
rect 14645 26364 14657 26367
rect 14608 26336 14657 26364
rect 14608 26324 14614 26336
rect 14645 26333 14657 26336
rect 14691 26333 14703 26367
rect 14645 26327 14703 26333
rect 14826 26324 14832 26376
rect 14884 26364 14890 26376
rect 14921 26367 14979 26373
rect 14921 26364 14933 26367
rect 14884 26336 14933 26364
rect 14884 26324 14890 26336
rect 14921 26333 14933 26336
rect 14967 26333 14979 26367
rect 14921 26327 14979 26333
rect 19705 26367 19763 26373
rect 19705 26333 19717 26367
rect 19751 26364 19763 26367
rect 20916 26364 20944 26392
rect 19751 26336 20944 26364
rect 19751 26333 19763 26336
rect 19705 26327 19763 26333
rect 20990 26324 20996 26376
rect 21048 26324 21054 26376
rect 25038 26324 25044 26376
rect 25096 26324 25102 26376
rect 25225 26367 25283 26373
rect 25225 26333 25237 26367
rect 25271 26333 25283 26367
rect 25225 26327 25283 26333
rect 10551 26268 11100 26296
rect 14277 26299 14335 26305
rect 10551 26265 10563 26268
rect 10505 26259 10563 26265
rect 14277 26265 14289 26299
rect 14323 26296 14335 26299
rect 14323 26268 14688 26296
rect 14323 26265 14335 26268
rect 14277 26259 14335 26265
rect 3605 26231 3663 26237
rect 3605 26197 3617 26231
rect 3651 26197 3663 26231
rect 3605 26191 3663 26197
rect 5534 26188 5540 26240
rect 5592 26188 5598 26240
rect 5902 26188 5908 26240
rect 5960 26188 5966 26240
rect 8662 26188 8668 26240
rect 8720 26188 8726 26240
rect 14660 26228 14688 26268
rect 14734 26256 14740 26308
rect 14792 26256 14798 26308
rect 15105 26299 15163 26305
rect 15105 26296 15117 26299
rect 15028 26268 15117 26296
rect 15028 26228 15056 26268
rect 15105 26265 15117 26268
rect 15151 26265 15163 26299
rect 15105 26259 15163 26265
rect 16574 26256 16580 26308
rect 16632 26256 16638 26308
rect 19797 26299 19855 26305
rect 19797 26265 19809 26299
rect 19843 26296 19855 26299
rect 20714 26296 20720 26308
rect 19843 26268 20720 26296
rect 19843 26265 19855 26268
rect 19797 26259 19855 26265
rect 20714 26256 20720 26268
rect 20772 26256 20778 26308
rect 23290 26296 23296 26308
rect 22770 26268 23296 26296
rect 23290 26256 23296 26268
rect 23348 26256 23354 26308
rect 23566 26256 23572 26308
rect 23624 26296 23630 26308
rect 24397 26299 24455 26305
rect 24397 26296 24409 26299
rect 23624 26268 24409 26296
rect 23624 26256 23630 26268
rect 24397 26265 24409 26268
rect 24443 26265 24455 26299
rect 25240 26296 25268 26327
rect 28074 26324 28080 26376
rect 28132 26364 28138 26376
rect 28169 26367 28227 26373
rect 28169 26364 28181 26367
rect 28132 26336 28181 26364
rect 28132 26324 28138 26336
rect 28169 26333 28181 26336
rect 28215 26333 28227 26367
rect 28169 26327 28227 26333
rect 28442 26324 28448 26376
rect 28500 26324 28506 26376
rect 28534 26324 28540 26376
rect 28592 26324 28598 26376
rect 28997 26367 29055 26373
rect 28997 26364 29009 26367
rect 28736 26336 29009 26364
rect 25240 26268 25452 26296
rect 24397 26259 24455 26265
rect 25424 26240 25452 26268
rect 25498 26256 25504 26308
rect 25556 26256 25562 26308
rect 27982 26296 27988 26308
rect 26726 26268 27988 26296
rect 27982 26256 27988 26268
rect 28040 26256 28046 26308
rect 28353 26299 28411 26305
rect 28353 26265 28365 26299
rect 28399 26296 28411 26299
rect 28626 26296 28632 26308
rect 28399 26268 28632 26296
rect 28399 26265 28411 26268
rect 28353 26259 28411 26265
rect 28626 26256 28632 26268
rect 28684 26256 28690 26308
rect 14660 26200 15056 26228
rect 23106 26188 23112 26240
rect 23164 26188 23170 26240
rect 25406 26188 25412 26240
rect 25464 26188 25470 26240
rect 28736 26237 28764 26336
rect 28997 26333 29009 26336
rect 29043 26333 29055 26367
rect 28997 26327 29055 26333
rect 29086 26324 29092 26376
rect 29144 26364 29150 26376
rect 29181 26367 29239 26373
rect 29181 26364 29193 26367
rect 29144 26336 29193 26364
rect 29144 26324 29150 26336
rect 29181 26333 29193 26336
rect 29227 26333 29239 26367
rect 29181 26327 29239 26333
rect 29273 26367 29331 26373
rect 29273 26333 29285 26367
rect 29319 26364 29331 26367
rect 29319 26336 29684 26364
rect 29319 26333 29331 26336
rect 29273 26327 29331 26333
rect 28721 26231 28779 26237
rect 28721 26197 28733 26231
rect 28767 26197 28779 26231
rect 29656 26228 29684 26336
rect 29748 26296 29776 26404
rect 30653 26401 30665 26404
rect 30699 26401 30711 26435
rect 31849 26435 31907 26441
rect 31849 26432 31861 26435
rect 30653 26395 30711 26401
rect 31220 26404 31861 26432
rect 29822 26324 29828 26376
rect 29880 26364 29886 26376
rect 31220 26373 31248 26404
rect 31849 26401 31861 26404
rect 31895 26401 31907 26435
rect 31849 26395 31907 26401
rect 33597 26435 33655 26441
rect 33597 26401 33609 26435
rect 33643 26401 33655 26435
rect 33597 26395 33655 26401
rect 30561 26367 30619 26373
rect 30561 26364 30573 26367
rect 29880 26336 30573 26364
rect 29880 26324 29886 26336
rect 30561 26333 30573 26336
rect 30607 26364 30619 26367
rect 31205 26367 31263 26373
rect 31205 26364 31217 26367
rect 30607 26336 31217 26364
rect 30607 26333 30619 26336
rect 30561 26327 30619 26333
rect 31205 26333 31217 26336
rect 31251 26333 31263 26367
rect 31481 26367 31539 26373
rect 31481 26364 31493 26367
rect 31205 26327 31263 26333
rect 31312 26336 31493 26364
rect 31312 26296 31340 26336
rect 31481 26333 31493 26336
rect 31527 26333 31539 26367
rect 31481 26327 31539 26333
rect 31570 26324 31576 26376
rect 31628 26324 31634 26376
rect 29748 26268 31340 26296
rect 31386 26256 31392 26308
rect 31444 26256 31450 26308
rect 32858 26256 32864 26308
rect 32916 26256 32922 26308
rect 33042 26256 33048 26308
rect 33100 26296 33106 26308
rect 33321 26299 33379 26305
rect 33321 26296 33333 26299
rect 33100 26268 33333 26296
rect 33100 26256 33106 26268
rect 33321 26265 33333 26268
rect 33367 26265 33379 26299
rect 33321 26259 33379 26265
rect 30101 26231 30159 26237
rect 30101 26228 30113 26231
rect 29656 26200 30113 26228
rect 28721 26191 28779 26197
rect 30101 26197 30113 26200
rect 30147 26197 30159 26231
rect 30101 26191 30159 26197
rect 30466 26188 30472 26240
rect 30524 26188 30530 26240
rect 31757 26231 31815 26237
rect 31757 26197 31769 26231
rect 31803 26228 31815 26231
rect 32306 26228 32312 26240
rect 31803 26200 32312 26228
rect 31803 26197 31815 26200
rect 31757 26191 31815 26197
rect 32306 26188 32312 26200
rect 32364 26188 32370 26240
rect 1104 26138 34840 26160
rect 1104 26086 9344 26138
rect 9396 26086 9408 26138
rect 9460 26086 9472 26138
rect 9524 26086 9536 26138
rect 9588 26086 9600 26138
rect 9652 26086 17738 26138
rect 17790 26086 17802 26138
rect 17854 26086 17866 26138
rect 17918 26086 17930 26138
rect 17982 26086 17994 26138
rect 18046 26086 26132 26138
rect 26184 26086 26196 26138
rect 26248 26086 26260 26138
rect 26312 26086 26324 26138
rect 26376 26086 26388 26138
rect 26440 26086 34526 26138
rect 34578 26086 34590 26138
rect 34642 26086 34654 26138
rect 34706 26086 34718 26138
rect 34770 26086 34782 26138
rect 34834 26086 34840 26138
rect 1104 26064 34840 26086
rect 3418 25984 3424 26036
rect 3476 26024 3482 26036
rect 3789 26027 3847 26033
rect 3789 26024 3801 26027
rect 3476 25996 3801 26024
rect 3476 25984 3482 25996
rect 3789 25993 3801 25996
rect 3835 25993 3847 26027
rect 3789 25987 3847 25993
rect 3970 25984 3976 26036
rect 4028 25984 4034 26036
rect 7190 25984 7196 26036
rect 7248 26024 7254 26036
rect 7377 26027 7435 26033
rect 7377 26024 7389 26027
rect 7248 25996 7389 26024
rect 7248 25984 7254 25996
rect 7377 25993 7389 25996
rect 7423 25993 7435 26027
rect 7377 25987 7435 25993
rect 7466 25984 7472 26036
rect 7524 25984 7530 26036
rect 20990 25984 20996 26036
rect 21048 26024 21054 26036
rect 21821 26027 21879 26033
rect 21821 26024 21833 26027
rect 21048 25996 21833 26024
rect 21048 25984 21054 25996
rect 21821 25993 21833 25996
rect 21867 25993 21879 26027
rect 21821 25987 21879 25993
rect 22189 26027 22247 26033
rect 22189 25993 22201 26027
rect 22235 26024 22247 26027
rect 23106 26024 23112 26036
rect 22235 25996 23112 26024
rect 22235 25993 22247 25996
rect 22189 25987 22247 25993
rect 23106 25984 23112 25996
rect 23164 25984 23170 26036
rect 25041 26027 25099 26033
rect 23308 25996 23796 26024
rect 5353 25959 5411 25965
rect 5353 25925 5365 25959
rect 5399 25956 5411 25959
rect 5534 25956 5540 25968
rect 5399 25928 5540 25956
rect 5399 25925 5411 25928
rect 5353 25919 5411 25925
rect 4154 25848 4160 25900
rect 4212 25888 4218 25900
rect 4341 25891 4399 25897
rect 4341 25888 4353 25891
rect 4212 25860 4353 25888
rect 4212 25848 4218 25860
rect 4341 25857 4353 25860
rect 4387 25857 4399 25891
rect 4341 25851 4399 25857
rect 4985 25891 5043 25897
rect 4985 25857 4997 25891
rect 5031 25888 5043 25891
rect 5368 25888 5396 25919
rect 5534 25916 5540 25928
rect 5592 25916 5598 25968
rect 6914 25916 6920 25968
rect 6972 25956 6978 25968
rect 7009 25959 7067 25965
rect 7009 25956 7021 25959
rect 6972 25928 7021 25956
rect 6972 25916 6978 25928
rect 7009 25925 7021 25928
rect 7055 25925 7067 25959
rect 7009 25919 7067 25925
rect 5718 25888 5724 25900
rect 5031 25860 5396 25888
rect 5460 25860 5724 25888
rect 5031 25857 5043 25860
rect 4985 25851 5043 25857
rect 4706 25780 4712 25832
rect 4764 25780 4770 25832
rect 4801 25823 4859 25829
rect 4801 25789 4813 25823
rect 4847 25789 4859 25823
rect 4801 25783 4859 25789
rect 4893 25823 4951 25829
rect 4893 25789 4905 25823
rect 4939 25820 4951 25823
rect 5460 25820 5488 25860
rect 5718 25848 5724 25860
rect 5776 25888 5782 25900
rect 5813 25891 5871 25897
rect 5813 25888 5825 25891
rect 5776 25860 5825 25888
rect 5776 25848 5782 25860
rect 5813 25857 5825 25860
rect 5859 25857 5871 25891
rect 5813 25851 5871 25857
rect 6549 25891 6607 25897
rect 6549 25857 6561 25891
rect 6595 25888 6607 25891
rect 7484 25888 7512 25984
rect 23308 25968 23336 25996
rect 12066 25916 12072 25968
rect 12124 25956 12130 25968
rect 12345 25959 12403 25965
rect 12345 25956 12357 25959
rect 12124 25928 12357 25956
rect 12124 25916 12130 25928
rect 12345 25925 12357 25928
rect 12391 25925 12403 25959
rect 12345 25919 12403 25925
rect 23290 25916 23296 25968
rect 23348 25916 23354 25968
rect 23385 25959 23443 25965
rect 23385 25925 23397 25959
rect 23431 25956 23443 25959
rect 23658 25956 23664 25968
rect 23431 25928 23664 25956
rect 23431 25925 23443 25928
rect 23385 25919 23443 25925
rect 23658 25916 23664 25928
rect 23716 25916 23722 25968
rect 23768 25956 23796 25996
rect 25041 25993 25053 26027
rect 25087 26024 25099 26027
rect 25498 26024 25504 26036
rect 25087 25996 25504 26024
rect 25087 25993 25099 25996
rect 25041 25987 25099 25993
rect 25498 25984 25504 25996
rect 25556 25984 25562 26036
rect 30377 26027 30435 26033
rect 30377 25993 30389 26027
rect 30423 26024 30435 26027
rect 30466 26024 30472 26036
rect 30423 25996 30472 26024
rect 30423 25993 30435 25996
rect 30377 25987 30435 25993
rect 30466 25984 30472 25996
rect 30524 25984 30530 26036
rect 32125 26027 32183 26033
rect 32125 25993 32137 26027
rect 32171 26024 32183 26027
rect 33042 26024 33048 26036
rect 32171 25996 33048 26024
rect 32171 25993 32183 25996
rect 32125 25987 32183 25993
rect 33042 25984 33048 25996
rect 33100 25984 33106 26036
rect 26329 25959 26387 25965
rect 26329 25956 26341 25959
rect 23768 25928 23874 25956
rect 24688 25928 26341 25956
rect 24688 25900 24716 25928
rect 26329 25925 26341 25928
rect 26375 25956 26387 25959
rect 28994 25956 29000 25968
rect 26375 25928 29000 25956
rect 26375 25925 26387 25928
rect 26329 25919 26387 25925
rect 28994 25916 29000 25928
rect 29052 25916 29058 25968
rect 7561 25891 7619 25897
rect 7561 25888 7573 25891
rect 6595 25860 6960 25888
rect 7484 25860 7573 25888
rect 6595 25857 6607 25860
rect 6549 25851 6607 25857
rect 6932 25832 6960 25860
rect 7561 25857 7573 25860
rect 7607 25857 7619 25891
rect 14369 25891 14427 25897
rect 14369 25888 14381 25891
rect 7561 25851 7619 25857
rect 12728 25860 14381 25888
rect 4939 25792 5488 25820
rect 5629 25823 5687 25829
rect 4939 25789 4951 25792
rect 4893 25783 4951 25789
rect 5629 25789 5641 25823
rect 5675 25789 5687 25823
rect 6641 25823 6699 25829
rect 6641 25820 6653 25823
rect 5629 25783 5687 25789
rect 6012 25792 6653 25820
rect 4816 25752 4844 25783
rect 4982 25752 4988 25764
rect 4816 25724 4988 25752
rect 4982 25712 4988 25724
rect 5040 25752 5046 25764
rect 5644 25752 5672 25783
rect 6012 25761 6040 25792
rect 6641 25789 6653 25792
rect 6687 25789 6699 25823
rect 6641 25783 6699 25789
rect 6914 25780 6920 25832
rect 6972 25780 6978 25832
rect 8757 25823 8815 25829
rect 8757 25820 8769 25823
rect 7852 25792 8769 25820
rect 5040 25724 5672 25752
rect 5997 25755 6055 25761
rect 5040 25712 5046 25724
rect 5997 25721 6009 25755
rect 6043 25721 6055 25755
rect 5997 25715 6055 25721
rect 7852 25696 7880 25792
rect 8757 25789 8769 25792
rect 8803 25789 8815 25823
rect 8757 25783 8815 25789
rect 12728 25764 12756 25860
rect 14369 25857 14381 25860
rect 14415 25888 14427 25891
rect 14734 25888 14740 25900
rect 14415 25860 14740 25888
rect 14415 25857 14427 25860
rect 14369 25851 14427 25857
rect 14734 25848 14740 25860
rect 14792 25848 14798 25900
rect 14826 25848 14832 25900
rect 14884 25848 14890 25900
rect 19978 25848 19984 25900
rect 20036 25888 20042 25900
rect 20990 25888 20996 25900
rect 20036 25860 20996 25888
rect 20036 25848 20042 25860
rect 20990 25848 20996 25860
rect 21048 25888 21054 25900
rect 21048 25860 22508 25888
rect 21048 25848 21054 25860
rect 14185 25823 14243 25829
rect 14185 25789 14197 25823
rect 14231 25820 14243 25823
rect 14844 25820 14872 25848
rect 14231 25792 14872 25820
rect 14231 25789 14243 25792
rect 14185 25783 14243 25789
rect 21634 25780 21640 25832
rect 21692 25820 21698 25832
rect 22480 25829 22508 25860
rect 23106 25848 23112 25900
rect 23164 25848 23170 25900
rect 24670 25848 24676 25900
rect 24728 25848 24734 25900
rect 25317 25891 25375 25897
rect 25317 25857 25329 25891
rect 25363 25857 25375 25891
rect 25317 25851 25375 25857
rect 22281 25823 22339 25829
rect 22281 25820 22293 25823
rect 21692 25792 22293 25820
rect 21692 25780 21698 25792
rect 22281 25789 22293 25792
rect 22327 25789 22339 25823
rect 22281 25783 22339 25789
rect 22465 25823 22523 25829
rect 22465 25789 22477 25823
rect 22511 25820 22523 25823
rect 22922 25820 22928 25832
rect 22511 25792 22928 25820
rect 22511 25789 22523 25792
rect 22465 25783 22523 25789
rect 22922 25780 22928 25792
rect 22980 25820 22986 25832
rect 22980 25792 24440 25820
rect 22980 25780 22986 25792
rect 12161 25755 12219 25761
rect 12161 25721 12173 25755
rect 12207 25752 12219 25755
rect 12526 25752 12532 25764
rect 12207 25724 12532 25752
rect 12207 25721 12219 25724
rect 12161 25715 12219 25721
rect 12526 25712 12532 25724
rect 12584 25712 12590 25764
rect 12710 25712 12716 25764
rect 12768 25712 12774 25764
rect 24412 25752 24440 25792
rect 25038 25780 25044 25832
rect 25096 25780 25102 25832
rect 25332 25820 25360 25851
rect 25590 25848 25596 25900
rect 25648 25848 25654 25900
rect 26421 25891 26479 25897
rect 26421 25857 26433 25891
rect 26467 25888 26479 25891
rect 26510 25888 26516 25900
rect 26467 25860 26516 25888
rect 26467 25857 26479 25860
rect 26421 25851 26479 25857
rect 26510 25848 26516 25860
rect 26568 25848 26574 25900
rect 26602 25848 26608 25900
rect 26660 25888 26666 25900
rect 27065 25891 27123 25897
rect 27065 25888 27077 25891
rect 26660 25860 27077 25888
rect 26660 25848 26666 25860
rect 27065 25857 27077 25860
rect 27111 25888 27123 25891
rect 27154 25888 27160 25900
rect 27111 25860 27160 25888
rect 27111 25857 27123 25860
rect 27065 25851 27123 25857
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 27246 25848 27252 25900
rect 27304 25848 27310 25900
rect 27433 25891 27491 25897
rect 27433 25857 27445 25891
rect 27479 25857 27491 25891
rect 27433 25851 27491 25857
rect 26620 25820 26648 25848
rect 25332 25792 26648 25820
rect 26789 25823 26847 25829
rect 26789 25789 26801 25823
rect 26835 25820 26847 25823
rect 27448 25820 27476 25851
rect 28166 25848 28172 25900
rect 28224 25848 28230 25900
rect 30006 25848 30012 25900
rect 30064 25848 30070 25900
rect 32306 25848 32312 25900
rect 32364 25848 32370 25900
rect 32490 25848 32496 25900
rect 32548 25848 32554 25900
rect 32582 25848 32588 25900
rect 32640 25848 32646 25900
rect 26835 25792 27476 25820
rect 26835 25789 26847 25792
rect 26789 25783 26847 25789
rect 25225 25755 25283 25761
rect 25225 25752 25237 25755
rect 24412 25724 25237 25752
rect 25225 25721 25237 25724
rect 25271 25752 25283 25755
rect 25682 25752 25688 25764
rect 25271 25724 25688 25752
rect 25271 25721 25283 25724
rect 25225 25715 25283 25721
rect 25682 25712 25688 25724
rect 25740 25712 25746 25764
rect 27154 25712 27160 25764
rect 27212 25752 27218 25764
rect 27249 25755 27307 25761
rect 27249 25752 27261 25755
rect 27212 25724 27261 25752
rect 27212 25712 27218 25724
rect 27249 25721 27261 25724
rect 27295 25752 27307 25755
rect 28184 25752 28212 25848
rect 30101 25823 30159 25829
rect 30101 25789 30113 25823
rect 30147 25820 30159 25823
rect 30650 25820 30656 25832
rect 30147 25792 30656 25820
rect 30147 25789 30159 25792
rect 30101 25783 30159 25789
rect 30650 25780 30656 25792
rect 30708 25780 30714 25832
rect 27295 25724 28212 25752
rect 27295 25721 27307 25724
rect 27249 25715 27307 25721
rect 3973 25687 4031 25693
rect 3973 25653 3985 25687
rect 4019 25684 4031 25687
rect 4525 25687 4583 25693
rect 4525 25684 4537 25687
rect 4019 25656 4537 25684
rect 4019 25653 4031 25656
rect 3973 25647 4031 25653
rect 4525 25653 4537 25656
rect 4571 25653 4583 25687
rect 4525 25647 4583 25653
rect 5810 25644 5816 25696
rect 5868 25644 5874 25696
rect 5902 25644 5908 25696
rect 5960 25684 5966 25696
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 5960 25656 6377 25684
rect 5960 25644 5966 25656
rect 6365 25653 6377 25656
rect 6411 25653 6423 25687
rect 6365 25647 6423 25653
rect 6917 25687 6975 25693
rect 6917 25653 6929 25687
rect 6963 25684 6975 25687
rect 7006 25684 7012 25696
rect 6963 25656 7012 25684
rect 6963 25653 6975 25656
rect 6917 25647 6975 25653
rect 7006 25644 7012 25656
rect 7064 25684 7070 25696
rect 7190 25684 7196 25696
rect 7064 25656 7196 25684
rect 7064 25644 7070 25656
rect 7190 25644 7196 25656
rect 7248 25644 7254 25696
rect 7834 25644 7840 25696
rect 7892 25644 7898 25696
rect 9122 25644 9128 25696
rect 9180 25684 9186 25696
rect 9401 25687 9459 25693
rect 9401 25684 9413 25687
rect 9180 25656 9413 25684
rect 9180 25644 9186 25656
rect 9401 25653 9413 25656
rect 9447 25653 9459 25687
rect 9401 25647 9459 25653
rect 9950 25644 9956 25696
rect 10008 25684 10014 25696
rect 12345 25687 12403 25693
rect 12345 25684 12357 25687
rect 10008 25656 12357 25684
rect 10008 25644 10014 25656
rect 12345 25653 12357 25656
rect 12391 25653 12403 25687
rect 12345 25647 12403 25653
rect 14550 25644 14556 25696
rect 14608 25644 14614 25696
rect 24854 25644 24860 25696
rect 24912 25644 24918 25696
rect 25314 25644 25320 25696
rect 25372 25684 25378 25696
rect 27709 25687 27767 25693
rect 27709 25684 27721 25687
rect 25372 25656 27721 25684
rect 25372 25644 25378 25656
rect 27709 25653 27721 25656
rect 27755 25684 27767 25687
rect 28442 25684 28448 25696
rect 27755 25656 28448 25684
rect 27755 25653 27767 25656
rect 27709 25647 27767 25653
rect 28442 25644 28448 25656
rect 28500 25644 28506 25696
rect 1104 25594 34684 25616
rect 1104 25542 5147 25594
rect 5199 25542 5211 25594
rect 5263 25542 5275 25594
rect 5327 25542 5339 25594
rect 5391 25542 5403 25594
rect 5455 25542 13541 25594
rect 13593 25542 13605 25594
rect 13657 25542 13669 25594
rect 13721 25542 13733 25594
rect 13785 25542 13797 25594
rect 13849 25542 21935 25594
rect 21987 25542 21999 25594
rect 22051 25542 22063 25594
rect 22115 25542 22127 25594
rect 22179 25542 22191 25594
rect 22243 25542 30329 25594
rect 30381 25542 30393 25594
rect 30445 25542 30457 25594
rect 30509 25542 30521 25594
rect 30573 25542 30585 25594
rect 30637 25542 34684 25594
rect 1104 25520 34684 25542
rect 4154 25440 4160 25492
rect 4212 25480 4218 25492
rect 4617 25483 4675 25489
rect 4617 25480 4629 25483
rect 4212 25452 4629 25480
rect 4212 25440 4218 25452
rect 4617 25449 4629 25452
rect 4663 25449 4675 25483
rect 4617 25443 4675 25449
rect 4801 25483 4859 25489
rect 4801 25449 4813 25483
rect 4847 25480 4859 25483
rect 5534 25480 5540 25492
rect 4847 25452 5540 25480
rect 4847 25449 4859 25452
rect 4801 25443 4859 25449
rect 5534 25440 5540 25452
rect 5592 25440 5598 25492
rect 7190 25440 7196 25492
rect 7248 25480 7254 25492
rect 7248 25452 7604 25480
rect 7248 25440 7254 25452
rect 4430 25304 4436 25356
rect 4488 25344 4494 25356
rect 4488 25316 5028 25344
rect 4488 25304 4494 25316
rect 3237 25279 3295 25285
rect 3237 25245 3249 25279
rect 3283 25276 3295 25279
rect 3326 25276 3332 25288
rect 3283 25248 3332 25276
rect 3283 25245 3295 25248
rect 3237 25239 3295 25245
rect 3326 25236 3332 25248
rect 3384 25236 3390 25288
rect 3418 25236 3424 25288
rect 3476 25236 3482 25288
rect 3513 25279 3571 25285
rect 3513 25245 3525 25279
rect 3559 25276 3571 25279
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 3559 25248 3801 25276
rect 3559 25245 3571 25248
rect 3513 25239 3571 25245
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 5000 25220 5028 25316
rect 5810 25304 5816 25356
rect 5868 25344 5874 25356
rect 7190 25344 7196 25356
rect 5868 25316 7196 25344
rect 5868 25304 5874 25316
rect 6656 25285 6684 25316
rect 7190 25304 7196 25316
rect 7248 25304 7254 25356
rect 7576 25344 7604 25452
rect 7834 25440 7840 25492
rect 7892 25440 7898 25492
rect 8662 25440 8668 25492
rect 8720 25480 8726 25492
rect 9033 25483 9091 25489
rect 9033 25480 9045 25483
rect 8720 25452 9045 25480
rect 8720 25440 8726 25452
rect 9033 25449 9045 25452
rect 9079 25449 9091 25483
rect 9033 25443 9091 25449
rect 9214 25440 9220 25492
rect 9272 25440 9278 25492
rect 15749 25483 15807 25489
rect 15749 25449 15761 25483
rect 15795 25480 15807 25483
rect 16025 25483 16083 25489
rect 16025 25480 16037 25483
rect 15795 25452 16037 25480
rect 15795 25449 15807 25452
rect 15749 25443 15807 25449
rect 16025 25449 16037 25452
rect 16071 25449 16083 25483
rect 16025 25443 16083 25449
rect 20714 25440 20720 25492
rect 20772 25480 20778 25492
rect 20993 25483 21051 25489
rect 20993 25480 21005 25483
rect 20772 25452 21005 25480
rect 20772 25440 20778 25452
rect 20993 25449 21005 25452
rect 21039 25449 21051 25483
rect 20993 25443 21051 25449
rect 26510 25440 26516 25492
rect 26568 25440 26574 25492
rect 28810 25440 28816 25492
rect 28868 25480 28874 25492
rect 29181 25483 29239 25489
rect 28868 25452 28994 25480
rect 28868 25440 28874 25452
rect 8680 25344 8708 25440
rect 9125 25415 9183 25421
rect 9125 25381 9137 25415
rect 9171 25381 9183 25415
rect 9232 25412 9260 25440
rect 9232 25384 9352 25412
rect 9125 25375 9183 25381
rect 9140 25344 9168 25375
rect 9324 25353 9352 25384
rect 10888 25384 12434 25412
rect 7576 25316 8708 25344
rect 8772 25316 9168 25344
rect 9217 25347 9275 25353
rect 7576 25285 7604 25316
rect 6641 25279 6699 25285
rect 6641 25245 6653 25279
rect 6687 25245 6699 25279
rect 6641 25239 6699 25245
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 7561 25279 7619 25285
rect 7561 25276 7573 25279
rect 6963 25248 7573 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 7561 25245 7573 25248
rect 7607 25245 7619 25279
rect 7742 25276 7748 25288
rect 7561 25239 7619 25245
rect 7668 25248 7748 25276
rect 4982 25168 4988 25220
rect 5040 25168 5046 25220
rect 7377 25211 7435 25217
rect 7377 25208 7389 25211
rect 6932 25180 7389 25208
rect 6932 25152 6960 25180
rect 7377 25177 7389 25180
rect 7423 25208 7435 25211
rect 7668 25208 7696 25248
rect 7742 25236 7748 25248
rect 7800 25276 7806 25288
rect 7929 25279 7987 25285
rect 7929 25276 7941 25279
rect 7800 25248 7941 25276
rect 7800 25236 7806 25248
rect 7929 25245 7941 25248
rect 7975 25245 7987 25279
rect 8772 25276 8800 25316
rect 9217 25313 9229 25347
rect 9263 25313 9275 25347
rect 9217 25307 9275 25313
rect 9309 25347 9367 25353
rect 9309 25313 9321 25347
rect 9355 25313 9367 25347
rect 9309 25307 9367 25313
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 7929 25239 7987 25245
rect 8496 25248 8800 25276
rect 8864 25248 8953 25276
rect 7423 25180 7696 25208
rect 7837 25211 7895 25217
rect 7423 25177 7435 25180
rect 7377 25171 7435 25177
rect 7837 25177 7849 25211
rect 7883 25208 7895 25211
rect 8496 25208 8524 25248
rect 8864 25208 8892 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 9232 25276 9260 25307
rect 10888 25288 10916 25384
rect 11057 25347 11115 25353
rect 11057 25313 11069 25347
rect 11103 25344 11115 25347
rect 11103 25316 11744 25344
rect 11103 25313 11115 25316
rect 11057 25307 11115 25313
rect 11716 25288 11744 25316
rect 10870 25276 10876 25288
rect 9232 25248 9352 25276
rect 10718 25248 10876 25276
rect 8941 25239 8999 25245
rect 7883 25180 8524 25208
rect 8588 25180 8892 25208
rect 7883 25177 7895 25180
rect 7837 25171 7895 25177
rect 2866 25100 2872 25152
rect 2924 25140 2930 25152
rect 4798 25149 4804 25152
rect 3053 25143 3111 25149
rect 3053 25140 3065 25143
rect 2924 25112 3065 25140
rect 2924 25100 2930 25112
rect 3053 25109 3065 25112
rect 3099 25109 3111 25143
rect 3053 25103 3111 25109
rect 4785 25143 4804 25149
rect 4785 25109 4797 25143
rect 4785 25103 4804 25109
rect 4798 25100 4804 25103
rect 4856 25100 4862 25152
rect 6454 25100 6460 25152
rect 6512 25100 6518 25152
rect 6825 25143 6883 25149
rect 6825 25109 6837 25143
rect 6871 25140 6883 25143
rect 6914 25140 6920 25152
rect 6871 25112 6920 25140
rect 6871 25109 6883 25112
rect 6825 25103 6883 25109
rect 6914 25100 6920 25112
rect 6972 25100 6978 25152
rect 7006 25100 7012 25152
rect 7064 25100 7070 25152
rect 7190 25149 7196 25152
rect 7177 25143 7196 25149
rect 7177 25109 7189 25143
rect 7177 25103 7196 25109
rect 7190 25100 7196 25103
rect 7248 25100 7254 25152
rect 8588 25149 8616 25180
rect 7653 25143 7711 25149
rect 7653 25109 7665 25143
rect 7699 25140 7711 25143
rect 8573 25143 8631 25149
rect 8573 25140 8585 25143
rect 7699 25112 8585 25140
rect 7699 25109 7711 25112
rect 7653 25103 7711 25109
rect 8573 25109 8585 25112
rect 8619 25109 8631 25143
rect 8573 25103 8631 25109
rect 9030 25100 9036 25152
rect 9088 25140 9094 25152
rect 9324 25140 9352 25248
rect 10870 25236 10876 25248
rect 10928 25236 10934 25288
rect 11330 25236 11336 25288
rect 11388 25236 11394 25288
rect 11698 25236 11704 25288
rect 11756 25236 11762 25288
rect 11885 25279 11943 25285
rect 11885 25245 11897 25279
rect 11931 25245 11943 25279
rect 11885 25239 11943 25245
rect 9585 25211 9643 25217
rect 9585 25177 9597 25211
rect 9631 25208 9643 25211
rect 9858 25208 9864 25220
rect 9631 25180 9864 25208
rect 9631 25177 9643 25180
rect 9585 25171 9643 25177
rect 9858 25168 9864 25180
rect 9916 25168 9922 25220
rect 11348 25208 11376 25236
rect 11900 25208 11928 25239
rect 11974 25236 11980 25288
rect 12032 25276 12038 25288
rect 12069 25279 12127 25285
rect 12069 25276 12081 25279
rect 12032 25248 12081 25276
rect 12032 25236 12038 25248
rect 12069 25245 12081 25248
rect 12115 25276 12127 25279
rect 12158 25276 12164 25288
rect 12115 25248 12164 25276
rect 12115 25245 12127 25248
rect 12069 25239 12127 25245
rect 12158 25236 12164 25248
rect 12216 25236 12222 25288
rect 12406 25276 12434 25384
rect 15580 25316 16528 25344
rect 12406 25248 12558 25276
rect 13906 25236 13912 25288
rect 13964 25236 13970 25288
rect 15580 25285 15608 25316
rect 16500 25288 16528 25316
rect 16758 25304 16764 25356
rect 16816 25344 16822 25356
rect 17313 25347 17371 25353
rect 17313 25344 17325 25347
rect 16816 25316 17325 25344
rect 16816 25304 16822 25316
rect 17313 25313 17325 25316
rect 17359 25344 17371 25347
rect 19245 25347 19303 25353
rect 19245 25344 19257 25347
rect 17359 25316 19257 25344
rect 17359 25313 17371 25316
rect 17313 25307 17371 25313
rect 19245 25313 19257 25316
rect 19291 25313 19303 25347
rect 26528 25344 26556 25440
rect 27157 25415 27215 25421
rect 27157 25381 27169 25415
rect 27203 25412 27215 25415
rect 27798 25412 27804 25424
rect 27203 25384 27804 25412
rect 27203 25381 27215 25384
rect 27157 25375 27215 25381
rect 27798 25372 27804 25384
rect 27856 25372 27862 25424
rect 19245 25307 19303 25313
rect 26252 25316 27016 25344
rect 15565 25279 15623 25285
rect 15565 25245 15577 25279
rect 15611 25245 15623 25279
rect 16301 25279 16359 25285
rect 16301 25276 16313 25279
rect 15565 25239 15623 25245
rect 15672 25248 16313 25276
rect 12250 25208 12256 25220
rect 11348 25180 12256 25208
rect 12250 25168 12256 25180
rect 12308 25168 12314 25220
rect 13630 25168 13636 25220
rect 13688 25168 13694 25220
rect 14550 25168 14556 25220
rect 14608 25208 14614 25220
rect 15381 25211 15439 25217
rect 15381 25208 15393 25211
rect 14608 25180 15393 25208
rect 14608 25168 14614 25180
rect 15381 25177 15393 25180
rect 15427 25208 15439 25211
rect 15672 25208 15700 25248
rect 16301 25245 16313 25248
rect 16347 25245 16359 25279
rect 16301 25239 16359 25245
rect 16482 25236 16488 25288
rect 16540 25236 16546 25288
rect 26252 25285 26280 25316
rect 26145 25279 26203 25285
rect 26145 25245 26157 25279
rect 26191 25245 26203 25279
rect 26145 25239 26203 25245
rect 26237 25279 26295 25285
rect 26237 25245 26249 25279
rect 26283 25245 26295 25279
rect 26602 25276 26608 25288
rect 26237 25239 26295 25245
rect 26344 25248 26608 25276
rect 15427 25180 15700 25208
rect 15427 25177 15439 25180
rect 15381 25171 15439 25177
rect 16206 25168 16212 25220
rect 16264 25208 16270 25220
rect 16574 25208 16580 25220
rect 16264 25180 16580 25208
rect 16264 25168 16270 25180
rect 16574 25168 16580 25180
rect 16632 25168 16638 25220
rect 16669 25211 16727 25217
rect 16669 25177 16681 25211
rect 16715 25208 16727 25211
rect 16942 25208 16948 25220
rect 16715 25180 16948 25208
rect 16715 25177 16727 25180
rect 16669 25171 16727 25177
rect 9950 25140 9956 25152
rect 9088 25112 9956 25140
rect 9088 25100 9094 25112
rect 9950 25100 9956 25112
rect 10008 25100 10014 25152
rect 11146 25100 11152 25152
rect 11204 25100 11210 25152
rect 11238 25100 11244 25152
rect 11296 25140 11302 25152
rect 11977 25143 12035 25149
rect 11977 25140 11989 25143
rect 11296 25112 11989 25140
rect 11296 25100 11302 25112
rect 11977 25109 11989 25112
rect 12023 25109 12035 25143
rect 11977 25103 12035 25109
rect 12158 25100 12164 25152
rect 12216 25100 12222 25152
rect 15838 25100 15844 25152
rect 15896 25100 15902 25152
rect 16009 25143 16067 25149
rect 16009 25109 16021 25143
rect 16055 25140 16067 25143
rect 16684 25140 16712 25171
rect 16942 25168 16948 25180
rect 17000 25168 17006 25220
rect 17589 25211 17647 25217
rect 17589 25177 17601 25211
rect 17635 25177 17647 25211
rect 18814 25180 19472 25208
rect 17589 25171 17647 25177
rect 16055 25112 16712 25140
rect 17604 25140 17632 25171
rect 18230 25140 18236 25152
rect 17604 25112 18236 25140
rect 16055 25109 16067 25112
rect 16009 25103 16067 25109
rect 18230 25100 18236 25112
rect 18288 25100 18294 25152
rect 19058 25100 19064 25152
rect 19116 25100 19122 25152
rect 19444 25140 19472 25180
rect 19518 25168 19524 25220
rect 19576 25168 19582 25220
rect 19978 25208 19984 25220
rect 19628 25180 19984 25208
rect 19628 25140 19656 25180
rect 19978 25168 19984 25180
rect 20036 25168 20042 25220
rect 20070 25168 20076 25220
rect 20128 25168 20134 25220
rect 23474 25168 23480 25220
rect 23532 25208 23538 25220
rect 24670 25208 24676 25220
rect 23532 25180 24676 25208
rect 23532 25168 23538 25180
rect 24670 25168 24676 25180
rect 24728 25168 24734 25220
rect 25406 25168 25412 25220
rect 25464 25168 25470 25220
rect 26160 25208 26188 25239
rect 26344 25208 26372 25248
rect 26602 25236 26608 25248
rect 26660 25236 26666 25288
rect 26988 25285 27016 25316
rect 26973 25279 27031 25285
rect 26973 25245 26985 25279
rect 27019 25245 27031 25279
rect 26973 25239 27031 25245
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25245 28779 25279
rect 28966 25276 28994 25452
rect 29181 25449 29193 25483
rect 29227 25480 29239 25483
rect 29227 25452 29776 25480
rect 29227 25449 29239 25452
rect 29181 25443 29239 25449
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 28966 25248 29561 25276
rect 28721 25239 28779 25245
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29748 25276 29776 25452
rect 29822 25440 29828 25492
rect 29880 25440 29886 25492
rect 30006 25440 30012 25492
rect 30064 25480 30070 25492
rect 30193 25483 30251 25489
rect 30193 25480 30205 25483
rect 30064 25452 30205 25480
rect 30064 25440 30070 25452
rect 30193 25449 30205 25452
rect 30239 25449 30251 25483
rect 30193 25443 30251 25449
rect 30208 25344 30236 25443
rect 32582 25440 32588 25492
rect 32640 25480 32646 25492
rect 32769 25483 32827 25489
rect 32769 25480 32781 25483
rect 32640 25452 32781 25480
rect 32640 25440 32646 25452
rect 32769 25449 32781 25452
rect 32815 25449 32827 25483
rect 32769 25443 32827 25449
rect 30208 25316 30512 25344
rect 30484 25285 30512 25316
rect 31386 25304 31392 25356
rect 31444 25344 31450 25356
rect 32033 25347 32091 25353
rect 32033 25344 32045 25347
rect 31444 25316 32045 25344
rect 31444 25304 31450 25316
rect 32033 25313 32045 25316
rect 32079 25313 32091 25347
rect 32033 25307 32091 25313
rect 33410 25304 33416 25356
rect 33468 25304 33474 25356
rect 30101 25279 30159 25285
rect 30101 25276 30113 25279
rect 29748 25248 30113 25276
rect 29549 25239 29607 25245
rect 30101 25245 30113 25248
rect 30147 25245 30159 25279
rect 30285 25279 30343 25285
rect 30285 25276 30297 25279
rect 30101 25239 30159 25245
rect 30208 25248 30297 25276
rect 26160 25180 26372 25208
rect 26421 25211 26479 25217
rect 26421 25177 26433 25211
rect 26467 25208 26479 25211
rect 27433 25211 27491 25217
rect 27433 25208 27445 25211
rect 26467 25180 27445 25208
rect 26467 25177 26479 25180
rect 26421 25171 26479 25177
rect 27433 25177 27445 25180
rect 27479 25177 27491 25211
rect 28736 25208 28764 25239
rect 29178 25208 29184 25220
rect 28736 25180 29184 25208
rect 27433 25171 27491 25177
rect 29178 25168 29184 25180
rect 29236 25208 29242 25220
rect 29822 25208 29828 25220
rect 29236 25180 29828 25208
rect 29236 25168 29242 25180
rect 29822 25168 29828 25180
rect 29880 25168 29886 25220
rect 30208 25152 30236 25248
rect 30285 25245 30297 25248
rect 30331 25245 30343 25279
rect 30285 25239 30343 25245
rect 30469 25279 30527 25285
rect 30469 25245 30481 25279
rect 30515 25245 30527 25279
rect 30469 25239 30527 25245
rect 30653 25279 30711 25285
rect 30653 25245 30665 25279
rect 30699 25276 30711 25279
rect 31846 25276 31852 25288
rect 30699 25248 31852 25276
rect 30699 25245 30711 25248
rect 30653 25239 30711 25245
rect 31846 25236 31852 25248
rect 31904 25276 31910 25288
rect 32125 25279 32183 25285
rect 32125 25276 32137 25279
rect 31904 25248 32137 25276
rect 31904 25236 31910 25248
rect 32125 25245 32137 25248
rect 32171 25245 32183 25279
rect 32125 25239 32183 25245
rect 32582 25168 32588 25220
rect 32640 25208 32646 25220
rect 33229 25211 33287 25217
rect 33229 25208 33241 25211
rect 32640 25180 33241 25208
rect 32640 25168 32646 25180
rect 33229 25177 33241 25180
rect 33275 25177 33287 25211
rect 33229 25171 33287 25177
rect 19444 25112 19656 25140
rect 26970 25100 26976 25152
rect 27028 25140 27034 25152
rect 27525 25143 27583 25149
rect 27525 25140 27537 25143
rect 27028 25112 27537 25140
rect 27028 25100 27034 25112
rect 27525 25109 27537 25112
rect 27571 25109 27583 25143
rect 27525 25103 27583 25109
rect 30009 25143 30067 25149
rect 30009 25109 30021 25143
rect 30055 25140 30067 25143
rect 30190 25140 30196 25152
rect 30055 25112 30196 25140
rect 30055 25109 30067 25112
rect 30009 25103 30067 25109
rect 30190 25100 30196 25112
rect 30248 25100 30254 25152
rect 30834 25100 30840 25152
rect 30892 25100 30898 25152
rect 32493 25143 32551 25149
rect 32493 25109 32505 25143
rect 32539 25140 32551 25143
rect 33137 25143 33195 25149
rect 33137 25140 33149 25143
rect 32539 25112 33149 25140
rect 32539 25109 32551 25112
rect 32493 25103 32551 25109
rect 33137 25109 33149 25112
rect 33183 25109 33195 25143
rect 33137 25103 33195 25109
rect 1104 25050 34840 25072
rect 1104 24998 9344 25050
rect 9396 24998 9408 25050
rect 9460 24998 9472 25050
rect 9524 24998 9536 25050
rect 9588 24998 9600 25050
rect 9652 24998 17738 25050
rect 17790 24998 17802 25050
rect 17854 24998 17866 25050
rect 17918 24998 17930 25050
rect 17982 24998 17994 25050
rect 18046 24998 26132 25050
rect 26184 24998 26196 25050
rect 26248 24998 26260 25050
rect 26312 24998 26324 25050
rect 26376 24998 26388 25050
rect 26440 24998 34526 25050
rect 34578 24998 34590 25050
rect 34642 24998 34654 25050
rect 34706 24998 34718 25050
rect 34770 24998 34782 25050
rect 34834 24998 34840 25050
rect 1104 24976 34840 24998
rect 3418 24896 3424 24948
rect 3476 24896 3482 24948
rect 3605 24939 3663 24945
rect 3605 24905 3617 24939
rect 3651 24936 3663 24939
rect 3881 24939 3939 24945
rect 3881 24936 3893 24939
rect 3651 24908 3893 24936
rect 3651 24905 3663 24908
rect 3605 24899 3663 24905
rect 3881 24905 3893 24908
rect 3927 24936 3939 24939
rect 4430 24936 4436 24948
rect 3927 24908 4436 24936
rect 3927 24905 3939 24908
rect 3881 24899 3939 24905
rect 4430 24896 4436 24908
rect 4488 24896 4494 24948
rect 4706 24896 4712 24948
rect 4764 24936 4770 24948
rect 4764 24908 5028 24936
rect 4764 24896 4770 24908
rect 3436 24800 3464 24896
rect 4798 24868 4804 24880
rect 3804 24840 4804 24868
rect 3804 24809 3832 24840
rect 4798 24828 4804 24840
rect 4856 24828 4862 24880
rect 5000 24868 5028 24908
rect 6454 24896 6460 24948
rect 6512 24936 6518 24948
rect 6549 24939 6607 24945
rect 6549 24936 6561 24939
rect 6512 24908 6561 24936
rect 6512 24896 6518 24908
rect 6549 24905 6561 24908
rect 6595 24905 6607 24939
rect 6549 24899 6607 24905
rect 7742 24896 7748 24948
rect 7800 24896 7806 24948
rect 9030 24936 9036 24948
rect 7852 24908 9036 24936
rect 7006 24868 7012 24880
rect 5000 24840 7012 24868
rect 3789 24803 3847 24809
rect 3789 24800 3801 24803
rect 1857 24735 1915 24741
rect 1857 24701 1869 24735
rect 1903 24701 1915 24735
rect 1857 24695 1915 24701
rect 2133 24735 2191 24741
rect 2133 24701 2145 24735
rect 2179 24732 2191 24735
rect 2866 24732 2872 24744
rect 2179 24704 2872 24732
rect 2179 24701 2191 24704
rect 2133 24695 2191 24701
rect 1872 24596 1900 24695
rect 2866 24692 2872 24704
rect 2924 24692 2930 24744
rect 3142 24596 3148 24608
rect 1872 24568 3148 24596
rect 3142 24556 3148 24568
rect 3200 24556 3206 24608
rect 3252 24596 3280 24786
rect 3436 24772 3801 24800
rect 3789 24769 3801 24772
rect 3835 24769 3847 24803
rect 3789 24763 3847 24769
rect 4065 24803 4123 24809
rect 4065 24769 4077 24803
rect 4111 24800 4123 24803
rect 4338 24800 4344 24812
rect 4111 24772 4344 24800
rect 4111 24769 4123 24772
rect 4065 24763 4123 24769
rect 4338 24760 4344 24772
rect 4396 24760 4402 24812
rect 5000 24809 5028 24840
rect 4985 24803 5043 24809
rect 4985 24769 4997 24803
rect 5031 24769 5043 24803
rect 4985 24763 5043 24769
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24800 5227 24803
rect 5718 24800 5724 24812
rect 5215 24772 5724 24800
rect 5215 24769 5227 24772
rect 5169 24763 5227 24769
rect 5718 24760 5724 24772
rect 5776 24760 5782 24812
rect 6932 24809 6960 24840
rect 7006 24828 7012 24840
rect 7064 24828 7070 24880
rect 6917 24803 6975 24809
rect 6917 24769 6929 24803
rect 6963 24769 6975 24803
rect 6917 24763 6975 24769
rect 3326 24692 3332 24744
rect 3384 24732 3390 24744
rect 7852 24732 7880 24908
rect 9030 24896 9036 24908
rect 9088 24896 9094 24948
rect 9214 24896 9220 24948
rect 9272 24896 9278 24948
rect 9858 24896 9864 24948
rect 9916 24936 9922 24948
rect 10229 24939 10287 24945
rect 10229 24936 10241 24939
rect 9916 24908 10241 24936
rect 9916 24896 9922 24908
rect 10229 24905 10241 24908
rect 10275 24905 10287 24939
rect 11146 24936 11152 24948
rect 10229 24899 10287 24905
rect 11072 24908 11152 24936
rect 9232 24868 9260 24896
rect 9232 24840 9536 24868
rect 9508 24809 9536 24840
rect 9493 24803 9551 24809
rect 3384 24704 4108 24732
rect 3384 24692 3390 24704
rect 4080 24673 4108 24704
rect 6840 24704 7880 24732
rect 8036 24772 8142 24800
rect 4065 24667 4123 24673
rect 4065 24633 4077 24667
rect 4111 24633 4123 24667
rect 4065 24627 4123 24633
rect 5626 24624 5632 24676
rect 5684 24664 5690 24676
rect 5684 24636 6592 24664
rect 5684 24624 5690 24636
rect 4522 24596 4528 24608
rect 3252 24568 4528 24596
rect 4522 24556 4528 24568
rect 4580 24556 4586 24608
rect 6362 24556 6368 24608
rect 6420 24556 6426 24608
rect 6564 24605 6592 24636
rect 6549 24599 6607 24605
rect 6549 24565 6561 24599
rect 6595 24596 6607 24599
rect 6840 24596 6868 24704
rect 8036 24664 8064 24772
rect 9493 24769 9505 24803
rect 9539 24769 9551 24803
rect 9493 24763 9551 24769
rect 10413 24803 10471 24809
rect 10413 24769 10425 24803
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 10689 24803 10747 24809
rect 10689 24769 10701 24803
rect 10735 24800 10747 24803
rect 11072 24800 11100 24908
rect 11146 24896 11152 24908
rect 11204 24896 11210 24948
rect 12066 24896 12072 24948
rect 12124 24896 12130 24948
rect 12250 24896 12256 24948
rect 12308 24936 12314 24948
rect 12361 24939 12419 24945
rect 12361 24936 12373 24939
rect 12308 24908 12373 24936
rect 12308 24896 12314 24908
rect 12361 24905 12373 24908
rect 12407 24905 12419 24939
rect 12361 24899 12419 24905
rect 12529 24939 12587 24945
rect 12529 24905 12541 24939
rect 12575 24936 12587 24939
rect 12710 24936 12716 24948
rect 12575 24908 12716 24936
rect 12575 24905 12587 24908
rect 12529 24899 12587 24905
rect 12710 24896 12716 24908
rect 12768 24896 12774 24948
rect 12897 24939 12955 24945
rect 12897 24905 12909 24939
rect 12943 24936 12955 24939
rect 13630 24936 13636 24948
rect 12943 24908 13636 24936
rect 12943 24905 12955 24908
rect 12897 24899 12955 24905
rect 13630 24896 13636 24908
rect 13688 24896 13694 24948
rect 15378 24896 15384 24948
rect 15436 24896 15442 24948
rect 16482 24896 16488 24948
rect 16540 24896 16546 24948
rect 18049 24939 18107 24945
rect 18049 24905 18061 24939
rect 18095 24905 18107 24939
rect 18049 24899 18107 24905
rect 12158 24868 12164 24880
rect 11624 24840 12164 24868
rect 10735 24772 11100 24800
rect 10735 24769 10747 24772
rect 10689 24763 10747 24769
rect 9122 24692 9128 24744
rect 9180 24732 9186 24744
rect 9217 24735 9275 24741
rect 9217 24732 9229 24735
rect 9180 24704 9229 24732
rect 9180 24692 9186 24704
rect 9217 24701 9229 24704
rect 9263 24701 9275 24735
rect 9217 24695 9275 24701
rect 7024 24636 8064 24664
rect 10428 24664 10456 24763
rect 11146 24760 11152 24812
rect 11204 24800 11210 24812
rect 11514 24800 11520 24812
rect 11204 24772 11520 24800
rect 11204 24760 11210 24772
rect 11514 24760 11520 24772
rect 11572 24760 11578 24812
rect 11624 24809 11652 24840
rect 12158 24828 12164 24840
rect 12216 24828 12222 24880
rect 15102 24828 15108 24880
rect 15160 24868 15166 24880
rect 15396 24868 15424 24896
rect 18064 24868 18092 24899
rect 18230 24896 18236 24948
rect 18288 24896 18294 24948
rect 19518 24896 19524 24948
rect 19576 24896 19582 24948
rect 21177 24939 21235 24945
rect 21177 24905 21189 24939
rect 21223 24936 21235 24939
rect 21223 24908 23428 24936
rect 21223 24905 21235 24908
rect 21177 24899 21235 24905
rect 22097 24871 22155 24877
rect 22097 24868 22109 24871
rect 15160 24840 15502 24868
rect 18064 24840 20116 24868
rect 15160 24828 15166 24840
rect 11609 24803 11667 24809
rect 11609 24769 11621 24803
rect 11655 24769 11667 24803
rect 11609 24763 11667 24769
rect 11698 24760 11704 24812
rect 11756 24760 11762 24812
rect 11808 24772 12388 24800
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24732 11023 24735
rect 11716 24732 11744 24760
rect 11808 24741 11836 24772
rect 11011 24704 11744 24732
rect 11793 24735 11851 24741
rect 11011 24701 11023 24704
rect 10965 24695 11023 24701
rect 11793 24701 11805 24735
rect 11839 24701 11851 24735
rect 11793 24695 11851 24701
rect 11885 24735 11943 24741
rect 11885 24701 11897 24735
rect 11931 24701 11943 24735
rect 11885 24695 11943 24701
rect 11238 24664 11244 24676
rect 10428 24636 11244 24664
rect 7024 24608 7052 24636
rect 6595 24568 6868 24596
rect 6595 24565 6607 24568
rect 6549 24559 6607 24565
rect 7006 24556 7012 24608
rect 7064 24556 7070 24608
rect 8036 24596 8064 24636
rect 11238 24624 11244 24636
rect 11296 24624 11302 24676
rect 11514 24624 11520 24676
rect 11572 24664 11578 24676
rect 11900 24664 11928 24695
rect 11572 24636 11928 24664
rect 11572 24624 11578 24636
rect 12360 24608 12388 24772
rect 12526 24760 12532 24812
rect 12584 24800 12590 24812
rect 12713 24803 12771 24809
rect 12713 24800 12725 24803
rect 12584 24772 12725 24800
rect 12584 24760 12590 24772
rect 12713 24769 12725 24772
rect 12759 24769 12771 24803
rect 12713 24763 12771 24769
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 14737 24803 14795 24809
rect 14737 24800 14749 24803
rect 13964 24772 14749 24800
rect 13964 24760 13970 24772
rect 14737 24769 14749 24772
rect 14783 24769 14795 24803
rect 14737 24763 14795 24769
rect 16942 24760 16948 24812
rect 17000 24760 17006 24812
rect 17034 24760 17040 24812
rect 17092 24800 17098 24812
rect 17497 24803 17555 24809
rect 17497 24800 17509 24803
rect 17092 24772 17509 24800
rect 17092 24760 17098 24772
rect 17497 24769 17509 24772
rect 17543 24769 17555 24803
rect 17497 24763 17555 24769
rect 18414 24760 18420 24812
rect 18472 24760 18478 24812
rect 19334 24760 19340 24812
rect 19392 24760 19398 24812
rect 15010 24692 15016 24744
rect 15068 24692 15074 24744
rect 20088 24732 20116 24840
rect 21836 24840 22109 24868
rect 20162 24760 20168 24812
rect 20220 24800 20226 24812
rect 21085 24803 21143 24809
rect 21085 24800 21097 24803
rect 20220 24772 21097 24800
rect 20220 24760 20226 24772
rect 21085 24769 21097 24772
rect 21131 24769 21143 24803
rect 21085 24763 21143 24769
rect 21266 24760 21272 24812
rect 21324 24800 21330 24812
rect 21836 24800 21864 24840
rect 22097 24837 22109 24840
rect 22143 24837 22155 24871
rect 22097 24831 22155 24837
rect 21324 24772 21864 24800
rect 23230 24772 23336 24800
rect 21324 24760 21330 24772
rect 23308 24744 23336 24772
rect 20990 24732 20996 24744
rect 20088 24704 20996 24732
rect 20990 24692 20996 24704
rect 21048 24692 21054 24744
rect 21821 24735 21879 24741
rect 21821 24701 21833 24735
rect 21867 24701 21879 24735
rect 21821 24695 21879 24701
rect 9766 24596 9772 24608
rect 8036 24568 9772 24596
rect 9766 24556 9772 24568
rect 9824 24556 9830 24608
rect 10597 24599 10655 24605
rect 10597 24565 10609 24599
rect 10643 24596 10655 24599
rect 11146 24596 11152 24608
rect 10643 24568 11152 24596
rect 10643 24565 10655 24568
rect 10597 24559 10655 24565
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 11330 24556 11336 24608
rect 11388 24556 11394 24608
rect 12342 24556 12348 24608
rect 12400 24556 12406 24608
rect 21542 24556 21548 24608
rect 21600 24556 21606 24608
rect 21836 24596 21864 24695
rect 23290 24692 23296 24744
rect 23348 24692 23354 24744
rect 23400 24608 23428 24908
rect 23658 24896 23664 24948
rect 23716 24896 23722 24948
rect 24305 24939 24363 24945
rect 24305 24905 24317 24939
rect 24351 24936 24363 24939
rect 24854 24936 24860 24948
rect 24351 24908 24860 24936
rect 24351 24905 24363 24908
rect 24305 24899 24363 24905
rect 24854 24896 24860 24908
rect 24912 24896 24918 24948
rect 30650 24896 30656 24948
rect 30708 24896 30714 24948
rect 31846 24896 31852 24948
rect 31904 24896 31910 24948
rect 25038 24828 25044 24880
rect 25096 24868 25102 24880
rect 25096 24840 27660 24868
rect 25096 24828 25102 24840
rect 23845 24803 23903 24809
rect 23845 24769 23857 24803
rect 23891 24800 23903 24803
rect 23891 24772 23980 24800
rect 23891 24769 23903 24772
rect 23845 24763 23903 24769
rect 23952 24673 23980 24772
rect 26970 24760 26976 24812
rect 27028 24760 27034 24812
rect 27154 24760 27160 24812
rect 27212 24760 27218 24812
rect 27249 24803 27307 24809
rect 27249 24769 27261 24803
rect 27295 24769 27307 24803
rect 27632 24800 27660 24840
rect 28994 24828 29000 24880
rect 29052 24868 29058 24880
rect 29052 24840 29500 24868
rect 29052 24828 29058 24840
rect 29472 24812 29500 24840
rect 30190 24828 30196 24880
rect 30248 24868 30254 24880
rect 30668 24868 30696 24896
rect 30248 24840 30604 24868
rect 30668 24840 30788 24868
rect 30248 24828 30254 24840
rect 27632 24772 28120 24800
rect 27249 24763 27307 24769
rect 24394 24692 24400 24744
rect 24452 24692 24458 24744
rect 24581 24735 24639 24741
rect 24581 24701 24593 24735
rect 24627 24732 24639 24735
rect 26510 24732 26516 24744
rect 24627 24704 26516 24732
rect 24627 24701 24639 24704
rect 24581 24695 24639 24701
rect 26510 24692 26516 24704
rect 26568 24732 26574 24744
rect 26988 24732 27016 24760
rect 26568 24704 27016 24732
rect 26568 24692 26574 24704
rect 27062 24692 27068 24744
rect 27120 24732 27126 24744
rect 27264 24732 27292 24763
rect 28092 24741 28120 24772
rect 28258 24760 28264 24812
rect 28316 24800 28322 24812
rect 28316 24772 29408 24800
rect 28316 24760 28322 24772
rect 27120 24704 27292 24732
rect 28077 24735 28135 24741
rect 27120 24692 27126 24704
rect 28077 24701 28089 24735
rect 28123 24732 28135 24735
rect 28626 24732 28632 24744
rect 28123 24704 28632 24732
rect 28123 24701 28135 24704
rect 28077 24695 28135 24701
rect 28626 24692 28632 24704
rect 28684 24692 28690 24744
rect 28810 24692 28816 24744
rect 28868 24692 28874 24744
rect 29380 24732 29408 24772
rect 29454 24760 29460 24812
rect 29512 24760 29518 24812
rect 30469 24803 30527 24809
rect 30469 24769 30481 24803
rect 30515 24769 30527 24803
rect 30576 24800 30604 24840
rect 30760 24809 30788 24840
rect 31312 24840 31892 24868
rect 31312 24812 31340 24840
rect 30653 24803 30711 24809
rect 30653 24800 30665 24803
rect 30576 24772 30665 24800
rect 30469 24763 30527 24769
rect 30653 24769 30665 24772
rect 30699 24769 30711 24803
rect 30653 24763 30711 24769
rect 30745 24803 30803 24809
rect 30745 24769 30757 24803
rect 30791 24800 30803 24803
rect 30929 24803 30987 24809
rect 30929 24800 30941 24803
rect 30791 24772 30941 24800
rect 30791 24769 30803 24772
rect 30745 24763 30803 24769
rect 30929 24769 30941 24772
rect 30975 24769 30987 24803
rect 30929 24763 30987 24769
rect 31113 24803 31171 24809
rect 31113 24769 31125 24803
rect 31159 24769 31171 24803
rect 31113 24763 31171 24769
rect 30193 24735 30251 24741
rect 30193 24732 30205 24735
rect 29380 24704 30205 24732
rect 30193 24701 30205 24704
rect 30239 24701 30251 24735
rect 30193 24695 30251 24701
rect 23937 24667 23995 24673
rect 23937 24633 23949 24667
rect 23983 24633 23995 24667
rect 23937 24627 23995 24633
rect 24854 24624 24860 24676
rect 24912 24664 24918 24676
rect 28828 24664 28856 24692
rect 24912 24636 28856 24664
rect 24912 24624 24918 24636
rect 29178 24624 29184 24676
rect 29236 24624 29242 24676
rect 29273 24667 29331 24673
rect 29273 24633 29285 24667
rect 29319 24664 29331 24667
rect 30006 24664 30012 24676
rect 29319 24636 30012 24664
rect 29319 24633 29331 24636
rect 29273 24627 29331 24633
rect 30006 24624 30012 24636
rect 30064 24664 30070 24676
rect 30484 24664 30512 24763
rect 31128 24732 31156 24763
rect 31294 24760 31300 24812
rect 31352 24760 31358 24812
rect 31386 24760 31392 24812
rect 31444 24760 31450 24812
rect 31481 24803 31539 24809
rect 31481 24769 31493 24803
rect 31527 24769 31539 24803
rect 31481 24763 31539 24769
rect 31573 24803 31631 24809
rect 31573 24769 31585 24803
rect 31619 24800 31631 24803
rect 31757 24803 31815 24809
rect 31757 24800 31769 24803
rect 31619 24772 31769 24800
rect 31619 24769 31631 24772
rect 31573 24763 31631 24769
rect 31757 24769 31769 24772
rect 31803 24769 31815 24803
rect 31864 24800 31892 24840
rect 31941 24803 31999 24809
rect 31941 24800 31953 24803
rect 31864 24772 31953 24800
rect 31757 24763 31815 24769
rect 31941 24769 31953 24772
rect 31987 24769 31999 24803
rect 31941 24763 31999 24769
rect 31496 24732 31524 24763
rect 31128 24704 31616 24732
rect 30064 24636 30512 24664
rect 30064 24624 30070 24636
rect 31588 24608 31616 24704
rect 23106 24596 23112 24608
rect 21836 24568 23112 24596
rect 23106 24556 23112 24568
rect 23164 24556 23170 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 23569 24599 23627 24605
rect 23569 24596 23581 24599
rect 23440 24568 23581 24596
rect 23440 24556 23446 24568
rect 23569 24565 23581 24568
rect 23615 24565 23627 24599
rect 23569 24559 23627 24565
rect 30469 24599 30527 24605
rect 30469 24565 30481 24599
rect 30515 24596 30527 24599
rect 30650 24596 30656 24608
rect 30515 24568 30656 24596
rect 30515 24565 30527 24568
rect 30469 24559 30527 24565
rect 30650 24556 30656 24568
rect 30708 24556 30714 24608
rect 31570 24556 31576 24608
rect 31628 24556 31634 24608
rect 1104 24506 34684 24528
rect 1104 24454 5147 24506
rect 5199 24454 5211 24506
rect 5263 24454 5275 24506
rect 5327 24454 5339 24506
rect 5391 24454 5403 24506
rect 5455 24454 13541 24506
rect 13593 24454 13605 24506
rect 13657 24454 13669 24506
rect 13721 24454 13733 24506
rect 13785 24454 13797 24506
rect 13849 24454 21935 24506
rect 21987 24454 21999 24506
rect 22051 24454 22063 24506
rect 22115 24454 22127 24506
rect 22179 24454 22191 24506
rect 22243 24454 30329 24506
rect 30381 24454 30393 24506
rect 30445 24454 30457 24506
rect 30509 24454 30521 24506
rect 30573 24454 30585 24506
rect 30637 24454 34684 24506
rect 1104 24432 34684 24454
rect 4338 24352 4344 24404
rect 4396 24352 4402 24404
rect 4706 24352 4712 24404
rect 4764 24352 4770 24404
rect 7190 24352 7196 24404
rect 7248 24392 7254 24404
rect 8021 24395 8079 24401
rect 8021 24392 8033 24395
rect 7248 24364 8033 24392
rect 7248 24352 7254 24364
rect 8021 24361 8033 24364
rect 8067 24361 8079 24395
rect 8021 24355 8079 24361
rect 11330 24352 11336 24404
rect 11388 24392 11394 24404
rect 11609 24395 11667 24401
rect 11609 24392 11621 24395
rect 11388 24364 11621 24392
rect 11388 24352 11394 24364
rect 11609 24361 11621 24364
rect 11655 24392 11667 24395
rect 11655 24364 12112 24392
rect 11655 24361 11667 24364
rect 11609 24355 11667 24361
rect 4356 24324 4384 24352
rect 11793 24327 11851 24333
rect 11793 24324 11805 24327
rect 4356 24296 5120 24324
rect 4985 24259 5043 24265
rect 4985 24256 4997 24259
rect 4540 24228 4997 24256
rect 4540 24197 4568 24228
rect 4985 24225 4997 24228
rect 5031 24225 5043 24259
rect 4985 24219 5043 24225
rect 5092 24200 5120 24296
rect 11440 24296 11805 24324
rect 5718 24216 5724 24268
rect 5776 24256 5782 24268
rect 5813 24259 5871 24265
rect 5813 24256 5825 24259
rect 5776 24228 5825 24256
rect 5776 24216 5782 24228
rect 5813 24225 5825 24228
rect 5859 24225 5871 24259
rect 5813 24219 5871 24225
rect 6273 24259 6331 24265
rect 6273 24225 6285 24259
rect 6319 24256 6331 24259
rect 8478 24256 8484 24268
rect 6319 24228 8484 24256
rect 6319 24225 6331 24228
rect 6273 24219 6331 24225
rect 8478 24216 8484 24228
rect 8536 24256 8542 24268
rect 9214 24256 9220 24268
rect 8536 24228 9220 24256
rect 8536 24216 8542 24228
rect 9214 24216 9220 24228
rect 9272 24216 9278 24268
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24157 4583 24191
rect 4525 24151 4583 24157
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 4816 24120 4844 24151
rect 4890 24148 4896 24200
rect 4948 24148 4954 24200
rect 5074 24148 5080 24200
rect 5132 24148 5138 24200
rect 11440 24197 11468 24296
rect 11793 24293 11805 24296
rect 11839 24293 11851 24327
rect 11793 24287 11851 24293
rect 12084 24197 12112 24364
rect 15010 24352 15016 24404
rect 15068 24392 15074 24404
rect 15473 24395 15531 24401
rect 15473 24392 15485 24395
rect 15068 24364 15485 24392
rect 15068 24352 15074 24364
rect 15473 24361 15485 24364
rect 15519 24361 15531 24395
rect 15473 24355 15531 24361
rect 17773 24395 17831 24401
rect 17773 24361 17785 24395
rect 17819 24392 17831 24395
rect 18414 24392 18420 24404
rect 17819 24364 18420 24392
rect 17819 24361 17831 24364
rect 17773 24355 17831 24361
rect 18414 24352 18420 24364
rect 18472 24352 18478 24404
rect 19245 24395 19303 24401
rect 19245 24361 19257 24395
rect 19291 24392 19303 24395
rect 19334 24392 19340 24404
rect 19291 24364 19340 24392
rect 19291 24361 19303 24364
rect 19245 24355 19303 24361
rect 19334 24352 19340 24364
rect 19392 24352 19398 24404
rect 21266 24352 21272 24404
rect 21324 24352 21330 24404
rect 21542 24352 21548 24404
rect 21600 24352 21606 24404
rect 31389 24395 31447 24401
rect 26528 24364 28580 24392
rect 16574 24284 16580 24336
rect 16632 24324 16638 24336
rect 17221 24327 17279 24333
rect 17221 24324 17233 24327
rect 16632 24296 17233 24324
rect 16632 24284 16638 24296
rect 17221 24293 17233 24296
rect 17267 24293 17279 24327
rect 19058 24324 19064 24336
rect 17221 24287 17279 24293
rect 18708 24296 19064 24324
rect 11425 24191 11483 24197
rect 11425 24157 11437 24191
rect 11471 24157 11483 24191
rect 11425 24151 11483 24157
rect 11701 24191 11759 24197
rect 11701 24157 11713 24191
rect 11747 24188 11759 24191
rect 12069 24191 12127 24197
rect 11747 24160 12020 24188
rect 11747 24157 11759 24160
rect 11701 24151 11759 24157
rect 5261 24123 5319 24129
rect 5261 24120 5273 24123
rect 4816 24092 5273 24120
rect 5261 24089 5273 24092
rect 5307 24089 5319 24123
rect 5261 24083 5319 24089
rect 6546 24080 6552 24132
rect 6604 24080 6610 24132
rect 6638 24080 6644 24132
rect 6696 24120 6702 24132
rect 7006 24120 7012 24132
rect 6696 24092 7012 24120
rect 6696 24080 6702 24092
rect 7006 24080 7012 24092
rect 7064 24080 7070 24132
rect 11793 24123 11851 24129
rect 11793 24089 11805 24123
rect 11839 24120 11851 24123
rect 11882 24120 11888 24132
rect 11839 24092 11888 24120
rect 11839 24089 11851 24092
rect 11793 24083 11851 24089
rect 11882 24080 11888 24092
rect 11940 24080 11946 24132
rect 4338 24012 4344 24064
rect 4396 24012 4402 24064
rect 11238 24012 11244 24064
rect 11296 24012 11302 24064
rect 11992 24061 12020 24160
rect 12069 24157 12081 24191
rect 12115 24157 12127 24191
rect 12069 24151 12127 24157
rect 15657 24191 15715 24197
rect 15657 24157 15669 24191
rect 15703 24188 15715 24191
rect 15838 24188 15844 24200
rect 15703 24160 15844 24188
rect 15703 24157 15715 24160
rect 15657 24151 15715 24157
rect 15838 24148 15844 24160
rect 15896 24148 15902 24200
rect 17494 24148 17500 24200
rect 17552 24188 17558 24200
rect 18708 24197 18736 24296
rect 19058 24284 19064 24296
rect 19116 24324 19122 24336
rect 19116 24296 20208 24324
rect 19116 24284 19122 24296
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 18831 24228 19564 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 19536 24200 19564 24228
rect 20180 24200 20208 24296
rect 18693 24191 18751 24197
rect 17552 24160 18460 24188
rect 17552 24148 17558 24160
rect 17589 24123 17647 24129
rect 17589 24089 17601 24123
rect 17635 24120 17647 24123
rect 18432 24120 18460 24160
rect 18693 24157 18705 24191
rect 18739 24157 18751 24191
rect 18693 24151 18751 24157
rect 19518 24148 19524 24200
rect 19576 24148 19582 24200
rect 20162 24148 20168 24200
rect 20220 24148 20226 24200
rect 21085 24191 21143 24197
rect 21085 24157 21097 24191
rect 21131 24188 21143 24191
rect 21560 24188 21588 24352
rect 23106 24216 23112 24268
rect 23164 24256 23170 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 23164 24228 24593 24256
rect 23164 24216 23170 24228
rect 24581 24225 24593 24228
rect 24627 24256 24639 24259
rect 25406 24256 25412 24268
rect 24627 24228 25412 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 25406 24216 25412 24228
rect 25464 24256 25470 24268
rect 25464 24228 25912 24256
rect 25464 24216 25470 24228
rect 25884 24200 25912 24228
rect 21131 24160 21588 24188
rect 21131 24157 21143 24160
rect 21085 24151 21143 24157
rect 25866 24148 25872 24200
rect 25924 24148 25930 24200
rect 26142 24148 26148 24200
rect 26200 24188 26206 24200
rect 26528 24188 26556 24364
rect 28552 24336 28580 24364
rect 31389 24361 31401 24395
rect 31435 24361 31447 24395
rect 31389 24355 31447 24361
rect 26605 24327 26663 24333
rect 26605 24293 26617 24327
rect 26651 24324 26663 24327
rect 26651 24296 27292 24324
rect 26651 24293 26663 24296
rect 26605 24287 26663 24293
rect 27062 24256 27068 24268
rect 26988 24228 27068 24256
rect 26988 24197 27016 24228
rect 27062 24216 27068 24228
rect 27120 24216 27126 24268
rect 27264 24265 27292 24296
rect 28534 24284 28540 24336
rect 28592 24284 28598 24336
rect 31404 24324 31432 24355
rect 31570 24352 31576 24404
rect 31628 24352 31634 24404
rect 32582 24352 32588 24404
rect 32640 24352 32646 24404
rect 31757 24327 31815 24333
rect 31757 24324 31769 24327
rect 28966 24296 30864 24324
rect 31404 24296 31769 24324
rect 27249 24259 27307 24265
rect 27249 24225 27261 24259
rect 27295 24225 27307 24259
rect 27249 24219 27307 24225
rect 26789 24191 26847 24197
rect 26789 24188 26801 24191
rect 26200 24160 26801 24188
rect 26200 24148 26206 24160
rect 26789 24157 26801 24160
rect 26835 24157 26847 24191
rect 26789 24151 26847 24157
rect 26973 24191 27031 24197
rect 26973 24157 26985 24191
rect 27019 24157 27031 24191
rect 26973 24151 27031 24157
rect 27154 24148 27160 24200
rect 27212 24148 27218 24200
rect 18782 24120 18788 24132
rect 17635 24092 18368 24120
rect 18432 24092 18788 24120
rect 17635 24089 17647 24092
rect 17589 24083 17647 24089
rect 11977 24055 12035 24061
rect 11977 24021 11989 24055
rect 12023 24052 12035 24055
rect 12066 24052 12072 24064
rect 12023 24024 12072 24052
rect 12023 24021 12035 24024
rect 11977 24015 12035 24021
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 17310 24012 17316 24064
rect 17368 24052 17374 24064
rect 18340 24061 18368 24092
rect 18782 24080 18788 24092
rect 18840 24120 18846 24132
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 18840 24092 19625 24120
rect 18840 24080 18846 24092
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 19613 24083 19671 24089
rect 19702 24080 19708 24132
rect 19760 24120 19766 24132
rect 19797 24123 19855 24129
rect 19797 24120 19809 24123
rect 19760 24092 19809 24120
rect 19760 24080 19766 24092
rect 19797 24089 19809 24092
rect 19843 24120 19855 24123
rect 22462 24120 22468 24132
rect 19843 24092 22468 24120
rect 19843 24089 19855 24092
rect 19797 24083 19855 24089
rect 22462 24080 22468 24092
rect 22520 24080 22526 24132
rect 24854 24080 24860 24132
rect 24912 24080 24918 24132
rect 25314 24080 25320 24132
rect 25372 24080 25378 24132
rect 26881 24123 26939 24129
rect 26881 24120 26893 24123
rect 26160 24092 26893 24120
rect 17405 24055 17463 24061
rect 17405 24052 17417 24055
rect 17368 24024 17417 24052
rect 17368 24012 17374 24024
rect 17405 24021 17417 24024
rect 17451 24021 17463 24055
rect 17405 24015 17463 24021
rect 18325 24055 18383 24061
rect 18325 24021 18337 24055
rect 18371 24021 18383 24055
rect 18325 24015 18383 24021
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 23382 24012 23388 24064
rect 23440 24052 23446 24064
rect 26160 24052 26188 24092
rect 26881 24089 26893 24092
rect 26927 24089 26939 24123
rect 28966 24120 28994 24296
rect 29454 24148 29460 24200
rect 29512 24188 29518 24200
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 29512 24160 29561 24188
rect 29512 24148 29518 24160
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 30836 24188 30864 24296
rect 31757 24293 31769 24296
rect 31803 24324 31815 24327
rect 32122 24324 32128 24336
rect 31803 24296 32128 24324
rect 31803 24293 31815 24296
rect 31757 24287 31815 24293
rect 32122 24284 32128 24296
rect 32180 24324 32186 24336
rect 32600 24324 32628 24352
rect 32180 24296 32628 24324
rect 32180 24284 32186 24296
rect 31481 24191 31539 24197
rect 31481 24188 31493 24191
rect 30836 24160 31493 24188
rect 29549 24151 29607 24157
rect 31481 24157 31493 24160
rect 31527 24188 31539 24191
rect 32033 24191 32091 24197
rect 32033 24188 32045 24191
rect 31527 24160 32045 24188
rect 31527 24157 31539 24160
rect 31481 24151 31539 24157
rect 32033 24157 32045 24160
rect 32079 24157 32091 24191
rect 32033 24151 32091 24157
rect 32950 24148 32956 24200
rect 33008 24148 33014 24200
rect 34330 24148 34336 24200
rect 34388 24148 34394 24200
rect 26881 24083 26939 24089
rect 26988 24092 28994 24120
rect 23440 24024 26188 24052
rect 26329 24055 26387 24061
rect 23440 24012 23446 24024
rect 26329 24021 26341 24055
rect 26375 24052 26387 24055
rect 26602 24052 26608 24064
rect 26375 24024 26608 24052
rect 26375 24021 26387 24024
rect 26329 24015 26387 24021
rect 26602 24012 26608 24024
rect 26660 24052 26666 24064
rect 26988 24052 27016 24092
rect 29822 24080 29828 24132
rect 29880 24120 29886 24132
rect 30285 24123 30343 24129
rect 30285 24120 30297 24123
rect 29880 24092 30297 24120
rect 29880 24080 29886 24092
rect 30285 24089 30297 24092
rect 30331 24089 30343 24123
rect 30285 24083 30343 24089
rect 34054 24080 34060 24132
rect 34112 24080 34118 24132
rect 26660 24024 27016 24052
rect 26660 24012 26666 24024
rect 27890 24012 27896 24064
rect 27948 24012 27954 24064
rect 30098 24012 30104 24064
rect 30156 24052 30162 24064
rect 31021 24055 31079 24061
rect 31021 24052 31033 24055
rect 30156 24024 31033 24052
rect 30156 24012 30162 24024
rect 31021 24021 31033 24024
rect 31067 24052 31079 24055
rect 31294 24052 31300 24064
rect 31067 24024 31300 24052
rect 31067 24021 31079 24024
rect 31021 24015 31079 24021
rect 31294 24012 31300 24024
rect 31352 24012 31358 24064
rect 1104 23962 34840 23984
rect 1104 23910 9344 23962
rect 9396 23910 9408 23962
rect 9460 23910 9472 23962
rect 9524 23910 9536 23962
rect 9588 23910 9600 23962
rect 9652 23910 17738 23962
rect 17790 23910 17802 23962
rect 17854 23910 17866 23962
rect 17918 23910 17930 23962
rect 17982 23910 17994 23962
rect 18046 23910 26132 23962
rect 26184 23910 26196 23962
rect 26248 23910 26260 23962
rect 26312 23910 26324 23962
rect 26376 23910 26388 23962
rect 26440 23910 34526 23962
rect 34578 23910 34590 23962
rect 34642 23910 34654 23962
rect 34706 23910 34718 23962
rect 34770 23910 34782 23962
rect 34834 23910 34840 23962
rect 1104 23888 34840 23910
rect 4338 23848 4344 23860
rect 4080 23820 4344 23848
rect 4080 23789 4108 23820
rect 4338 23808 4344 23820
rect 4396 23808 4402 23860
rect 5537 23851 5595 23857
rect 5537 23817 5549 23851
rect 5583 23848 5595 23851
rect 5718 23848 5724 23860
rect 5583 23820 5724 23848
rect 5583 23817 5595 23820
rect 5537 23811 5595 23817
rect 5718 23808 5724 23820
rect 5776 23808 5782 23860
rect 6362 23808 6368 23860
rect 6420 23808 6426 23860
rect 6546 23808 6552 23860
rect 6604 23808 6610 23860
rect 12066 23808 12072 23860
rect 12124 23808 12130 23860
rect 13906 23848 13912 23860
rect 12912 23820 13912 23848
rect 4065 23783 4123 23789
rect 4065 23749 4077 23783
rect 4111 23749 4123 23783
rect 4065 23743 4123 23749
rect 4522 23740 4528 23792
rect 4580 23740 4586 23792
rect 3142 23672 3148 23724
rect 3200 23712 3206 23724
rect 3789 23715 3847 23721
rect 3789 23712 3801 23715
rect 3200 23684 3801 23712
rect 3200 23672 3206 23684
rect 3789 23681 3801 23684
rect 3835 23681 3847 23715
rect 6380 23712 6408 23808
rect 9766 23740 9772 23792
rect 9824 23740 9830 23792
rect 6733 23715 6791 23721
rect 6733 23712 6745 23715
rect 6380 23684 6745 23712
rect 3789 23675 3847 23681
rect 6733 23681 6745 23684
rect 6779 23681 6791 23715
rect 6733 23675 6791 23681
rect 8478 23672 8484 23724
rect 8536 23672 8542 23724
rect 12342 23672 12348 23724
rect 12400 23712 12406 23724
rect 12912 23721 12940 23820
rect 13906 23808 13912 23820
rect 13964 23808 13970 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 19426 23848 19432 23860
rect 19383 23820 19432 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 19426 23808 19432 23820
rect 19484 23808 19490 23860
rect 19518 23808 19524 23860
rect 19576 23808 19582 23860
rect 20714 23808 20720 23860
rect 20772 23808 20778 23860
rect 23014 23808 23020 23860
rect 23072 23808 23078 23860
rect 23290 23808 23296 23860
rect 23348 23848 23354 23860
rect 24765 23851 24823 23857
rect 23348 23820 23980 23848
rect 23348 23808 23354 23820
rect 13170 23740 13176 23792
rect 13228 23740 13234 23792
rect 14458 23780 14464 23792
rect 14398 23752 14464 23780
rect 14458 23740 14464 23752
rect 14516 23780 14522 23792
rect 15102 23780 15108 23792
rect 14516 23752 15108 23780
rect 14516 23740 14522 23752
rect 15102 23740 15108 23752
rect 15160 23780 15166 23792
rect 16758 23780 16764 23792
rect 15160 23752 16764 23780
rect 15160 23740 15166 23752
rect 16758 23740 16764 23752
rect 16816 23740 16822 23792
rect 18969 23783 19027 23789
rect 18969 23749 18981 23783
rect 19015 23780 19027 23783
rect 19015 23752 19288 23780
rect 19015 23749 19027 23752
rect 18969 23743 19027 23749
rect 19260 23724 19288 23752
rect 12621 23715 12679 23721
rect 12621 23712 12633 23715
rect 12400 23684 12633 23712
rect 12400 23672 12406 23684
rect 12621 23681 12633 23684
rect 12667 23681 12679 23715
rect 12621 23675 12679 23681
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23681 12955 23715
rect 12897 23675 12955 23681
rect 19153 23715 19211 23721
rect 19153 23681 19165 23715
rect 19199 23681 19211 23715
rect 19153 23675 19211 23681
rect 8202 23604 8208 23656
rect 8260 23644 8266 23656
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 8260 23616 8769 23644
rect 8260 23604 8266 23616
rect 8757 23613 8769 23616
rect 8803 23613 8815 23647
rect 19168 23644 19196 23675
rect 19242 23672 19248 23724
rect 19300 23712 19306 23724
rect 19429 23715 19487 23721
rect 19429 23712 19441 23715
rect 19300 23684 19441 23712
rect 19300 23672 19306 23684
rect 19429 23681 19441 23684
rect 19475 23681 19487 23715
rect 19429 23675 19487 23681
rect 19613 23715 19671 23721
rect 19613 23681 19625 23715
rect 19659 23712 19671 23715
rect 20732 23712 20760 23808
rect 23032 23780 23060 23808
rect 23952 23780 23980 23820
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 26602 23848 26608 23860
rect 24811 23820 26608 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 26602 23808 26608 23820
rect 26660 23808 26666 23860
rect 27154 23808 27160 23860
rect 27212 23808 27218 23860
rect 27617 23851 27675 23857
rect 27617 23817 27629 23851
rect 27663 23848 27675 23851
rect 27706 23848 27712 23860
rect 27663 23820 27712 23848
rect 27663 23817 27675 23820
rect 27617 23811 27675 23817
rect 27706 23808 27712 23820
rect 27764 23808 27770 23860
rect 27890 23808 27896 23860
rect 27948 23808 27954 23860
rect 32677 23851 32735 23857
rect 32677 23817 32689 23851
rect 32723 23817 32735 23851
rect 32677 23811 32735 23817
rect 33229 23851 33287 23857
rect 33229 23817 33241 23851
rect 33275 23848 33287 23851
rect 34054 23848 34060 23860
rect 33275 23820 34060 23848
rect 33275 23817 33287 23820
rect 33229 23811 33287 23817
rect 25222 23780 25228 23792
rect 22388 23752 23060 23780
rect 23874 23752 25228 23780
rect 19659 23684 20760 23712
rect 22097 23715 22155 23721
rect 19659 23681 19671 23684
rect 19613 23675 19671 23681
rect 22097 23681 22109 23715
rect 22143 23712 22155 23715
rect 22278 23712 22284 23724
rect 22143 23684 22284 23712
rect 22143 23681 22155 23684
rect 22097 23675 22155 23681
rect 19628 23644 19656 23675
rect 22278 23672 22284 23684
rect 22336 23672 22342 23724
rect 22388 23721 22416 23752
rect 25222 23740 25228 23752
rect 25280 23740 25286 23792
rect 25869 23783 25927 23789
rect 25869 23749 25881 23783
rect 25915 23780 25927 23783
rect 25958 23780 25964 23792
rect 25915 23752 25964 23780
rect 25915 23749 25927 23752
rect 25869 23743 25927 23749
rect 25958 23740 25964 23752
rect 26016 23740 26022 23792
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23681 22431 23715
rect 25317 23715 25375 23721
rect 25317 23712 25329 23715
rect 22373 23675 22431 23681
rect 24596 23684 25329 23712
rect 24596 23653 24624 23684
rect 25317 23681 25329 23684
rect 25363 23712 25375 23715
rect 26510 23712 26516 23724
rect 25363 23684 26516 23712
rect 25363 23681 25375 23684
rect 25317 23675 25375 23681
rect 26510 23672 26516 23684
rect 26568 23672 26574 23724
rect 22649 23647 22707 23653
rect 22649 23644 22661 23647
rect 19168 23616 19656 23644
rect 22296 23616 22661 23644
rect 8757 23607 8815 23613
rect 22296 23585 22324 23616
rect 22649 23613 22661 23616
rect 22695 23613 22707 23647
rect 22649 23607 22707 23613
rect 24581 23647 24639 23653
rect 24581 23613 24593 23647
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 24670 23604 24676 23656
rect 24728 23604 24734 23656
rect 27172 23644 27200 23808
rect 27908 23780 27936 23808
rect 27448 23752 27936 23780
rect 27448 23721 27476 23752
rect 28626 23740 28632 23792
rect 28684 23780 28690 23792
rect 31478 23780 31484 23792
rect 28684 23752 31484 23780
rect 28684 23740 28690 23752
rect 31478 23740 31484 23752
rect 31536 23780 31542 23792
rect 32309 23783 32367 23789
rect 32309 23780 32321 23783
rect 31536 23752 32321 23780
rect 31536 23740 31542 23752
rect 32309 23749 32321 23752
rect 32355 23749 32367 23783
rect 32692 23780 32720 23811
rect 34054 23808 34060 23820
rect 34112 23808 34118 23860
rect 32692 23752 33088 23780
rect 32309 23743 32367 23749
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23681 27491 23715
rect 27433 23675 27491 23681
rect 27709 23715 27767 23721
rect 27709 23681 27721 23715
rect 27755 23712 27767 23715
rect 28350 23712 28356 23724
rect 27755 23684 28356 23712
rect 27755 23681 27767 23684
rect 27709 23675 27767 23681
rect 28350 23672 28356 23684
rect 28408 23672 28414 23724
rect 29730 23672 29736 23724
rect 29788 23672 29794 23724
rect 29914 23672 29920 23724
rect 29972 23672 29978 23724
rect 30006 23672 30012 23724
rect 30064 23672 30070 23724
rect 30098 23672 30104 23724
rect 30156 23672 30162 23724
rect 30282 23672 30288 23724
rect 30340 23672 30346 23724
rect 32122 23672 32128 23724
rect 32180 23672 32186 23724
rect 32401 23715 32459 23721
rect 32401 23681 32413 23715
rect 32447 23681 32459 23715
rect 32401 23675 32459 23681
rect 32493 23715 32551 23721
rect 32493 23681 32505 23715
rect 32539 23681 32551 23715
rect 32493 23675 32551 23681
rect 27893 23647 27951 23653
rect 27893 23644 27905 23647
rect 27172 23616 27905 23644
rect 27893 23613 27905 23616
rect 27939 23613 27951 23647
rect 27893 23607 27951 23613
rect 28534 23604 28540 23656
rect 28592 23604 28598 23656
rect 22281 23579 22339 23585
rect 22281 23545 22293 23579
rect 22327 23545 22339 23579
rect 22281 23539 22339 23545
rect 24118 23536 24124 23588
rect 24176 23576 24182 23588
rect 32416 23576 32444 23675
rect 24176 23548 32444 23576
rect 24176 23536 24182 23548
rect 10226 23468 10232 23520
rect 10284 23468 10290 23520
rect 14645 23511 14703 23517
rect 14645 23477 14657 23511
rect 14691 23508 14703 23511
rect 14918 23508 14924 23520
rect 14691 23480 14924 23508
rect 14691 23477 14703 23480
rect 14645 23471 14703 23477
rect 14918 23468 14924 23480
rect 14976 23468 14982 23520
rect 25130 23468 25136 23520
rect 25188 23468 25194 23520
rect 27246 23468 27252 23520
rect 27304 23468 27310 23520
rect 29549 23511 29607 23517
rect 29549 23477 29561 23511
rect 29595 23508 29607 23511
rect 31294 23508 31300 23520
rect 29595 23480 31300 23508
rect 29595 23477 29607 23480
rect 29549 23471 29607 23477
rect 31294 23468 31300 23480
rect 31352 23468 31358 23520
rect 31662 23468 31668 23520
rect 31720 23508 31726 23520
rect 32508 23508 32536 23675
rect 32582 23672 32588 23724
rect 32640 23672 32646 23724
rect 32766 23672 32772 23724
rect 32824 23672 32830 23724
rect 33060 23721 33088 23752
rect 32861 23715 32919 23721
rect 32861 23681 32873 23715
rect 32907 23681 32919 23715
rect 32861 23675 32919 23681
rect 33045 23715 33103 23721
rect 33045 23681 33057 23715
rect 33091 23681 33103 23715
rect 33045 23675 33103 23681
rect 32600 23644 32628 23672
rect 32876 23644 32904 23675
rect 32600 23616 32904 23644
rect 31720 23480 32536 23508
rect 31720 23468 31726 23480
rect 1104 23418 34684 23440
rect 1104 23366 5147 23418
rect 5199 23366 5211 23418
rect 5263 23366 5275 23418
rect 5327 23366 5339 23418
rect 5391 23366 5403 23418
rect 5455 23366 13541 23418
rect 13593 23366 13605 23418
rect 13657 23366 13669 23418
rect 13721 23366 13733 23418
rect 13785 23366 13797 23418
rect 13849 23366 21935 23418
rect 21987 23366 21999 23418
rect 22051 23366 22063 23418
rect 22115 23366 22127 23418
rect 22179 23366 22191 23418
rect 22243 23366 30329 23418
rect 30381 23366 30393 23418
rect 30445 23366 30457 23418
rect 30509 23366 30521 23418
rect 30573 23366 30585 23418
rect 30637 23366 34684 23418
rect 1104 23344 34684 23366
rect 12342 23264 12348 23316
rect 12400 23264 12406 23316
rect 19242 23304 19248 23316
rect 18432 23276 19248 23304
rect 5902 23168 5908 23180
rect 5276 23140 5908 23168
rect 4982 23060 4988 23112
rect 5040 23100 5046 23112
rect 5276 23109 5304 23140
rect 5902 23128 5908 23140
rect 5960 23128 5966 23180
rect 10597 23171 10655 23177
rect 10597 23168 10609 23171
rect 9232 23140 10609 23168
rect 9232 23112 9260 23140
rect 10597 23137 10609 23140
rect 10643 23137 10655 23171
rect 10597 23131 10655 23137
rect 10873 23171 10931 23177
rect 10873 23137 10885 23171
rect 10919 23168 10931 23171
rect 11238 23168 11244 23180
rect 10919 23140 11244 23168
rect 10919 23137 10931 23140
rect 10873 23131 10931 23137
rect 11238 23128 11244 23140
rect 11296 23128 11302 23180
rect 18432 23177 18460 23276
rect 19242 23264 19248 23276
rect 19300 23264 19306 23316
rect 21634 23264 21640 23316
rect 21692 23264 21698 23316
rect 22278 23264 22284 23316
rect 22336 23304 22342 23316
rect 22465 23307 22523 23313
rect 22465 23304 22477 23307
rect 22336 23276 22477 23304
rect 22336 23264 22342 23276
rect 22465 23273 22477 23276
rect 22511 23273 22523 23307
rect 22465 23267 22523 23273
rect 24765 23307 24823 23313
rect 24765 23273 24777 23307
rect 24811 23304 24823 23307
rect 24854 23304 24860 23316
rect 24811 23276 24860 23304
rect 24811 23273 24823 23276
rect 24765 23267 24823 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 28350 23264 28356 23316
rect 28408 23264 28414 23316
rect 29012 23276 30420 23304
rect 19061 23239 19119 23245
rect 19061 23205 19073 23239
rect 19107 23205 19119 23239
rect 28261 23239 28319 23245
rect 19061 23199 19119 23205
rect 22066 23208 23336 23236
rect 18417 23171 18475 23177
rect 18417 23137 18429 23171
rect 18463 23137 18475 23171
rect 18417 23131 18475 23137
rect 18782 23128 18788 23180
rect 18840 23128 18846 23180
rect 5077 23103 5135 23109
rect 5077 23100 5089 23103
rect 5040 23072 5089 23100
rect 5040 23060 5046 23072
rect 5077 23069 5089 23072
rect 5123 23069 5135 23103
rect 5077 23063 5135 23069
rect 5261 23103 5319 23109
rect 5261 23069 5273 23103
rect 5307 23069 5319 23103
rect 5261 23063 5319 23069
rect 5442 23060 5448 23112
rect 5500 23100 5506 23112
rect 5629 23103 5687 23109
rect 5629 23100 5641 23103
rect 5500 23072 5641 23100
rect 5500 23060 5506 23072
rect 5629 23069 5641 23072
rect 5675 23069 5687 23103
rect 5629 23063 5687 23069
rect 5994 23060 6000 23112
rect 6052 23060 6058 23112
rect 9214 23060 9220 23112
rect 9272 23060 9278 23112
rect 10137 23103 10195 23109
rect 10137 23069 10149 23103
rect 10183 23100 10195 23103
rect 10226 23100 10232 23112
rect 10183 23072 10232 23100
rect 10183 23069 10195 23072
rect 10137 23063 10195 23069
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 15933 23103 15991 23109
rect 15933 23069 15945 23103
rect 15979 23100 15991 23103
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15979 23072 16037 23100
rect 15979 23069 15991 23072
rect 15933 23063 15991 23069
rect 16025 23069 16037 23072
rect 16071 23069 16083 23103
rect 16025 23063 16083 23069
rect 4522 22992 4528 23044
rect 4580 23032 4586 23044
rect 4580 23004 5764 23032
rect 4580 22992 4586 23004
rect 4890 22924 4896 22976
rect 4948 22964 4954 22976
rect 5169 22967 5227 22973
rect 5169 22964 5181 22967
rect 4948 22936 5181 22964
rect 4948 22924 4954 22936
rect 5169 22933 5181 22936
rect 5215 22933 5227 22967
rect 5736 22964 5764 23004
rect 6288 23004 6394 23032
rect 11072 23004 11362 23032
rect 6288 22964 6316 23004
rect 11072 22976 11100 23004
rect 15102 22992 15108 23044
rect 15160 22992 15166 23044
rect 15654 22992 15660 23044
rect 15712 22992 15718 23044
rect 15948 23032 15976 23063
rect 16390 23060 16396 23112
rect 16448 23060 16454 23112
rect 19076 23100 19104 23199
rect 20622 23128 20628 23180
rect 20680 23168 20686 23180
rect 22066 23168 22094 23208
rect 23308 23180 23336 23208
rect 28261 23205 28273 23239
rect 28307 23236 28319 23239
rect 28534 23236 28540 23248
rect 28307 23208 28540 23236
rect 28307 23205 28319 23208
rect 28261 23199 28319 23205
rect 28534 23196 28540 23208
rect 28592 23236 28598 23248
rect 29012 23236 29040 23276
rect 28592 23208 29040 23236
rect 28592 23196 28598 23208
rect 29914 23196 29920 23248
rect 29972 23196 29978 23248
rect 20680 23140 22094 23168
rect 20680 23128 20686 23140
rect 22922 23128 22928 23180
rect 22980 23168 22986 23180
rect 23017 23171 23075 23177
rect 23017 23168 23029 23171
rect 22980 23140 23029 23168
rect 22980 23128 22986 23140
rect 23017 23137 23029 23140
rect 23063 23168 23075 23171
rect 23106 23168 23112 23180
rect 23063 23140 23112 23168
rect 23063 23137 23075 23140
rect 23017 23131 23075 23137
rect 23106 23128 23112 23140
rect 23164 23128 23170 23180
rect 23290 23128 23296 23180
rect 23348 23128 23354 23180
rect 25866 23128 25872 23180
rect 25924 23168 25930 23180
rect 26513 23171 26571 23177
rect 26513 23168 26525 23171
rect 25924 23140 26525 23168
rect 25924 23128 25930 23140
rect 26513 23137 26525 23140
rect 26559 23137 26571 23171
rect 26513 23131 26571 23137
rect 26789 23171 26847 23177
rect 26789 23137 26801 23171
rect 26835 23168 26847 23171
rect 27246 23168 27252 23180
rect 26835 23140 27252 23168
rect 26835 23137 26847 23140
rect 26789 23131 26847 23137
rect 27246 23128 27252 23140
rect 27304 23128 27310 23180
rect 27982 23128 27988 23180
rect 28040 23128 28046 23180
rect 28902 23128 28908 23180
rect 28960 23128 28966 23180
rect 29932 23168 29960 23196
rect 30392 23177 30420 23276
rect 30650 23264 30656 23316
rect 30708 23264 30714 23316
rect 30668 23236 30696 23264
rect 30484 23208 30696 23236
rect 29288 23140 29960 23168
rect 30009 23171 30067 23177
rect 19613 23103 19671 23109
rect 19613 23100 19625 23103
rect 19076 23072 19625 23100
rect 19613 23069 19625 23072
rect 19659 23069 19671 23103
rect 19613 23063 19671 23069
rect 19886 23060 19892 23112
rect 19944 23060 19950 23112
rect 22189 23103 22247 23109
rect 22189 23069 22201 23103
rect 22235 23100 22247 23103
rect 22646 23100 22652 23112
rect 22235 23072 22652 23100
rect 22235 23069 22247 23072
rect 22189 23063 22247 23069
rect 22646 23060 22652 23072
rect 22704 23060 22710 23112
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 24118 23100 24124 23112
rect 22879 23072 24124 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 24118 23060 24124 23072
rect 24176 23060 24182 23112
rect 24670 23060 24676 23112
rect 24728 23060 24734 23112
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 25130 23100 25136 23112
rect 24995 23072 25136 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 25130 23060 25136 23072
rect 25188 23060 25194 23112
rect 28000 23100 28028 23128
rect 27922 23072 28028 23100
rect 28813 23103 28871 23109
rect 28813 23069 28825 23103
rect 28859 23100 28871 23103
rect 29086 23100 29092 23112
rect 28859 23072 29092 23100
rect 28859 23069 28871 23072
rect 28813 23063 28871 23069
rect 29086 23060 29092 23072
rect 29144 23100 29150 23112
rect 29288 23100 29316 23140
rect 30009 23137 30021 23171
rect 30055 23168 30067 23171
rect 30377 23171 30435 23177
rect 30055 23140 30144 23168
rect 30055 23137 30067 23140
rect 30009 23131 30067 23137
rect 29144 23072 29316 23100
rect 29917 23103 29975 23109
rect 29144 23060 29150 23072
rect 29917 23069 29929 23103
rect 29963 23100 29975 23103
rect 30116 23100 30144 23140
rect 30377 23137 30389 23171
rect 30423 23137 30435 23171
rect 30377 23131 30435 23137
rect 30484 23100 30512 23208
rect 30653 23171 30711 23177
rect 30653 23137 30665 23171
rect 30699 23168 30711 23171
rect 31205 23171 31263 23177
rect 31205 23168 31217 23171
rect 30699 23140 31217 23168
rect 30699 23137 30711 23140
rect 30653 23131 30711 23137
rect 31205 23137 31217 23140
rect 31251 23137 31263 23171
rect 31205 23131 31263 23137
rect 29963 23072 30052 23100
rect 30116 23072 30512 23100
rect 29963 23069 29975 23072
rect 29917 23063 29975 23069
rect 15856 23004 15976 23032
rect 15856 22976 15884 23004
rect 16758 22992 16764 23044
rect 16816 22992 16822 23044
rect 17865 23035 17923 23041
rect 17865 23001 17877 23035
rect 17911 23032 17923 23035
rect 18230 23032 18236 23044
rect 17911 23004 18236 23032
rect 17911 23001 17923 23004
rect 17865 22995 17923 23001
rect 18230 22992 18236 23004
rect 18288 22992 18294 23044
rect 18874 22992 18880 23044
rect 18932 23041 18938 23044
rect 18932 23035 18960 23041
rect 18948 23001 18960 23035
rect 20165 23035 20223 23041
rect 20165 23032 20177 23035
rect 18932 22995 18960 23001
rect 19812 23004 20177 23032
rect 18932 22992 18938 22995
rect 6638 22964 6644 22976
rect 5736 22936 6644 22964
rect 5169 22927 5227 22933
rect 6638 22924 6644 22936
rect 6696 22924 6702 22976
rect 7423 22967 7481 22973
rect 7423 22933 7435 22967
rect 7469 22964 7481 22967
rect 7742 22964 7748 22976
rect 7469 22936 7748 22964
rect 7469 22933 7481 22936
rect 7423 22927 7481 22933
rect 7742 22924 7748 22936
rect 7800 22924 7806 22976
rect 8754 22924 8760 22976
rect 8812 22964 8818 22976
rect 9493 22967 9551 22973
rect 9493 22964 9505 22967
rect 8812 22936 9505 22964
rect 8812 22924 8818 22936
rect 9493 22933 9505 22936
rect 9539 22933 9551 22967
rect 9493 22927 9551 22933
rect 11054 22924 11060 22976
rect 11112 22964 11118 22976
rect 12526 22964 12532 22976
rect 11112 22936 12532 22964
rect 11112 22924 11118 22936
rect 12526 22924 12532 22936
rect 12584 22924 12590 22976
rect 14185 22967 14243 22973
rect 14185 22933 14197 22967
rect 14231 22964 14243 22967
rect 15378 22964 15384 22976
rect 14231 22936 15384 22964
rect 14231 22933 14243 22936
rect 14185 22927 14243 22933
rect 15378 22924 15384 22936
rect 15436 22924 15442 22976
rect 15838 22924 15844 22976
rect 15896 22924 15902 22976
rect 17310 22924 17316 22976
rect 17368 22964 17374 22976
rect 18693 22967 18751 22973
rect 18693 22964 18705 22967
rect 17368 22936 18705 22964
rect 17368 22924 17374 22936
rect 18693 22933 18705 22936
rect 18739 22964 18751 22967
rect 19702 22964 19708 22976
rect 18739 22936 19708 22964
rect 18739 22933 18751 22936
rect 18693 22927 18751 22933
rect 19702 22924 19708 22936
rect 19760 22924 19766 22976
rect 19812 22973 19840 23004
rect 20165 23001 20177 23004
rect 20211 23001 20223 23035
rect 20622 23032 20628 23044
rect 20165 22995 20223 23001
rect 20272 23004 20628 23032
rect 19797 22967 19855 22973
rect 19797 22933 19809 22967
rect 19843 22933 19855 22967
rect 19797 22927 19855 22933
rect 20070 22924 20076 22976
rect 20128 22964 20134 22976
rect 20272 22964 20300 23004
rect 20622 22992 20628 23004
rect 20680 22992 20686 23044
rect 22281 23035 22339 23041
rect 22281 23001 22293 23035
rect 22327 23032 22339 23035
rect 24688 23032 24716 23060
rect 22327 23004 24716 23032
rect 28721 23035 28779 23041
rect 22327 23001 22339 23004
rect 22281 22995 22339 23001
rect 28721 23001 28733 23035
rect 28767 23032 28779 23035
rect 28767 23004 29592 23032
rect 28767 23001 28779 23004
rect 28721 22995 28779 23001
rect 20128 22936 20300 22964
rect 20128 22924 20134 22936
rect 22922 22924 22928 22976
rect 22980 22924 22986 22976
rect 29564 22973 29592 23004
rect 30024 22976 30052 23072
rect 31110 23060 31116 23112
rect 31168 23060 31174 23112
rect 31294 23060 31300 23112
rect 31352 23060 31358 23112
rect 30834 22992 30840 23044
rect 30892 23041 30898 23044
rect 30892 23035 30920 23041
rect 30908 23001 30920 23035
rect 30892 22995 30920 23001
rect 30892 22992 30898 22995
rect 29549 22967 29607 22973
rect 29549 22933 29561 22967
rect 29595 22933 29607 22967
rect 29549 22927 29607 22933
rect 30006 22924 30012 22976
rect 30064 22924 30070 22976
rect 30742 22924 30748 22976
rect 30800 22924 30806 22976
rect 31021 22967 31079 22973
rect 31021 22933 31033 22967
rect 31067 22964 31079 22967
rect 31110 22964 31116 22976
rect 31067 22936 31116 22964
rect 31067 22933 31079 22936
rect 31021 22927 31079 22933
rect 31110 22924 31116 22936
rect 31168 22924 31174 22976
rect 1104 22874 34840 22896
rect 1104 22822 9344 22874
rect 9396 22822 9408 22874
rect 9460 22822 9472 22874
rect 9524 22822 9536 22874
rect 9588 22822 9600 22874
rect 9652 22822 17738 22874
rect 17790 22822 17802 22874
rect 17854 22822 17866 22874
rect 17918 22822 17930 22874
rect 17982 22822 17994 22874
rect 18046 22822 26132 22874
rect 26184 22822 26196 22874
rect 26248 22822 26260 22874
rect 26312 22822 26324 22874
rect 26376 22822 26388 22874
rect 26440 22822 34526 22874
rect 34578 22822 34590 22874
rect 34642 22822 34654 22874
rect 34706 22822 34718 22874
rect 34770 22822 34782 22874
rect 34834 22822 34840 22874
rect 1104 22800 34840 22822
rect 13170 22760 13176 22772
rect 11992 22732 13176 22760
rect 6638 22652 6644 22704
rect 6696 22692 6702 22704
rect 6696 22664 7774 22692
rect 6696 22652 6702 22664
rect 5442 22584 5448 22636
rect 5500 22624 5506 22636
rect 11992 22633 12020 22732
rect 13170 22720 13176 22732
rect 13228 22720 13234 22772
rect 15654 22720 15660 22772
rect 15712 22720 15718 22772
rect 16390 22720 16396 22772
rect 16448 22760 16454 22772
rect 16669 22763 16727 22769
rect 16669 22760 16681 22763
rect 16448 22732 16681 22760
rect 16448 22720 16454 22732
rect 16669 22729 16681 22732
rect 16715 22729 16727 22763
rect 16669 22723 16727 22729
rect 16853 22763 16911 22769
rect 16853 22729 16865 22763
rect 16899 22760 16911 22763
rect 17405 22763 17463 22769
rect 17405 22760 17417 22763
rect 16899 22732 17417 22760
rect 16899 22729 16911 22732
rect 16853 22723 16911 22729
rect 17405 22729 17417 22732
rect 17451 22729 17463 22763
rect 17405 22723 17463 22729
rect 17494 22720 17500 22772
rect 17552 22720 17558 22772
rect 18785 22763 18843 22769
rect 18785 22729 18797 22763
rect 18831 22760 18843 22763
rect 18874 22760 18880 22772
rect 18831 22732 18880 22760
rect 18831 22729 18843 22732
rect 18785 22723 18843 22729
rect 18874 22720 18880 22732
rect 18932 22720 18938 22772
rect 19242 22720 19248 22772
rect 19300 22720 19306 22772
rect 29365 22763 29423 22769
rect 29365 22729 29377 22763
rect 29411 22760 29423 22763
rect 29730 22760 29736 22772
rect 29411 22732 29736 22760
rect 29411 22729 29423 22732
rect 29365 22723 29423 22729
rect 29730 22720 29736 22732
rect 29788 22720 29794 22772
rect 29914 22720 29920 22772
rect 29972 22720 29978 22772
rect 30009 22763 30067 22769
rect 30009 22729 30021 22763
rect 30055 22760 30067 22763
rect 30742 22760 30748 22772
rect 30055 22732 30748 22760
rect 30055 22729 30067 22732
rect 30009 22723 30067 22729
rect 30742 22720 30748 22732
rect 30800 22720 30806 22772
rect 31110 22720 31116 22772
rect 31168 22720 31174 22772
rect 14366 22692 14372 22704
rect 13478 22664 14372 22692
rect 14366 22652 14372 22664
rect 14424 22652 14430 22704
rect 7009 22627 7067 22633
rect 7009 22624 7021 22627
rect 5500 22596 7021 22624
rect 5500 22584 5506 22596
rect 7009 22593 7021 22596
rect 7055 22593 7067 22627
rect 7009 22587 7067 22593
rect 11977 22627 12035 22633
rect 11977 22593 11989 22627
rect 12023 22593 12035 22627
rect 11977 22587 12035 22593
rect 7024 22420 7052 22587
rect 7282 22516 7288 22568
rect 7340 22516 7346 22568
rect 7650 22516 7656 22568
rect 7708 22556 7714 22568
rect 9033 22559 9091 22565
rect 9033 22556 9045 22559
rect 7708 22528 9045 22556
rect 7708 22516 7714 22528
rect 9033 22525 9045 22528
rect 9079 22525 9091 22559
rect 9033 22519 9091 22525
rect 12250 22516 12256 22568
rect 12308 22516 12314 22568
rect 12802 22516 12808 22568
rect 12860 22556 12866 22568
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 12860 22528 14013 22556
rect 12860 22516 12866 22528
rect 14001 22525 14013 22528
rect 14047 22525 14059 22559
rect 14001 22519 14059 22525
rect 8294 22420 8300 22432
rect 7024 22392 8300 22420
rect 8294 22380 8300 22392
rect 8352 22420 8358 22432
rect 9306 22420 9312 22432
rect 8352 22392 9312 22420
rect 8352 22380 8358 22392
rect 9306 22380 9312 22392
rect 9364 22380 9370 22432
rect 15672 22420 15700 22720
rect 16942 22652 16948 22704
rect 17000 22692 17006 22704
rect 17310 22692 17316 22704
rect 17000 22664 17316 22692
rect 17000 22652 17006 22664
rect 17310 22652 17316 22664
rect 17368 22652 17374 22704
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 16669 22627 16727 22633
rect 16669 22624 16681 22627
rect 16632 22596 16681 22624
rect 16632 22584 16638 22596
rect 16669 22593 16681 22596
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22624 17095 22627
rect 17512 22624 17540 22720
rect 19153 22695 19211 22701
rect 19153 22692 19165 22695
rect 18156 22664 19165 22692
rect 18156 22636 18184 22664
rect 19153 22661 19165 22664
rect 19199 22661 19211 22695
rect 21634 22692 21640 22704
rect 19153 22655 19211 22661
rect 19628 22664 21640 22692
rect 17083 22596 17540 22624
rect 17083 22593 17095 22596
rect 17037 22587 17095 22593
rect 18138 22584 18144 22636
rect 18196 22584 18202 22636
rect 18969 22627 19027 22633
rect 18969 22593 18981 22627
rect 19015 22624 19027 22627
rect 19168 22624 19196 22655
rect 19628 22633 19656 22664
rect 21634 22652 21640 22664
rect 21692 22652 21698 22704
rect 19429 22627 19487 22633
rect 19429 22624 19441 22627
rect 19015 22596 19104 22624
rect 19168 22596 19441 22624
rect 19015 22593 19027 22596
rect 18969 22587 19027 22593
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22556 18107 22559
rect 18230 22556 18236 22568
rect 18095 22528 18236 22556
rect 18095 22525 18107 22528
rect 18049 22519 18107 22525
rect 18230 22516 18236 22528
rect 18288 22556 18294 22568
rect 19076 22556 19104 22596
rect 19429 22593 19441 22596
rect 19475 22593 19487 22627
rect 19429 22587 19487 22593
rect 19613 22627 19671 22633
rect 19613 22593 19625 22627
rect 19659 22593 19671 22627
rect 19613 22587 19671 22593
rect 19628 22556 19656 22587
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 20809 22627 20867 22633
rect 20809 22624 20821 22627
rect 20772 22596 20821 22624
rect 20772 22584 20778 22596
rect 20809 22593 20821 22596
rect 20855 22593 20867 22627
rect 20990 22624 20996 22636
rect 20809 22587 20867 22593
rect 20916 22596 20996 22624
rect 20916 22565 20944 22596
rect 20990 22584 20996 22596
rect 21048 22624 21054 22636
rect 24394 22624 24400 22636
rect 21048 22596 24400 22624
rect 21048 22584 21054 22596
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 28626 22584 28632 22636
rect 28684 22624 28690 22636
rect 29273 22627 29331 22633
rect 29273 22624 29285 22627
rect 28684 22596 29285 22624
rect 28684 22584 28690 22596
rect 29273 22593 29285 22596
rect 29319 22593 29331 22627
rect 29748 22624 29776 22720
rect 29932 22692 29960 22720
rect 31128 22692 31156 22720
rect 31205 22695 31263 22701
rect 31205 22692 31217 22695
rect 29932 22664 30144 22692
rect 31128 22664 31217 22692
rect 30116 22633 30144 22664
rect 31205 22661 31217 22664
rect 31251 22661 31263 22695
rect 31205 22655 31263 22661
rect 29917 22627 29975 22633
rect 29917 22624 29929 22627
rect 29748 22596 29929 22624
rect 29273 22587 29331 22593
rect 29917 22593 29929 22596
rect 29963 22593 29975 22627
rect 29917 22587 29975 22593
rect 30101 22627 30159 22633
rect 30101 22593 30113 22627
rect 30147 22593 30159 22627
rect 32950 22624 32956 22636
rect 32890 22596 32956 22624
rect 30101 22587 30159 22593
rect 32950 22584 32956 22596
rect 33008 22584 33014 22636
rect 18288 22528 19012 22556
rect 19076 22528 19656 22556
rect 20901 22559 20959 22565
rect 18288 22516 18294 22528
rect 18984 22500 19012 22528
rect 20901 22525 20913 22559
rect 20947 22525 20959 22559
rect 20901 22519 20959 22525
rect 24765 22559 24823 22565
rect 24765 22525 24777 22559
rect 24811 22556 24823 22559
rect 24946 22556 24952 22568
rect 24811 22528 24952 22556
rect 24811 22525 24823 22528
rect 24765 22519 24823 22525
rect 24946 22516 24952 22528
rect 25004 22516 25010 22568
rect 28721 22559 28779 22565
rect 28721 22525 28733 22559
rect 28767 22556 28779 22559
rect 29086 22556 29092 22568
rect 28767 22528 29092 22556
rect 28767 22525 28779 22528
rect 28721 22519 28779 22525
rect 29086 22516 29092 22528
rect 29144 22516 29150 22568
rect 30006 22516 30012 22568
rect 30064 22516 30070 22568
rect 32214 22516 32220 22568
rect 32272 22556 32278 22568
rect 33965 22559 34023 22565
rect 33965 22556 33977 22559
rect 32272 22528 33977 22556
rect 32272 22516 32278 22528
rect 33965 22525 33977 22528
rect 34011 22525 34023 22559
rect 34241 22559 34299 22565
rect 34241 22556 34253 22559
rect 33965 22519 34023 22525
rect 34164 22528 34253 22556
rect 18966 22448 18972 22500
rect 19024 22448 19030 22500
rect 21174 22448 21180 22500
rect 21232 22448 21238 22500
rect 28997 22491 29055 22497
rect 28997 22457 29009 22491
rect 29043 22488 29055 22491
rect 30024 22488 30052 22516
rect 29043 22460 30052 22488
rect 31389 22491 31447 22497
rect 29043 22457 29055 22460
rect 28997 22451 29055 22457
rect 31389 22457 31401 22491
rect 31435 22488 31447 22491
rect 32122 22488 32128 22500
rect 31435 22460 32128 22488
rect 31435 22457 31447 22460
rect 31389 22451 31447 22457
rect 32122 22448 32128 22460
rect 32180 22448 32186 22500
rect 32416 22460 32996 22488
rect 23566 22420 23572 22432
rect 15672 22392 23572 22420
rect 23566 22380 23572 22392
rect 23624 22380 23630 22432
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 24121 22423 24179 22429
rect 24121 22420 24133 22423
rect 23716 22392 24133 22420
rect 23716 22380 23722 22392
rect 24121 22389 24133 22392
rect 24167 22389 24179 22423
rect 24121 22383 24179 22389
rect 29730 22380 29736 22432
rect 29788 22420 29794 22432
rect 32416 22420 32444 22460
rect 29788 22392 32444 22420
rect 29788 22380 29794 22392
rect 32490 22380 32496 22432
rect 32548 22380 32554 22432
rect 32968 22420 32996 22460
rect 34164 22420 34192 22528
rect 34241 22525 34253 22528
rect 34287 22525 34299 22559
rect 34241 22519 34299 22525
rect 34330 22420 34336 22432
rect 32968 22392 34336 22420
rect 34330 22380 34336 22392
rect 34388 22380 34394 22432
rect 1104 22330 34684 22352
rect 1104 22278 5147 22330
rect 5199 22278 5211 22330
rect 5263 22278 5275 22330
rect 5327 22278 5339 22330
rect 5391 22278 5403 22330
rect 5455 22278 13541 22330
rect 13593 22278 13605 22330
rect 13657 22278 13669 22330
rect 13721 22278 13733 22330
rect 13785 22278 13797 22330
rect 13849 22278 21935 22330
rect 21987 22278 21999 22330
rect 22051 22278 22063 22330
rect 22115 22278 22127 22330
rect 22179 22278 22191 22330
rect 22243 22278 30329 22330
rect 30381 22278 30393 22330
rect 30445 22278 30457 22330
rect 30509 22278 30521 22330
rect 30573 22278 30585 22330
rect 30637 22278 34684 22330
rect 1104 22256 34684 22278
rect 5994 22176 6000 22228
rect 6052 22216 6058 22228
rect 6181 22219 6239 22225
rect 6181 22216 6193 22219
rect 6052 22188 6193 22216
rect 6052 22176 6058 22188
rect 6181 22185 6193 22188
rect 6227 22185 6239 22219
rect 6181 22179 6239 22185
rect 12161 22219 12219 22225
rect 12161 22185 12173 22219
rect 12207 22216 12219 22219
rect 12250 22216 12256 22228
rect 12207 22188 12256 22216
rect 12207 22185 12219 22188
rect 12161 22179 12219 22185
rect 12250 22176 12256 22188
rect 12308 22176 12314 22228
rect 15583 22219 15641 22225
rect 15583 22185 15595 22219
rect 15629 22216 15641 22219
rect 24302 22216 24308 22228
rect 15629 22188 24308 22216
rect 15629 22185 15641 22188
rect 15583 22179 15641 22185
rect 24302 22176 24308 22188
rect 24360 22176 24366 22228
rect 24946 22176 24952 22228
rect 25004 22216 25010 22228
rect 25004 22188 26234 22216
rect 25004 22176 25010 22188
rect 12526 22108 12532 22160
rect 12584 22148 12590 22160
rect 14366 22148 14372 22160
rect 12584 22120 14372 22148
rect 12584 22108 12590 22120
rect 14366 22108 14372 22120
rect 14424 22108 14430 22160
rect 6549 22083 6607 22089
rect 6549 22080 6561 22083
rect 5460 22052 6561 22080
rect 5460 22024 5488 22052
rect 6549 22049 6561 22052
rect 6595 22080 6607 22083
rect 6595 22052 8156 22080
rect 6595 22049 6607 22052
rect 6549 22043 6607 22049
rect 1946 21972 1952 22024
rect 2004 22012 2010 22024
rect 3789 22015 3847 22021
rect 3789 22012 3801 22015
rect 2004 21984 3801 22012
rect 2004 21972 2010 21984
rect 3789 21981 3801 21984
rect 3835 21981 3847 22015
rect 3789 21975 3847 21981
rect 5442 21972 5448 22024
rect 5500 21972 5506 22024
rect 6362 21972 6368 22024
rect 6420 21972 6426 22024
rect 6641 22015 6699 22021
rect 6641 21981 6653 22015
rect 6687 22012 6699 22015
rect 7101 22015 7159 22021
rect 7101 22012 7113 22015
rect 6687 21984 7113 22012
rect 6687 21981 6699 21984
rect 6641 21975 6699 21981
rect 7101 21981 7113 21984
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 7742 21972 7748 22024
rect 7800 21972 7806 22024
rect 8128 22012 8156 22052
rect 8202 22040 8208 22092
rect 8260 22040 8266 22092
rect 8665 22083 8723 22089
rect 8665 22080 8677 22083
rect 8312 22052 8677 22080
rect 8312 22012 8340 22052
rect 8665 22049 8677 22052
rect 8711 22049 8723 22083
rect 8665 22043 8723 22049
rect 9306 22040 9312 22092
rect 9364 22040 9370 22092
rect 12713 22083 12771 22089
rect 12713 22080 12725 22083
rect 12406 22052 12725 22080
rect 8128 21984 8340 22012
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 8541 22015 8599 22021
rect 8444 21984 8489 22012
rect 8444 21972 8450 21984
rect 8541 21981 8553 22015
rect 8587 22012 8599 22015
rect 8587 21984 8708 22012
rect 8587 21981 8599 21984
rect 8541 21975 8599 21981
rect 2682 21904 2688 21956
rect 2740 21904 2746 21956
rect 4065 21947 4123 21953
rect 4065 21913 4077 21947
rect 4111 21944 4123 21947
rect 4338 21944 4344 21956
rect 4111 21916 4344 21944
rect 4111 21913 4123 21916
rect 4065 21907 4123 21913
rect 4338 21904 4344 21916
rect 4396 21904 4402 21956
rect 4522 21944 4528 21956
rect 4448 21916 4528 21944
rect 2700 21876 2728 21904
rect 4448 21876 4476 21916
rect 4522 21904 4528 21916
rect 4580 21904 4586 21956
rect 5350 21904 5356 21956
rect 5408 21944 5414 21956
rect 5810 21944 5816 21956
rect 5408 21916 5816 21944
rect 5408 21904 5414 21916
rect 5810 21904 5816 21916
rect 5868 21904 5874 21956
rect 2700 21848 4476 21876
rect 8680 21876 8708 21984
rect 8754 21972 8760 22024
rect 8812 21972 8818 22024
rect 11054 22012 11060 22024
rect 10718 21984 11060 22012
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 22012 12035 22015
rect 12406 22012 12434 22052
rect 12713 22049 12725 22052
rect 12759 22049 12771 22083
rect 12713 22043 12771 22049
rect 23106 22040 23112 22092
rect 23164 22040 23170 22092
rect 24854 22080 24860 22092
rect 23400 22052 24860 22080
rect 12023 21984 12434 22012
rect 12621 22015 12679 22021
rect 12023 21981 12035 21984
rect 11977 21975 12035 21981
rect 12621 21981 12633 22015
rect 12667 22012 12679 22015
rect 12897 22015 12955 22021
rect 12897 22012 12909 22015
rect 12667 21984 12909 22012
rect 12667 21981 12679 21984
rect 12621 21975 12679 21981
rect 12897 21981 12909 21984
rect 12943 21981 12955 22015
rect 12897 21975 12955 21981
rect 12986 21972 12992 22024
rect 13044 21972 13050 22024
rect 14274 21972 14280 22024
rect 14332 22012 14338 22024
rect 14332 21998 14490 22012
rect 14332 21984 14504 21998
rect 14332 21972 14338 21984
rect 9214 21904 9220 21956
rect 9272 21944 9278 21956
rect 9585 21947 9643 21953
rect 9585 21944 9597 21947
rect 9272 21916 9597 21944
rect 9272 21904 9278 21916
rect 9585 21913 9597 21916
rect 9631 21913 9643 21947
rect 9585 21907 9643 21913
rect 11330 21904 11336 21956
rect 11388 21904 11394 21956
rect 12253 21947 12311 21953
rect 12253 21913 12265 21947
rect 12299 21913 12311 21947
rect 12253 21907 12311 21913
rect 12437 21947 12495 21953
rect 12437 21913 12449 21947
rect 12483 21944 12495 21947
rect 12802 21944 12808 21956
rect 12483 21916 12808 21944
rect 12483 21913 12495 21916
rect 12437 21907 12495 21913
rect 9950 21876 9956 21888
rect 8680 21848 9956 21876
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 12268 21876 12296 21907
rect 12802 21904 12808 21916
rect 12860 21904 12866 21956
rect 12710 21876 12716 21888
rect 12268 21848 12716 21876
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 14090 21836 14096 21888
rect 14148 21836 14154 21888
rect 14476 21876 14504 21984
rect 15838 21972 15844 22024
rect 15896 21972 15902 22024
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 18969 22015 19027 22021
rect 18969 22012 18981 22015
rect 18288 21984 18981 22012
rect 18288 21972 18294 21984
rect 18969 21981 18981 21984
rect 19015 21981 19027 22015
rect 18969 21975 19027 21981
rect 23014 21972 23020 22024
rect 23072 22012 23078 22024
rect 23400 22012 23428 22052
rect 24854 22040 24860 22052
rect 24912 22040 24918 22092
rect 26206 22080 26234 22188
rect 32214 22176 32220 22228
rect 32272 22176 32278 22228
rect 33410 22108 33416 22160
rect 33468 22148 33474 22160
rect 33468 22120 33548 22148
rect 33468 22108 33474 22120
rect 28261 22083 28319 22089
rect 28261 22080 28273 22083
rect 26206 22052 28273 22080
rect 28261 22049 28273 22052
rect 28307 22049 28319 22083
rect 32490 22080 32496 22092
rect 28261 22043 28319 22049
rect 31312 22052 32496 22080
rect 23072 21984 23428 22012
rect 23072 21972 23078 21984
rect 23658 21972 23664 22024
rect 23716 21972 23722 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 17494 21904 17500 21956
rect 17552 21944 17558 21956
rect 23385 21947 23443 21953
rect 17552 21916 22094 21944
rect 17552 21904 17558 21916
rect 14734 21876 14740 21888
rect 14476 21848 14740 21876
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 18598 21836 18604 21888
rect 18656 21876 18662 21888
rect 18785 21879 18843 21885
rect 18785 21876 18797 21879
rect 18656 21848 18797 21876
rect 18656 21836 18662 21848
rect 18785 21845 18797 21848
rect 18831 21845 18843 21879
rect 18785 21839 18843 21845
rect 19702 21836 19708 21888
rect 19760 21876 19766 21888
rect 20622 21876 20628 21888
rect 19760 21848 20628 21876
rect 19760 21836 19766 21848
rect 20622 21836 20628 21848
rect 20680 21836 20686 21888
rect 22066 21876 22094 21916
rect 23385 21913 23397 21947
rect 23431 21944 23443 21947
rect 23676 21944 23704 21972
rect 24044 21944 24072 21975
rect 24578 21972 24584 22024
rect 24636 21972 24642 22024
rect 30282 21972 30288 22024
rect 30340 22012 30346 22024
rect 31312 22021 31340 22052
rect 32490 22040 32496 22052
rect 32548 22080 32554 22092
rect 33520 22089 33548 22120
rect 33321 22083 33379 22089
rect 33321 22080 33333 22083
rect 32548 22052 33333 22080
rect 32548 22040 32554 22052
rect 33321 22049 33333 22052
rect 33367 22049 33379 22083
rect 33321 22043 33379 22049
rect 33505 22083 33563 22089
rect 33505 22049 33517 22083
rect 33551 22080 33563 22083
rect 33551 22052 33585 22080
rect 33551 22049 33563 22052
rect 33505 22043 33563 22049
rect 31297 22015 31355 22021
rect 31297 22012 31309 22015
rect 30340 21984 31309 22012
rect 30340 21972 30346 21984
rect 31297 21981 31309 21984
rect 31343 21981 31355 22015
rect 31297 21975 31355 21981
rect 31662 21972 31668 22024
rect 31720 21972 31726 22024
rect 32401 22015 32459 22021
rect 32401 21981 32413 22015
rect 32447 21981 32459 22015
rect 32401 21975 32459 21981
rect 25133 21947 25191 21953
rect 25133 21944 25145 21947
rect 23431 21916 23704 21944
rect 23768 21916 24072 21944
rect 24780 21916 25145 21944
rect 23431 21913 23443 21916
rect 23385 21907 23443 21913
rect 23198 21876 23204 21888
rect 22066 21848 23204 21876
rect 23198 21836 23204 21848
rect 23256 21836 23262 21888
rect 23290 21836 23296 21888
rect 23348 21836 23354 21888
rect 23768 21885 23796 21916
rect 23753 21879 23811 21885
rect 23753 21845 23765 21879
rect 23799 21845 23811 21879
rect 23753 21839 23811 21845
rect 23842 21836 23848 21888
rect 23900 21836 23906 21888
rect 24780 21885 24808 21916
rect 25133 21913 25145 21916
rect 25179 21913 25191 21947
rect 25133 21907 25191 21913
rect 25332 21916 25622 21944
rect 25332 21888 25360 21916
rect 31478 21904 31484 21956
rect 31536 21904 31542 21956
rect 31573 21947 31631 21953
rect 31573 21913 31585 21947
rect 31619 21913 31631 21947
rect 31573 21907 31631 21913
rect 24765 21879 24823 21885
rect 24765 21845 24777 21879
rect 24811 21845 24823 21879
rect 24765 21839 24823 21845
rect 25314 21836 25320 21888
rect 25372 21836 25378 21888
rect 26602 21836 26608 21888
rect 26660 21876 26666 21888
rect 28626 21876 28632 21888
rect 26660 21848 28632 21876
rect 26660 21836 26666 21848
rect 28626 21836 28632 21848
rect 28684 21836 28690 21888
rect 28905 21879 28963 21885
rect 28905 21845 28917 21879
rect 28951 21876 28963 21879
rect 31588 21876 31616 21907
rect 28951 21848 31616 21876
rect 31849 21879 31907 21885
rect 28951 21845 28963 21848
rect 28905 21839 28963 21845
rect 31849 21845 31861 21879
rect 31895 21876 31907 21879
rect 32416 21876 32444 21975
rect 32674 21972 32680 22024
rect 32732 21972 32738 22024
rect 31895 21848 32444 21876
rect 31895 21845 31907 21848
rect 31849 21839 31907 21845
rect 32582 21836 32588 21888
rect 32640 21836 32646 21888
rect 32766 21836 32772 21888
rect 32824 21876 32830 21888
rect 32861 21879 32919 21885
rect 32861 21876 32873 21879
rect 32824 21848 32873 21876
rect 32824 21836 32830 21848
rect 32861 21845 32873 21848
rect 32907 21845 32919 21879
rect 32861 21839 32919 21845
rect 33226 21836 33232 21888
rect 33284 21836 33290 21888
rect 1104 21786 34840 21808
rect 1104 21734 9344 21786
rect 9396 21734 9408 21786
rect 9460 21734 9472 21786
rect 9524 21734 9536 21786
rect 9588 21734 9600 21786
rect 9652 21734 17738 21786
rect 17790 21734 17802 21786
rect 17854 21734 17866 21786
rect 17918 21734 17930 21786
rect 17982 21734 17994 21786
rect 18046 21734 26132 21786
rect 26184 21734 26196 21786
rect 26248 21734 26260 21786
rect 26312 21734 26324 21786
rect 26376 21734 26388 21786
rect 26440 21734 34526 21786
rect 34578 21734 34590 21786
rect 34642 21734 34654 21786
rect 34706 21734 34718 21786
rect 34770 21734 34782 21786
rect 34834 21734 34840 21786
rect 1104 21712 34840 21734
rect 4338 21632 4344 21684
rect 4396 21672 4402 21684
rect 4801 21675 4859 21681
rect 4801 21672 4813 21675
rect 4396 21644 4813 21672
rect 4396 21632 4402 21644
rect 4801 21641 4813 21644
rect 4847 21641 4859 21675
rect 4801 21635 4859 21641
rect 7193 21675 7251 21681
rect 7193 21641 7205 21675
rect 7239 21672 7251 21675
rect 7282 21672 7288 21684
rect 7239 21644 7288 21672
rect 7239 21641 7251 21644
rect 7193 21635 7251 21641
rect 7282 21632 7288 21644
rect 7340 21632 7346 21684
rect 8386 21672 8392 21684
rect 7392 21644 8392 21672
rect 7392 21604 7420 21644
rect 8386 21632 8392 21644
rect 8444 21672 8450 21684
rect 8444 21644 9168 21672
rect 8444 21632 8450 21644
rect 7929 21607 7987 21613
rect 7929 21604 7941 21607
rect 4724 21576 7420 21604
rect 4724 21548 4752 21576
rect 4706 21496 4712 21548
rect 4764 21496 4770 21548
rect 5092 21545 5120 21576
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21505 5043 21539
rect 4985 21499 5043 21505
rect 5077 21539 5135 21545
rect 5077 21505 5089 21539
rect 5123 21505 5135 21539
rect 5077 21499 5135 21505
rect 5000 21468 5028 21499
rect 5350 21496 5356 21548
rect 5408 21496 5414 21548
rect 5534 21496 5540 21548
rect 5592 21496 5598 21548
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21505 5779 21539
rect 5721 21499 5779 21505
rect 5629 21471 5687 21477
rect 5629 21468 5641 21471
rect 5000 21440 5641 21468
rect 5629 21437 5641 21440
rect 5675 21437 5687 21471
rect 5629 21431 5687 21437
rect 5736 21400 5764 21499
rect 7282 21496 7288 21548
rect 7340 21536 7346 21548
rect 7392 21545 7420 21576
rect 7484 21576 7941 21604
rect 7484 21545 7512 21576
rect 7929 21573 7941 21576
rect 7975 21573 7987 21607
rect 7929 21567 7987 21573
rect 7377 21539 7435 21545
rect 7377 21536 7389 21539
rect 7340 21508 7389 21536
rect 7340 21496 7346 21508
rect 7377 21505 7389 21508
rect 7423 21505 7435 21539
rect 7377 21499 7435 21505
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21505 7527 21539
rect 7745 21539 7803 21545
rect 7745 21536 7757 21539
rect 7469 21499 7527 21505
rect 7576 21508 7757 21536
rect 7576 21480 7604 21508
rect 7745 21505 7757 21508
rect 7791 21505 7803 21539
rect 7745 21499 7803 21505
rect 7834 21496 7840 21548
rect 7892 21496 7898 21548
rect 8021 21539 8079 21545
rect 8021 21505 8033 21539
rect 8067 21505 8079 21539
rect 8021 21499 8079 21505
rect 7558 21428 7564 21480
rect 7616 21428 7622 21480
rect 5994 21400 6000 21412
rect 5736 21372 6000 21400
rect 5994 21360 6000 21372
rect 6052 21400 6058 21412
rect 8036 21400 8064 21499
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 9140 21468 9168 21644
rect 9214 21632 9220 21684
rect 9272 21672 9278 21684
rect 9585 21675 9643 21681
rect 9585 21672 9597 21675
rect 9272 21644 9597 21672
rect 9272 21632 9278 21644
rect 9585 21641 9597 21644
rect 9631 21641 9643 21675
rect 9585 21635 9643 21641
rect 9950 21632 9956 21684
rect 10008 21672 10014 21684
rect 10045 21675 10103 21681
rect 10045 21672 10057 21675
rect 10008 21644 10057 21672
rect 10008 21632 10014 21644
rect 10045 21641 10057 21644
rect 10091 21641 10103 21675
rect 12897 21675 12955 21681
rect 12897 21672 12909 21675
rect 10045 21635 10103 21641
rect 12360 21644 12909 21672
rect 12360 21613 12388 21644
rect 12897 21641 12909 21644
rect 12943 21672 12955 21675
rect 12986 21672 12992 21684
rect 12943 21644 12992 21672
rect 12943 21641 12955 21644
rect 12897 21635 12955 21641
rect 12986 21632 12992 21644
rect 13044 21632 13050 21684
rect 14090 21632 14096 21684
rect 14148 21672 14154 21684
rect 14148 21644 15332 21672
rect 14148 21632 14154 21644
rect 15304 21613 15332 21644
rect 15838 21632 15844 21684
rect 15896 21672 15902 21684
rect 19886 21672 19892 21684
rect 15896 21644 19892 21672
rect 15896 21632 15902 21644
rect 9769 21607 9827 21613
rect 9769 21604 9781 21607
rect 9324 21576 9781 21604
rect 9324 21545 9352 21576
rect 9769 21573 9781 21576
rect 9815 21573 9827 21607
rect 12345 21607 12403 21613
rect 9769 21567 9827 21573
rect 9876 21576 10180 21604
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21505 9367 21539
rect 9309 21499 9367 21505
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21505 9459 21539
rect 9401 21499 9459 21505
rect 9416 21468 9444 21499
rect 9674 21496 9680 21548
rect 9732 21496 9738 21548
rect 9876 21545 9904 21576
rect 10152 21545 10180 21576
rect 12345 21573 12357 21607
rect 12391 21573 12403 21607
rect 12345 21567 12403 21573
rect 12437 21607 12495 21613
rect 12437 21573 12449 21607
rect 12483 21604 12495 21607
rect 15289 21607 15347 21613
rect 12483 21576 12664 21604
rect 12483 21573 12495 21576
rect 12437 21567 12495 21573
rect 12636 21548 12664 21576
rect 15289 21573 15301 21607
rect 15335 21573 15347 21607
rect 15289 21567 15347 21573
rect 17494 21564 17500 21616
rect 17552 21564 17558 21616
rect 17862 21564 17868 21616
rect 17920 21564 17926 21616
rect 18138 21564 18144 21616
rect 18196 21564 18202 21616
rect 18230 21564 18236 21616
rect 18288 21564 18294 21616
rect 9861 21539 9919 21545
rect 9861 21505 9873 21539
rect 9907 21505 9919 21539
rect 9861 21499 9919 21505
rect 9953 21539 10011 21545
rect 9953 21505 9965 21539
rect 9999 21505 10011 21539
rect 9953 21499 10011 21505
rect 10137 21539 10195 21545
rect 10137 21505 10149 21539
rect 10183 21505 10195 21539
rect 10137 21499 10195 21505
rect 9140 21440 9444 21468
rect 9876 21400 9904 21499
rect 9968 21468 9996 21499
rect 10962 21496 10968 21548
rect 11020 21496 11026 21548
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 12529 21539 12587 21545
rect 12207 21508 12480 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 10980 21468 11008 21496
rect 9968 21440 11008 21468
rect 6052 21372 9904 21400
rect 6052 21360 6058 21372
rect 4798 21292 4804 21344
rect 4856 21332 4862 21344
rect 5261 21335 5319 21341
rect 5261 21332 5273 21335
rect 4856 21304 5273 21332
rect 4856 21292 4862 21304
rect 5261 21301 5273 21304
rect 5307 21332 5319 21335
rect 5442 21332 5448 21344
rect 5307 21304 5448 21332
rect 5307 21301 5319 21304
rect 5261 21295 5319 21301
rect 5442 21292 5448 21304
rect 5500 21332 5506 21344
rect 7653 21335 7711 21341
rect 7653 21332 7665 21335
rect 5500 21304 7665 21332
rect 5500 21292 5506 21304
rect 7653 21301 7665 21304
rect 7699 21332 7711 21335
rect 9125 21335 9183 21341
rect 9125 21332 9137 21335
rect 7699 21304 9137 21332
rect 7699 21301 7711 21304
rect 7653 21295 7711 21301
rect 9125 21301 9137 21304
rect 9171 21301 9183 21335
rect 9876 21332 9904 21372
rect 12452 21344 12480 21508
rect 12529 21505 12541 21539
rect 12575 21505 12587 21539
rect 12529 21499 12587 21505
rect 12544 21468 12572 21499
rect 12618 21496 12624 21548
rect 12676 21496 12682 21548
rect 12710 21496 12716 21548
rect 12768 21496 12774 21548
rect 12802 21496 12808 21548
rect 12860 21496 12866 21548
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 12728 21468 12756 21496
rect 13004 21468 13032 21499
rect 16298 21496 16304 21548
rect 16356 21496 16362 21548
rect 14829 21471 14887 21477
rect 14829 21468 14841 21471
rect 12544 21440 14841 21468
rect 14829 21437 14841 21440
rect 14875 21437 14887 21471
rect 14829 21431 14887 21437
rect 12713 21403 12771 21409
rect 12713 21369 12725 21403
rect 12759 21400 12771 21403
rect 13262 21400 13268 21412
rect 12759 21372 13268 21400
rect 12759 21369 12771 21372
rect 12713 21363 12771 21369
rect 13262 21360 13268 21372
rect 13320 21360 13326 21412
rect 15013 21403 15071 21409
rect 15013 21369 15025 21403
rect 15059 21400 15071 21403
rect 17512 21400 17540 21564
rect 17589 21539 17647 21545
rect 17589 21505 17601 21539
rect 17635 21536 17647 21539
rect 18156 21536 18184 21564
rect 17635 21508 18184 21536
rect 17635 21505 17647 21508
rect 17589 21499 17647 21505
rect 17954 21428 17960 21480
rect 18012 21428 18018 21480
rect 18046 21428 18052 21480
rect 18104 21477 18110 21480
rect 18104 21471 18132 21477
rect 18120 21437 18132 21471
rect 18104 21431 18132 21437
rect 18104 21428 18110 21431
rect 18248 21409 18276 21564
rect 18340 21545 18368 21644
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 20073 21675 20131 21681
rect 20073 21641 20085 21675
rect 20119 21672 20131 21675
rect 22922 21672 22928 21684
rect 20119 21644 22928 21672
rect 20119 21641 20131 21644
rect 20073 21635 20131 21641
rect 18598 21564 18604 21616
rect 18656 21564 18662 21616
rect 18325 21539 18383 21545
rect 18325 21505 18337 21539
rect 18371 21505 18383 21539
rect 18325 21499 18383 21505
rect 19702 21496 19708 21548
rect 19760 21496 19766 21548
rect 19242 21428 19248 21480
rect 19300 21468 19306 21480
rect 20088 21468 20116 21635
rect 22922 21632 22928 21644
rect 22980 21632 22986 21684
rect 24857 21675 24915 21681
rect 24857 21641 24869 21675
rect 24903 21672 24915 21675
rect 24946 21672 24952 21684
rect 24903 21644 24952 21672
rect 24903 21641 24915 21644
rect 24857 21635 24915 21641
rect 24946 21632 24952 21644
rect 25004 21632 25010 21684
rect 25317 21675 25375 21681
rect 25317 21641 25329 21675
rect 25363 21672 25375 21675
rect 26602 21672 26608 21684
rect 25363 21644 26608 21672
rect 25363 21641 25375 21644
rect 25317 21635 25375 21641
rect 26602 21632 26608 21644
rect 26660 21632 26666 21684
rect 30377 21675 30435 21681
rect 30377 21641 30389 21675
rect 30423 21672 30435 21675
rect 30650 21672 30656 21684
rect 30423 21644 30656 21672
rect 30423 21641 30435 21644
rect 30377 21635 30435 21641
rect 30650 21632 30656 21644
rect 30708 21632 30714 21684
rect 31021 21675 31079 21681
rect 31021 21641 31033 21675
rect 31067 21672 31079 21675
rect 31202 21672 31208 21684
rect 31067 21644 31208 21672
rect 31067 21641 31079 21644
rect 31021 21635 31079 21641
rect 31202 21632 31208 21644
rect 31260 21632 31266 21684
rect 33226 21632 33232 21684
rect 33284 21632 33290 21684
rect 21174 21564 21180 21616
rect 21232 21604 21238 21616
rect 21478 21607 21536 21613
rect 21478 21604 21490 21607
rect 21232 21576 21490 21604
rect 21232 21564 21238 21576
rect 21478 21573 21490 21576
rect 21524 21573 21536 21607
rect 21478 21567 21536 21573
rect 21634 21564 21640 21616
rect 21692 21604 21698 21616
rect 22005 21607 22063 21613
rect 22005 21604 22017 21607
rect 21692 21576 22017 21604
rect 21692 21564 21698 21576
rect 22005 21573 22017 21576
rect 22051 21573 22063 21607
rect 22005 21567 22063 21573
rect 25130 21564 25136 21616
rect 25188 21604 25194 21616
rect 25409 21607 25467 21613
rect 25409 21604 25421 21607
rect 25188 21576 25421 21604
rect 25188 21564 25194 21576
rect 25409 21573 25421 21576
rect 25455 21573 25467 21607
rect 25409 21567 25467 21573
rect 27706 21564 27712 21616
rect 27764 21564 27770 21616
rect 31386 21564 31392 21616
rect 31444 21564 31450 21616
rect 31496 21576 32352 21604
rect 20349 21539 20407 21545
rect 20349 21505 20361 21539
rect 20395 21536 20407 21539
rect 20714 21536 20720 21548
rect 20395 21508 20720 21536
rect 20395 21505 20407 21508
rect 20349 21499 20407 21505
rect 20714 21496 20720 21508
rect 20772 21496 20778 21548
rect 21361 21539 21419 21545
rect 21361 21505 21373 21539
rect 21407 21536 21419 21539
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21407 21508 21833 21536
rect 21407 21505 21419 21508
rect 21361 21499 21419 21505
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 22189 21539 22247 21545
rect 22189 21505 22201 21539
rect 22235 21536 22247 21539
rect 22646 21536 22652 21548
rect 22235 21508 22652 21536
rect 22235 21505 22247 21508
rect 22189 21499 22247 21505
rect 22646 21496 22652 21508
rect 22704 21496 22710 21548
rect 25038 21536 25044 21548
rect 24518 21508 25044 21536
rect 25038 21496 25044 21508
rect 25096 21536 25102 21548
rect 25314 21536 25320 21548
rect 25096 21508 25320 21536
rect 25096 21496 25102 21508
rect 25314 21496 25320 21508
rect 25372 21496 25378 21548
rect 26602 21496 26608 21548
rect 26660 21496 26666 21548
rect 26970 21496 26976 21548
rect 27028 21496 27034 21548
rect 29914 21536 29920 21548
rect 29380 21508 29920 21536
rect 19300 21440 20116 21468
rect 20625 21471 20683 21477
rect 19300 21428 19306 21440
rect 20625 21437 20637 21471
rect 20671 21468 20683 21471
rect 20993 21471 21051 21477
rect 20993 21468 21005 21471
rect 20671 21440 21005 21468
rect 20671 21437 20683 21440
rect 20625 21431 20683 21437
rect 20993 21437 21005 21440
rect 21039 21437 21051 21471
rect 20993 21431 21051 21437
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21437 21327 21471
rect 21269 21431 21327 21437
rect 15059 21372 17540 21400
rect 18233 21403 18291 21409
rect 15059 21369 15071 21372
rect 15013 21363 15071 21369
rect 18233 21369 18245 21403
rect 18279 21369 18291 21403
rect 18233 21363 18291 21369
rect 20640 21344 20668 21431
rect 20806 21360 20812 21412
rect 20864 21400 20870 21412
rect 21284 21400 21312 21431
rect 23014 21428 23020 21480
rect 23072 21468 23078 21480
rect 23109 21471 23167 21477
rect 23109 21468 23121 21471
rect 23072 21440 23121 21468
rect 23072 21428 23078 21440
rect 23109 21437 23121 21440
rect 23155 21437 23167 21471
rect 23109 21431 23167 21437
rect 23385 21471 23443 21477
rect 23385 21437 23397 21471
rect 23431 21468 23443 21471
rect 23842 21468 23848 21480
rect 23431 21440 23848 21468
rect 23431 21437 23443 21440
rect 23385 21431 23443 21437
rect 23842 21428 23848 21440
rect 23900 21428 23906 21480
rect 24578 21428 24584 21480
rect 24636 21428 24642 21480
rect 25222 21428 25228 21480
rect 25280 21428 25286 21480
rect 29380 21477 29408 21508
rect 29914 21496 29920 21508
rect 29972 21496 29978 21548
rect 30469 21539 30527 21545
rect 30469 21505 30481 21539
rect 30515 21536 30527 21539
rect 30926 21536 30932 21548
rect 30515 21508 30932 21536
rect 30515 21505 30527 21508
rect 30469 21499 30527 21505
rect 30926 21496 30932 21508
rect 30984 21536 30990 21548
rect 31297 21539 31355 21545
rect 31297 21536 31309 21539
rect 30984 21508 31309 21536
rect 30984 21496 30990 21508
rect 31297 21505 31309 21508
rect 31343 21505 31355 21539
rect 31297 21499 31355 21505
rect 25593 21471 25651 21477
rect 25593 21437 25605 21471
rect 25639 21437 25651 21471
rect 27249 21471 27307 21477
rect 27249 21468 27261 21471
rect 25593 21431 25651 21437
rect 26804 21440 27261 21468
rect 20864 21372 21312 21400
rect 24596 21400 24624 21428
rect 24949 21403 25007 21409
rect 24949 21400 24961 21403
rect 24596 21372 24961 21400
rect 20864 21360 20870 21372
rect 24949 21369 24961 21372
rect 24995 21369 25007 21403
rect 24949 21363 25007 21369
rect 11146 21332 11152 21344
rect 9876 21304 11152 21332
rect 9125 21295 9183 21301
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 12434 21292 12440 21344
rect 12492 21292 12498 21344
rect 15930 21292 15936 21344
rect 15988 21332 15994 21344
rect 16117 21335 16175 21341
rect 16117 21332 16129 21335
rect 15988 21304 16129 21332
rect 15988 21292 15994 21304
rect 16117 21301 16129 21304
rect 16163 21301 16175 21335
rect 16117 21295 16175 21301
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 17862 21332 17868 21344
rect 17000 21304 17868 21332
rect 17000 21292 17006 21304
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 20622 21292 20628 21344
rect 20680 21292 20686 21344
rect 20714 21292 20720 21344
rect 20772 21292 20778 21344
rect 20898 21292 20904 21344
rect 20956 21292 20962 21344
rect 21634 21292 21640 21344
rect 21692 21292 21698 21344
rect 23198 21292 23204 21344
rect 23256 21332 23262 21344
rect 25240 21332 25268 21428
rect 23256 21304 25268 21332
rect 25608 21332 25636 21431
rect 26804 21409 26832 21440
rect 27249 21437 27261 21440
rect 27295 21437 27307 21471
rect 27249 21431 27307 21437
rect 28721 21471 28779 21477
rect 28721 21437 28733 21471
rect 28767 21468 28779 21471
rect 29365 21471 29423 21477
rect 29365 21468 29377 21471
rect 28767 21440 29377 21468
rect 28767 21437 28779 21440
rect 28721 21431 28779 21437
rect 29365 21437 29377 21440
rect 29411 21437 29423 21471
rect 29365 21431 29423 21437
rect 30742 21428 30748 21480
rect 30800 21428 30806 21480
rect 31110 21428 31116 21480
rect 31168 21468 31174 21480
rect 31496 21477 31524 21576
rect 32324 21545 32352 21576
rect 31665 21539 31723 21545
rect 31665 21505 31677 21539
rect 31711 21505 31723 21539
rect 31665 21499 31723 21505
rect 32309 21539 32367 21545
rect 32309 21505 32321 21539
rect 32355 21505 32367 21539
rect 32309 21499 32367 21505
rect 31481 21471 31539 21477
rect 31481 21468 31493 21471
rect 31168 21440 31493 21468
rect 31168 21428 31174 21440
rect 31481 21437 31493 21440
rect 31527 21437 31539 21471
rect 31680 21468 31708 21499
rect 32217 21471 32275 21477
rect 32217 21468 32229 21471
rect 31680 21440 32229 21468
rect 31481 21431 31539 21437
rect 26789 21403 26847 21409
rect 26789 21369 26801 21403
rect 26835 21369 26847 21403
rect 26789 21363 26847 21369
rect 29840 21372 30420 21400
rect 29840 21344 29868 21372
rect 26510 21332 26516 21344
rect 25608 21304 26516 21332
rect 23256 21292 23262 21304
rect 26510 21292 26516 21304
rect 26568 21332 26574 21344
rect 26878 21332 26884 21344
rect 26568 21304 26884 21332
rect 26568 21292 26574 21304
rect 26878 21292 26884 21304
rect 26936 21292 26942 21344
rect 28810 21292 28816 21344
rect 28868 21292 28874 21344
rect 29822 21292 29828 21344
rect 29880 21292 29886 21344
rect 30098 21292 30104 21344
rect 30156 21332 30162 21344
rect 30193 21335 30251 21341
rect 30193 21332 30205 21335
rect 30156 21304 30205 21332
rect 30156 21292 30162 21304
rect 30193 21301 30205 21304
rect 30239 21332 30251 21335
rect 30282 21332 30288 21344
rect 30239 21304 30288 21332
rect 30239 21301 30251 21304
rect 30193 21295 30251 21301
rect 30282 21292 30288 21304
rect 30340 21292 30346 21344
rect 30392 21332 30420 21372
rect 30558 21332 30564 21344
rect 30392 21304 30564 21332
rect 30558 21292 30564 21304
rect 30616 21292 30622 21344
rect 30834 21292 30840 21344
rect 30892 21332 30898 21344
rect 31294 21332 31300 21344
rect 30892 21304 31300 21332
rect 30892 21292 30898 21304
rect 31294 21292 31300 21304
rect 31352 21292 31358 21344
rect 31478 21292 31484 21344
rect 31536 21332 31542 21344
rect 31726 21332 31754 21440
rect 32217 21437 32229 21440
rect 32263 21437 32275 21471
rect 32217 21431 32275 21437
rect 32677 21471 32735 21477
rect 32677 21437 32689 21471
rect 32723 21468 32735 21471
rect 33244 21468 33272 21632
rect 34333 21539 34391 21545
rect 34333 21505 34345 21539
rect 34379 21536 34391 21539
rect 34790 21536 34796 21548
rect 34379 21508 34796 21536
rect 34379 21505 34391 21508
rect 34333 21499 34391 21505
rect 34790 21496 34796 21508
rect 34848 21496 34854 21548
rect 32723 21440 33272 21468
rect 32723 21437 32735 21440
rect 32677 21431 32735 21437
rect 31536 21304 31754 21332
rect 34149 21335 34207 21341
rect 31536 21292 31542 21304
rect 34149 21301 34161 21335
rect 34195 21332 34207 21335
rect 34195 21304 34744 21332
rect 34195 21301 34207 21304
rect 34149 21295 34207 21301
rect 1104 21242 34684 21264
rect 1104 21190 5147 21242
rect 5199 21190 5211 21242
rect 5263 21190 5275 21242
rect 5327 21190 5339 21242
rect 5391 21190 5403 21242
rect 5455 21190 13541 21242
rect 13593 21190 13605 21242
rect 13657 21190 13669 21242
rect 13721 21190 13733 21242
rect 13785 21190 13797 21242
rect 13849 21190 21935 21242
rect 21987 21190 21999 21242
rect 22051 21190 22063 21242
rect 22115 21190 22127 21242
rect 22179 21190 22191 21242
rect 22243 21190 30329 21242
rect 30381 21190 30393 21242
rect 30445 21190 30457 21242
rect 30509 21190 30521 21242
rect 30573 21190 30585 21242
rect 30637 21190 34684 21242
rect 1104 21168 34684 21190
rect 9674 21088 9680 21140
rect 9732 21128 9738 21140
rect 9861 21131 9919 21137
rect 9861 21128 9873 21131
rect 9732 21100 9873 21128
rect 9732 21088 9738 21100
rect 9861 21097 9873 21100
rect 9907 21128 9919 21131
rect 12342 21128 12348 21140
rect 9907 21100 12348 21128
rect 9907 21097 9919 21100
rect 9861 21091 9919 21097
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 13262 21088 13268 21140
rect 13320 21128 13326 21140
rect 13645 21131 13703 21137
rect 13645 21128 13657 21131
rect 13320 21100 13657 21128
rect 13320 21088 13326 21100
rect 13645 21097 13657 21100
rect 13691 21097 13703 21131
rect 13645 21091 13703 21097
rect 15828 21131 15886 21137
rect 15828 21097 15840 21131
rect 15874 21128 15886 21131
rect 15930 21128 15936 21140
rect 15874 21100 15936 21128
rect 15874 21097 15886 21100
rect 15828 21091 15886 21097
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 16298 21088 16304 21140
rect 16356 21128 16362 21140
rect 17497 21131 17555 21137
rect 17497 21128 17509 21131
rect 16356 21100 17509 21128
rect 16356 21088 16362 21100
rect 17497 21097 17509 21100
rect 17543 21097 17555 21131
rect 17497 21091 17555 21097
rect 18046 21088 18052 21140
rect 18104 21128 18110 21140
rect 18969 21131 19027 21137
rect 18969 21128 18981 21131
rect 18104 21100 18981 21128
rect 18104 21088 18110 21100
rect 18969 21097 18981 21100
rect 19015 21097 19027 21131
rect 18969 21091 19027 21097
rect 20441 21131 20499 21137
rect 20441 21097 20453 21131
rect 20487 21128 20499 21131
rect 20622 21128 20628 21140
rect 20487 21100 20628 21128
rect 20487 21097 20499 21100
rect 20441 21091 20499 21097
rect 20622 21088 20628 21100
rect 20680 21088 20686 21140
rect 20806 21088 20812 21140
rect 20864 21088 20870 21140
rect 20898 21088 20904 21140
rect 20956 21088 20962 21140
rect 21726 21088 21732 21140
rect 21784 21088 21790 21140
rect 22097 21131 22155 21137
rect 22097 21097 22109 21131
rect 22143 21128 22155 21131
rect 22462 21128 22468 21140
rect 22143 21100 22468 21128
rect 22143 21097 22155 21100
rect 22097 21091 22155 21097
rect 22462 21088 22468 21100
rect 22520 21088 22526 21140
rect 26602 21088 26608 21140
rect 26660 21128 26666 21140
rect 26697 21131 26755 21137
rect 26697 21128 26709 21131
rect 26660 21100 26709 21128
rect 26660 21088 26666 21100
rect 26697 21097 26709 21100
rect 26743 21097 26755 21131
rect 26697 21091 26755 21097
rect 28810 21088 28816 21140
rect 28868 21088 28874 21140
rect 29914 21088 29920 21140
rect 29972 21128 29978 21140
rect 30193 21131 30251 21137
rect 30193 21128 30205 21131
rect 29972 21100 30205 21128
rect 29972 21088 29978 21100
rect 30193 21097 30205 21100
rect 30239 21097 30251 21131
rect 30193 21091 30251 21097
rect 30653 21131 30711 21137
rect 30653 21097 30665 21131
rect 30699 21128 30711 21131
rect 30742 21128 30748 21140
rect 30699 21100 30748 21128
rect 30699 21097 30711 21100
rect 30653 21091 30711 21097
rect 30742 21088 30748 21100
rect 30800 21088 30806 21140
rect 30834 21088 30840 21140
rect 30892 21088 30898 21140
rect 30926 21088 30932 21140
rect 30984 21088 30990 21140
rect 31110 21088 31116 21140
rect 31168 21128 31174 21140
rect 31205 21131 31263 21137
rect 31205 21128 31217 21131
rect 31168 21100 31217 21128
rect 31168 21088 31174 21100
rect 31205 21097 31217 21100
rect 31251 21097 31263 21131
rect 34716 21128 34744 21304
rect 31205 21091 31263 21097
rect 34256 21100 34744 21128
rect 20257 21063 20315 21069
rect 20257 21029 20269 21063
rect 20303 21060 20315 21063
rect 20824 21060 20852 21088
rect 20303 21032 20852 21060
rect 20303 21029 20315 21032
rect 20257 21023 20315 21029
rect 11885 20995 11943 21001
rect 11885 20961 11897 20995
rect 11931 20992 11943 20995
rect 12434 20992 12440 21004
rect 11931 20964 12440 20992
rect 11931 20961 11943 20964
rect 11885 20955 11943 20961
rect 12434 20952 12440 20964
rect 12492 20952 12498 21004
rect 13170 20952 13176 21004
rect 13228 20992 13234 21004
rect 13909 20995 13967 21001
rect 13909 20992 13921 20995
rect 13228 20964 13921 20992
rect 13228 20952 13234 20964
rect 13909 20961 13921 20964
rect 13955 20992 13967 20995
rect 15565 20995 15623 21001
rect 15565 20992 15577 20995
rect 13955 20964 15577 20992
rect 13955 20961 13967 20964
rect 13909 20955 13967 20961
rect 15565 20961 15577 20964
rect 15611 20992 15623 20995
rect 15838 20992 15844 21004
rect 15611 20964 15844 20992
rect 15611 20961 15623 20964
rect 15565 20955 15623 20961
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 20824 21001 20852 21032
rect 20809 20995 20867 21001
rect 20180 20964 20668 20992
rect 20180 20936 20208 20964
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 6730 20924 6736 20936
rect 5592 20896 6736 20924
rect 5592 20884 5598 20896
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 7098 20884 7104 20936
rect 7156 20924 7162 20936
rect 7285 20927 7343 20933
rect 7285 20924 7297 20927
rect 7156 20896 7297 20924
rect 7156 20884 7162 20896
rect 7285 20893 7297 20896
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 11330 20884 11336 20936
rect 11388 20884 11394 20936
rect 11514 20884 11520 20936
rect 11572 20884 11578 20936
rect 12526 20884 12532 20936
rect 12584 20884 12590 20936
rect 14734 20884 14740 20936
rect 14792 20884 14798 20936
rect 17494 20884 17500 20936
rect 17552 20924 17558 20936
rect 17656 20927 17714 20933
rect 17656 20924 17668 20927
rect 17552 20896 17668 20924
rect 17552 20884 17558 20896
rect 17656 20893 17668 20896
rect 17702 20893 17714 20927
rect 17656 20887 17714 20893
rect 18141 20927 18199 20933
rect 18141 20893 18153 20927
rect 18187 20924 18199 20927
rect 18230 20924 18236 20936
rect 18187 20896 18236 20924
rect 18187 20893 18199 20896
rect 18141 20887 18199 20893
rect 18230 20884 18236 20896
rect 18288 20924 18294 20936
rect 18601 20927 18659 20933
rect 18601 20924 18613 20927
rect 18288 20896 18613 20924
rect 18288 20884 18294 20896
rect 18601 20893 18613 20896
rect 18647 20893 18659 20927
rect 18601 20887 18659 20893
rect 20162 20884 20168 20936
rect 20220 20884 20226 20936
rect 20640 20933 20668 20964
rect 20809 20961 20821 20995
rect 20855 20961 20867 20995
rect 20916 20992 20944 21088
rect 20993 20995 21051 21001
rect 20993 20992 21005 20995
rect 20916 20964 21005 20992
rect 20809 20955 20867 20961
rect 20993 20961 21005 20964
rect 21039 20961 21051 20995
rect 21744 20992 21772 21088
rect 22833 21063 22891 21069
rect 22833 21029 22845 21063
rect 22879 21060 22891 21063
rect 23106 21060 23112 21072
rect 22879 21032 23112 21060
rect 22879 21029 22891 21032
rect 22833 21023 22891 21029
rect 23106 21020 23112 21032
rect 23164 21020 23170 21072
rect 23293 20995 23351 21001
rect 21744 20964 22094 20992
rect 20993 20955 21051 20961
rect 20349 20927 20407 20933
rect 20349 20893 20361 20927
rect 20395 20924 20407 20927
rect 20441 20927 20499 20933
rect 20441 20924 20453 20927
rect 20395 20896 20453 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 20441 20893 20453 20896
rect 20487 20893 20499 20927
rect 20441 20887 20499 20893
rect 20625 20927 20683 20933
rect 20625 20893 20637 20927
rect 20671 20893 20683 20927
rect 20625 20887 20683 20893
rect 21177 20927 21235 20933
rect 21177 20893 21189 20927
rect 21223 20893 21235 20927
rect 21177 20887 21235 20893
rect 4982 20816 4988 20868
rect 5040 20816 5046 20868
rect 6270 20816 6276 20868
rect 6328 20856 6334 20868
rect 7466 20856 7472 20868
rect 6328 20828 7472 20856
rect 6328 20816 6334 20828
rect 7466 20816 7472 20828
rect 7524 20816 7530 20868
rect 14752 20856 14780 20884
rect 17862 20856 17868 20868
rect 14752 20828 16330 20856
rect 17604 20828 17868 20856
rect 17604 20800 17632 20828
rect 17862 20816 17868 20828
rect 17920 20816 17926 20868
rect 18782 20816 18788 20868
rect 18840 20856 18846 20868
rect 19242 20856 19248 20868
rect 18840 20828 19248 20856
rect 18840 20816 18846 20828
rect 19242 20816 19248 20828
rect 19300 20816 19306 20868
rect 20364 20800 20392 20887
rect 21192 20856 21220 20887
rect 21542 20884 21548 20936
rect 21600 20924 21606 20936
rect 21637 20927 21695 20933
rect 21637 20924 21649 20927
rect 21600 20896 21649 20924
rect 21600 20884 21606 20896
rect 21637 20893 21649 20896
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 21729 20927 21787 20933
rect 21729 20893 21741 20927
rect 21775 20924 21787 20927
rect 21818 20924 21824 20936
rect 21775 20896 21824 20924
rect 21775 20893 21787 20896
rect 21729 20887 21787 20893
rect 21818 20884 21824 20896
rect 21876 20884 21882 20936
rect 22066 20924 22094 20964
rect 22756 20964 23152 20992
rect 22756 20936 22784 20964
rect 22281 20927 22339 20933
rect 22281 20924 22293 20927
rect 22066 20896 22293 20924
rect 22281 20893 22293 20896
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 22649 20927 22707 20933
rect 22649 20893 22661 20927
rect 22695 20924 22707 20927
rect 22738 20924 22744 20936
rect 22695 20896 22744 20924
rect 22695 20893 22707 20896
rect 22649 20887 22707 20893
rect 22738 20884 22744 20896
rect 22796 20884 22802 20936
rect 22922 20884 22928 20936
rect 22980 20884 22986 20936
rect 23124 20933 23152 20964
rect 23293 20961 23305 20995
rect 23339 20992 23351 20995
rect 23339 20964 25728 20992
rect 23339 20961 23351 20964
rect 23293 20955 23351 20961
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20924 23167 20927
rect 23201 20927 23259 20933
rect 23201 20924 23213 20927
rect 23155 20896 23213 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 23201 20893 23213 20896
rect 23247 20893 23259 20927
rect 23201 20887 23259 20893
rect 25041 20927 25099 20933
rect 25041 20893 25053 20927
rect 25087 20924 25099 20927
rect 25087 20896 25544 20924
rect 25087 20893 25099 20896
rect 25041 20887 25099 20893
rect 22370 20856 22376 20868
rect 21192 20828 22376 20856
rect 22370 20816 22376 20828
rect 22428 20816 22434 20868
rect 22465 20859 22523 20865
rect 22465 20825 22477 20859
rect 22511 20825 22523 20859
rect 22465 20819 22523 20825
rect 22557 20859 22615 20865
rect 22557 20825 22569 20859
rect 22603 20856 22615 20859
rect 22940 20856 22968 20884
rect 22603 20828 22968 20856
rect 22603 20825 22615 20828
rect 22557 20819 22615 20825
rect 4798 20748 4804 20800
rect 4856 20788 4862 20800
rect 4893 20791 4951 20797
rect 4893 20788 4905 20791
rect 4856 20760 4905 20788
rect 4856 20748 4862 20760
rect 4893 20757 4905 20760
rect 4939 20757 4951 20791
rect 4893 20751 4951 20757
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 7101 20791 7159 20797
rect 7101 20788 7113 20791
rect 5592 20760 7113 20788
rect 5592 20748 5598 20760
rect 7101 20757 7113 20760
rect 7147 20757 7159 20791
rect 7101 20751 7159 20757
rect 17310 20748 17316 20800
rect 17368 20748 17374 20800
rect 17586 20748 17592 20800
rect 17644 20748 17650 20800
rect 17773 20791 17831 20797
rect 17773 20757 17785 20791
rect 17819 20788 17831 20791
rect 17954 20788 17960 20800
rect 17819 20760 17960 20788
rect 17819 20757 17831 20760
rect 17773 20751 17831 20757
rect 17954 20748 17960 20760
rect 18012 20788 18018 20800
rect 18506 20788 18512 20800
rect 18012 20760 18512 20788
rect 18012 20748 18018 20760
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 20346 20748 20352 20800
rect 20404 20748 20410 20800
rect 22480 20788 22508 20819
rect 22646 20788 22652 20800
rect 22480 20760 22652 20788
rect 22646 20748 22652 20760
rect 22704 20748 22710 20800
rect 22922 20748 22928 20800
rect 22980 20788 22986 20800
rect 23017 20791 23075 20797
rect 23017 20788 23029 20791
rect 22980 20760 23029 20788
rect 22980 20748 22986 20760
rect 23017 20757 23029 20760
rect 23063 20757 23075 20791
rect 23017 20751 23075 20757
rect 24394 20748 24400 20800
rect 24452 20748 24458 20800
rect 25406 20748 25412 20800
rect 25464 20748 25470 20800
rect 25516 20788 25544 20896
rect 25590 20884 25596 20936
rect 25648 20884 25654 20936
rect 25700 20856 25728 20964
rect 26878 20952 26884 21004
rect 26936 20992 26942 21004
rect 27249 20995 27307 21001
rect 27249 20992 27261 20995
rect 26936 20964 27261 20992
rect 26936 20952 26942 20964
rect 27249 20961 27261 20964
rect 27295 20961 27307 20995
rect 28828 20992 28856 21088
rect 30098 21020 30104 21072
rect 30156 21020 30162 21072
rect 30561 21063 30619 21069
rect 30561 21029 30573 21063
rect 30607 21060 30619 21063
rect 30944 21060 30972 21088
rect 30607 21032 31248 21060
rect 30607 21029 30619 21032
rect 30561 21023 30619 21029
rect 27249 20955 27307 20961
rect 27908 20964 28856 20992
rect 27065 20927 27123 20933
rect 27065 20893 27077 20927
rect 27111 20924 27123 20927
rect 27908 20924 27936 20964
rect 27111 20896 27936 20924
rect 27111 20893 27123 20896
rect 27065 20887 27123 20893
rect 28718 20884 28724 20936
rect 28776 20884 28782 20936
rect 30116 20933 30144 21020
rect 30650 20952 30656 21004
rect 30708 20992 30714 21004
rect 30708 20964 31156 20992
rect 30708 20952 30714 20964
rect 30101 20927 30159 20933
rect 30101 20893 30113 20927
rect 30147 20893 30159 20927
rect 30101 20887 30159 20893
rect 30852 20865 30880 20964
rect 31128 20933 31156 20964
rect 31113 20927 31171 20933
rect 31113 20893 31125 20927
rect 31159 20893 31171 20927
rect 31220 20924 31248 21032
rect 34057 20995 34115 21001
rect 34057 20961 34069 20995
rect 34103 20992 34115 20995
rect 34256 20992 34284 21100
rect 34103 20964 34284 20992
rect 34103 20961 34115 20964
rect 34057 20955 34115 20961
rect 34330 20952 34336 21004
rect 34388 20952 34394 21004
rect 31297 20927 31355 20933
rect 31297 20924 31309 20927
rect 31220 20896 31309 20924
rect 31113 20887 31171 20893
rect 31297 20893 31309 20896
rect 31343 20893 31355 20927
rect 31297 20887 31355 20893
rect 32030 20884 32036 20936
rect 32088 20924 32094 20936
rect 32582 20924 32588 20936
rect 32088 20896 32588 20924
rect 32088 20884 32094 20896
rect 32582 20884 32588 20896
rect 32640 20884 32646 20936
rect 32950 20884 32956 20936
rect 33008 20884 33014 20936
rect 27157 20859 27215 20865
rect 27157 20856 27169 20859
rect 25700 20828 27169 20856
rect 27157 20825 27169 20828
rect 27203 20825 27215 20859
rect 30821 20859 30880 20865
rect 27157 20819 27215 20825
rect 28092 20828 28396 20856
rect 28092 20788 28120 20828
rect 25516 20760 28120 20788
rect 28166 20748 28172 20800
rect 28224 20748 28230 20800
rect 28368 20788 28396 20828
rect 30821 20825 30833 20859
rect 30867 20828 30880 20859
rect 30867 20825 30879 20828
rect 30821 20819 30879 20825
rect 30926 20816 30932 20868
rect 30984 20856 30990 20868
rect 31021 20859 31079 20865
rect 31021 20856 31033 20859
rect 30984 20828 31033 20856
rect 30984 20816 30990 20828
rect 31021 20825 31033 20828
rect 31067 20825 31079 20859
rect 31021 20819 31079 20825
rect 31128 20828 31754 20856
rect 31128 20788 31156 20828
rect 28368 20760 31156 20788
rect 31726 20788 31754 20828
rect 32585 20791 32643 20797
rect 32585 20788 32597 20791
rect 31726 20760 32597 20788
rect 32585 20757 32597 20760
rect 32631 20757 32643 20791
rect 32585 20751 32643 20757
rect 1104 20698 34840 20720
rect 1104 20646 9344 20698
rect 9396 20646 9408 20698
rect 9460 20646 9472 20698
rect 9524 20646 9536 20698
rect 9588 20646 9600 20698
rect 9652 20646 17738 20698
rect 17790 20646 17802 20698
rect 17854 20646 17866 20698
rect 17918 20646 17930 20698
rect 17982 20646 17994 20698
rect 18046 20646 26132 20698
rect 26184 20646 26196 20698
rect 26248 20646 26260 20698
rect 26312 20646 26324 20698
rect 26376 20646 26388 20698
rect 26440 20646 34526 20698
rect 34578 20646 34590 20698
rect 34642 20646 34654 20698
rect 34706 20646 34718 20698
rect 34770 20646 34782 20698
rect 34834 20646 34840 20698
rect 1104 20624 34840 20646
rect 4982 20544 4988 20596
rect 5040 20544 5046 20596
rect 6362 20544 6368 20596
rect 6420 20584 6426 20596
rect 6733 20587 6791 20593
rect 6733 20584 6745 20587
rect 6420 20556 6745 20584
rect 6420 20544 6426 20556
rect 6733 20553 6745 20556
rect 6779 20553 6791 20587
rect 6733 20547 6791 20553
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 8662 20584 8668 20596
rect 6972 20556 8668 20584
rect 6972 20544 6978 20556
rect 8662 20544 8668 20556
rect 8720 20544 8726 20596
rect 10594 20584 10600 20596
rect 10244 20556 10600 20584
rect 10244 20528 10272 20556
rect 10594 20544 10600 20556
rect 10652 20544 10658 20596
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 11609 20587 11667 20593
rect 11609 20584 11621 20587
rect 11572 20556 11621 20584
rect 11572 20544 11578 20556
rect 11609 20553 11621 20556
rect 11655 20553 11667 20587
rect 11609 20547 11667 20553
rect 15838 20544 15844 20596
rect 15896 20544 15902 20596
rect 17494 20544 17500 20596
rect 17552 20544 17558 20596
rect 18138 20544 18144 20596
rect 18196 20544 18202 20596
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 21600 20556 22017 20584
rect 21600 20544 21606 20556
rect 2682 20476 2688 20528
rect 2740 20476 2746 20528
rect 4890 20476 4896 20528
rect 4948 20516 4954 20528
rect 5353 20519 5411 20525
rect 5353 20516 5365 20519
rect 4948 20488 5365 20516
rect 4948 20476 4954 20488
rect 5353 20485 5365 20488
rect 5399 20485 5411 20519
rect 5902 20516 5908 20528
rect 5353 20479 5411 20485
rect 5552 20488 5908 20516
rect 4065 20451 4123 20457
rect 4065 20417 4077 20451
rect 4111 20448 4123 20451
rect 4522 20448 4528 20460
rect 4111 20420 4528 20448
rect 4111 20417 4123 20420
rect 4065 20411 4123 20417
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 5552 20457 5580 20488
rect 5902 20476 5908 20488
rect 5960 20516 5966 20528
rect 7742 20516 7748 20528
rect 5960 20488 6497 20516
rect 5960 20476 5966 20488
rect 5169 20451 5227 20457
rect 5169 20417 5181 20451
rect 5215 20417 5227 20451
rect 5169 20411 5227 20417
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 1394 20340 1400 20392
rect 1452 20380 1458 20392
rect 1946 20380 1952 20392
rect 1452 20352 1952 20380
rect 1452 20340 1458 20352
rect 1946 20340 1952 20352
rect 2004 20340 2010 20392
rect 2314 20340 2320 20392
rect 2372 20340 2378 20392
rect 4614 20340 4620 20392
rect 4672 20340 4678 20392
rect 4798 20340 4804 20392
rect 4856 20340 4862 20392
rect 5184 20380 5212 20411
rect 5626 20408 5632 20460
rect 5684 20408 5690 20460
rect 5718 20408 5724 20460
rect 5776 20408 5782 20460
rect 5810 20408 5816 20460
rect 5868 20448 5874 20460
rect 6270 20448 6276 20460
rect 5868 20420 6276 20448
rect 5868 20408 5874 20420
rect 6270 20408 6276 20420
rect 6328 20448 6334 20460
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 6328 20420 6377 20448
rect 6328 20408 6334 20420
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 5736 20380 5764 20408
rect 5184 20352 5764 20380
rect 6469 20380 6497 20488
rect 6656 20488 7748 20516
rect 6546 20408 6552 20460
rect 6604 20408 6610 20460
rect 6656 20457 6684 20488
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20417 6699 20451
rect 6641 20411 6699 20417
rect 6914 20408 6920 20460
rect 6972 20408 6978 20460
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20417 7067 20451
rect 7009 20411 7067 20417
rect 7024 20380 7052 20411
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 7156 20420 7205 20448
rect 7156 20408 7162 20420
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 7282 20408 7288 20460
rect 7340 20408 7346 20460
rect 7392 20457 7420 20488
rect 7742 20476 7748 20488
rect 7800 20516 7806 20528
rect 7800 20488 9352 20516
rect 7800 20476 7806 20488
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 7466 20408 7472 20460
rect 7524 20408 7530 20460
rect 8021 20451 8079 20457
rect 8021 20417 8033 20451
rect 8067 20448 8079 20451
rect 8386 20448 8392 20460
rect 8067 20420 8392 20448
rect 8067 20417 8079 20420
rect 8021 20411 8079 20417
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 8938 20408 8944 20460
rect 8996 20408 9002 20460
rect 9324 20457 9352 20488
rect 9674 20476 9680 20528
rect 9732 20516 9738 20528
rect 9953 20519 10011 20525
rect 9953 20516 9965 20519
rect 9732 20488 9965 20516
rect 9732 20476 9738 20488
rect 9953 20485 9965 20488
rect 9999 20516 10011 20519
rect 10226 20516 10232 20528
rect 9999 20488 10232 20516
rect 9999 20485 10011 20488
rect 9953 20479 10011 20485
rect 10226 20476 10232 20488
rect 10284 20476 10290 20528
rect 10781 20519 10839 20525
rect 10781 20516 10793 20519
rect 10428 20488 10793 20516
rect 10428 20460 10456 20488
rect 10781 20485 10793 20488
rect 10827 20485 10839 20519
rect 15856 20516 15884 20544
rect 17129 20519 17187 20525
rect 15856 20488 16160 20516
rect 10781 20479 10839 20485
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20417 9367 20451
rect 9309 20411 9367 20417
rect 10137 20451 10195 20457
rect 10137 20417 10149 20451
rect 10183 20448 10195 20451
rect 10183 20420 10364 20448
rect 10183 20417 10195 20420
rect 10137 20411 10195 20417
rect 7929 20383 7987 20389
rect 7929 20380 7941 20383
rect 6469 20352 7941 20380
rect 7929 20349 7941 20352
rect 7975 20349 7987 20383
rect 7929 20343 7987 20349
rect 9401 20383 9459 20389
rect 9401 20349 9413 20383
rect 9447 20380 9459 20383
rect 9769 20383 9827 20389
rect 9769 20380 9781 20383
rect 9447 20352 9781 20380
rect 9447 20349 9459 20352
rect 9401 20343 9459 20349
rect 9769 20349 9781 20352
rect 9815 20380 9827 20383
rect 9858 20380 9864 20392
rect 9815 20352 9864 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 9858 20340 9864 20352
rect 9916 20380 9922 20392
rect 10229 20383 10287 20389
rect 10229 20380 10241 20383
rect 9916 20352 10241 20380
rect 9916 20340 9922 20352
rect 10229 20349 10241 20352
rect 10275 20349 10287 20383
rect 10336 20380 10364 20420
rect 10410 20408 10416 20460
rect 10468 20408 10474 20460
rect 10594 20408 10600 20460
rect 10652 20448 10658 20460
rect 10689 20451 10747 20457
rect 10689 20448 10701 20451
rect 10652 20420 10701 20448
rect 10652 20408 10658 20420
rect 10689 20417 10701 20420
rect 10735 20417 10747 20451
rect 10689 20411 10747 20417
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 10502 20380 10508 20392
rect 10336 20352 10508 20380
rect 10229 20343 10287 20349
rect 10502 20340 10508 20352
rect 10560 20380 10566 20392
rect 10888 20380 10916 20411
rect 10560 20352 10916 20380
rect 10560 20340 10566 20352
rect 4982 20272 4988 20324
rect 5040 20312 5046 20324
rect 5040 20284 6500 20312
rect 5040 20272 5046 20284
rect 4154 20204 4160 20256
rect 4212 20204 4218 20256
rect 5537 20247 5595 20253
rect 5537 20213 5549 20247
rect 5583 20244 5595 20247
rect 5994 20244 6000 20256
rect 5583 20216 6000 20244
rect 5583 20213 5595 20216
rect 5537 20207 5595 20213
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 6472 20253 6500 20284
rect 8662 20272 8668 20324
rect 8720 20312 8726 20324
rect 8757 20315 8815 20321
rect 8757 20312 8769 20315
rect 8720 20284 8769 20312
rect 8720 20272 8726 20284
rect 8757 20281 8769 20284
rect 8803 20281 8815 20315
rect 11716 20312 11744 20411
rect 12250 20408 12256 20460
rect 12308 20408 12314 20460
rect 12434 20408 12440 20460
rect 12492 20457 12498 20460
rect 12492 20451 12507 20457
rect 12495 20448 12507 20451
rect 12894 20448 12900 20460
rect 12495 20420 12900 20448
rect 12495 20417 12507 20420
rect 12492 20411 12507 20417
rect 12492 20408 12498 20411
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 14734 20408 14740 20460
rect 14792 20408 14798 20460
rect 16132 20457 16160 20488
rect 17129 20485 17141 20519
rect 17175 20516 17187 20519
rect 17218 20516 17224 20528
rect 17175 20488 17224 20516
rect 17175 20485 17187 20488
rect 17129 20479 17187 20485
rect 17218 20476 17224 20488
rect 17276 20516 17282 20528
rect 18293 20519 18351 20525
rect 18293 20516 18305 20519
rect 17276 20488 18305 20516
rect 17276 20476 17282 20488
rect 18293 20485 18305 20488
rect 18339 20485 18351 20519
rect 18293 20479 18351 20485
rect 18509 20519 18567 20525
rect 18509 20485 18521 20519
rect 18555 20516 18567 20519
rect 18782 20516 18788 20528
rect 18555 20488 18788 20516
rect 18555 20485 18567 20488
rect 18509 20479 18567 20485
rect 18782 20476 18788 20488
rect 18840 20476 18846 20528
rect 21634 20476 21640 20528
rect 21692 20476 21698 20528
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20417 16175 20451
rect 16117 20411 16175 20417
rect 17034 20408 17040 20460
rect 17092 20448 17098 20460
rect 17310 20448 17316 20460
rect 17092 20420 17316 20448
rect 17092 20408 17098 20420
rect 17310 20408 17316 20420
rect 17368 20448 17374 20460
rect 17862 20448 17868 20460
rect 17368 20420 17868 20448
rect 17368 20408 17374 20420
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 15841 20383 15899 20389
rect 15841 20349 15853 20383
rect 15887 20380 15899 20383
rect 21652 20380 21680 20476
rect 21744 20460 21772 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 26970 20544 26976 20596
rect 27028 20584 27034 20596
rect 29730 20584 29736 20596
rect 27028 20556 29736 20584
rect 27028 20544 27034 20556
rect 22204 20488 22784 20516
rect 21726 20408 21732 20460
rect 21784 20408 21790 20460
rect 22204 20457 22232 20488
rect 21821 20451 21879 20457
rect 21821 20417 21833 20451
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 22189 20451 22247 20457
rect 22189 20417 22201 20451
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 21836 20380 21864 20411
rect 22462 20408 22468 20460
rect 22520 20408 22526 20460
rect 22756 20457 22784 20488
rect 23106 20476 23112 20528
rect 23164 20476 23170 20528
rect 25317 20519 25375 20525
rect 25317 20485 25329 20519
rect 25363 20516 25375 20519
rect 25406 20516 25412 20528
rect 25363 20488 25412 20516
rect 25363 20485 25375 20488
rect 25317 20479 25375 20485
rect 25406 20476 25412 20488
rect 25464 20476 25470 20528
rect 27706 20516 27712 20528
rect 26542 20488 27712 20516
rect 27706 20476 27712 20488
rect 27764 20476 27770 20528
rect 22557 20451 22615 20457
rect 22557 20417 22569 20451
rect 22603 20417 22615 20451
rect 22557 20411 22615 20417
rect 22741 20451 22799 20457
rect 22741 20417 22753 20451
rect 22787 20448 22799 20451
rect 23124 20448 23152 20476
rect 22787 20420 23152 20448
rect 22787 20417 22799 20420
rect 22741 20411 22799 20417
rect 22572 20380 22600 20411
rect 24854 20408 24860 20460
rect 24912 20448 24918 20460
rect 25041 20451 25099 20457
rect 25041 20448 25053 20451
rect 24912 20420 25053 20448
rect 24912 20408 24918 20420
rect 25041 20417 25053 20420
rect 25087 20417 25099 20451
rect 27816 20448 27844 20556
rect 29730 20544 29736 20556
rect 29788 20544 29794 20596
rect 30469 20587 30527 20593
rect 30469 20553 30481 20587
rect 30515 20584 30527 20587
rect 30926 20584 30932 20596
rect 30515 20556 30932 20584
rect 30515 20553 30527 20556
rect 30469 20547 30527 20553
rect 30926 20544 30932 20556
rect 30984 20584 30990 20596
rect 31386 20584 31392 20596
rect 30984 20556 31392 20584
rect 30984 20544 30990 20556
rect 31386 20544 31392 20556
rect 31444 20544 31450 20596
rect 32674 20544 32680 20596
rect 32732 20584 32738 20596
rect 32769 20587 32827 20593
rect 32769 20584 32781 20587
rect 32732 20556 32781 20584
rect 32732 20544 32738 20556
rect 32769 20553 32781 20556
rect 32815 20553 32827 20587
rect 32769 20547 32827 20553
rect 28074 20476 28080 20528
rect 28132 20516 28138 20528
rect 28132 20488 28658 20516
rect 28132 20476 28138 20488
rect 30742 20476 30748 20528
rect 30800 20516 30806 20528
rect 31110 20516 31116 20528
rect 30800 20488 31116 20516
rect 30800 20476 30806 20488
rect 31110 20476 31116 20488
rect 31168 20476 31174 20528
rect 27893 20451 27951 20457
rect 27893 20448 27905 20451
rect 27816 20420 27905 20448
rect 25041 20411 25099 20417
rect 27893 20417 27905 20420
rect 27939 20417 27951 20451
rect 29998 20449 30056 20455
rect 29998 20446 30010 20449
rect 27893 20411 27951 20417
rect 29932 20418 30010 20446
rect 29932 20380 29960 20418
rect 29998 20415 30010 20418
rect 30044 20415 30056 20449
rect 29998 20409 30056 20415
rect 33042 20408 33048 20460
rect 33100 20448 33106 20460
rect 33137 20451 33195 20457
rect 33137 20448 33149 20451
rect 33100 20420 33149 20448
rect 33100 20408 33106 20420
rect 33137 20417 33149 20420
rect 33183 20417 33195 20451
rect 33137 20411 33195 20417
rect 33229 20383 33287 20389
rect 33229 20380 33241 20383
rect 15887 20352 19012 20380
rect 21652 20352 21864 20380
rect 15887 20349 15899 20352
rect 15841 20343 15899 20349
rect 8757 20275 8815 20281
rect 10336 20284 11744 20312
rect 18984 20312 19012 20352
rect 21542 20312 21548 20324
rect 18984 20284 21548 20312
rect 10336 20256 10364 20284
rect 21542 20272 21548 20284
rect 21600 20272 21606 20324
rect 6457 20247 6515 20253
rect 6457 20213 6469 20247
rect 6503 20213 6515 20247
rect 6457 20207 6515 20213
rect 7282 20204 7288 20256
rect 7340 20244 7346 20256
rect 7558 20244 7564 20256
rect 7340 20216 7564 20244
rect 7340 20204 7346 20216
rect 7558 20204 7564 20216
rect 7616 20204 7622 20256
rect 7742 20204 7748 20256
rect 7800 20204 7806 20256
rect 10318 20204 10324 20256
rect 10376 20204 10382 20256
rect 10597 20247 10655 20253
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 10962 20244 10968 20256
rect 10643 20216 10968 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 12437 20247 12495 20253
rect 12437 20213 12449 20247
rect 12483 20244 12495 20247
rect 12618 20244 12624 20256
rect 12483 20216 12624 20244
rect 12483 20213 12495 20216
rect 12437 20207 12495 20213
rect 12618 20204 12624 20216
rect 12676 20204 12682 20256
rect 14366 20204 14372 20256
rect 14424 20204 14430 20256
rect 17862 20204 17868 20256
rect 17920 20244 17926 20256
rect 18325 20247 18383 20253
rect 18325 20244 18337 20247
rect 17920 20216 18337 20244
rect 17920 20204 17926 20216
rect 18325 20213 18337 20216
rect 18371 20244 18383 20247
rect 21174 20244 21180 20256
rect 18371 20216 21180 20244
rect 18371 20213 18383 20216
rect 18325 20207 18383 20213
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 21836 20244 21864 20352
rect 22204 20352 22600 20380
rect 26804 20352 29960 20380
rect 22204 20244 22232 20352
rect 22296 20284 22968 20312
rect 22296 20253 22324 20284
rect 22940 20256 22968 20284
rect 21836 20216 22232 20244
rect 22281 20247 22339 20253
rect 22281 20213 22293 20247
rect 22327 20213 22339 20247
rect 22281 20207 22339 20213
rect 22370 20204 22376 20256
rect 22428 20244 22434 20256
rect 22649 20247 22707 20253
rect 22649 20244 22661 20247
rect 22428 20216 22661 20244
rect 22428 20204 22434 20216
rect 22649 20213 22661 20216
rect 22695 20213 22707 20247
rect 22649 20207 22707 20213
rect 22922 20204 22928 20256
rect 22980 20204 22986 20256
rect 25682 20204 25688 20256
rect 25740 20244 25746 20256
rect 26804 20253 26832 20352
rect 29932 20312 29960 20352
rect 31726 20352 33241 20380
rect 30006 20312 30012 20324
rect 29932 20284 30012 20312
rect 30006 20272 30012 20284
rect 30064 20272 30070 20324
rect 31726 20312 31754 20352
rect 33229 20349 33241 20352
rect 33275 20349 33287 20383
rect 33229 20343 33287 20349
rect 33410 20340 33416 20392
rect 33468 20340 33474 20392
rect 30300 20284 31754 20312
rect 26789 20247 26847 20253
rect 26789 20244 26801 20247
rect 25740 20216 26801 20244
rect 25740 20204 25746 20216
rect 26789 20213 26801 20216
rect 26835 20213 26847 20247
rect 26789 20207 26847 20213
rect 27706 20204 27712 20256
rect 27764 20244 27770 20256
rect 27982 20244 27988 20256
rect 27764 20216 27988 20244
rect 27764 20204 27770 20216
rect 27982 20204 27988 20216
rect 28040 20204 28046 20256
rect 28166 20253 28172 20256
rect 28156 20247 28172 20253
rect 28156 20213 28168 20247
rect 28156 20207 28172 20213
rect 28166 20204 28172 20207
rect 28224 20204 28230 20256
rect 29641 20247 29699 20253
rect 29641 20213 29653 20247
rect 29687 20244 29699 20247
rect 29914 20244 29920 20256
rect 29687 20216 29920 20244
rect 29687 20213 29699 20216
rect 29641 20207 29699 20213
rect 29914 20204 29920 20216
rect 29972 20244 29978 20256
rect 30300 20253 30328 20284
rect 30285 20247 30343 20253
rect 30285 20244 30297 20247
rect 29972 20216 30297 20244
rect 29972 20204 29978 20216
rect 30285 20213 30297 20216
rect 30331 20213 30343 20247
rect 30285 20207 30343 20213
rect 1104 20154 34684 20176
rect 1104 20102 5147 20154
rect 5199 20102 5211 20154
rect 5263 20102 5275 20154
rect 5327 20102 5339 20154
rect 5391 20102 5403 20154
rect 5455 20102 13541 20154
rect 13593 20102 13605 20154
rect 13657 20102 13669 20154
rect 13721 20102 13733 20154
rect 13785 20102 13797 20154
rect 13849 20102 21935 20154
rect 21987 20102 21999 20154
rect 22051 20102 22063 20154
rect 22115 20102 22127 20154
rect 22179 20102 22191 20154
rect 22243 20102 30329 20154
rect 30381 20102 30393 20154
rect 30445 20102 30457 20154
rect 30509 20102 30521 20154
rect 30573 20102 30585 20154
rect 30637 20102 34684 20154
rect 1104 20080 34684 20102
rect 2314 20000 2320 20052
rect 2372 20040 2378 20052
rect 2685 20043 2743 20049
rect 2685 20040 2697 20043
rect 2372 20012 2697 20040
rect 2372 20000 2378 20012
rect 2685 20009 2697 20012
rect 2731 20009 2743 20043
rect 2685 20003 2743 20009
rect 4154 20000 4160 20052
rect 4212 20000 4218 20052
rect 4341 20043 4399 20049
rect 4341 20009 4353 20043
rect 4387 20009 4399 20043
rect 4341 20003 4399 20009
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 4614 20040 4620 20052
rect 4571 20012 4620 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 4172 19904 4200 20000
rect 4356 19972 4384 20003
rect 4614 20000 4620 20012
rect 4672 20000 4678 20052
rect 4706 20000 4712 20052
rect 4764 20040 4770 20052
rect 5077 20043 5135 20049
rect 5077 20040 5089 20043
rect 4764 20012 5089 20040
rect 4764 20000 4770 20012
rect 5077 20009 5089 20012
rect 5123 20009 5135 20043
rect 5077 20003 5135 20009
rect 5534 20000 5540 20052
rect 5592 20000 5598 20052
rect 7098 20000 7104 20052
rect 7156 20000 7162 20052
rect 7285 20043 7343 20049
rect 7285 20009 7297 20043
rect 7331 20040 7343 20043
rect 7742 20040 7748 20052
rect 7331 20012 7748 20040
rect 7331 20009 7343 20012
rect 7285 20003 7343 20009
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 9858 20000 9864 20052
rect 9916 20000 9922 20052
rect 10410 20000 10416 20052
rect 10468 20000 10474 20052
rect 12250 20000 12256 20052
rect 12308 20040 12314 20052
rect 12526 20040 12532 20052
rect 12308 20012 12532 20040
rect 12308 20000 12314 20012
rect 12526 20000 12532 20012
rect 12584 20040 12590 20052
rect 13357 20043 13415 20049
rect 13357 20040 13369 20043
rect 12584 20012 13369 20040
rect 12584 20000 12590 20012
rect 13357 20009 13369 20012
rect 13403 20009 13415 20043
rect 13357 20003 13415 20009
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 5552 19972 5580 20000
rect 4356 19944 5580 19972
rect 2884 19876 4200 19904
rect 4908 19876 5764 19904
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 2884 19845 2912 19876
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 2869 19839 2927 19845
rect 2869 19805 2881 19839
rect 2915 19805 2927 19839
rect 2869 19799 2927 19805
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19836 4031 19839
rect 4341 19839 4399 19845
rect 4019 19808 4200 19836
rect 4019 19805 4031 19808
rect 3973 19799 4031 19805
rect 4172 19780 4200 19808
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 4614 19836 4620 19848
rect 4387 19808 4620 19836
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4798 19836 4804 19848
rect 4755 19808 4804 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 4908 19845 4936 19876
rect 5736 19848 5764 19876
rect 6638 19864 6644 19916
rect 6696 19904 6702 19916
rect 7282 19904 7288 19916
rect 6696 19876 7288 19904
rect 6696 19864 6702 19876
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 8588 19876 9536 19904
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19805 4951 19839
rect 5261 19839 5319 19845
rect 5261 19836 5273 19839
rect 4893 19799 4951 19805
rect 5000 19808 5273 19836
rect 4154 19728 4160 19780
rect 4212 19728 4218 19780
rect 1578 19660 1584 19712
rect 1636 19660 1642 19712
rect 3602 19660 3608 19712
rect 3660 19700 3666 19712
rect 4801 19703 4859 19709
rect 4801 19700 4813 19703
rect 3660 19672 4813 19700
rect 3660 19660 3666 19672
rect 4801 19669 4813 19672
rect 4847 19700 4859 19703
rect 5000 19700 5028 19808
rect 5261 19805 5273 19808
rect 5307 19805 5319 19839
rect 5261 19799 5319 19805
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19838 5595 19839
rect 5583 19810 5672 19838
rect 5583 19805 5595 19810
rect 5537 19799 5595 19805
rect 5644 19768 5672 19810
rect 5718 19796 5724 19848
rect 5776 19796 5782 19848
rect 5902 19796 5908 19848
rect 5960 19796 5966 19848
rect 7009 19839 7067 19845
rect 7009 19836 7021 19839
rect 6840 19808 7021 19836
rect 6840 19780 6868 19808
rect 7009 19805 7021 19808
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7190 19796 7196 19848
rect 7248 19796 7254 19848
rect 7396 19839 7454 19845
rect 7396 19805 7408 19839
rect 7442 19836 7454 19839
rect 7561 19839 7619 19845
rect 7442 19808 7512 19836
rect 7442 19805 7454 19808
rect 7396 19799 7454 19805
rect 5994 19768 6000 19780
rect 5644 19740 6000 19768
rect 5994 19728 6000 19740
rect 6052 19728 6058 19780
rect 6822 19728 6828 19780
rect 6880 19728 6886 19780
rect 7484 19768 7512 19808
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 8386 19836 8392 19848
rect 7607 19808 8392 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 8588 19845 8616 19876
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19805 8631 19839
rect 8573 19799 8631 19805
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19836 8815 19839
rect 9030 19836 9036 19848
rect 8803 19808 9036 19836
rect 8803 19805 8815 19808
rect 8757 19799 8815 19805
rect 9030 19796 9036 19808
rect 9088 19836 9094 19848
rect 9508 19845 9536 19876
rect 9493 19839 9551 19845
rect 9088 19808 9352 19836
rect 9088 19796 9094 19808
rect 9324 19777 9352 19808
rect 9493 19805 9505 19839
rect 9539 19836 9551 19839
rect 9674 19836 9680 19848
rect 9539 19808 9680 19836
rect 9539 19805 9551 19808
rect 9493 19799 9551 19805
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 9876 19845 9904 20000
rect 10045 19975 10103 19981
rect 10045 19941 10057 19975
rect 10091 19972 10103 19975
rect 10226 19972 10232 19984
rect 10091 19944 10232 19972
rect 10091 19941 10103 19944
rect 10045 19935 10103 19941
rect 10226 19932 10232 19944
rect 10284 19932 10290 19984
rect 10428 19904 10456 20000
rect 11054 19904 11060 19916
rect 10152 19876 10456 19904
rect 10520 19876 11060 19904
rect 10152 19845 10180 19876
rect 9861 19839 9919 19845
rect 9861 19805 9873 19839
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 10318 19796 10324 19848
rect 10376 19796 10382 19848
rect 10520 19845 10548 19876
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 10965 19839 11023 19845
rect 10965 19805 10977 19839
rect 11011 19836 11023 19839
rect 11330 19836 11336 19848
rect 11011 19808 11336 19836
rect 11011 19805 11023 19808
rect 10965 19799 11023 19805
rect 9309 19771 9367 19777
rect 7484 19740 9168 19768
rect 9140 19712 9168 19740
rect 9309 19737 9321 19771
rect 9355 19737 9367 19771
rect 10980 19768 11008 19799
rect 11330 19796 11336 19808
rect 11388 19796 11394 19848
rect 13265 19839 13323 19845
rect 13265 19805 13277 19839
rect 13311 19836 13323 19839
rect 17144 19836 17172 20003
rect 17218 20000 17224 20052
rect 17276 20000 17282 20052
rect 17313 20043 17371 20049
rect 17313 20009 17325 20043
rect 17359 20040 17371 20043
rect 18230 20040 18236 20052
rect 17359 20012 18236 20040
rect 17359 20009 17371 20012
rect 17313 20003 17371 20009
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 22462 20000 22468 20052
rect 22520 20040 22526 20052
rect 22557 20043 22615 20049
rect 22557 20040 22569 20043
rect 22520 20012 22569 20040
rect 22520 20000 22526 20012
rect 22557 20009 22569 20012
rect 22603 20009 22615 20043
rect 22557 20003 22615 20009
rect 25317 20043 25375 20049
rect 25317 20009 25329 20043
rect 25363 20040 25375 20043
rect 25590 20040 25596 20052
rect 25363 20012 25596 20040
rect 25363 20009 25375 20012
rect 25317 20003 25375 20009
rect 25590 20000 25596 20012
rect 25648 20000 25654 20052
rect 28077 20043 28135 20049
rect 28077 20009 28089 20043
rect 28123 20040 28135 20043
rect 28718 20040 28724 20052
rect 28123 20012 28724 20040
rect 28123 20009 28135 20012
rect 28077 20003 28135 20009
rect 28718 20000 28724 20012
rect 28776 20000 28782 20052
rect 29914 20000 29920 20052
rect 29972 20000 29978 20052
rect 30006 20000 30012 20052
rect 30064 20000 30070 20052
rect 17236 19904 17264 20000
rect 21174 19932 21180 19984
rect 21232 19972 21238 19984
rect 21232 19944 23152 19972
rect 21232 19932 21238 19944
rect 17405 19907 17463 19913
rect 17405 19904 17417 19907
rect 17236 19876 17417 19904
rect 17405 19873 17417 19876
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 20809 19907 20867 19913
rect 20809 19904 20821 19907
rect 19668 19876 20821 19904
rect 19668 19864 19674 19876
rect 20809 19873 20821 19876
rect 20855 19873 20867 19907
rect 20809 19867 20867 19873
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 23014 19904 23020 19916
rect 21131 19876 23020 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 23014 19864 23020 19876
rect 23072 19864 23078 19916
rect 17773 19839 17831 19845
rect 13311 19808 13492 19836
rect 17144 19808 17356 19836
rect 13311 19805 13323 19808
rect 13265 19799 13323 19805
rect 13464 19780 13492 19808
rect 9309 19731 9367 19737
rect 9876 19740 11008 19768
rect 4847 19672 5028 19700
rect 4847 19669 4859 19672
rect 4801 19663 4859 19669
rect 5442 19660 5448 19712
rect 5500 19660 5506 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 8665 19703 8723 19709
rect 8665 19700 8677 19703
rect 5592 19672 8677 19700
rect 5592 19660 5598 19672
rect 8665 19669 8677 19672
rect 8711 19669 8723 19703
rect 8665 19663 8723 19669
rect 9122 19660 9128 19712
rect 9180 19660 9186 19712
rect 9324 19700 9352 19731
rect 9876 19700 9904 19740
rect 13446 19728 13452 19780
rect 13504 19728 13510 19780
rect 16945 19771 17003 19777
rect 16945 19737 16957 19771
rect 16991 19768 17003 19771
rect 17034 19768 17040 19780
rect 16991 19740 17040 19768
rect 16991 19737 17003 19740
rect 16945 19731 17003 19737
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 17328 19712 17356 19808
rect 17773 19805 17785 19839
rect 17819 19836 17831 19839
rect 18506 19836 18512 19848
rect 17819 19808 18512 19836
rect 17819 19805 17831 19808
rect 17773 19799 17831 19805
rect 18506 19796 18512 19808
rect 18564 19796 18570 19848
rect 19702 19796 19708 19848
rect 19760 19796 19766 19848
rect 22554 19796 22560 19848
rect 22612 19796 22618 19848
rect 22738 19796 22744 19848
rect 22796 19836 22802 19848
rect 23124 19836 23152 19944
rect 23750 19932 23756 19984
rect 23808 19932 23814 19984
rect 27433 19975 27491 19981
rect 27433 19972 27445 19975
rect 23860 19944 27445 19972
rect 23198 19864 23204 19916
rect 23256 19904 23262 19916
rect 23569 19907 23627 19913
rect 23569 19904 23581 19907
rect 23256 19876 23581 19904
rect 23256 19864 23262 19876
rect 23569 19873 23581 19876
rect 23615 19904 23627 19907
rect 23768 19904 23796 19932
rect 23615 19876 23796 19904
rect 23615 19873 23627 19876
rect 23569 19867 23627 19873
rect 23290 19836 23296 19848
rect 22796 19808 23296 19836
rect 22796 19796 22802 19808
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 23750 19796 23756 19848
rect 23808 19796 23814 19848
rect 23860 19845 23888 19944
rect 27433 19941 27445 19944
rect 27479 19941 27491 19975
rect 27433 19935 27491 19941
rect 25961 19907 26019 19913
rect 23952 19876 24716 19904
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19805 23903 19839
rect 23845 19799 23903 19805
rect 17586 19728 17592 19780
rect 17644 19768 17650 19780
rect 17890 19771 17948 19777
rect 17890 19768 17902 19771
rect 17644 19740 17902 19768
rect 17644 19728 17650 19740
rect 17890 19737 17902 19740
rect 17936 19737 17948 19771
rect 23768 19768 23796 19796
rect 23952 19768 23980 19876
rect 24688 19845 24716 19876
rect 25961 19873 25973 19907
rect 26007 19904 26019 19907
rect 26878 19904 26884 19916
rect 26007 19876 26884 19904
rect 26007 19873 26019 19876
rect 25961 19867 26019 19873
rect 26878 19864 26884 19876
rect 26936 19864 26942 19916
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 23768 19740 23980 19768
rect 24228 19808 24593 19836
rect 17890 19731 17948 19737
rect 9324 19672 9904 19700
rect 10502 19660 10508 19712
rect 10560 19660 10566 19712
rect 10873 19703 10931 19709
rect 10873 19669 10885 19703
rect 10919 19700 10931 19703
rect 11054 19700 11060 19712
rect 10919 19672 11060 19700
rect 10919 19669 10931 19672
rect 10873 19663 10931 19669
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 17126 19660 17132 19712
rect 17184 19709 17190 19712
rect 17184 19703 17203 19709
rect 17191 19669 17203 19703
rect 17184 19663 17203 19669
rect 17184 19660 17190 19663
rect 17310 19660 17316 19712
rect 17368 19660 17374 19712
rect 17494 19660 17500 19712
rect 17552 19700 17558 19712
rect 17681 19703 17739 19709
rect 17681 19700 17693 19703
rect 17552 19672 17693 19700
rect 17552 19660 17558 19672
rect 17681 19669 17693 19672
rect 17727 19669 17739 19703
rect 17681 19663 17739 19669
rect 18049 19703 18107 19709
rect 18049 19669 18061 19703
rect 18095 19700 18107 19703
rect 18138 19700 18144 19712
rect 18095 19672 18144 19700
rect 18095 19669 18107 19672
rect 18049 19663 18107 19669
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 22278 19700 22284 19712
rect 19392 19672 22284 19700
rect 19392 19660 19398 19672
rect 22278 19660 22284 19672
rect 22336 19700 22342 19712
rect 23658 19700 23664 19712
rect 22336 19672 23664 19700
rect 22336 19660 22342 19672
rect 23658 19660 23664 19672
rect 23716 19700 23722 19712
rect 24228 19709 24256 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 24673 19839 24731 19845
rect 24673 19805 24685 19839
rect 24719 19805 24731 19839
rect 24673 19799 24731 19805
rect 25682 19796 25688 19848
rect 25740 19796 25746 19848
rect 26786 19796 26792 19848
rect 26844 19796 26850 19848
rect 27448 19836 27476 19935
rect 27798 19864 27804 19916
rect 27856 19904 27862 19916
rect 28442 19904 28448 19916
rect 27856 19876 28448 19904
rect 27856 19864 27862 19876
rect 28442 19864 28448 19876
rect 28500 19864 28506 19916
rect 28537 19907 28595 19913
rect 28537 19873 28549 19907
rect 28583 19904 28595 19907
rect 29932 19904 29960 20000
rect 28583 19876 29960 19904
rect 28583 19873 28595 19876
rect 28537 19867 28595 19873
rect 28261 19839 28319 19845
rect 28261 19836 28273 19839
rect 27448 19808 28273 19836
rect 28261 19805 28273 19808
rect 28307 19805 28319 19839
rect 28261 19799 28319 19805
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19805 28687 19839
rect 28629 19799 28687 19805
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19836 28871 19839
rect 29362 19836 29368 19848
rect 28859 19808 29368 19836
rect 28859 19805 28871 19808
rect 28813 19799 28871 19805
rect 24765 19771 24823 19777
rect 24765 19737 24777 19771
rect 24811 19768 24823 19771
rect 25777 19771 25835 19777
rect 25777 19768 25789 19771
rect 24811 19740 25789 19768
rect 24811 19737 24823 19740
rect 24765 19731 24823 19737
rect 25777 19737 25789 19740
rect 25823 19737 25835 19771
rect 25777 19731 25835 19737
rect 28166 19728 28172 19780
rect 28224 19768 28230 19780
rect 28644 19768 28672 19799
rect 29362 19796 29368 19808
rect 29420 19796 29426 19848
rect 29932 19845 29960 19876
rect 29917 19839 29975 19845
rect 29917 19805 29929 19839
rect 29963 19805 29975 19839
rect 29917 19799 29975 19805
rect 28224 19740 28672 19768
rect 28224 19728 28230 19740
rect 23753 19703 23811 19709
rect 23753 19700 23765 19703
rect 23716 19672 23765 19700
rect 23716 19660 23722 19672
rect 23753 19669 23765 19672
rect 23799 19669 23811 19703
rect 23753 19663 23811 19669
rect 24213 19703 24271 19709
rect 24213 19669 24225 19703
rect 24259 19669 24271 19703
rect 24213 19663 24271 19669
rect 24394 19660 24400 19712
rect 24452 19660 24458 19712
rect 30374 19660 30380 19712
rect 30432 19660 30438 19712
rect 1104 19610 34840 19632
rect 1104 19558 9344 19610
rect 9396 19558 9408 19610
rect 9460 19558 9472 19610
rect 9524 19558 9536 19610
rect 9588 19558 9600 19610
rect 9652 19558 17738 19610
rect 17790 19558 17802 19610
rect 17854 19558 17866 19610
rect 17918 19558 17930 19610
rect 17982 19558 17994 19610
rect 18046 19558 26132 19610
rect 26184 19558 26196 19610
rect 26248 19558 26260 19610
rect 26312 19558 26324 19610
rect 26376 19558 26388 19610
rect 26440 19558 34526 19610
rect 34578 19558 34590 19610
rect 34642 19558 34654 19610
rect 34706 19558 34718 19610
rect 34770 19558 34782 19610
rect 34834 19558 34840 19610
rect 1104 19536 34840 19558
rect 3142 19456 3148 19508
rect 3200 19456 3206 19508
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 4706 19496 4712 19508
rect 4212 19468 4712 19496
rect 4212 19456 4218 19468
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 4798 19456 4804 19508
rect 4856 19456 4862 19508
rect 4982 19456 4988 19508
rect 5040 19496 5046 19508
rect 5169 19499 5227 19505
rect 5169 19496 5181 19499
rect 5040 19468 5181 19496
rect 5040 19456 5046 19468
rect 5169 19465 5181 19468
rect 5215 19465 5227 19499
rect 5169 19459 5227 19465
rect 5626 19456 5632 19508
rect 5684 19496 5690 19508
rect 6822 19496 6828 19508
rect 5684 19468 6828 19496
rect 5684 19456 5690 19468
rect 6822 19456 6828 19468
rect 6880 19496 6886 19508
rect 12802 19496 12808 19508
rect 6880 19468 12808 19496
rect 6880 19456 6886 19468
rect 12802 19456 12808 19468
rect 12860 19496 12866 19508
rect 13446 19496 13452 19508
rect 12860 19468 13452 19496
rect 12860 19456 12866 19468
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 15197 19499 15255 19505
rect 15197 19465 15209 19499
rect 15243 19496 15255 19499
rect 15286 19496 15292 19508
rect 15243 19468 15292 19496
rect 15243 19465 15255 19468
rect 15197 19459 15255 19465
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 17218 19456 17224 19508
rect 17276 19456 17282 19508
rect 17405 19499 17463 19505
rect 17405 19465 17417 19499
rect 17451 19496 17463 19499
rect 17586 19496 17592 19508
rect 17451 19468 17592 19496
rect 17451 19465 17463 19468
rect 17405 19459 17463 19465
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 19334 19456 19340 19508
rect 19392 19456 19398 19508
rect 22066 19468 31064 19496
rect 1578 19388 1584 19440
rect 1636 19428 1642 19440
rect 1673 19431 1731 19437
rect 1673 19428 1685 19431
rect 1636 19400 1685 19428
rect 1636 19388 1642 19400
rect 1673 19397 1685 19400
rect 1719 19397 1731 19431
rect 1673 19391 1731 19397
rect 2682 19388 2688 19440
rect 2740 19388 2746 19440
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 3878 19320 3884 19372
rect 3936 19360 3942 19372
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 3936 19332 4261 19360
rect 3936 19320 3942 19332
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19360 4491 19363
rect 4816 19360 4844 19456
rect 5353 19431 5411 19437
rect 5353 19397 5365 19431
rect 5399 19428 5411 19431
rect 7098 19428 7104 19440
rect 5399 19400 7104 19428
rect 5399 19397 5411 19400
rect 5353 19391 5411 19397
rect 7098 19388 7104 19400
rect 7156 19388 7162 19440
rect 8386 19388 8392 19440
rect 8444 19388 8450 19440
rect 9125 19431 9183 19437
rect 9125 19397 9137 19431
rect 9171 19428 9183 19431
rect 13725 19431 13783 19437
rect 13725 19428 13737 19431
rect 9171 19400 13737 19428
rect 9171 19397 9183 19400
rect 9125 19391 9183 19397
rect 13725 19397 13737 19400
rect 13771 19397 13783 19431
rect 13725 19391 13783 19397
rect 14734 19388 14740 19440
rect 14792 19388 14798 19440
rect 17236 19428 17264 19456
rect 17497 19431 17555 19437
rect 17497 19428 17509 19431
rect 17236 19400 17509 19428
rect 17497 19397 17509 19400
rect 17543 19397 17555 19431
rect 17497 19391 17555 19397
rect 17604 19400 17908 19428
rect 4479 19332 4844 19360
rect 4479 19329 4491 19332
rect 4433 19323 4491 19329
rect 4890 19320 4896 19372
rect 4948 19360 4954 19372
rect 5445 19363 5503 19369
rect 5445 19360 5457 19363
rect 4948 19332 5457 19360
rect 4948 19320 4954 19332
rect 5445 19329 5457 19332
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 5902 19320 5908 19372
rect 5960 19320 5966 19372
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7193 19363 7251 19369
rect 7193 19360 7205 19363
rect 6972 19332 7205 19360
rect 6972 19320 6978 19332
rect 7193 19329 7205 19332
rect 7239 19329 7251 19363
rect 7193 19323 7251 19329
rect 7374 19320 7380 19372
rect 7432 19320 7438 19372
rect 8404 19360 8432 19388
rect 11698 19360 11704 19372
rect 8404 19332 11704 19360
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 11790 19320 11796 19372
rect 11848 19320 11854 19372
rect 11974 19320 11980 19372
rect 12032 19360 12038 19372
rect 12437 19363 12495 19369
rect 12437 19360 12449 19363
rect 12032 19332 12449 19360
rect 12032 19320 12038 19332
rect 12437 19329 12449 19332
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12618 19320 12624 19372
rect 12676 19320 12682 19372
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 4617 19295 4675 19301
rect 4617 19261 4629 19295
rect 4663 19261 4675 19295
rect 4617 19255 4675 19261
rect 4632 19156 4660 19255
rect 4706 19252 4712 19304
rect 4764 19292 4770 19304
rect 4801 19295 4859 19301
rect 4801 19292 4813 19295
rect 4764 19264 4813 19292
rect 4764 19252 4770 19264
rect 4801 19261 4813 19264
rect 4847 19261 4859 19295
rect 4801 19255 4859 19261
rect 4985 19295 5043 19301
rect 4985 19261 4997 19295
rect 5031 19261 5043 19295
rect 4985 19255 5043 19261
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5166 19292 5172 19304
rect 5123 19264 5172 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5000 19224 5028 19255
rect 5166 19252 5172 19264
rect 5224 19292 5230 19304
rect 5718 19292 5724 19304
rect 5224 19264 5724 19292
rect 5224 19252 5230 19264
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 5920 19224 5948 19320
rect 8478 19252 8484 19304
rect 8536 19252 8542 19304
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 9824 19264 12265 19292
rect 9824 19252 9830 19264
rect 12253 19261 12265 19264
rect 12299 19292 12311 19295
rect 13096 19292 13124 19323
rect 13170 19320 13176 19372
rect 13228 19360 13234 19372
rect 13449 19363 13507 19369
rect 13449 19360 13461 19363
rect 13228 19332 13461 19360
rect 13228 19320 13234 19332
rect 13449 19329 13461 19332
rect 13495 19329 13507 19363
rect 13449 19323 13507 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19360 17279 19363
rect 17310 19360 17316 19372
rect 17267 19332 17316 19360
rect 17267 19329 17279 19332
rect 17221 19323 17279 19329
rect 17052 19292 17080 19323
rect 17310 19320 17316 19332
rect 17368 19360 17374 19372
rect 17604 19360 17632 19400
rect 17880 19369 17908 19400
rect 17368 19332 17632 19360
rect 17681 19363 17739 19369
rect 17368 19320 17374 19332
rect 17681 19329 17693 19363
rect 17727 19329 17739 19363
rect 17681 19323 17739 19329
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19360 17923 19363
rect 19352 19360 19380 19456
rect 19705 19431 19763 19437
rect 19705 19397 19717 19431
rect 19751 19428 19763 19431
rect 22066 19428 22094 19468
rect 31036 19440 31064 19468
rect 31386 19456 31392 19508
rect 31444 19496 31450 19508
rect 31444 19468 31800 19496
rect 31444 19456 31450 19468
rect 19751 19400 22094 19428
rect 19751 19397 19763 19400
rect 19705 19391 19763 19397
rect 22554 19388 22560 19440
rect 22612 19428 22618 19440
rect 23750 19428 23756 19440
rect 22612 19400 23756 19428
rect 22612 19388 22618 19400
rect 23750 19388 23756 19400
rect 23808 19388 23814 19440
rect 25038 19428 25044 19440
rect 24978 19400 25044 19428
rect 25038 19388 25044 19400
rect 25096 19388 25102 19440
rect 26786 19428 26792 19440
rect 25240 19400 26792 19428
rect 17911 19332 19380 19360
rect 17911 19329 17923 19332
rect 17865 19323 17923 19329
rect 17126 19292 17132 19304
rect 12299 19264 12388 19292
rect 13096 19264 13308 19292
rect 17052 19264 17132 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12360 19236 12388 19264
rect 5000 19196 5948 19224
rect 12342 19184 12348 19236
rect 12400 19184 12406 19236
rect 13280 19168 13308 19264
rect 17126 19252 17132 19264
rect 17184 19292 17190 19304
rect 17696 19292 17724 19323
rect 20254 19320 20260 19372
rect 20312 19360 20318 19372
rect 20533 19363 20591 19369
rect 20533 19360 20545 19363
rect 20312 19332 20545 19360
rect 20312 19320 20318 19332
rect 20533 19329 20545 19332
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 17184 19264 17724 19292
rect 17184 19252 17190 19264
rect 17586 19184 17592 19236
rect 17644 19224 17650 19236
rect 17696 19224 17724 19264
rect 20346 19252 20352 19304
rect 20404 19252 20410 19304
rect 20548 19292 20576 19323
rect 20622 19320 20628 19372
rect 20680 19360 20686 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20680 19332 20729 19360
rect 20680 19320 20686 19332
rect 20717 19329 20729 19332
rect 20763 19360 20775 19363
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20763 19332 20821 19360
rect 20763 19329 20775 19332
rect 20717 19323 20775 19329
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20809 19323 20867 19329
rect 20916 19332 21005 19360
rect 20916 19304 20944 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 20898 19292 20904 19304
rect 20548 19264 20904 19292
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 23474 19252 23480 19304
rect 23532 19252 23538 19304
rect 23753 19295 23811 19301
rect 23753 19261 23765 19295
rect 23799 19292 23811 19295
rect 24394 19292 24400 19304
rect 23799 19264 24400 19292
rect 23799 19261 23811 19264
rect 23753 19255 23811 19261
rect 24394 19252 24400 19264
rect 24452 19252 24458 19304
rect 25240 19301 25268 19400
rect 26786 19388 26792 19400
rect 26844 19388 26850 19440
rect 27338 19428 27344 19440
rect 26896 19400 27344 19428
rect 26510 19320 26516 19372
rect 26568 19320 26574 19372
rect 26896 19360 26924 19400
rect 27338 19388 27344 19400
rect 27396 19428 27402 19440
rect 27396 19400 27738 19428
rect 27396 19388 27402 19400
rect 30374 19388 30380 19440
rect 30432 19388 30438 19440
rect 31018 19388 31024 19440
rect 31076 19388 31082 19440
rect 31128 19400 31616 19428
rect 26620 19332 26924 19360
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19261 25283 19295
rect 25225 19255 25283 19261
rect 23382 19224 23388 19236
rect 17644 19196 17724 19224
rect 18248 19196 23388 19224
rect 17644 19184 17650 19196
rect 5626 19156 5632 19168
rect 4632 19128 5632 19156
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 7558 19116 7564 19168
rect 7616 19116 7622 19168
rect 13262 19116 13268 19168
rect 13320 19116 13326 19168
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 18248 19165 18276 19196
rect 23382 19184 23388 19196
rect 23440 19184 23446 19236
rect 24946 19184 24952 19236
rect 25004 19224 25010 19236
rect 26620 19224 26648 19332
rect 26970 19320 26976 19372
rect 27028 19320 27034 19372
rect 30009 19363 30067 19369
rect 30009 19360 30021 19363
rect 28736 19332 30021 19360
rect 28736 19304 28764 19332
rect 30009 19329 30021 19332
rect 30055 19360 30067 19363
rect 30392 19360 30420 19388
rect 31128 19360 31156 19400
rect 31588 19369 31616 19400
rect 31772 19369 31800 19468
rect 33042 19456 33048 19508
rect 33100 19496 33106 19508
rect 33137 19499 33195 19505
rect 33137 19496 33149 19499
rect 33100 19468 33149 19496
rect 33100 19456 33106 19468
rect 33137 19465 33149 19468
rect 33183 19465 33195 19499
rect 33137 19459 33195 19465
rect 30055 19332 30328 19360
rect 30392 19332 31156 19360
rect 31205 19363 31263 19369
rect 30055 19329 30067 19332
rect 30009 19323 30067 19329
rect 27249 19295 27307 19301
rect 27249 19292 27261 19295
rect 26712 19264 27261 19292
rect 26712 19233 26740 19264
rect 27249 19261 27261 19264
rect 27295 19261 27307 19295
rect 27249 19255 27307 19261
rect 28718 19252 28724 19304
rect 28776 19252 28782 19304
rect 30300 19292 30328 19332
rect 31036 19301 31064 19332
rect 31205 19329 31217 19363
rect 31251 19360 31263 19363
rect 31481 19363 31539 19369
rect 31481 19360 31493 19363
rect 31251 19332 31340 19360
rect 31251 19329 31263 19332
rect 31205 19323 31263 19329
rect 31021 19295 31079 19301
rect 30300 19264 30696 19292
rect 30668 19236 30696 19264
rect 31021 19261 31033 19295
rect 31067 19261 31079 19295
rect 31021 19255 31079 19261
rect 25004 19196 26648 19224
rect 25004 19184 25010 19196
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 13964 19128 18245 19156
rect 13964 19116 13970 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18233 19119 18291 19125
rect 20809 19159 20867 19165
rect 20809 19125 20821 19159
rect 20855 19156 20867 19159
rect 25130 19156 25136 19168
rect 20855 19128 25136 19156
rect 20855 19125 20867 19128
rect 20809 19119 20867 19125
rect 25130 19116 25136 19128
rect 25188 19116 25194 19168
rect 26620 19156 26648 19196
rect 26697 19227 26755 19233
rect 26697 19193 26709 19227
rect 26743 19193 26755 19227
rect 26697 19187 26755 19193
rect 30650 19184 30656 19236
rect 30708 19184 30714 19236
rect 31312 19224 31340 19332
rect 31404 19332 31493 19360
rect 31404 19304 31432 19332
rect 31481 19329 31493 19332
rect 31527 19329 31539 19363
rect 31481 19323 31539 19329
rect 31573 19363 31631 19369
rect 31573 19329 31585 19363
rect 31619 19329 31631 19363
rect 31573 19323 31631 19329
rect 31757 19363 31815 19369
rect 31757 19329 31769 19363
rect 31803 19329 31815 19363
rect 31757 19323 31815 19329
rect 32490 19320 32496 19372
rect 32548 19360 32554 19372
rect 32769 19363 32827 19369
rect 32769 19360 32781 19363
rect 32548 19332 32781 19360
rect 32548 19320 32554 19332
rect 32769 19329 32781 19332
rect 32815 19329 32827 19363
rect 32769 19323 32827 19329
rect 31386 19252 31392 19304
rect 31444 19252 31450 19304
rect 31665 19295 31723 19301
rect 31665 19261 31677 19295
rect 31711 19292 31723 19295
rect 32508 19292 32536 19320
rect 31711 19264 32536 19292
rect 31711 19261 31723 19264
rect 31665 19255 31723 19261
rect 32674 19252 32680 19304
rect 32732 19252 32738 19304
rect 32122 19224 32128 19236
rect 31312 19196 32128 19224
rect 32122 19184 32128 19196
rect 32180 19184 32186 19236
rect 26786 19156 26792 19168
rect 26620 19128 26792 19156
rect 26786 19116 26792 19128
rect 26844 19116 26850 19168
rect 30190 19116 30196 19168
rect 30248 19116 30254 19168
rect 30469 19159 30527 19165
rect 30469 19125 30481 19159
rect 30515 19156 30527 19159
rect 31570 19156 31576 19168
rect 30515 19128 31576 19156
rect 30515 19125 30527 19128
rect 30469 19119 30527 19125
rect 31570 19116 31576 19128
rect 31628 19116 31634 19168
rect 1104 19066 34684 19088
rect 1104 19014 5147 19066
rect 5199 19014 5211 19066
rect 5263 19014 5275 19066
rect 5327 19014 5339 19066
rect 5391 19014 5403 19066
rect 5455 19014 13541 19066
rect 13593 19014 13605 19066
rect 13657 19014 13669 19066
rect 13721 19014 13733 19066
rect 13785 19014 13797 19066
rect 13849 19014 21935 19066
rect 21987 19014 21999 19066
rect 22051 19014 22063 19066
rect 22115 19014 22127 19066
rect 22179 19014 22191 19066
rect 22243 19014 30329 19066
rect 30381 19014 30393 19066
rect 30445 19014 30457 19066
rect 30509 19014 30521 19066
rect 30573 19014 30585 19066
rect 30637 19014 34684 19066
rect 1104 18992 34684 19014
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 9766 18952 9772 18964
rect 1912 18924 9772 18952
rect 1912 18912 1918 18924
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 12986 18912 12992 18964
rect 13044 18912 13050 18964
rect 18601 18955 18659 18961
rect 18601 18921 18613 18955
rect 18647 18952 18659 18955
rect 19610 18952 19616 18964
rect 18647 18924 19616 18952
rect 18647 18921 18659 18924
rect 18601 18915 18659 18921
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 20548 18924 23152 18952
rect 6362 18844 6368 18896
rect 6420 18884 6426 18896
rect 7282 18884 7288 18896
rect 6420 18856 7288 18884
rect 6420 18844 6426 18856
rect 7282 18844 7288 18856
rect 7340 18884 7346 18896
rect 8573 18887 8631 18893
rect 7340 18856 8524 18884
rect 7340 18844 7346 18856
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 1581 18819 1639 18825
rect 1581 18816 1593 18819
rect 1452 18788 1593 18816
rect 1452 18776 1458 18788
rect 1581 18785 1593 18788
rect 1627 18816 1639 18819
rect 8294 18816 8300 18828
rect 1627 18788 8300 18816
rect 1627 18785 1639 18788
rect 1581 18779 1639 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 2958 18708 2964 18760
rect 3016 18708 3022 18760
rect 5258 18708 5264 18760
rect 5316 18748 5322 18760
rect 5718 18748 5724 18760
rect 5316 18720 5724 18748
rect 5316 18708 5322 18720
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18748 6883 18751
rect 6914 18748 6920 18760
rect 6871 18720 6920 18748
rect 6871 18717 6883 18720
rect 6825 18711 6883 18717
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 7374 18708 7380 18760
rect 7432 18708 7438 18760
rect 7558 18708 7564 18760
rect 7616 18748 7622 18760
rect 7745 18751 7803 18757
rect 7745 18748 7757 18751
rect 7616 18720 7757 18748
rect 7616 18708 7622 18720
rect 7745 18717 7757 18720
rect 7791 18717 7803 18751
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 7745 18711 7803 18717
rect 7852 18720 8401 18748
rect 1854 18640 1860 18692
rect 1912 18640 1918 18692
rect 3605 18683 3663 18689
rect 3605 18649 3617 18683
rect 3651 18680 3663 18683
rect 3694 18680 3700 18692
rect 3651 18652 3700 18680
rect 3651 18649 3663 18652
rect 3605 18643 3663 18649
rect 3694 18640 3700 18652
rect 3752 18640 3758 18692
rect 7392 18680 7420 18708
rect 7852 18680 7880 18720
rect 8389 18717 8401 18720
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 7392 18652 7880 18680
rect 8021 18683 8079 18689
rect 8021 18649 8033 18683
rect 8067 18680 8079 18683
rect 8294 18680 8300 18692
rect 8067 18652 8300 18680
rect 8067 18649 8079 18652
rect 8021 18643 8079 18649
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 8496 18680 8524 18856
rect 8573 18853 8585 18887
rect 8619 18884 8631 18887
rect 9582 18884 9588 18896
rect 8619 18856 9588 18884
rect 8619 18853 8631 18856
rect 8573 18847 8631 18853
rect 9582 18844 9588 18856
rect 9640 18844 9646 18896
rect 9858 18844 9864 18896
rect 9916 18884 9922 18896
rect 10318 18884 10324 18896
rect 9916 18856 10324 18884
rect 9916 18844 9922 18856
rect 10318 18844 10324 18856
rect 10376 18884 10382 18896
rect 10376 18856 10732 18884
rect 10376 18844 10382 18856
rect 8754 18776 8760 18828
rect 8812 18816 8818 18828
rect 9033 18819 9091 18825
rect 9033 18816 9045 18819
rect 8812 18788 9045 18816
rect 8812 18776 8818 18788
rect 9033 18785 9045 18788
rect 9079 18816 9091 18819
rect 9079 18788 9996 18816
rect 9079 18785 9091 18788
rect 9033 18779 9091 18785
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 9674 18748 9680 18760
rect 8628 18720 9680 18748
rect 8628 18708 8634 18720
rect 9646 18716 9680 18720
rect 9674 18708 9680 18716
rect 9732 18708 9738 18760
rect 9766 18708 9772 18760
rect 9824 18757 9830 18760
rect 9968 18757 9996 18788
rect 10704 18757 10732 18856
rect 12161 18819 12219 18825
rect 12161 18785 12173 18819
rect 12207 18785 12219 18819
rect 13004 18816 13032 18912
rect 15565 18887 15623 18893
rect 15565 18853 15577 18887
rect 15611 18884 15623 18887
rect 20254 18884 20260 18896
rect 15611 18856 20260 18884
rect 15611 18853 15623 18856
rect 15565 18847 15623 18853
rect 20254 18844 20260 18856
rect 20312 18844 20318 18896
rect 13004 18788 15148 18816
rect 12161 18779 12219 18785
rect 9824 18751 9845 18757
rect 9833 18717 9845 18751
rect 9824 18711 9845 18717
rect 9953 18751 10011 18757
rect 9953 18717 9965 18751
rect 9999 18717 10011 18751
rect 9953 18711 10011 18717
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 9824 18708 9830 18711
rect 11054 18708 11060 18760
rect 11112 18708 11118 18760
rect 11330 18708 11336 18760
rect 11388 18748 11394 18760
rect 12176 18748 12204 18779
rect 12802 18748 12808 18760
rect 11388 18720 12204 18748
rect 12268 18720 12808 18748
rect 11388 18708 11394 18720
rect 9309 18683 9367 18689
rect 9309 18680 9321 18683
rect 8496 18652 9321 18680
rect 9309 18649 9321 18652
rect 9355 18649 9367 18683
rect 9309 18643 9367 18649
rect 10042 18640 10048 18692
rect 10100 18680 10106 18692
rect 10100 18652 10272 18680
rect 10100 18640 10106 18652
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7377 18615 7435 18621
rect 7377 18612 7389 18615
rect 7156 18584 7389 18612
rect 7156 18572 7162 18584
rect 7377 18581 7389 18584
rect 7423 18612 7435 18615
rect 7834 18612 7840 18624
rect 7423 18584 7840 18612
rect 7423 18581 7435 18584
rect 7377 18575 7435 18581
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 9217 18615 9275 18621
rect 9217 18612 9229 18615
rect 8628 18584 9229 18612
rect 8628 18572 8634 18584
rect 9217 18581 9229 18584
rect 9263 18581 9275 18615
rect 9217 18575 9275 18581
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 9766 18612 9772 18624
rect 9723 18584 9772 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 9766 18572 9772 18584
rect 9824 18572 9830 18624
rect 10134 18572 10140 18624
rect 10192 18572 10198 18624
rect 10244 18612 10272 18652
rect 12066 18640 12072 18692
rect 12124 18680 12130 18692
rect 12268 18680 12296 18720
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18748 13415 18751
rect 13446 18748 13452 18760
rect 13403 18720 13452 18748
rect 13403 18717 13415 18720
rect 13357 18711 13415 18717
rect 13446 18708 13452 18720
rect 13504 18708 13510 18760
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18748 13783 18751
rect 14090 18748 14096 18760
rect 13771 18720 14096 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 12124 18652 12296 18680
rect 12621 18683 12679 18689
rect 12124 18640 12130 18652
rect 12621 18649 12633 18683
rect 12667 18680 12679 18683
rect 13262 18680 13268 18692
rect 12667 18652 13268 18680
rect 12667 18649 12679 18652
rect 12621 18643 12679 18649
rect 13262 18640 13268 18652
rect 13320 18640 13326 18692
rect 13740 18612 13768 18711
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 15120 18680 15148 18788
rect 15764 18788 16528 18816
rect 15764 18760 15792 18788
rect 15746 18708 15752 18760
rect 15804 18708 15810 18760
rect 16500 18757 16528 18788
rect 18138 18776 18144 18828
rect 18196 18776 18202 18828
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18748 16083 18751
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 16071 18720 16313 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 16301 18717 16313 18720
rect 16347 18717 16359 18751
rect 16301 18711 16359 18717
rect 16485 18751 16543 18757
rect 16485 18717 16497 18751
rect 16531 18717 16543 18751
rect 18156 18748 18184 18776
rect 18417 18751 18475 18757
rect 18417 18748 18429 18751
rect 18156 18720 18429 18748
rect 16485 18711 16543 18717
rect 18417 18717 18429 18720
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 16040 18680 16068 18711
rect 18690 18708 18696 18760
rect 18748 18708 18754 18760
rect 20548 18757 20576 18924
rect 21818 18844 21824 18896
rect 21876 18844 21882 18896
rect 22462 18884 22468 18896
rect 22020 18856 22468 18884
rect 22020 18757 22048 18856
rect 22462 18844 22468 18856
rect 22520 18884 22526 18896
rect 23124 18884 23152 18924
rect 23198 18912 23204 18964
rect 23256 18912 23262 18964
rect 26329 18955 26387 18961
rect 26329 18921 26341 18955
rect 26375 18952 26387 18955
rect 26510 18952 26516 18964
rect 26375 18924 26516 18952
rect 26375 18921 26387 18924
rect 26329 18915 26387 18921
rect 26510 18912 26516 18924
rect 26568 18912 26574 18964
rect 29362 18912 29368 18964
rect 29420 18952 29426 18964
rect 29917 18955 29975 18961
rect 29917 18952 29929 18955
rect 29420 18924 29929 18952
rect 29420 18912 29426 18924
rect 29917 18921 29929 18924
rect 29963 18921 29975 18955
rect 29917 18915 29975 18921
rect 30834 18912 30840 18964
rect 30892 18952 30898 18964
rect 31205 18955 31263 18961
rect 31205 18952 31217 18955
rect 30892 18924 31217 18952
rect 30892 18912 30898 18924
rect 31205 18921 31217 18924
rect 31251 18921 31263 18955
rect 31205 18915 31263 18921
rect 31312 18924 32628 18952
rect 24946 18884 24952 18896
rect 22520 18856 22968 18884
rect 23124 18856 24952 18884
rect 22520 18844 22526 18856
rect 22940 18816 22968 18856
rect 24946 18844 24952 18856
rect 25004 18844 25010 18896
rect 30929 18887 30987 18893
rect 30929 18884 30941 18887
rect 30208 18856 30941 18884
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 22112 18788 22876 18816
rect 22940 18788 23121 18816
rect 22112 18757 22140 18788
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18717 20591 18751
rect 20533 18711 20591 18717
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 22097 18751 22155 18757
rect 22097 18717 22109 18751
rect 22143 18717 22155 18751
rect 22097 18711 22155 18717
rect 22186 18708 22192 18760
rect 22244 18708 22250 18760
rect 22554 18708 22560 18760
rect 22612 18708 22618 18760
rect 22738 18708 22744 18760
rect 22796 18708 22802 18760
rect 22848 18757 22876 18788
rect 23109 18785 23121 18788
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 23661 18819 23719 18825
rect 23661 18785 23673 18819
rect 23707 18816 23719 18819
rect 26789 18819 26847 18825
rect 26789 18816 26801 18819
rect 23707 18788 26801 18816
rect 23707 18785 23719 18788
rect 23661 18779 23719 18785
rect 26789 18785 26801 18788
rect 26835 18785 26847 18819
rect 26789 18779 26847 18785
rect 26878 18776 26884 18828
rect 26936 18776 26942 18828
rect 28445 18819 28503 18825
rect 28445 18785 28457 18819
rect 28491 18816 28503 18819
rect 28718 18816 28724 18828
rect 28491 18788 28724 18816
rect 28491 18785 28503 18788
rect 28445 18779 28503 18785
rect 28718 18776 28724 18788
rect 28776 18776 28782 18828
rect 22833 18751 22891 18757
rect 22833 18717 22845 18751
rect 22879 18748 22891 18751
rect 23569 18751 23627 18757
rect 22879 18720 23060 18748
rect 22879 18717 22891 18720
rect 22833 18711 22891 18717
rect 15120 18652 16068 18680
rect 16669 18683 16727 18689
rect 16669 18649 16681 18683
rect 16715 18680 16727 18683
rect 16715 18652 19334 18680
rect 16715 18649 16727 18652
rect 16669 18643 16727 18649
rect 10244 18584 13768 18612
rect 18874 18572 18880 18624
rect 18932 18572 18938 18624
rect 19306 18612 19334 18652
rect 19610 18640 19616 18692
rect 19668 18680 19674 18692
rect 19981 18683 20039 18689
rect 19981 18680 19993 18683
rect 19668 18652 19993 18680
rect 19668 18640 19674 18652
rect 19981 18649 19993 18652
rect 20027 18649 20039 18683
rect 19981 18643 20039 18649
rect 21821 18683 21879 18689
rect 21821 18649 21833 18683
rect 21867 18680 21879 18683
rect 21867 18652 22094 18680
rect 21867 18649 21879 18652
rect 21821 18643 21879 18649
rect 20438 18612 20444 18624
rect 19306 18584 20444 18612
rect 20438 18572 20444 18584
rect 20496 18572 20502 18624
rect 22066 18612 22094 18652
rect 22278 18640 22284 18692
rect 22336 18680 22342 18692
rect 22373 18683 22431 18689
rect 22373 18680 22385 18683
rect 22336 18652 22385 18680
rect 22336 18640 22342 18652
rect 22373 18649 22385 18652
rect 22419 18649 22431 18683
rect 22373 18643 22431 18649
rect 22465 18683 22523 18689
rect 22465 18649 22477 18683
rect 22511 18680 22523 18683
rect 22756 18680 22784 18708
rect 22511 18652 22784 18680
rect 22511 18649 22523 18652
rect 22465 18643 22523 18649
rect 23032 18624 23060 18720
rect 23569 18717 23581 18751
rect 23615 18717 23627 18751
rect 23569 18711 23627 18717
rect 23584 18680 23612 18711
rect 24394 18708 24400 18760
rect 24452 18708 24458 18760
rect 28626 18708 28632 18760
rect 28684 18708 28690 18760
rect 28994 18708 29000 18760
rect 29052 18748 29058 18760
rect 30055 18751 30113 18757
rect 30055 18748 30067 18751
rect 29052 18720 30067 18748
rect 29052 18708 29058 18720
rect 30055 18717 30067 18720
rect 30101 18717 30113 18751
rect 30055 18711 30113 18717
rect 30208 18692 30236 18856
rect 30929 18853 30941 18856
rect 30975 18853 30987 18887
rect 30929 18847 30987 18853
rect 30300 18788 30788 18816
rect 30300 18757 30328 18788
rect 30285 18751 30343 18757
rect 30285 18717 30297 18751
rect 30331 18717 30343 18751
rect 30468 18751 30526 18757
rect 30468 18748 30480 18751
rect 30285 18711 30343 18717
rect 30392 18720 30480 18748
rect 23124 18652 23612 18680
rect 26697 18683 26755 18689
rect 23124 18624 23152 18652
rect 26697 18649 26709 18683
rect 26743 18680 26755 18683
rect 27801 18683 27859 18689
rect 27801 18680 27813 18683
rect 26743 18652 27813 18680
rect 26743 18649 26755 18652
rect 26697 18643 26755 18649
rect 27801 18649 27813 18652
rect 27847 18649 27859 18683
rect 27801 18643 27859 18649
rect 28258 18640 28264 18692
rect 28316 18680 28322 18692
rect 30190 18680 30196 18692
rect 28316 18652 30196 18680
rect 28316 18640 28322 18652
rect 30190 18640 30196 18652
rect 30248 18640 30254 18692
rect 22741 18615 22799 18621
rect 22741 18612 22753 18615
rect 22066 18584 22753 18612
rect 22741 18581 22753 18584
rect 22787 18612 22799 18615
rect 22922 18612 22928 18624
rect 22787 18584 22928 18612
rect 22787 18581 22799 18584
rect 22741 18575 22799 18581
rect 22922 18572 22928 18584
rect 22980 18572 22986 18624
rect 23014 18572 23020 18624
rect 23072 18572 23078 18624
rect 23106 18572 23112 18624
rect 23164 18572 23170 18624
rect 23290 18572 23296 18624
rect 23348 18612 23354 18624
rect 23385 18615 23443 18621
rect 23385 18612 23397 18615
rect 23348 18584 23397 18612
rect 23348 18572 23354 18584
rect 23385 18581 23397 18584
rect 23431 18581 23443 18615
rect 23385 18575 23443 18581
rect 24578 18572 24584 18624
rect 24636 18572 24642 18624
rect 29181 18615 29239 18621
rect 29181 18581 29193 18615
rect 29227 18612 29239 18615
rect 29362 18612 29368 18624
rect 29227 18584 29368 18612
rect 29227 18581 29239 18584
rect 29181 18575 29239 18581
rect 29362 18572 29368 18584
rect 29420 18572 29426 18624
rect 30392 18612 30420 18720
rect 30468 18717 30480 18720
rect 30514 18717 30526 18751
rect 30468 18711 30526 18717
rect 30558 18708 30564 18760
rect 30616 18708 30622 18760
rect 30650 18708 30656 18760
rect 30708 18708 30714 18760
rect 30760 18748 30788 18788
rect 31312 18748 31340 18924
rect 32306 18884 32312 18896
rect 31404 18856 32312 18884
rect 31404 18757 31432 18856
rect 32306 18844 32312 18856
rect 32364 18844 32370 18896
rect 32401 18887 32459 18893
rect 32401 18853 32413 18887
rect 32447 18853 32459 18887
rect 32600 18884 32628 18924
rect 32674 18912 32680 18964
rect 32732 18952 32738 18964
rect 32769 18955 32827 18961
rect 32769 18952 32781 18955
rect 32732 18924 32781 18952
rect 32732 18912 32738 18924
rect 32769 18921 32781 18924
rect 32815 18921 32827 18955
rect 32769 18915 32827 18921
rect 33689 18887 33747 18893
rect 33689 18884 33701 18887
rect 32600 18856 33701 18884
rect 32401 18847 32459 18853
rect 33689 18853 33701 18856
rect 33735 18853 33747 18887
rect 33689 18847 33747 18853
rect 32416 18816 32444 18847
rect 31496 18788 32444 18816
rect 32692 18788 33272 18816
rect 30760 18720 31340 18748
rect 31389 18751 31447 18757
rect 31389 18717 31401 18751
rect 31435 18717 31447 18751
rect 31389 18711 31447 18717
rect 31496 18680 31524 18788
rect 31570 18708 31576 18760
rect 31628 18708 31634 18760
rect 31662 18708 31668 18760
rect 31720 18708 31726 18760
rect 31757 18751 31815 18757
rect 31757 18717 31769 18751
rect 31803 18717 31815 18751
rect 31757 18711 31815 18717
rect 31036 18652 31524 18680
rect 31588 18680 31616 18708
rect 31772 18680 31800 18711
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32401 18751 32459 18757
rect 32401 18748 32413 18751
rect 32272 18720 32413 18748
rect 32272 18708 32278 18720
rect 32401 18717 32413 18720
rect 32447 18717 32459 18751
rect 32692 18735 32720 18788
rect 32401 18711 32459 18717
rect 32673 18729 32731 18735
rect 32673 18695 32685 18729
rect 32719 18695 32731 18729
rect 32950 18708 32956 18760
rect 33008 18708 33014 18760
rect 33244 18757 33272 18788
rect 33229 18751 33287 18757
rect 33229 18717 33241 18751
rect 33275 18748 33287 18751
rect 33321 18751 33379 18757
rect 33321 18748 33333 18751
rect 33275 18720 33333 18748
rect 33275 18717 33287 18720
rect 33229 18711 33287 18717
rect 33321 18717 33333 18720
rect 33367 18717 33379 18751
rect 33321 18711 33379 18717
rect 32673 18692 32731 18695
rect 32673 18689 32680 18692
rect 31588 18652 31800 18680
rect 31036 18612 31064 18652
rect 32674 18640 32680 18689
rect 32732 18640 32738 18692
rect 33505 18683 33563 18689
rect 33505 18649 33517 18683
rect 33551 18649 33563 18683
rect 33505 18643 33563 18649
rect 30392 18584 31064 18612
rect 31113 18615 31171 18621
rect 31113 18581 31125 18615
rect 31159 18612 31171 18615
rect 31386 18612 31392 18624
rect 31159 18584 31392 18612
rect 31159 18581 31171 18584
rect 31113 18575 31171 18581
rect 31386 18572 31392 18584
rect 31444 18612 31450 18624
rect 31570 18612 31576 18624
rect 31444 18584 31576 18612
rect 31444 18572 31450 18584
rect 31570 18572 31576 18584
rect 31628 18572 31634 18624
rect 31846 18572 31852 18624
rect 31904 18572 31910 18624
rect 32585 18615 32643 18621
rect 32585 18581 32597 18615
rect 32631 18612 32643 18615
rect 32858 18612 32864 18624
rect 32631 18584 32864 18612
rect 32631 18581 32643 18584
rect 32585 18575 32643 18581
rect 32858 18572 32864 18584
rect 32916 18612 32922 18624
rect 33137 18615 33195 18621
rect 33137 18612 33149 18615
rect 32916 18584 33149 18612
rect 32916 18572 32922 18584
rect 33137 18581 33149 18584
rect 33183 18612 33195 18615
rect 33520 18612 33548 18643
rect 33183 18584 33548 18612
rect 33183 18581 33195 18584
rect 33137 18575 33195 18581
rect 1104 18522 34840 18544
rect 1104 18470 9344 18522
rect 9396 18470 9408 18522
rect 9460 18470 9472 18522
rect 9524 18470 9536 18522
rect 9588 18470 9600 18522
rect 9652 18470 17738 18522
rect 17790 18470 17802 18522
rect 17854 18470 17866 18522
rect 17918 18470 17930 18522
rect 17982 18470 17994 18522
rect 18046 18470 26132 18522
rect 26184 18470 26196 18522
rect 26248 18470 26260 18522
rect 26312 18470 26324 18522
rect 26376 18470 26388 18522
rect 26440 18470 34526 18522
rect 34578 18470 34590 18522
rect 34642 18470 34654 18522
rect 34706 18470 34718 18522
rect 34770 18470 34782 18522
rect 34834 18470 34840 18522
rect 1104 18448 34840 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 3421 18411 3479 18417
rect 3421 18408 3433 18411
rect 1912 18380 3433 18408
rect 1912 18368 1918 18380
rect 3421 18377 3433 18380
rect 3467 18377 3479 18411
rect 3421 18371 3479 18377
rect 3694 18368 3700 18420
rect 3752 18408 3758 18420
rect 3752 18380 4752 18408
rect 3752 18368 3758 18380
rect 3602 18232 3608 18284
rect 3660 18232 3666 18284
rect 3712 18281 3740 18368
rect 3789 18343 3847 18349
rect 3789 18309 3801 18343
rect 3835 18340 3847 18343
rect 3878 18340 3884 18352
rect 3835 18312 3884 18340
rect 3835 18309 3847 18312
rect 3789 18303 3847 18309
rect 3878 18300 3884 18312
rect 3936 18300 3942 18352
rect 3697 18275 3755 18281
rect 3697 18241 3709 18275
rect 3743 18241 3755 18275
rect 3697 18235 3755 18241
rect 3970 18232 3976 18284
rect 4028 18232 4034 18284
rect 4522 18232 4528 18284
rect 4580 18232 4586 18284
rect 4724 18272 4752 18380
rect 4982 18368 4988 18420
rect 5040 18408 5046 18420
rect 5369 18411 5427 18417
rect 5369 18408 5381 18411
rect 5040 18380 5381 18408
rect 5040 18368 5046 18380
rect 5369 18377 5381 18380
rect 5415 18408 5427 18411
rect 5718 18408 5724 18420
rect 5415 18380 5724 18408
rect 5415 18377 5427 18380
rect 5369 18371 5427 18377
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 6089 18411 6147 18417
rect 6089 18377 6101 18411
rect 6135 18408 6147 18411
rect 6914 18408 6920 18420
rect 6135 18380 6920 18408
rect 6135 18377 6147 18380
rect 6089 18371 6147 18377
rect 6914 18368 6920 18380
rect 6972 18368 6978 18420
rect 9401 18411 9459 18417
rect 9401 18408 9413 18411
rect 7576 18380 9413 18408
rect 4798 18300 4804 18352
rect 4856 18340 4862 18352
rect 5169 18343 5227 18349
rect 5169 18340 5181 18343
rect 4856 18312 5181 18340
rect 4856 18300 4862 18312
rect 5169 18309 5181 18312
rect 5215 18309 5227 18343
rect 5169 18303 5227 18309
rect 5552 18312 6500 18340
rect 5552 18284 5580 18312
rect 5534 18272 5540 18284
rect 4724 18244 5540 18272
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 5629 18275 5687 18281
rect 5629 18241 5641 18275
rect 5675 18272 5687 18275
rect 5810 18272 5816 18284
rect 5675 18244 5816 18272
rect 5675 18241 5687 18244
rect 5629 18235 5687 18241
rect 5810 18232 5816 18244
rect 5868 18232 5874 18284
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 6362 18272 6368 18284
rect 5951 18244 6368 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 6472 18281 6500 18312
rect 7576 18281 7604 18380
rect 9401 18377 9413 18380
rect 9447 18408 9459 18411
rect 9858 18408 9864 18420
rect 9447 18380 9864 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 9858 18368 9864 18380
rect 9916 18368 9922 18420
rect 12342 18368 12348 18420
rect 12400 18408 12406 18420
rect 15473 18411 15531 18417
rect 12400 18380 14412 18408
rect 12400 18368 12406 18380
rect 8110 18300 8116 18352
rect 8168 18300 8174 18352
rect 8294 18300 8300 18352
rect 8352 18340 8358 18352
rect 8352 18312 8800 18340
rect 8352 18300 8358 18312
rect 6457 18275 6515 18281
rect 6457 18241 6469 18275
rect 6503 18241 6515 18275
rect 6457 18235 6515 18241
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 7561 18275 7619 18281
rect 7561 18241 7573 18275
rect 7607 18241 7619 18275
rect 7561 18235 7619 18241
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18272 7895 18275
rect 8662 18272 8668 18284
rect 7883 18244 8668 18272
rect 7883 18241 7895 18244
rect 7837 18235 7895 18241
rect 4540 18204 4568 18232
rect 5994 18204 6000 18216
rect 4540 18176 6000 18204
rect 5994 18164 6000 18176
rect 6052 18204 6058 18216
rect 6840 18204 6868 18235
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 8772 18272 8800 18312
rect 8846 18300 8852 18352
rect 8904 18340 8910 18352
rect 8941 18343 8999 18349
rect 8941 18340 8953 18343
rect 8904 18312 8953 18340
rect 8904 18300 8910 18312
rect 8941 18309 8953 18312
rect 8987 18309 8999 18343
rect 8941 18303 8999 18309
rect 9585 18343 9643 18349
rect 9585 18309 9597 18343
rect 9631 18340 9643 18343
rect 11793 18343 11851 18349
rect 9631 18312 10272 18340
rect 9631 18309 9643 18312
rect 9585 18303 9643 18309
rect 9033 18275 9091 18281
rect 9033 18272 9045 18275
rect 8772 18244 9045 18272
rect 9033 18241 9045 18244
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 9122 18232 9128 18284
rect 9180 18232 9186 18284
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 9766 18272 9772 18284
rect 9364 18244 9772 18272
rect 9364 18232 9370 18244
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18272 9919 18275
rect 10134 18272 10140 18284
rect 9907 18244 10140 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 10134 18232 10140 18244
rect 10192 18232 10198 18284
rect 10244 18272 10272 18312
rect 11793 18309 11805 18343
rect 11839 18340 11851 18343
rect 14384 18340 14412 18380
rect 15473 18377 15485 18411
rect 15519 18408 15531 18411
rect 15746 18408 15752 18420
rect 15519 18380 15752 18408
rect 15519 18377 15531 18380
rect 15473 18371 15531 18377
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 17494 18368 17500 18420
rect 17552 18408 17558 18420
rect 17865 18411 17923 18417
rect 17865 18408 17877 18411
rect 17552 18380 17877 18408
rect 17552 18368 17558 18380
rect 17865 18377 17877 18380
rect 17911 18377 17923 18411
rect 17865 18371 17923 18377
rect 18233 18411 18291 18417
rect 18233 18377 18245 18411
rect 18279 18408 18291 18411
rect 18690 18408 18696 18420
rect 18279 18380 18696 18408
rect 18279 18377 18291 18380
rect 18233 18371 18291 18377
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 18874 18408 18880 18420
rect 18800 18380 18880 18408
rect 16117 18343 16175 18349
rect 16117 18340 16129 18343
rect 11839 18312 14320 18340
rect 14384 18312 16129 18340
rect 11839 18309 11851 18312
rect 11793 18303 11851 18309
rect 11146 18272 11152 18284
rect 10244 18244 11152 18272
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 12529 18275 12587 18281
rect 11563 18244 11744 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 6052 18176 6868 18204
rect 7929 18207 7987 18213
rect 6052 18164 6058 18176
rect 7929 18173 7941 18207
rect 7975 18204 7987 18207
rect 8478 18204 8484 18216
rect 7975 18176 8484 18204
rect 7975 18173 7987 18176
rect 7929 18167 7987 18173
rect 8478 18164 8484 18176
rect 8536 18164 8542 18216
rect 8680 18204 8708 18232
rect 9324 18204 9352 18232
rect 8680 18176 9352 18204
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 11609 18207 11667 18213
rect 11609 18204 11621 18207
rect 9732 18176 11621 18204
rect 9732 18164 9738 18176
rect 11609 18173 11621 18176
rect 11655 18173 11667 18207
rect 11609 18167 11667 18173
rect 5721 18139 5779 18145
rect 5721 18105 5733 18139
rect 5767 18136 5779 18139
rect 5810 18136 5816 18148
rect 5767 18108 5816 18136
rect 5767 18105 5779 18108
rect 5721 18099 5779 18105
rect 5810 18096 5816 18108
rect 5868 18096 5874 18148
rect 8662 18096 8668 18148
rect 8720 18136 8726 18148
rect 11716 18136 11744 18244
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 11793 18207 11851 18213
rect 11793 18173 11805 18207
rect 11839 18204 11851 18207
rect 11974 18204 11980 18216
rect 11839 18176 11980 18204
rect 11839 18173 11851 18176
rect 11793 18167 11851 18173
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 12544 18204 12572 18235
rect 12710 18232 12716 18284
rect 12768 18232 12774 18284
rect 12802 18232 12808 18284
rect 12860 18232 12866 18284
rect 12894 18232 12900 18284
rect 12952 18232 12958 18284
rect 13262 18232 13268 18284
rect 13320 18232 13326 18284
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18241 13691 18275
rect 13633 18235 13691 18241
rect 12820 18204 12848 18232
rect 12986 18204 12992 18216
rect 12544 18176 12756 18204
rect 12820 18176 12992 18204
rect 8720 18108 12020 18136
rect 8720 18096 8726 18108
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 5258 18068 5264 18080
rect 5040 18040 5264 18068
rect 5040 18028 5046 18040
rect 5258 18028 5264 18040
rect 5316 18068 5322 18080
rect 5353 18071 5411 18077
rect 5353 18068 5365 18071
rect 5316 18040 5365 18068
rect 5316 18028 5322 18040
rect 5353 18037 5365 18040
rect 5399 18037 5411 18071
rect 5353 18031 5411 18037
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 5537 18071 5595 18077
rect 5537 18068 5549 18071
rect 5500 18040 5549 18068
rect 5500 18028 5506 18040
rect 5537 18037 5549 18040
rect 5583 18068 5595 18071
rect 8938 18068 8944 18080
rect 5583 18040 8944 18068
rect 5583 18037 5595 18040
rect 5537 18031 5595 18037
rect 8938 18028 8944 18040
rect 8996 18028 9002 18080
rect 9232 18077 9260 18108
rect 11992 18080 12020 18108
rect 12728 18080 12756 18176
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 12805 18139 12863 18145
rect 12805 18105 12817 18139
rect 12851 18136 12863 18139
rect 13648 18136 13676 18235
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 14185 18275 14243 18281
rect 14185 18272 14197 18275
rect 13780 18244 14197 18272
rect 13780 18232 13786 18244
rect 14185 18241 14197 18244
rect 14231 18241 14243 18275
rect 14292 18272 14320 18312
rect 16117 18309 16129 18312
rect 16163 18309 16175 18343
rect 16117 18303 16175 18309
rect 17957 18343 18015 18349
rect 17957 18309 17969 18343
rect 18003 18340 18015 18343
rect 18506 18340 18512 18352
rect 18003 18312 18512 18340
rect 18003 18309 18015 18312
rect 17957 18303 18015 18309
rect 18506 18300 18512 18312
rect 18564 18300 18570 18352
rect 18800 18349 18828 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 23290 18368 23296 18420
rect 23348 18368 23354 18420
rect 24578 18408 24584 18420
rect 24504 18380 24584 18408
rect 18785 18343 18843 18349
rect 18785 18309 18797 18343
rect 18831 18309 18843 18343
rect 18785 18303 18843 18309
rect 19518 18300 19524 18352
rect 19576 18300 19582 18352
rect 21726 18300 21732 18352
rect 21784 18340 21790 18352
rect 21784 18312 22784 18340
rect 21784 18300 21790 18312
rect 14550 18272 14556 18284
rect 14292 18244 14556 18272
rect 14185 18235 14243 18241
rect 14550 18232 14556 18244
rect 14608 18272 14614 18284
rect 14645 18275 14703 18281
rect 14645 18272 14657 18275
rect 14608 18244 14657 18272
rect 14608 18232 14614 18244
rect 14645 18241 14657 18244
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 15102 18232 15108 18284
rect 15160 18232 15166 18284
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18272 15255 18275
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15243 18244 15424 18272
rect 15243 18241 15255 18244
rect 15197 18235 15255 18241
rect 14461 18207 14519 18213
rect 14461 18173 14473 18207
rect 14507 18204 14519 18207
rect 14734 18204 14740 18216
rect 14507 18176 14740 18204
rect 14507 18173 14519 18176
rect 14461 18167 14519 18173
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 14826 18164 14832 18216
rect 14884 18204 14890 18216
rect 15013 18207 15071 18213
rect 15013 18204 15025 18207
rect 14884 18176 15025 18204
rect 14884 18164 14890 18176
rect 15013 18173 15025 18176
rect 15059 18173 15071 18207
rect 15013 18167 15071 18173
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18173 15347 18207
rect 15289 18167 15347 18173
rect 12851 18108 13676 18136
rect 14369 18139 14427 18145
rect 12851 18105 12863 18108
rect 12805 18099 12863 18105
rect 14369 18105 14381 18139
rect 14415 18136 14427 18139
rect 15304 18136 15332 18167
rect 14415 18108 15332 18136
rect 15396 18136 15424 18244
rect 15856 18244 15945 18272
rect 15856 18148 15884 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18272 17647 18275
rect 17678 18272 17684 18284
rect 17635 18244 17684 18272
rect 17635 18241 17647 18244
rect 17589 18235 17647 18241
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 22462 18232 22468 18284
rect 22520 18232 22526 18284
rect 22756 18281 22784 18312
rect 22741 18275 22799 18281
rect 22741 18241 22753 18275
rect 22787 18241 22799 18275
rect 22741 18235 22799 18241
rect 22922 18232 22928 18284
rect 22980 18232 22986 18284
rect 23308 18281 23336 18368
rect 24504 18349 24532 18380
rect 24578 18368 24584 18380
rect 24636 18368 24642 18420
rect 26786 18368 26792 18420
rect 26844 18408 26850 18420
rect 32769 18411 32827 18417
rect 26844 18380 29868 18408
rect 26844 18368 26850 18380
rect 24489 18343 24547 18349
rect 23492 18312 24256 18340
rect 23492 18284 23520 18312
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 23474 18232 23480 18284
rect 23532 18232 23538 18284
rect 23569 18275 23627 18281
rect 23569 18241 23581 18275
rect 23615 18241 23627 18275
rect 23569 18235 23627 18241
rect 18046 18164 18052 18216
rect 18104 18213 18110 18216
rect 18104 18207 18132 18213
rect 18120 18173 18132 18207
rect 18104 18167 18132 18173
rect 18104 18164 18110 18167
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18288 18176 18521 18204
rect 18288 18164 18294 18176
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 23014 18164 23020 18216
rect 23072 18204 23078 18216
rect 23385 18207 23443 18213
rect 23385 18204 23397 18207
rect 23072 18176 23397 18204
rect 23072 18164 23078 18176
rect 23385 18173 23397 18176
rect 23431 18173 23443 18207
rect 23385 18167 23443 18173
rect 15470 18136 15476 18148
rect 15396 18108 15476 18136
rect 14415 18105 14427 18108
rect 14369 18099 14427 18105
rect 15120 18080 15148 18108
rect 15470 18096 15476 18108
rect 15528 18136 15534 18148
rect 15838 18136 15844 18148
rect 15528 18108 15844 18136
rect 15528 18096 15534 18108
rect 15838 18096 15844 18108
rect 15896 18096 15902 18148
rect 20254 18096 20260 18148
rect 20312 18136 20318 18148
rect 20312 18108 22094 18136
rect 20312 18096 20318 18108
rect 9217 18071 9275 18077
rect 9217 18037 9229 18071
rect 9263 18037 9275 18071
rect 9217 18031 9275 18037
rect 9585 18071 9643 18077
rect 9585 18037 9597 18071
rect 9631 18068 9643 18071
rect 9950 18068 9956 18080
rect 9631 18040 9956 18068
rect 9631 18037 9643 18040
rect 9585 18031 9643 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 11974 18028 11980 18080
rect 12032 18028 12038 18080
rect 12710 18028 12716 18080
rect 12768 18028 12774 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 14829 18071 14887 18077
rect 14829 18068 14841 18071
rect 14792 18040 14841 18068
rect 14792 18028 14798 18040
rect 14829 18037 14841 18040
rect 14875 18037 14887 18071
rect 14829 18031 14887 18037
rect 15102 18028 15108 18080
rect 15160 18028 15166 18080
rect 15194 18028 15200 18080
rect 15252 18068 15258 18080
rect 15562 18068 15568 18080
rect 15252 18040 15568 18068
rect 15252 18028 15258 18040
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 16298 18028 16304 18080
rect 16356 18028 16362 18080
rect 18506 18028 18512 18080
rect 18564 18068 18570 18080
rect 21913 18071 21971 18077
rect 21913 18068 21925 18071
rect 18564 18040 21925 18068
rect 18564 18028 18570 18040
rect 21913 18037 21925 18040
rect 21959 18037 21971 18071
rect 22066 18068 22094 18108
rect 22278 18096 22284 18148
rect 22336 18136 22342 18148
rect 23106 18136 23112 18148
rect 22336 18108 23112 18136
rect 22336 18096 22342 18108
rect 23106 18096 23112 18108
rect 23164 18136 23170 18148
rect 23584 18136 23612 18235
rect 23658 18232 23664 18284
rect 23716 18232 23722 18284
rect 23937 18275 23995 18281
rect 23937 18272 23949 18275
rect 23768 18244 23949 18272
rect 23164 18108 23612 18136
rect 23164 18096 23170 18108
rect 23474 18068 23480 18080
rect 22066 18040 23480 18068
rect 21913 18031 21971 18037
rect 23474 18028 23480 18040
rect 23532 18068 23538 18080
rect 23768 18068 23796 18244
rect 23937 18241 23949 18244
rect 23983 18241 23995 18275
rect 23937 18235 23995 18241
rect 24118 18164 24124 18216
rect 24176 18204 24182 18216
rect 24228 18213 24256 18312
rect 24489 18309 24501 18343
rect 24535 18309 24547 18343
rect 24489 18303 24547 18309
rect 24946 18300 24952 18352
rect 25004 18300 25010 18352
rect 28350 18232 28356 18284
rect 28408 18232 28414 18284
rect 29730 18232 29736 18284
rect 29788 18232 29794 18284
rect 29840 18272 29868 18380
rect 32769 18377 32781 18411
rect 32815 18408 32827 18411
rect 32858 18408 32864 18420
rect 32815 18380 32864 18408
rect 32815 18377 32827 18380
rect 32769 18371 32827 18377
rect 32858 18368 32864 18380
rect 32916 18368 32922 18420
rect 31570 18300 31576 18352
rect 31628 18340 31634 18352
rect 32950 18340 32956 18352
rect 31628 18312 32956 18340
rect 31628 18300 31634 18312
rect 29917 18275 29975 18281
rect 29917 18272 29929 18275
rect 29840 18244 29929 18272
rect 29917 18241 29929 18244
rect 29963 18241 29975 18275
rect 29917 18235 29975 18241
rect 31846 18232 31852 18284
rect 31904 18272 31910 18284
rect 32582 18272 32588 18284
rect 31904 18244 32588 18272
rect 31904 18232 31910 18244
rect 32582 18232 32588 18244
rect 32640 18272 32646 18284
rect 32876 18281 32904 18312
rect 32950 18300 32956 18312
rect 33008 18300 33014 18352
rect 32677 18275 32735 18281
rect 32677 18272 32689 18275
rect 32640 18244 32689 18272
rect 32640 18232 32646 18244
rect 32677 18241 32689 18244
rect 32723 18241 32735 18275
rect 32677 18235 32735 18241
rect 32861 18275 32919 18281
rect 32861 18241 32873 18275
rect 32907 18241 32919 18275
rect 32861 18235 32919 18241
rect 24213 18207 24271 18213
rect 24213 18204 24225 18207
rect 24176 18176 24225 18204
rect 24176 18164 24182 18176
rect 24213 18173 24225 18176
rect 24259 18173 24271 18207
rect 24213 18167 24271 18173
rect 25961 18207 26019 18213
rect 25961 18173 25973 18207
rect 26007 18204 26019 18207
rect 27157 18207 27215 18213
rect 27157 18204 27169 18207
rect 26007 18176 27169 18204
rect 26007 18173 26019 18176
rect 25961 18167 26019 18173
rect 27157 18173 27169 18176
rect 27203 18173 27215 18207
rect 28368 18204 28396 18232
rect 30193 18207 30251 18213
rect 30193 18204 30205 18207
rect 28368 18176 30205 18204
rect 27157 18167 27215 18173
rect 30193 18173 30205 18176
rect 30239 18173 30251 18207
rect 30193 18167 30251 18173
rect 23532 18040 23796 18068
rect 23532 18028 23538 18040
rect 23842 18028 23848 18080
rect 23900 18028 23906 18080
rect 27798 18028 27804 18080
rect 27856 18028 27862 18080
rect 27985 18071 28043 18077
rect 27985 18037 27997 18071
rect 28031 18068 28043 18071
rect 28258 18068 28264 18080
rect 28031 18040 28264 18068
rect 28031 18037 28043 18040
rect 27985 18031 28043 18037
rect 28258 18028 28264 18040
rect 28316 18028 28322 18080
rect 29362 18028 29368 18080
rect 29420 18068 29426 18080
rect 29469 18071 29527 18077
rect 29469 18068 29481 18071
rect 29420 18040 29481 18068
rect 29420 18028 29426 18040
rect 29469 18037 29481 18040
rect 29515 18037 29527 18071
rect 29469 18031 29527 18037
rect 32214 18028 32220 18080
rect 32272 18068 32278 18080
rect 32858 18068 32864 18080
rect 32272 18040 32864 18068
rect 32272 18028 32278 18040
rect 32858 18028 32864 18040
rect 32916 18028 32922 18080
rect 1104 17978 34684 18000
rect 1104 17926 5147 17978
rect 5199 17926 5211 17978
rect 5263 17926 5275 17978
rect 5327 17926 5339 17978
rect 5391 17926 5403 17978
rect 5455 17926 13541 17978
rect 13593 17926 13605 17978
rect 13657 17926 13669 17978
rect 13721 17926 13733 17978
rect 13785 17926 13797 17978
rect 13849 17926 21935 17978
rect 21987 17926 21999 17978
rect 22051 17926 22063 17978
rect 22115 17926 22127 17978
rect 22179 17926 22191 17978
rect 22243 17926 30329 17978
rect 30381 17926 30393 17978
rect 30445 17926 30457 17978
rect 30509 17926 30521 17978
rect 30573 17926 30585 17978
rect 30637 17926 34684 17978
rect 1104 17904 34684 17926
rect 3878 17824 3884 17876
rect 3936 17824 3942 17876
rect 3970 17824 3976 17876
rect 4028 17864 4034 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4028 17836 4537 17864
rect 4028 17824 4034 17836
rect 4525 17833 4537 17836
rect 4571 17833 4583 17867
rect 9766 17864 9772 17876
rect 4525 17827 4583 17833
rect 8220 17836 9772 17864
rect 3418 17756 3424 17808
rect 3476 17796 3482 17808
rect 3896 17796 3924 17824
rect 3476 17768 4384 17796
rect 3476 17756 3482 17768
rect 3513 17731 3571 17737
rect 3513 17697 3525 17731
rect 3559 17728 3571 17731
rect 3559 17700 4200 17728
rect 3559 17697 3571 17700
rect 3513 17691 3571 17697
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17629 3479 17663
rect 3421 17623 3479 17629
rect 3436 17592 3464 17623
rect 3602 17620 3608 17672
rect 3660 17620 3666 17672
rect 3694 17620 3700 17672
rect 3752 17660 3758 17672
rect 4172 17669 4200 17700
rect 4356 17669 4384 17768
rect 7374 17756 7380 17808
rect 7432 17756 7438 17808
rect 4706 17688 4712 17740
rect 4764 17688 4770 17740
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 4985 17731 5043 17737
rect 4985 17728 4997 17731
rect 4856 17700 4997 17728
rect 4856 17688 4862 17700
rect 4985 17697 4997 17700
rect 5031 17697 5043 17731
rect 5534 17728 5540 17740
rect 4985 17691 5043 17697
rect 5276 17700 5540 17728
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3752 17632 3985 17660
rect 3752 17620 3758 17632
rect 3973 17629 3985 17632
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 4341 17663 4399 17669
rect 4341 17629 4353 17663
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 3510 17592 3516 17604
rect 3436 17564 3516 17592
rect 3510 17552 3516 17564
rect 3568 17592 3574 17604
rect 4065 17595 4123 17601
rect 3568 17564 3924 17592
rect 3568 17552 3574 17564
rect 3786 17484 3792 17536
rect 3844 17484 3850 17536
rect 3896 17524 3924 17564
rect 4065 17561 4077 17595
rect 4111 17592 4123 17595
rect 4246 17592 4252 17604
rect 4111 17564 4252 17592
rect 4111 17561 4123 17564
rect 4065 17555 4123 17561
rect 4246 17552 4252 17564
rect 4304 17552 4310 17604
rect 4448 17592 4476 17623
rect 4522 17620 4528 17672
rect 4580 17660 4586 17672
rect 4617 17663 4675 17669
rect 4617 17660 4629 17663
rect 4580 17632 4629 17660
rect 4580 17620 4586 17632
rect 4617 17629 4629 17632
rect 4663 17629 4675 17663
rect 4617 17623 4675 17629
rect 4724 17592 4752 17688
rect 5276 17669 5304 17700
rect 5534 17688 5540 17700
rect 5592 17728 5598 17740
rect 5592 17700 5948 17728
rect 5592 17688 5598 17700
rect 5920 17672 5948 17700
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 6972 17700 7941 17728
rect 6972 17688 6978 17700
rect 7929 17697 7941 17700
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 5261 17663 5319 17669
rect 5261 17629 5273 17663
rect 5307 17629 5319 17663
rect 5261 17623 5319 17629
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 5902 17620 5908 17672
rect 5960 17660 5966 17672
rect 6270 17660 6276 17672
rect 5960 17632 6276 17660
rect 5960 17620 5966 17632
rect 6270 17620 6276 17632
rect 6328 17660 6334 17672
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 6328 17632 6653 17660
rect 6328 17620 6334 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 7282 17620 7288 17672
rect 7340 17620 7346 17672
rect 7469 17663 7527 17669
rect 7469 17629 7481 17663
rect 7515 17629 7527 17663
rect 7469 17623 7527 17629
rect 4448 17564 4752 17592
rect 5828 17592 5856 17620
rect 7484 17592 7512 17623
rect 7650 17592 7656 17604
rect 5828 17564 7656 17592
rect 4448 17524 4476 17564
rect 7650 17552 7656 17564
rect 7708 17552 7714 17604
rect 3896 17496 4476 17524
rect 5905 17527 5963 17533
rect 5905 17493 5917 17527
rect 5951 17524 5963 17527
rect 8110 17524 8116 17536
rect 5951 17496 8116 17524
rect 5951 17493 5963 17496
rect 5905 17487 5963 17493
rect 8110 17484 8116 17496
rect 8168 17524 8174 17536
rect 8220 17524 8248 17836
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 10873 17867 10931 17873
rect 10873 17833 10885 17867
rect 10919 17864 10931 17867
rect 10919 17836 12756 17864
rect 10919 17833 10931 17836
rect 10873 17827 10931 17833
rect 8938 17756 8944 17808
rect 8996 17796 9002 17808
rect 8996 17768 9674 17796
rect 8996 17756 9002 17768
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 9122 17728 9128 17740
rect 8352 17700 9128 17728
rect 8352 17688 8358 17700
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 9646 17672 9674 17768
rect 12728 17740 12756 17836
rect 14826 17824 14832 17876
rect 14884 17824 14890 17876
rect 16301 17867 16359 17873
rect 16301 17833 16313 17867
rect 16347 17864 16359 17867
rect 18325 17867 18383 17873
rect 16347 17836 18276 17864
rect 16347 17833 16359 17836
rect 16301 17827 16359 17833
rect 16390 17796 16396 17808
rect 16132 17768 16396 17796
rect 10318 17688 10324 17740
rect 10376 17728 10382 17740
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 10376 17700 10977 17728
rect 10376 17688 10382 17700
rect 10965 17697 10977 17700
rect 11011 17728 11023 17731
rect 12342 17728 12348 17740
rect 11011 17700 12348 17728
rect 11011 17697 11023 17700
rect 10965 17691 11023 17697
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 12710 17688 12716 17740
rect 12768 17688 12774 17740
rect 13170 17688 13176 17740
rect 13228 17688 13234 17740
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17660 8815 17663
rect 8846 17660 8852 17672
rect 8803 17632 8852 17660
rect 8803 17629 8815 17632
rect 8757 17623 8815 17629
rect 8846 17620 8852 17632
rect 8904 17620 8910 17672
rect 8938 17620 8944 17672
rect 8996 17620 9002 17672
rect 9030 17620 9036 17672
rect 9088 17660 9094 17672
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 9088 17632 9229 17660
rect 9088 17620 9094 17632
rect 9217 17629 9229 17632
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17660 9459 17663
rect 9493 17663 9551 17669
rect 9493 17660 9505 17663
rect 9447 17632 9505 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 9493 17629 9505 17632
rect 9539 17629 9551 17663
rect 9646 17632 9680 17672
rect 9493 17623 9551 17629
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 10686 17620 10692 17672
rect 10744 17620 10750 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 11057 17663 11115 17669
rect 11057 17660 11069 17663
rect 10827 17632 11069 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 11057 17629 11069 17632
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17660 11299 17663
rect 11330 17660 11336 17672
rect 11287 17632 11336 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 11422 17620 11428 17672
rect 11480 17620 11486 17672
rect 11514 17620 11520 17672
rect 11572 17620 11578 17672
rect 11606 17620 11612 17672
rect 11664 17620 11670 17672
rect 13354 17660 13360 17672
rect 11808 17632 13360 17660
rect 8864 17592 8892 17620
rect 11808 17592 11836 17632
rect 12169 17626 12205 17632
rect 13354 17620 13360 17632
rect 13412 17660 13418 17672
rect 13906 17660 13912 17672
rect 13412 17632 13912 17660
rect 13412 17620 13418 17632
rect 13906 17620 13912 17632
rect 13964 17620 13970 17672
rect 14550 17620 14556 17672
rect 14608 17620 14614 17672
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17660 14887 17663
rect 15470 17660 15476 17672
rect 14875 17632 15476 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 16132 17669 16160 17768
rect 16390 17756 16396 17768
rect 16448 17796 16454 17808
rect 16942 17796 16948 17808
rect 16448 17768 16948 17796
rect 16448 17756 16454 17768
rect 16942 17756 16948 17768
rect 17000 17756 17006 17808
rect 17678 17756 17684 17808
rect 17736 17796 17742 17808
rect 18141 17799 18199 17805
rect 18141 17796 18153 17799
rect 17736 17768 18153 17796
rect 17736 17756 17742 17768
rect 18141 17765 18153 17768
rect 18187 17765 18199 17799
rect 18248 17796 18276 17836
rect 18325 17833 18337 17867
rect 18371 17864 18383 17867
rect 19334 17864 19340 17876
rect 18371 17836 19340 17864
rect 18371 17833 18383 17836
rect 18325 17827 18383 17833
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 20349 17867 20407 17873
rect 20349 17833 20361 17867
rect 20395 17864 20407 17867
rect 20622 17864 20628 17876
rect 20395 17836 20628 17864
rect 20395 17833 20407 17836
rect 20349 17827 20407 17833
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 21361 17867 21419 17873
rect 21361 17833 21373 17867
rect 21407 17864 21419 17867
rect 22278 17864 22284 17876
rect 21407 17836 22284 17864
rect 21407 17833 21419 17836
rect 21361 17827 21419 17833
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 22554 17824 22560 17876
rect 22612 17824 22618 17876
rect 23198 17824 23204 17876
rect 23256 17864 23262 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 23256 17836 23305 17864
rect 23256 17824 23262 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23566 17864 23572 17876
rect 23293 17827 23351 17833
rect 23400 17836 23572 17864
rect 19886 17796 19892 17808
rect 18248 17768 19892 17796
rect 18141 17759 18199 17765
rect 19886 17756 19892 17768
rect 19944 17796 19950 17808
rect 21545 17799 21603 17805
rect 21545 17796 21557 17799
rect 19944 17768 20024 17796
rect 19944 17756 19950 17768
rect 19996 17737 20024 17768
rect 21192 17768 21557 17796
rect 19981 17731 20039 17737
rect 19981 17697 19993 17731
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 20180 17700 21118 17728
rect 20180 17672 20208 17700
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 16117 17663 16175 17669
rect 16117 17629 16129 17663
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 8864 17564 11836 17592
rect 11885 17595 11943 17601
rect 11885 17561 11897 17595
rect 11931 17592 11943 17595
rect 12066 17592 12072 17604
rect 11931 17564 12072 17592
rect 11931 17561 11943 17564
rect 11885 17555 11943 17561
rect 12066 17552 12072 17564
rect 12124 17552 12130 17604
rect 15856 17592 15884 17623
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16485 17663 16543 17669
rect 16485 17660 16497 17663
rect 16356 17632 16497 17660
rect 16356 17620 16362 17632
rect 16485 17629 16497 17632
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 16316 17592 16344 17620
rect 15856 17564 16344 17592
rect 8168 17496 8248 17524
rect 8168 17484 8174 17496
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 8812 17496 9045 17524
rect 8812 17484 8818 17496
rect 9033 17493 9045 17496
rect 9079 17493 9091 17527
rect 9033 17487 9091 17493
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 9585 17527 9643 17533
rect 9585 17524 9597 17527
rect 9272 17496 9597 17524
rect 9272 17484 9278 17496
rect 9585 17493 9597 17496
rect 9631 17493 9643 17527
rect 9585 17487 9643 17493
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 13078 17524 13084 17536
rect 11204 17496 13084 17524
rect 11204 17484 11210 17496
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 14642 17484 14648 17536
rect 14700 17484 14706 17536
rect 15933 17527 15991 17533
rect 15933 17493 15945 17527
rect 15979 17524 15991 17527
rect 16022 17524 16028 17536
rect 15979 17496 16028 17524
rect 15979 17493 15991 17496
rect 15933 17487 15991 17493
rect 16022 17484 16028 17496
rect 16080 17524 16086 17536
rect 16776 17524 16804 17623
rect 16942 17620 16948 17672
rect 17000 17660 17006 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 17000 17632 17325 17660
rect 17000 17620 17006 17632
rect 17313 17629 17325 17632
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 18046 17620 18052 17672
rect 18104 17620 18110 17672
rect 20162 17620 20168 17672
rect 20220 17620 20226 17672
rect 20898 17620 20904 17672
rect 20956 17620 20962 17672
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17629 21051 17663
rect 20993 17623 21051 17629
rect 17586 17552 17592 17604
rect 17644 17592 17650 17604
rect 17681 17595 17739 17601
rect 17681 17592 17693 17595
rect 17644 17564 17693 17592
rect 17644 17552 17650 17564
rect 17681 17561 17693 17564
rect 17727 17561 17739 17595
rect 17681 17555 17739 17561
rect 17865 17595 17923 17601
rect 17865 17561 17877 17595
rect 17911 17592 17923 17595
rect 18509 17595 18567 17601
rect 18509 17592 18521 17595
rect 17911 17564 18521 17592
rect 17911 17561 17923 17564
rect 17865 17555 17923 17561
rect 18509 17561 18521 17564
rect 18555 17592 18567 17595
rect 20254 17592 20260 17604
rect 18555 17564 20260 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 20254 17552 20260 17564
rect 20312 17552 20318 17604
rect 21008 17536 21036 17623
rect 21090 17592 21118 17700
rect 21192 17669 21220 17768
rect 21545 17765 21557 17768
rect 21591 17765 21603 17799
rect 23400 17796 23428 17836
rect 23566 17824 23572 17836
rect 23624 17824 23630 17876
rect 23934 17824 23940 17876
rect 23992 17864 23998 17876
rect 23992 17836 24348 17864
rect 23992 17824 23998 17836
rect 21545 17759 21603 17765
rect 22756 17768 23428 17796
rect 21284 17700 21680 17728
rect 21177 17663 21235 17669
rect 21177 17629 21189 17663
rect 21223 17629 21235 17663
rect 21177 17623 21235 17629
rect 21284 17592 21312 17700
rect 21652 17672 21680 17700
rect 21453 17663 21511 17669
rect 21453 17629 21465 17663
rect 21499 17629 21511 17663
rect 21453 17623 21511 17629
rect 21090 17564 21312 17592
rect 16080 17496 16804 17524
rect 17405 17527 17463 17533
rect 16080 17484 16086 17496
rect 17405 17493 17417 17527
rect 17451 17524 17463 17527
rect 18138 17524 18144 17536
rect 17451 17496 18144 17524
rect 17451 17493 17463 17496
rect 17405 17487 17463 17493
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 18309 17527 18367 17533
rect 18309 17493 18321 17527
rect 18355 17524 18367 17527
rect 18690 17524 18696 17536
rect 18355 17496 18696 17524
rect 18355 17493 18367 17496
rect 18309 17487 18367 17493
rect 18690 17484 18696 17496
rect 18748 17484 18754 17536
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 21468 17524 21496 17623
rect 21634 17620 21640 17672
rect 21692 17620 21698 17672
rect 22756 17669 22784 17768
rect 23474 17756 23480 17808
rect 23532 17796 23538 17808
rect 24320 17796 24348 17836
rect 24394 17824 24400 17876
rect 24452 17824 24458 17876
rect 28534 17824 28540 17876
rect 28592 17824 28598 17876
rect 28626 17824 28632 17876
rect 28684 17864 28690 17876
rect 28721 17867 28779 17873
rect 28721 17864 28733 17867
rect 28684 17836 28733 17864
rect 28684 17824 28690 17836
rect 28721 17833 28733 17836
rect 28767 17833 28779 17867
rect 28721 17827 28779 17833
rect 31478 17824 31484 17876
rect 31536 17864 31542 17876
rect 31665 17867 31723 17873
rect 31665 17864 31677 17867
rect 31536 17836 31677 17864
rect 31536 17824 31542 17836
rect 31665 17833 31677 17836
rect 31711 17833 31723 17867
rect 31665 17827 31723 17833
rect 32582 17824 32588 17876
rect 32640 17864 32646 17876
rect 33137 17867 33195 17873
rect 33137 17864 33149 17867
rect 32640 17836 33149 17864
rect 32640 17824 32646 17836
rect 33137 17833 33149 17836
rect 33183 17833 33195 17867
rect 33137 17827 33195 17833
rect 24762 17796 24768 17808
rect 23532 17768 23980 17796
rect 24320 17768 24768 17796
rect 23532 17756 23538 17768
rect 23952 17728 23980 17768
rect 24762 17756 24768 17768
rect 24820 17796 24826 17808
rect 26878 17796 26884 17808
rect 24820 17768 24992 17796
rect 24820 17756 24826 17768
rect 24964 17737 24992 17768
rect 26436 17768 26884 17796
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 23058 17700 23880 17728
rect 23952 17700 24869 17728
rect 23058 17669 23086 17700
rect 23852 17672 23880 17700
rect 24857 17697 24869 17700
rect 24903 17697 24915 17731
rect 24857 17691 24915 17697
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17697 25007 17731
rect 24949 17691 25007 17697
rect 26053 17731 26111 17737
rect 26053 17697 26065 17731
rect 26099 17728 26111 17731
rect 26436 17728 26464 17768
rect 26878 17756 26884 17768
rect 26936 17756 26942 17808
rect 28552 17796 28580 17824
rect 30006 17796 30012 17808
rect 28552 17768 30012 17796
rect 30006 17756 30012 17768
rect 30064 17796 30070 17808
rect 30650 17796 30656 17808
rect 30064 17768 30656 17796
rect 30064 17756 30070 17768
rect 30650 17756 30656 17768
rect 30708 17756 30714 17808
rect 27798 17728 27804 17740
rect 26099 17700 26464 17728
rect 26528 17700 27804 17728
rect 26099 17697 26111 17700
rect 26053 17691 26111 17697
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 22572 17632 22753 17660
rect 22572 17536 22600 17632
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 23043 17663 23101 17669
rect 23043 17629 23055 17663
rect 23089 17629 23101 17663
rect 23043 17623 23101 17629
rect 23201 17663 23259 17669
rect 23201 17629 23213 17663
rect 23247 17660 23259 17663
rect 23474 17660 23480 17672
rect 23247 17632 23480 17660
rect 23247 17629 23259 17632
rect 23201 17623 23259 17629
rect 23474 17620 23480 17632
rect 23532 17620 23538 17672
rect 23566 17620 23572 17672
rect 23624 17620 23630 17672
rect 23842 17620 23848 17672
rect 23900 17620 23906 17672
rect 24765 17663 24823 17669
rect 24765 17629 24777 17663
rect 24811 17660 24823 17663
rect 26528 17660 26556 17700
rect 27798 17688 27804 17700
rect 27856 17728 27862 17740
rect 27856 17700 28580 17728
rect 27856 17688 27862 17700
rect 24811 17632 26556 17660
rect 24811 17629 24823 17632
rect 24765 17623 24823 17629
rect 26602 17620 26608 17672
rect 26660 17660 26666 17672
rect 26881 17663 26939 17669
rect 26881 17660 26893 17663
rect 26660 17632 26893 17660
rect 26660 17620 26666 17632
rect 26881 17629 26893 17632
rect 26927 17629 26939 17663
rect 26881 17623 26939 17629
rect 27982 17620 27988 17672
rect 28040 17620 28046 17672
rect 28166 17620 28172 17672
rect 28224 17620 28230 17672
rect 28258 17620 28264 17672
rect 28316 17620 28322 17672
rect 28353 17663 28411 17669
rect 28353 17629 28365 17663
rect 28399 17660 28411 17663
rect 28442 17660 28448 17672
rect 28399 17632 28448 17660
rect 28399 17629 28411 17632
rect 28353 17623 28411 17629
rect 22833 17595 22891 17601
rect 22833 17561 22845 17595
rect 22879 17561 22891 17595
rect 22833 17555 22891 17561
rect 21048 17496 21496 17524
rect 21048 17484 21054 17496
rect 22554 17484 22560 17536
rect 22612 17484 22618 17536
rect 22848 17524 22876 17555
rect 22922 17552 22928 17604
rect 22980 17592 22986 17604
rect 23293 17595 23351 17601
rect 23293 17592 23305 17595
rect 22980 17564 23305 17592
rect 22980 17552 22986 17564
rect 23293 17561 23305 17564
rect 23339 17592 23351 17595
rect 23339 17564 23612 17592
rect 23339 17561 23351 17564
rect 23293 17555 23351 17561
rect 23474 17524 23480 17536
rect 22848 17496 23480 17524
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 23584 17524 23612 17564
rect 23658 17552 23664 17604
rect 23716 17592 23722 17604
rect 23852 17592 23880 17620
rect 23716 17564 23880 17592
rect 23937 17595 23995 17601
rect 23716 17552 23722 17564
rect 23937 17561 23949 17595
rect 23983 17592 23995 17595
rect 26145 17595 26203 17601
rect 26145 17592 26157 17595
rect 23983 17564 26157 17592
rect 23983 17561 23995 17564
rect 23937 17555 23995 17561
rect 26145 17561 26157 17564
rect 26191 17561 26203 17595
rect 26145 17555 26203 17561
rect 26237 17595 26295 17601
rect 26237 17561 26249 17595
rect 26283 17592 26295 17595
rect 27614 17592 27620 17604
rect 26283 17564 27620 17592
rect 26283 17561 26295 17564
rect 26237 17555 26295 17561
rect 27614 17552 27620 17564
rect 27672 17552 27678 17604
rect 27890 17552 27896 17604
rect 27948 17592 27954 17604
rect 28368 17592 28396 17623
rect 28442 17620 28448 17632
rect 28500 17620 28506 17672
rect 28552 17669 28580 17700
rect 31110 17688 31116 17740
rect 31168 17728 31174 17740
rect 31570 17728 31576 17740
rect 31168 17700 31576 17728
rect 31168 17688 31174 17700
rect 31570 17688 31576 17700
rect 31628 17728 31634 17740
rect 32677 17731 32735 17737
rect 32677 17728 32689 17731
rect 31628 17700 32689 17728
rect 31628 17688 31634 17700
rect 32677 17697 32689 17700
rect 32723 17728 32735 17731
rect 32723 17700 33180 17728
rect 32723 17697 32735 17700
rect 32677 17691 32735 17697
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 31846 17620 31852 17672
rect 31904 17660 31910 17672
rect 31941 17663 31999 17669
rect 31941 17660 31953 17663
rect 31904 17632 31953 17660
rect 31904 17620 31910 17632
rect 31941 17629 31953 17632
rect 31987 17629 31999 17663
rect 31941 17623 31999 17629
rect 32033 17663 32091 17669
rect 32033 17629 32045 17663
rect 32079 17629 32091 17663
rect 32033 17623 32091 17629
rect 27948 17564 28396 17592
rect 32048 17592 32076 17623
rect 32122 17620 32128 17672
rect 32180 17620 32186 17672
rect 32309 17663 32367 17669
rect 32309 17629 32321 17663
rect 32355 17660 32367 17663
rect 32355 17632 32444 17660
rect 32355 17629 32367 17632
rect 32309 17623 32367 17629
rect 32048 17564 32260 17592
rect 27948 17552 27954 17564
rect 32232 17536 32260 17564
rect 24854 17524 24860 17536
rect 23584 17496 24860 17524
rect 24854 17484 24860 17496
rect 24912 17484 24918 17536
rect 26602 17484 26608 17536
rect 26660 17484 26666 17536
rect 26694 17484 26700 17536
rect 26752 17484 26758 17536
rect 29546 17484 29552 17536
rect 29604 17524 29610 17536
rect 30926 17524 30932 17536
rect 29604 17496 30932 17524
rect 29604 17484 29610 17496
rect 30926 17484 30932 17496
rect 30984 17484 30990 17536
rect 32214 17484 32220 17536
rect 32272 17484 32278 17536
rect 32416 17533 32444 17632
rect 32490 17620 32496 17672
rect 32548 17660 32554 17672
rect 33152 17669 33180 17700
rect 32585 17663 32643 17669
rect 32585 17660 32597 17663
rect 32548 17632 32597 17660
rect 32548 17620 32554 17632
rect 32585 17629 32597 17632
rect 32631 17660 32643 17663
rect 33137 17663 33195 17669
rect 32631 17632 32720 17660
rect 32631 17629 32643 17632
rect 32585 17623 32643 17629
rect 32401 17527 32459 17533
rect 32401 17493 32413 17527
rect 32447 17493 32459 17527
rect 32692 17524 32720 17632
rect 33137 17629 33149 17663
rect 33183 17629 33195 17663
rect 33137 17623 33195 17629
rect 33229 17663 33287 17669
rect 33229 17629 33241 17663
rect 33275 17629 33287 17663
rect 33229 17623 33287 17629
rect 32766 17552 32772 17604
rect 32824 17592 32830 17604
rect 33045 17595 33103 17601
rect 33045 17592 33057 17595
rect 32824 17564 33057 17592
rect 32824 17552 32830 17564
rect 33045 17561 33057 17564
rect 33091 17561 33103 17595
rect 33045 17555 33103 17561
rect 33244 17524 33272 17623
rect 32692 17496 33272 17524
rect 32401 17487 32459 17493
rect 33502 17484 33508 17536
rect 33560 17484 33566 17536
rect 1104 17434 34840 17456
rect 1104 17382 9344 17434
rect 9396 17382 9408 17434
rect 9460 17382 9472 17434
rect 9524 17382 9536 17434
rect 9588 17382 9600 17434
rect 9652 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 17930 17434
rect 17982 17382 17994 17434
rect 18046 17382 26132 17434
rect 26184 17382 26196 17434
rect 26248 17382 26260 17434
rect 26312 17382 26324 17434
rect 26376 17382 26388 17434
rect 26440 17382 34526 17434
rect 34578 17382 34590 17434
rect 34642 17382 34654 17434
rect 34706 17382 34718 17434
rect 34770 17382 34782 17434
rect 34834 17382 34840 17434
rect 1104 17360 34840 17382
rect 3418 17280 3424 17332
rect 3476 17280 3482 17332
rect 3602 17280 3608 17332
rect 3660 17320 3666 17332
rect 4246 17320 4252 17332
rect 3660 17292 4252 17320
rect 3660 17280 3666 17292
rect 4246 17280 4252 17292
rect 4304 17320 4310 17332
rect 7837 17323 7895 17329
rect 4304 17292 6500 17320
rect 4304 17280 4310 17292
rect 2958 17184 2964 17196
rect 2806 17156 2964 17184
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 3436 17193 3464 17280
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 3510 17144 3516 17196
rect 3568 17144 3574 17196
rect 3602 17144 3608 17196
rect 3660 17144 3666 17196
rect 3694 17144 3700 17196
rect 3752 17193 3758 17196
rect 5000 17193 5028 17292
rect 5074 17212 5080 17264
rect 5132 17252 5138 17264
rect 5132 17224 5212 17252
rect 5132 17212 5138 17224
rect 5184 17193 5212 17224
rect 3752 17187 3801 17193
rect 3752 17153 3755 17187
rect 3789 17153 3801 17187
rect 3752 17147 3801 17153
rect 4985 17187 5043 17193
rect 4985 17153 4997 17187
rect 5031 17153 5043 17187
rect 4985 17147 5043 17153
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 5261 17190 5319 17193
rect 5261 17187 5396 17190
rect 5261 17153 5273 17187
rect 5307 17184 5396 17187
rect 5718 17184 5724 17196
rect 5307 17162 5724 17184
rect 5307 17153 5319 17162
rect 5368 17156 5724 17162
rect 5261 17147 5319 17153
rect 3752 17146 3766 17147
rect 3752 17144 3758 17146
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 1394 17076 1400 17128
rect 1452 17076 1458 17128
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 3237 17119 3295 17125
rect 3237 17116 3249 17119
rect 1719 17088 3249 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 3237 17085 3249 17088
rect 3283 17085 3295 17119
rect 3237 17079 3295 17085
rect 3878 17076 3884 17128
rect 3936 17076 3942 17128
rect 4798 17076 4804 17128
rect 4856 17076 4862 17128
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17085 5135 17119
rect 5077 17079 5135 17085
rect 4816 17048 4844 17076
rect 5092 17048 5120 17079
rect 4816 17020 5120 17048
rect 3142 16940 3148 16992
rect 3200 16940 3206 16992
rect 4982 16940 4988 16992
rect 5040 16980 5046 16992
rect 5445 16983 5503 16989
rect 5445 16980 5457 16983
rect 5040 16952 5457 16980
rect 5040 16940 5046 16952
rect 5445 16949 5457 16952
rect 5491 16949 5503 16983
rect 6472 16980 6500 17292
rect 7837 17289 7849 17323
rect 7883 17320 7895 17323
rect 9030 17320 9036 17332
rect 7883 17292 9036 17320
rect 7883 17289 7895 17292
rect 7837 17283 7895 17289
rect 9030 17280 9036 17292
rect 9088 17280 9094 17332
rect 9232 17292 11192 17320
rect 7576 17224 8340 17252
rect 7374 17144 7380 17196
rect 7432 17144 7438 17196
rect 7576 17193 7604 17224
rect 8312 17196 8340 17224
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7650 17144 7656 17196
rect 7708 17144 7714 17196
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7800 17156 8033 17184
rect 7800 17144 7806 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8294 17144 8300 17196
rect 8352 17144 8358 17196
rect 9232 17193 9260 17292
rect 9674 17252 9680 17264
rect 9508 17224 9680 17252
rect 9508 17193 9536 17224
rect 9674 17212 9680 17224
rect 9732 17212 9738 17264
rect 9766 17212 9772 17264
rect 9824 17252 9830 17264
rect 9824 17224 11100 17252
rect 9824 17212 9830 17224
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17116 7527 17119
rect 7760 17116 7788 17144
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 7515 17088 7788 17116
rect 7852 17088 8125 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 7650 17008 7656 17060
rect 7708 17048 7714 17060
rect 7852 17048 7880 17088
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 9232 17116 9260 17147
rect 8113 17079 8171 17085
rect 8220 17088 9260 17116
rect 8220 17048 8248 17088
rect 7708 17020 7880 17048
rect 7944 17020 8248 17048
rect 7708 17008 7714 17020
rect 7742 16980 7748 16992
rect 6472 16952 7748 16980
rect 5445 16943 5503 16949
rect 7742 16940 7748 16952
rect 7800 16980 7806 16992
rect 7944 16980 7972 17020
rect 8478 17008 8484 17060
rect 8536 17048 8542 17060
rect 9600 17048 9628 17147
rect 8536 17020 9628 17048
rect 9692 17048 9720 17212
rect 11072 17193 11100 17224
rect 11164 17193 11192 17292
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 12154 17323 12212 17329
rect 12154 17320 12166 17323
rect 11572 17292 12166 17320
rect 11572 17280 11578 17292
rect 12154 17289 12166 17292
rect 12200 17289 12212 17323
rect 12154 17283 12212 17289
rect 11238 17212 11244 17264
rect 11296 17252 11302 17264
rect 12069 17255 12127 17261
rect 12069 17252 12081 17255
rect 11296 17224 12081 17252
rect 11296 17212 11302 17224
rect 12069 17221 12081 17224
rect 12115 17221 12127 17255
rect 12169 17252 12197 17283
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 13541 17323 13599 17329
rect 12492 17292 12756 17320
rect 12492 17280 12498 17292
rect 12169 17224 12664 17252
rect 12069 17215 12127 17221
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 9784 17156 10885 17184
rect 9784 17128 9812 17156
rect 10873 17153 10885 17156
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 11057 17187 11115 17193
rect 11057 17153 11069 17187
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17153 11207 17187
rect 11606 17184 11612 17196
rect 11149 17147 11207 17153
rect 11348 17156 11612 17184
rect 9766 17076 9772 17128
rect 9824 17076 9830 17128
rect 10888 17048 10916 17147
rect 11072 17116 11100 17147
rect 11348 17116 11376 17156
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 11882 17144 11888 17196
rect 11940 17144 11946 17196
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 11072 17088 11376 17116
rect 11333 17051 11391 17057
rect 9692 17020 10456 17048
rect 10888 17020 11008 17048
rect 8536 17008 8542 17020
rect 10428 16992 10456 17020
rect 7800 16952 7972 16980
rect 8205 16983 8263 16989
rect 7800 16940 7806 16952
rect 8205 16949 8217 16983
rect 8251 16980 8263 16983
rect 8294 16980 8300 16992
rect 8251 16952 8300 16980
rect 8251 16949 8263 16952
rect 8205 16943 8263 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 8389 16983 8447 16989
rect 8389 16949 8401 16983
rect 8435 16980 8447 16983
rect 9122 16980 9128 16992
rect 8435 16952 9128 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 9214 16940 9220 16992
rect 9272 16980 9278 16992
rect 9309 16983 9367 16989
rect 9309 16980 9321 16983
rect 9272 16952 9321 16980
rect 9272 16940 9278 16952
rect 9309 16949 9321 16952
rect 9355 16949 9367 16983
rect 9309 16943 9367 16949
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 9732 16952 9781 16980
rect 9732 16940 9738 16952
rect 9769 16949 9781 16952
rect 9815 16949 9827 16983
rect 9769 16943 9827 16949
rect 10410 16940 10416 16992
rect 10468 16940 10474 16992
rect 10870 16940 10876 16992
rect 10928 16940 10934 16992
rect 10980 16980 11008 17020
rect 11333 17017 11345 17051
rect 11379 17048 11391 17051
rect 11992 17048 12020 17147
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 12636 17193 12664 17224
rect 12728 17193 12756 17292
rect 13541 17289 13553 17323
rect 13587 17320 13599 17323
rect 14642 17320 14648 17332
rect 13587 17292 14648 17320
rect 13587 17289 13599 17292
rect 13541 17283 13599 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 17957 17323 18015 17329
rect 17957 17320 17969 17323
rect 17552 17292 17969 17320
rect 17552 17280 17558 17292
rect 17957 17289 17969 17292
rect 18003 17289 18015 17323
rect 17957 17283 18015 17289
rect 18138 17280 18144 17332
rect 18196 17320 18202 17332
rect 18196 17292 18828 17320
rect 18196 17280 18202 17292
rect 18800 17264 18828 17292
rect 27982 17280 27988 17332
rect 28040 17320 28046 17332
rect 28261 17323 28319 17329
rect 28261 17320 28273 17323
rect 28040 17292 28273 17320
rect 28040 17280 28046 17292
rect 28261 17289 28273 17292
rect 28307 17289 28319 17323
rect 28994 17320 29000 17332
rect 28261 17283 28319 17289
rect 28460 17292 29000 17320
rect 12897 17255 12955 17261
rect 12897 17221 12909 17255
rect 12943 17252 12955 17255
rect 12943 17224 13952 17252
rect 12943 17221 12955 17224
rect 12897 17215 12955 17221
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12400 17156 12449 17184
rect 12400 17144 12406 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 12713 17187 12771 17193
rect 12713 17153 12725 17187
rect 12759 17153 12771 17187
rect 12713 17147 12771 17153
rect 11379 17020 12020 17048
rect 11379 17017 11391 17020
rect 11333 17011 11391 17017
rect 11606 16980 11612 16992
rect 10980 16952 11612 16980
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 11793 16983 11851 16989
rect 11793 16949 11805 16983
rect 11839 16980 11851 16983
rect 11974 16980 11980 16992
rect 11839 16952 11980 16980
rect 11839 16949 11851 16952
rect 11793 16943 11851 16949
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12452 16980 12480 17147
rect 12986 17144 12992 17196
rect 13044 17144 13050 17196
rect 13078 17144 13084 17196
rect 13136 17144 13142 17196
rect 13262 17144 13268 17196
rect 13320 17144 13326 17196
rect 13446 17144 13452 17196
rect 13504 17144 13510 17196
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 13924 17193 13952 17224
rect 17586 17212 17592 17264
rect 17644 17252 17650 17264
rect 18417 17255 18475 17261
rect 18417 17252 18429 17255
rect 17644 17224 17724 17252
rect 17644 17212 17650 17224
rect 13633 17187 13691 17193
rect 13633 17184 13645 17187
rect 13596 17156 13645 17184
rect 13596 17144 13602 17156
rect 13633 17153 13645 17156
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 13817 17187 13875 17193
rect 13817 17153 13829 17187
rect 13863 17153 13875 17187
rect 13817 17147 13875 17153
rect 13909 17187 13967 17193
rect 13909 17153 13921 17187
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 13004 17116 13032 17144
rect 13173 17119 13231 17125
rect 13173 17116 13185 17119
rect 13004 17088 13185 17116
rect 13173 17085 13185 17088
rect 13219 17085 13231 17119
rect 13173 17079 13231 17085
rect 13357 17119 13415 17125
rect 13357 17085 13369 17119
rect 13403 17085 13415 17119
rect 13357 17079 13415 17085
rect 12526 17008 12532 17060
rect 12584 17008 12590 17060
rect 12710 17008 12716 17060
rect 12768 17048 12774 17060
rect 13372 17048 13400 17079
rect 12768 17020 13400 17048
rect 13464 17048 13492 17144
rect 13633 17051 13691 17057
rect 13633 17048 13645 17051
rect 13464 17020 13645 17048
rect 12768 17008 12774 17020
rect 13633 17017 13645 17020
rect 13679 17017 13691 17051
rect 13832 17048 13860 17147
rect 14918 17144 14924 17196
rect 14976 17144 14982 17196
rect 17696 17193 17724 17224
rect 17788 17224 18429 17252
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 15304 17156 15577 17184
rect 15194 17076 15200 17128
rect 15252 17076 15258 17128
rect 13906 17048 13912 17060
rect 13832 17020 13912 17048
rect 13633 17011 13691 17017
rect 13906 17008 13912 17020
rect 13964 17008 13970 17060
rect 15304 16992 15332 17156
rect 15565 17153 15577 17156
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 17405 17187 17463 17193
rect 17405 17153 17417 17187
rect 17451 17153 17463 17187
rect 17405 17147 17463 17153
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 17221 17119 17279 17125
rect 17221 17085 17233 17119
rect 17267 17085 17279 17119
rect 17420 17116 17448 17147
rect 17788 17116 17816 17224
rect 18417 17221 18429 17224
rect 18463 17252 18475 17255
rect 18463 17224 18736 17252
rect 18463 17221 18475 17224
rect 18417 17215 18475 17221
rect 18708 17196 18736 17224
rect 18782 17212 18788 17264
rect 18840 17212 18846 17264
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17184 18107 17187
rect 18506 17184 18512 17196
rect 18095 17156 18512 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 17420 17088 17816 17116
rect 18166 17119 18224 17125
rect 17221 17079 17279 17085
rect 18166 17085 18178 17119
rect 18212 17116 18224 17119
rect 18322 17116 18328 17128
rect 18212 17088 18328 17116
rect 18212 17085 18224 17088
rect 18166 17079 18224 17085
rect 17236 17048 17264 17079
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 18616 17116 18644 17147
rect 18690 17144 18696 17196
rect 18748 17144 18754 17196
rect 18800 17184 18828 17212
rect 20990 17184 20996 17196
rect 18800 17156 20996 17184
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17184 21235 17187
rect 21634 17184 21640 17196
rect 21223 17156 21640 17184
rect 21223 17153 21235 17156
rect 21177 17147 21235 17153
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 28460 17193 28488 17292
rect 28994 17280 29000 17292
rect 29052 17280 29058 17332
rect 31573 17323 31631 17329
rect 29656 17292 30144 17320
rect 29546 17252 29552 17264
rect 28736 17224 29552 17252
rect 28736 17193 28764 17224
rect 29546 17212 29552 17224
rect 29604 17212 29610 17264
rect 28445 17187 28503 17193
rect 28445 17153 28457 17187
rect 28491 17153 28503 17187
rect 28445 17147 28503 17153
rect 28537 17187 28595 17193
rect 28537 17153 28549 17187
rect 28583 17153 28595 17187
rect 28537 17147 28595 17153
rect 28721 17187 28779 17193
rect 28721 17153 28733 17187
rect 28767 17153 28779 17187
rect 28721 17147 28779 17153
rect 19334 17116 19340 17128
rect 18616 17088 19340 17116
rect 18616 17048 18644 17088
rect 19334 17076 19340 17088
rect 19392 17116 19398 17128
rect 19978 17116 19984 17128
rect 19392 17088 19984 17116
rect 19392 17076 19398 17088
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 21008 17116 21036 17144
rect 22278 17116 22284 17128
rect 21008 17088 22284 17116
rect 22278 17076 22284 17088
rect 22336 17076 22342 17128
rect 28552 17116 28580 17147
rect 28810 17144 28816 17196
rect 28868 17144 28874 17196
rect 28902 17144 28908 17196
rect 28960 17144 28966 17196
rect 29270 17144 29276 17196
rect 29328 17184 29334 17196
rect 29656 17184 29684 17292
rect 29733 17187 29791 17193
rect 29733 17184 29745 17187
rect 29328 17156 29745 17184
rect 29328 17144 29334 17156
rect 29733 17153 29745 17156
rect 29779 17153 29791 17187
rect 29917 17187 29975 17193
rect 29917 17184 29929 17187
rect 29733 17147 29791 17153
rect 29840 17156 29929 17184
rect 28920 17116 28948 17144
rect 28552 17088 28948 17116
rect 29840 17116 29868 17156
rect 29917 17153 29929 17156
rect 29963 17153 29975 17187
rect 30116 17184 30144 17292
rect 31573 17289 31585 17323
rect 31619 17320 31631 17323
rect 31662 17320 31668 17332
rect 31619 17292 31668 17320
rect 31619 17289 31631 17292
rect 31573 17283 31631 17289
rect 31662 17280 31668 17292
rect 31720 17280 31726 17332
rect 32674 17280 32680 17332
rect 32732 17320 32738 17332
rect 32861 17323 32919 17329
rect 32861 17320 32873 17323
rect 32732 17292 32873 17320
rect 32732 17280 32738 17292
rect 32861 17289 32873 17292
rect 32907 17289 32919 17323
rect 32861 17283 32919 17289
rect 33410 17280 33416 17332
rect 33468 17320 33474 17332
rect 33468 17292 33916 17320
rect 33468 17280 33474 17292
rect 30926 17212 30932 17264
rect 30984 17252 30990 17264
rect 33781 17255 33839 17261
rect 33781 17252 33793 17255
rect 30984 17224 33793 17252
rect 30984 17212 30990 17224
rect 33781 17221 33793 17224
rect 33827 17221 33839 17255
rect 33781 17215 33839 17221
rect 30193 17187 30251 17193
rect 30193 17184 30205 17187
rect 30116 17156 30205 17184
rect 29917 17147 29975 17153
rect 30193 17153 30205 17156
rect 30239 17153 30251 17187
rect 30193 17147 30251 17153
rect 30377 17187 30435 17193
rect 30377 17153 30389 17187
rect 30423 17153 30435 17187
rect 31018 17184 31024 17196
rect 30377 17147 30435 17153
rect 30944 17156 31024 17184
rect 30392 17116 30420 17147
rect 29840 17088 30420 17116
rect 30944 17116 30972 17156
rect 31018 17144 31024 17156
rect 31076 17144 31082 17196
rect 31110 17144 31116 17196
rect 31168 17144 31174 17196
rect 31202 17144 31208 17196
rect 31260 17184 31266 17196
rect 31297 17187 31355 17193
rect 31297 17184 31309 17187
rect 31260 17156 31309 17184
rect 31260 17144 31266 17156
rect 31297 17153 31309 17156
rect 31343 17153 31355 17187
rect 31297 17147 31355 17153
rect 31389 17187 31447 17193
rect 31389 17153 31401 17187
rect 31435 17184 31447 17187
rect 31570 17184 31576 17196
rect 31435 17156 31576 17184
rect 31435 17153 31447 17156
rect 31389 17147 31447 17153
rect 31570 17144 31576 17156
rect 31628 17144 31634 17196
rect 32677 17187 32735 17193
rect 32677 17153 32689 17187
rect 32723 17184 32735 17187
rect 32766 17184 32772 17196
rect 32723 17156 32772 17184
rect 32723 17153 32735 17156
rect 32677 17147 32735 17153
rect 32692 17116 32720 17147
rect 32766 17144 32772 17156
rect 32824 17144 32830 17196
rect 32950 17144 32956 17196
rect 33008 17144 33014 17196
rect 33134 17144 33140 17196
rect 33192 17144 33198 17196
rect 33686 17144 33692 17196
rect 33744 17144 33750 17196
rect 33888 17193 33916 17292
rect 33873 17187 33931 17193
rect 33873 17153 33885 17187
rect 33919 17153 33931 17187
rect 33873 17147 33931 17153
rect 30944 17088 32720 17116
rect 17236 17020 18644 17048
rect 27614 17008 27620 17060
rect 27672 17048 27678 17060
rect 29840 17048 29868 17088
rect 27672 17020 29868 17048
rect 30101 17051 30159 17057
rect 27672 17008 27678 17020
rect 30101 17017 30113 17051
rect 30147 17048 30159 17051
rect 30926 17048 30932 17060
rect 30147 17020 30932 17048
rect 30147 17017 30159 17020
rect 30101 17011 30159 17017
rect 30926 17008 30932 17020
rect 30984 17008 30990 17060
rect 14182 16980 14188 16992
rect 12452 16952 14188 16980
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 15286 16940 15292 16992
rect 15344 16940 15350 16992
rect 15470 16940 15476 16992
rect 15528 16940 15534 16992
rect 15654 16940 15660 16992
rect 15712 16940 15718 16992
rect 18138 16940 18144 16992
rect 18196 16980 18202 16992
rect 18325 16983 18383 16989
rect 18325 16980 18337 16983
rect 18196 16952 18337 16980
rect 18196 16940 18202 16952
rect 18325 16949 18337 16952
rect 18371 16949 18383 16983
rect 18325 16943 18383 16949
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 18785 16983 18843 16989
rect 18785 16980 18797 16983
rect 18472 16952 18797 16980
rect 18472 16940 18478 16952
rect 18785 16949 18797 16952
rect 18831 16949 18843 16983
rect 18785 16943 18843 16949
rect 21174 16940 21180 16992
rect 21232 16940 21238 16992
rect 30285 16983 30343 16989
rect 30285 16949 30297 16983
rect 30331 16980 30343 16983
rect 30650 16980 30656 16992
rect 30331 16952 30656 16980
rect 30331 16949 30343 16952
rect 30285 16943 30343 16949
rect 30650 16940 30656 16952
rect 30708 16940 30714 16992
rect 1104 16890 34684 16912
rect 1104 16838 5147 16890
rect 5199 16838 5211 16890
rect 5263 16838 5275 16890
rect 5327 16838 5339 16890
rect 5391 16838 5403 16890
rect 5455 16838 13541 16890
rect 13593 16838 13605 16890
rect 13657 16838 13669 16890
rect 13721 16838 13733 16890
rect 13785 16838 13797 16890
rect 13849 16838 21935 16890
rect 21987 16838 21999 16890
rect 22051 16838 22063 16890
rect 22115 16838 22127 16890
rect 22179 16838 22191 16890
rect 22243 16838 30329 16890
rect 30381 16838 30393 16890
rect 30445 16838 30457 16890
rect 30509 16838 30521 16890
rect 30573 16838 30585 16890
rect 30637 16838 34684 16890
rect 1104 16816 34684 16838
rect 3970 16736 3976 16788
rect 4028 16776 4034 16788
rect 5626 16785 5632 16788
rect 5610 16779 5632 16785
rect 5610 16776 5622 16779
rect 4028 16748 5622 16776
rect 4028 16736 4034 16748
rect 5610 16745 5622 16748
rect 5610 16739 5632 16745
rect 5626 16736 5632 16739
rect 5684 16736 5690 16788
rect 5810 16736 5816 16788
rect 5868 16776 5874 16788
rect 5905 16779 5963 16785
rect 5905 16776 5917 16779
rect 5868 16748 5917 16776
rect 5868 16736 5874 16748
rect 5905 16745 5917 16748
rect 5951 16745 5963 16779
rect 5905 16739 5963 16745
rect 6917 16779 6975 16785
rect 6917 16745 6929 16779
rect 6963 16776 6975 16779
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 6963 16748 7481 16776
rect 6963 16745 6975 16748
rect 6917 16739 6975 16745
rect 7469 16745 7481 16748
rect 7515 16745 7527 16779
rect 7469 16739 7527 16745
rect 5721 16711 5779 16717
rect 5721 16708 5733 16711
rect 3896 16680 5733 16708
rect 3142 16532 3148 16584
rect 3200 16572 3206 16584
rect 3329 16575 3387 16581
rect 3329 16572 3341 16575
rect 3200 16544 3341 16572
rect 3200 16532 3206 16544
rect 3329 16541 3341 16544
rect 3375 16541 3387 16575
rect 3329 16535 3387 16541
rect 3896 16516 3924 16680
rect 5721 16677 5733 16680
rect 5767 16677 5779 16711
rect 5721 16671 5779 16677
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 5813 16643 5871 16649
rect 5813 16640 5825 16643
rect 4120 16612 5825 16640
rect 4120 16600 4126 16612
rect 5813 16609 5825 16612
rect 5859 16609 5871 16643
rect 5920 16640 5948 16739
rect 7834 16736 7840 16788
rect 7892 16776 7898 16788
rect 9766 16776 9772 16788
rect 7892 16748 9772 16776
rect 7892 16736 7898 16748
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 9876 16748 13553 16776
rect 6733 16711 6791 16717
rect 6733 16677 6745 16711
rect 6779 16708 6791 16711
rect 7377 16711 7435 16717
rect 6779 16680 7052 16708
rect 6779 16677 6791 16680
rect 6733 16671 6791 16677
rect 7024 16640 7052 16680
rect 7377 16677 7389 16711
rect 7423 16708 7435 16711
rect 9876 16708 9904 16748
rect 13541 16745 13553 16748
rect 13587 16745 13599 16779
rect 13541 16739 13599 16745
rect 13906 16736 13912 16788
rect 13964 16736 13970 16788
rect 15102 16736 15108 16788
rect 15160 16736 15166 16788
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 15378 16776 15384 16788
rect 15335 16748 15384 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 15378 16736 15384 16748
rect 15436 16776 15442 16788
rect 15746 16776 15752 16788
rect 15436 16748 15752 16776
rect 15436 16736 15442 16748
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16022 16736 16028 16788
rect 16080 16776 16086 16788
rect 16117 16779 16175 16785
rect 16117 16776 16129 16779
rect 16080 16748 16129 16776
rect 16080 16736 16086 16748
rect 16117 16745 16129 16748
rect 16163 16745 16175 16779
rect 16117 16739 16175 16745
rect 21174 16736 21180 16788
rect 21232 16776 21238 16788
rect 21453 16779 21511 16785
rect 21453 16776 21465 16779
rect 21232 16748 21465 16776
rect 21232 16736 21238 16748
rect 21453 16745 21465 16748
rect 21499 16745 21511 16779
rect 21453 16739 21511 16745
rect 21821 16779 21879 16785
rect 21821 16745 21833 16779
rect 21867 16776 21879 16779
rect 22738 16776 22744 16788
rect 21867 16748 22744 16776
rect 21867 16745 21879 16748
rect 21821 16739 21879 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 22925 16779 22983 16785
rect 22925 16745 22937 16779
rect 22971 16776 22983 16779
rect 23658 16776 23664 16788
rect 22971 16748 23664 16776
rect 22971 16745 22983 16748
rect 22925 16739 22983 16745
rect 23658 16736 23664 16748
rect 23716 16736 23722 16788
rect 24762 16736 24768 16788
rect 24820 16736 24826 16788
rect 26132 16779 26190 16785
rect 26132 16745 26144 16779
rect 26178 16776 26190 16779
rect 26694 16776 26700 16788
rect 26178 16748 26700 16776
rect 26178 16745 26190 16748
rect 26132 16739 26190 16745
rect 26694 16736 26700 16748
rect 26752 16736 26758 16788
rect 27614 16736 27620 16788
rect 27672 16736 27678 16788
rect 29270 16736 29276 16788
rect 29328 16736 29334 16788
rect 30745 16779 30803 16785
rect 30745 16745 30757 16779
rect 30791 16776 30803 16779
rect 31018 16776 31024 16788
rect 30791 16748 31024 16776
rect 30791 16745 30803 16748
rect 30745 16739 30803 16745
rect 31018 16736 31024 16748
rect 31076 16736 31082 16788
rect 31113 16779 31171 16785
rect 31113 16745 31125 16779
rect 31159 16776 31171 16779
rect 31202 16776 31208 16788
rect 31159 16748 31208 16776
rect 31159 16745 31171 16748
rect 31113 16739 31171 16745
rect 31202 16736 31208 16748
rect 31260 16736 31266 16788
rect 31294 16736 31300 16788
rect 31352 16736 31358 16788
rect 31665 16779 31723 16785
rect 31665 16745 31677 16779
rect 31711 16776 31723 16779
rect 32401 16779 32459 16785
rect 32401 16776 32413 16779
rect 31711 16748 32413 16776
rect 31711 16745 31723 16748
rect 31665 16739 31723 16745
rect 32401 16745 32413 16748
rect 32447 16776 32459 16779
rect 33134 16776 33140 16788
rect 32447 16748 33140 16776
rect 32447 16745 32459 16748
rect 32401 16739 32459 16745
rect 33134 16736 33140 16748
rect 33192 16736 33198 16788
rect 33502 16736 33508 16788
rect 33560 16736 33566 16788
rect 33686 16736 33692 16788
rect 33744 16776 33750 16788
rect 33781 16779 33839 16785
rect 33781 16776 33793 16779
rect 33744 16748 33793 16776
rect 33744 16736 33750 16748
rect 33781 16745 33793 16748
rect 33827 16745 33839 16779
rect 33781 16739 33839 16745
rect 7423 16680 9904 16708
rect 7423 16677 7435 16680
rect 7377 16671 7435 16677
rect 10870 16668 10876 16720
rect 10928 16708 10934 16720
rect 11882 16708 11888 16720
rect 10928 16680 11888 16708
rect 10928 16668 10934 16680
rect 11882 16668 11888 16680
rect 11940 16668 11946 16720
rect 15120 16708 15148 16736
rect 12452 16680 13860 16708
rect 15120 16680 15884 16708
rect 12452 16652 12480 16680
rect 8113 16643 8171 16649
rect 8113 16640 8125 16643
rect 5920 16612 6776 16640
rect 7024 16612 7144 16640
rect 5813 16603 5871 16609
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16572 5503 16575
rect 5534 16572 5540 16584
rect 5491 16544 5540 16572
rect 5491 16541 5503 16544
rect 5445 16535 5503 16541
rect 5534 16532 5540 16544
rect 5592 16572 5598 16584
rect 5994 16572 6000 16584
rect 5592 16544 6000 16572
rect 5592 16532 5598 16544
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 6270 16532 6276 16584
rect 6328 16572 6334 16584
rect 6748 16581 6776 16612
rect 6549 16575 6607 16581
rect 6549 16572 6561 16575
rect 6328 16544 6561 16572
rect 6328 16532 6334 16544
rect 6549 16541 6561 16544
rect 6595 16541 6607 16575
rect 6549 16535 6607 16541
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16541 6791 16575
rect 6733 16535 6791 16541
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 3878 16504 3884 16516
rect 3108 16476 3884 16504
rect 3108 16464 3114 16476
rect 3878 16464 3884 16476
rect 3936 16464 3942 16516
rect 6362 16396 6368 16448
rect 6420 16396 6426 16448
rect 6748 16436 6776 16535
rect 6822 16532 6828 16584
rect 6880 16532 6886 16584
rect 7116 16581 7144 16612
rect 7208 16612 8125 16640
rect 7208 16581 7236 16612
rect 8113 16609 8125 16612
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 8662 16640 8668 16652
rect 8619 16612 8668 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 12434 16600 12440 16652
rect 12492 16600 12498 16652
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16640 12679 16643
rect 13538 16640 13544 16652
rect 12667 16612 13544 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 13832 16649 13860 16680
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16609 13875 16643
rect 13817 16603 13875 16609
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15286 16640 15292 16652
rect 15151 16612 15292 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15856 16640 15884 16680
rect 20162 16668 20168 16720
rect 20220 16668 20226 16720
rect 24780 16708 24808 16736
rect 33520 16708 33548 16736
rect 24780 16680 24992 16708
rect 15856 16612 15976 16640
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16541 7251 16575
rect 7193 16535 7251 16541
rect 7374 16532 7380 16584
rect 7432 16572 7438 16584
rect 7650 16572 7656 16584
rect 7432 16544 7656 16572
rect 7432 16532 7438 16544
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 7742 16532 7748 16584
rect 7800 16532 7806 16584
rect 7834 16532 7840 16584
rect 7892 16532 7898 16584
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 8297 16575 8355 16581
rect 8297 16572 8309 16575
rect 7929 16535 7987 16541
rect 8220 16544 8309 16572
rect 7558 16464 7564 16516
rect 7616 16504 7622 16516
rect 7944 16504 7972 16535
rect 8220 16504 8248 16544
rect 8297 16541 8309 16544
rect 8343 16541 8355 16575
rect 8297 16535 8355 16541
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16572 8539 16575
rect 8527 16544 8708 16572
rect 8527 16541 8539 16544
rect 8481 16535 8539 16541
rect 7616 16476 7972 16504
rect 8129 16476 8248 16504
rect 7616 16464 7622 16476
rect 8129 16436 8157 16476
rect 6748 16408 8157 16436
rect 8680 16436 8708 16544
rect 9398 16532 9404 16584
rect 9456 16572 9462 16584
rect 9493 16575 9551 16581
rect 9493 16572 9505 16575
rect 9456 16544 9505 16572
rect 9456 16532 9462 16544
rect 9493 16541 9505 16544
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 9585 16575 9643 16581
rect 9585 16541 9597 16575
rect 9631 16572 9643 16575
rect 9674 16572 9680 16584
rect 9631 16544 9680 16572
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 9769 16575 9827 16581
rect 9769 16541 9781 16575
rect 9815 16572 9827 16575
rect 11238 16572 11244 16584
rect 9815 16544 11244 16572
rect 9815 16541 9827 16544
rect 9769 16535 9827 16541
rect 9306 16464 9312 16516
rect 9364 16504 9370 16516
rect 9784 16504 9812 16535
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 13449 16575 13507 16581
rect 13449 16572 13461 16575
rect 12308 16544 13461 16572
rect 12308 16532 12314 16544
rect 13449 16541 13461 16544
rect 13495 16541 13507 16575
rect 13449 16535 13507 16541
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16541 13783 16575
rect 13725 16535 13783 16541
rect 9364 16476 9812 16504
rect 9364 16464 9370 16476
rect 13354 16464 13360 16516
rect 13412 16464 13418 16516
rect 9766 16436 9772 16448
rect 8680 16408 9772 16436
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 9953 16439 10011 16445
rect 9953 16405 9965 16439
rect 9999 16436 10011 16439
rect 10686 16436 10692 16448
rect 9999 16408 10692 16436
rect 9999 16405 10011 16408
rect 9953 16399 10011 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 13464 16436 13492 16535
rect 13538 16464 13544 16516
rect 13596 16504 13602 16516
rect 13740 16504 13768 16535
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 15010 16572 15016 16584
rect 14424 16544 15016 16572
rect 14424 16532 14430 16544
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 15194 16532 15200 16584
rect 15252 16532 15258 16584
rect 15381 16575 15439 16581
rect 15381 16541 15393 16575
rect 15427 16572 15439 16575
rect 15470 16572 15476 16584
rect 15427 16544 15476 16572
rect 15427 16541 15439 16544
rect 15381 16535 15439 16541
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16572 15807 16575
rect 15838 16572 15844 16584
rect 15795 16544 15844 16572
rect 15795 16541 15807 16544
rect 15749 16535 15807 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 15948 16581 15976 16612
rect 19886 16600 19892 16652
rect 19944 16640 19950 16652
rect 20180 16640 20208 16668
rect 19944 16612 20024 16640
rect 19944 16600 19950 16612
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16541 15991 16575
rect 15933 16535 15991 16541
rect 16114 16532 16120 16584
rect 16172 16532 16178 16584
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16572 18107 16575
rect 18138 16572 18144 16584
rect 18095 16544 18144 16572
rect 18095 16541 18107 16544
rect 18049 16535 18107 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18230 16532 18236 16584
rect 18288 16532 18294 16584
rect 19996 16581 20024 16612
rect 20134 16612 20208 16640
rect 20349 16643 20407 16649
rect 20134 16581 20162 16612
rect 20349 16609 20361 16643
rect 20395 16640 20407 16643
rect 21361 16643 21419 16649
rect 21361 16640 21373 16643
rect 20395 16612 21373 16640
rect 20395 16609 20407 16612
rect 20349 16603 20407 16609
rect 21361 16609 21373 16612
rect 21407 16640 21419 16643
rect 22557 16643 22615 16649
rect 22557 16640 22569 16643
rect 21407 16612 22569 16640
rect 21407 16609 21419 16612
rect 21361 16603 21419 16609
rect 22557 16609 22569 16612
rect 22603 16609 22615 16643
rect 22557 16603 22615 16609
rect 24854 16600 24860 16652
rect 24912 16600 24918 16652
rect 24964 16649 24992 16680
rect 30668 16680 31754 16708
rect 30668 16652 30696 16680
rect 24949 16643 25007 16649
rect 24949 16609 24961 16643
rect 24995 16609 25007 16643
rect 24949 16603 25007 16609
rect 25869 16643 25927 16649
rect 25869 16609 25881 16643
rect 25915 16640 25927 16643
rect 26878 16640 26884 16652
rect 25915 16612 26884 16640
rect 25915 16609 25927 16612
rect 25869 16603 25927 16609
rect 26878 16600 26884 16612
rect 26936 16600 26942 16652
rect 30561 16643 30619 16649
rect 30561 16609 30573 16643
rect 30607 16640 30619 16643
rect 30650 16640 30656 16652
rect 30607 16612 30656 16640
rect 30607 16609 30619 16612
rect 30561 16603 30619 16609
rect 30650 16600 30656 16612
rect 30708 16600 30714 16652
rect 31726 16640 31754 16680
rect 32508 16680 33548 16708
rect 32508 16649 32536 16680
rect 32493 16643 32551 16649
rect 30944 16612 31616 16640
rect 31726 16612 31800 16640
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 20119 16575 20177 16581
rect 20119 16541 20131 16575
rect 20165 16541 20177 16575
rect 20119 16535 20177 16541
rect 20254 16532 20260 16584
rect 20312 16532 20318 16584
rect 20438 16532 20444 16584
rect 20496 16532 20502 16584
rect 21634 16532 21640 16584
rect 21692 16532 21698 16584
rect 22741 16575 22799 16581
rect 22741 16541 22753 16575
rect 22787 16572 22799 16575
rect 22922 16572 22928 16584
rect 22787 16544 22928 16572
rect 22787 16541 22799 16544
rect 22741 16535 22799 16541
rect 22922 16532 22928 16544
rect 22980 16532 22986 16584
rect 28258 16532 28264 16584
rect 28316 16532 28322 16584
rect 29181 16575 29239 16581
rect 29181 16572 29193 16575
rect 28920 16544 29193 16572
rect 13596 16476 13768 16504
rect 13596 16464 13602 16476
rect 14274 16436 14280 16448
rect 13464 16408 14280 16436
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 14829 16439 14887 16445
rect 14829 16405 14841 16439
rect 14875 16436 14887 16439
rect 15212 16436 15240 16532
rect 15289 16507 15347 16513
rect 15289 16473 15301 16507
rect 15335 16504 15347 16507
rect 15562 16504 15568 16516
rect 15335 16476 15568 16504
rect 15335 16473 15347 16476
rect 15289 16467 15347 16473
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 18248 16504 18276 16532
rect 24118 16504 24124 16516
rect 18248 16476 24124 16504
rect 24118 16464 24124 16476
rect 24176 16464 24182 16516
rect 26786 16464 26792 16516
rect 26844 16464 26850 16516
rect 28920 16448 28948 16544
rect 29181 16541 29193 16544
rect 29227 16541 29239 16575
rect 29181 16535 29239 16541
rect 30668 16504 30696 16600
rect 30944 16584 30972 16612
rect 30926 16532 30932 16584
rect 30984 16532 30990 16584
rect 31018 16532 31024 16584
rect 31076 16532 31082 16584
rect 31588 16581 31616 16612
rect 31772 16581 31800 16612
rect 32493 16609 32505 16643
rect 32539 16609 32551 16643
rect 32493 16603 32551 16609
rect 33505 16643 33563 16649
rect 33505 16609 33517 16643
rect 33551 16640 33563 16643
rect 33965 16643 34023 16649
rect 33965 16640 33977 16643
rect 33551 16612 33977 16640
rect 33551 16609 33563 16612
rect 33505 16603 33563 16609
rect 33965 16609 33977 16612
rect 34011 16609 34023 16643
rect 33965 16603 34023 16609
rect 31573 16575 31631 16581
rect 31573 16541 31585 16575
rect 31619 16541 31631 16575
rect 31573 16535 31631 16541
rect 31757 16575 31815 16581
rect 31757 16541 31769 16575
rect 31803 16541 31815 16575
rect 31757 16535 31815 16541
rect 32585 16575 32643 16581
rect 32585 16541 32597 16575
rect 32631 16541 32643 16575
rect 32585 16535 32643 16541
rect 31265 16507 31323 16513
rect 31265 16504 31277 16507
rect 30668 16476 31277 16504
rect 31265 16473 31277 16476
rect 31311 16473 31323 16507
rect 31481 16507 31539 16513
rect 31481 16504 31493 16507
rect 31265 16467 31323 16473
rect 31404 16476 31493 16504
rect 31404 16448 31432 16476
rect 31481 16473 31493 16476
rect 31527 16473 31539 16507
rect 31481 16467 31539 16473
rect 32600 16448 32628 16535
rect 33134 16532 33140 16584
rect 33192 16572 33198 16584
rect 33413 16575 33471 16581
rect 33413 16572 33425 16575
rect 33192 16544 33425 16572
rect 33192 16532 33198 16544
rect 33413 16541 33425 16544
rect 33459 16541 33471 16575
rect 33413 16535 33471 16541
rect 33873 16575 33931 16581
rect 33873 16541 33885 16575
rect 33919 16541 33931 16575
rect 33873 16535 33931 16541
rect 34057 16575 34115 16581
rect 34057 16541 34069 16575
rect 34103 16541 34115 16575
rect 34057 16535 34115 16541
rect 32766 16464 32772 16516
rect 32824 16504 32830 16516
rect 33888 16504 33916 16535
rect 32824 16476 33916 16504
rect 32824 16464 32830 16476
rect 14875 16408 15240 16436
rect 14875 16405 14887 16408
rect 14829 16399 14887 16405
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 15654 16436 15660 16448
rect 15436 16408 15660 16436
rect 15436 16396 15442 16408
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 18233 16439 18291 16445
rect 18233 16405 18245 16439
rect 18279 16436 18291 16439
rect 18414 16436 18420 16448
rect 18279 16408 18420 16436
rect 18279 16405 18291 16408
rect 18233 16399 18291 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 24394 16396 24400 16448
rect 24452 16396 24458 16448
rect 24762 16396 24768 16448
rect 24820 16396 24826 16448
rect 27706 16396 27712 16448
rect 27764 16396 27770 16448
rect 28902 16396 28908 16448
rect 28960 16396 28966 16448
rect 31386 16396 31392 16448
rect 31444 16396 31450 16448
rect 31846 16396 31852 16448
rect 31904 16436 31910 16448
rect 32217 16439 32275 16445
rect 32217 16436 32229 16439
rect 31904 16408 32229 16436
rect 31904 16396 31910 16408
rect 32217 16405 32229 16408
rect 32263 16405 32275 16439
rect 32217 16399 32275 16405
rect 32582 16396 32588 16448
rect 32640 16396 32646 16448
rect 32950 16396 32956 16448
rect 33008 16436 33014 16448
rect 34072 16436 34100 16535
rect 33008 16408 34100 16436
rect 33008 16396 33014 16408
rect 1104 16346 34840 16368
rect 1104 16294 9344 16346
rect 9396 16294 9408 16346
rect 9460 16294 9472 16346
rect 9524 16294 9536 16346
rect 9588 16294 9600 16346
rect 9652 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 17930 16346
rect 17982 16294 17994 16346
rect 18046 16294 26132 16346
rect 26184 16294 26196 16346
rect 26248 16294 26260 16346
rect 26312 16294 26324 16346
rect 26376 16294 26388 16346
rect 26440 16294 34526 16346
rect 34578 16294 34590 16346
rect 34642 16294 34654 16346
rect 34706 16294 34718 16346
rect 34770 16294 34782 16346
rect 34834 16294 34840 16346
rect 1104 16272 34840 16294
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3602 16232 3608 16244
rect 3283 16204 3608 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 3602 16192 3608 16204
rect 3660 16192 3666 16244
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 5166 16232 5172 16244
rect 4856 16204 5172 16232
rect 4856 16192 4862 16204
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 5445 16235 5503 16241
rect 5445 16201 5457 16235
rect 5491 16232 5503 16235
rect 7926 16232 7932 16244
rect 5491 16204 7932 16232
rect 5491 16201 5503 16204
rect 5445 16195 5503 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 8294 16232 8300 16244
rect 8260 16204 8300 16232
rect 8260 16192 8266 16204
rect 8294 16192 8300 16204
rect 8352 16232 8358 16244
rect 8352 16204 8432 16232
rect 8352 16192 8358 16204
rect 4614 16124 4620 16176
rect 4672 16164 4678 16176
rect 5184 16164 5212 16192
rect 8404 16173 8432 16204
rect 8570 16192 8576 16244
rect 8628 16192 8634 16244
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 9493 16235 9551 16241
rect 9493 16232 9505 16235
rect 9180 16204 9505 16232
rect 9180 16192 9186 16204
rect 9493 16201 9505 16204
rect 9539 16232 9551 16235
rect 11146 16232 11152 16244
rect 9539 16204 11152 16232
rect 9539 16201 9551 16204
rect 9493 16195 9551 16201
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 13265 16235 13323 16241
rect 13265 16232 13277 16235
rect 12584 16204 13277 16232
rect 12584 16192 12590 16204
rect 13265 16201 13277 16204
rect 13311 16201 13323 16235
rect 13265 16195 13323 16201
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 18472 16204 18552 16232
rect 18472 16192 18478 16204
rect 18524 16173 18552 16204
rect 19978 16192 19984 16244
rect 20036 16192 20042 16244
rect 22189 16235 22247 16241
rect 22189 16201 22201 16235
rect 22235 16232 22247 16235
rect 22278 16232 22284 16244
rect 22235 16204 22284 16232
rect 22235 16201 22247 16204
rect 22189 16195 22247 16201
rect 22278 16192 22284 16204
rect 22336 16232 22342 16244
rect 23198 16232 23204 16244
rect 22336 16204 23204 16232
rect 22336 16192 22342 16204
rect 23198 16192 23204 16204
rect 23256 16232 23262 16244
rect 23477 16235 23535 16241
rect 23256 16204 23428 16232
rect 23256 16192 23262 16204
rect 5813 16167 5871 16173
rect 5813 16164 5825 16167
rect 4672 16136 5028 16164
rect 5184 16136 5825 16164
rect 4672 16124 4678 16136
rect 1486 16056 1492 16108
rect 1544 16096 1550 16108
rect 2869 16099 2927 16105
rect 2869 16096 2881 16099
rect 1544 16068 2881 16096
rect 1544 16056 1550 16068
rect 2869 16065 2881 16068
rect 2915 16096 2927 16099
rect 4062 16096 4068 16108
rect 2915 16068 4068 16096
rect 2915 16065 2927 16068
rect 2869 16059 2927 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4157 16059 4215 16065
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16096 4399 16099
rect 4706 16096 4712 16108
rect 4387 16068 4712 16096
rect 4387 16065 4399 16068
rect 4341 16059 4399 16065
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 16028 3019 16031
rect 3050 16028 3056 16040
rect 3007 16000 3056 16028
rect 3007 15997 3019 16000
rect 2961 15991 3019 15997
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 4172 16028 4200 16059
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 5000 16105 5028 16136
rect 5813 16133 5825 16136
rect 5859 16133 5871 16167
rect 8389 16167 8447 16173
rect 5813 16127 5871 16133
rect 7024 16136 8340 16164
rect 4985 16099 5043 16105
rect 4985 16065 4997 16099
rect 5031 16096 5043 16099
rect 5261 16099 5319 16105
rect 5031 16068 5212 16096
rect 5031 16065 5043 16068
rect 4985 16059 5043 16065
rect 4798 16028 4804 16040
rect 4172 16000 4804 16028
rect 4798 15988 4804 16000
rect 4856 16028 4862 16040
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 4856 16000 5089 16028
rect 4856 15988 4862 16000
rect 5077 15997 5089 16000
rect 5123 15997 5135 16031
rect 5184 16028 5212 16068
rect 5261 16065 5273 16099
rect 5307 16096 5319 16099
rect 5442 16096 5448 16108
rect 5307 16068 5448 16096
rect 5307 16065 5319 16068
rect 5261 16059 5319 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 7024 16028 7052 16136
rect 8312 16108 8340 16136
rect 8389 16133 8401 16167
rect 8435 16133 8447 16167
rect 18509 16167 18567 16173
rect 8389 16127 8447 16133
rect 15028 16136 15516 16164
rect 15028 16108 15056 16136
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 8220 16028 8248 16059
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 8352 16068 9413 16096
rect 8352 16056 8358 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9674 16056 9680 16108
rect 9732 16056 9738 16108
rect 9858 16056 9864 16108
rect 9916 16056 9922 16108
rect 10318 16056 10324 16108
rect 10376 16056 10382 16108
rect 10502 16056 10508 16108
rect 10560 16056 10566 16108
rect 10686 16056 10692 16108
rect 10744 16056 10750 16108
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16096 10931 16099
rect 11330 16096 11336 16108
rect 10919 16068 11336 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 13173 16099 13231 16105
rect 13173 16096 13185 16099
rect 12860 16068 13185 16096
rect 12860 16056 12866 16068
rect 13173 16065 13185 16068
rect 13219 16065 13231 16099
rect 13173 16059 13231 16065
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 5184 16000 7052 16028
rect 8036 16000 8248 16028
rect 5077 15991 5135 15997
rect 8036 15972 8064 16000
rect 8846 15988 8852 16040
rect 8904 16028 8910 16040
rect 9692 16028 9720 16056
rect 8904 16000 9720 16028
rect 8904 15988 8910 16000
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 10597 16031 10655 16037
rect 10597 16028 10609 16031
rect 10468 16000 10609 16028
rect 10468 15988 10474 16000
rect 10597 15997 10609 16000
rect 10643 16028 10655 16031
rect 11882 16028 11888 16040
rect 10643 16000 11888 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 11882 15988 11888 16000
rect 11940 16028 11946 16040
rect 13372 16028 13400 16059
rect 15010 16056 15016 16108
rect 15068 16056 15074 16108
rect 15194 16056 15200 16108
rect 15252 16056 15258 16108
rect 15378 16056 15384 16108
rect 15436 16056 15442 16108
rect 15488 16105 15516 16136
rect 18509 16133 18521 16167
rect 18555 16133 18567 16167
rect 19996 16164 20024 16192
rect 22738 16164 22744 16176
rect 19996 16136 22744 16164
rect 18509 16127 18567 16133
rect 22738 16124 22744 16136
rect 22796 16124 22802 16176
rect 23400 16164 23428 16204
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 23750 16232 23756 16244
rect 23523 16204 23756 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 24394 16192 24400 16244
rect 24452 16192 24458 16244
rect 24762 16192 24768 16244
rect 24820 16232 24826 16244
rect 26786 16232 26792 16244
rect 24820 16204 26792 16232
rect 24820 16192 24826 16204
rect 26786 16192 26792 16204
rect 26844 16192 26850 16244
rect 27706 16232 27712 16244
rect 27448 16204 27712 16232
rect 24412 16164 24440 16192
rect 23400 16136 23796 16164
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 15562 16056 15568 16108
rect 15620 16096 15626 16108
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 15620 16068 15669 16096
rect 15620 16056 15626 16068
rect 15657 16065 15669 16068
rect 15703 16096 15715 16099
rect 16206 16096 16212 16108
rect 15703 16068 16212 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 19610 16056 19616 16108
rect 19668 16056 19674 16108
rect 22833 16099 22891 16105
rect 22833 16065 22845 16099
rect 22879 16096 22891 16099
rect 22922 16096 22928 16108
rect 22879 16068 22928 16096
rect 22879 16065 22891 16068
rect 22833 16059 22891 16065
rect 22922 16056 22928 16068
rect 22980 16056 22986 16108
rect 23017 16099 23075 16105
rect 23017 16065 23029 16099
rect 23063 16065 23075 16099
rect 23017 16059 23075 16065
rect 11940 16000 13400 16028
rect 15289 16031 15347 16037
rect 11940 15988 11946 16000
rect 15289 15997 15301 16031
rect 15335 16028 15347 16031
rect 15746 16028 15752 16040
rect 15335 16000 15752 16028
rect 15335 15997 15347 16000
rect 15289 15991 15347 15997
rect 15746 15988 15752 16000
rect 15804 15988 15810 16040
rect 18230 15988 18236 16040
rect 18288 15988 18294 16040
rect 22278 15988 22284 16040
rect 22336 15988 22342 16040
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 16028 22523 16031
rect 22738 16028 22744 16040
rect 22511 16000 22744 16028
rect 22511 15997 22523 16000
rect 22465 15991 22523 15997
rect 22738 15988 22744 16000
rect 22796 15988 22802 16040
rect 1946 15920 1952 15972
rect 2004 15960 2010 15972
rect 6914 15960 6920 15972
rect 2004 15932 6920 15960
rect 2004 15920 2010 15932
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 8018 15920 8024 15972
rect 8076 15920 8082 15972
rect 8110 15920 8116 15972
rect 8168 15960 8174 15972
rect 10778 15960 10784 15972
rect 8168 15932 10784 15960
rect 8168 15920 8174 15932
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 11698 15960 11704 15972
rect 10888 15932 11704 15960
rect 4522 15852 4528 15904
rect 4580 15852 4586 15904
rect 5166 15852 5172 15904
rect 5224 15852 5230 15904
rect 5721 15895 5779 15901
rect 5721 15861 5733 15895
rect 5767 15892 5779 15895
rect 6086 15892 6092 15904
rect 5767 15864 6092 15892
rect 5767 15861 5779 15864
rect 5721 15855 5779 15861
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 10888 15892 10916 15932
rect 11698 15920 11704 15932
rect 11756 15920 11762 15972
rect 13262 15920 13268 15972
rect 13320 15960 13326 15972
rect 13538 15960 13544 15972
rect 13320 15932 13544 15960
rect 13320 15920 13326 15932
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 21821 15963 21879 15969
rect 21821 15929 21833 15963
rect 21867 15960 21879 15963
rect 22646 15960 22652 15972
rect 21867 15932 22652 15960
rect 21867 15929 21879 15932
rect 21821 15923 21879 15929
rect 22646 15920 22652 15932
rect 22704 15920 22710 15972
rect 23032 15960 23060 16059
rect 23106 16056 23112 16108
rect 23164 16056 23170 16108
rect 23201 16099 23259 16105
rect 23201 16065 23213 16099
rect 23247 16065 23259 16099
rect 23201 16059 23259 16065
rect 23216 16028 23244 16059
rect 23290 16056 23296 16108
rect 23348 16096 23354 16108
rect 23768 16105 23796 16136
rect 23860 16136 24440 16164
rect 23860 16105 23888 16136
rect 26694 16124 26700 16176
rect 26752 16124 26758 16176
rect 27448 16173 27476 16204
rect 27706 16192 27712 16204
rect 27764 16192 27770 16244
rect 30006 16192 30012 16244
rect 30064 16192 30070 16244
rect 31481 16235 31539 16241
rect 31481 16201 31493 16235
rect 31527 16232 31539 16235
rect 31527 16204 31754 16232
rect 31527 16201 31539 16204
rect 31481 16195 31539 16201
rect 27433 16167 27491 16173
rect 27433 16133 27445 16167
rect 27479 16133 27491 16167
rect 27433 16127 27491 16133
rect 28166 16124 28172 16176
rect 28224 16124 28230 16176
rect 29733 16167 29791 16173
rect 29733 16164 29745 16167
rect 29380 16136 29745 16164
rect 23569 16099 23627 16105
rect 23569 16096 23581 16099
rect 23348 16068 23581 16096
rect 23348 16056 23354 16068
rect 23569 16065 23581 16068
rect 23615 16065 23627 16099
rect 23569 16059 23627 16065
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16065 23811 16099
rect 23753 16059 23811 16065
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16065 23903 16099
rect 23845 16059 23903 16065
rect 24118 16056 24124 16108
rect 24176 16056 24182 16108
rect 26712 16096 26740 16124
rect 29380 16108 29408 16136
rect 29733 16133 29745 16136
rect 29779 16133 29791 16167
rect 30024 16164 30052 16192
rect 31726 16164 31754 16204
rect 32582 16192 32588 16244
rect 32640 16192 32646 16244
rect 32309 16167 32367 16173
rect 32309 16164 32321 16167
rect 30024 16136 30144 16164
rect 31726 16136 32321 16164
rect 29733 16127 29791 16133
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 23216 16000 23673 16028
rect 23661 15997 23673 16000
rect 23707 15997 23719 16031
rect 24397 16031 24455 16037
rect 24397 16028 24409 16031
rect 23661 15991 23719 15997
rect 24044 16000 24409 16028
rect 23474 15960 23480 15972
rect 23032 15932 23480 15960
rect 23474 15920 23480 15932
rect 23532 15920 23538 15972
rect 24044 15969 24072 16000
rect 24397 15997 24409 16000
rect 24443 15997 24455 16031
rect 25516 16028 25544 16082
rect 25700 16068 26740 16096
rect 25590 16028 25596 16040
rect 25516 16000 25596 16028
rect 24397 15991 24455 15997
rect 25590 15988 25596 16000
rect 25648 16028 25654 16040
rect 25700 16028 25728 16068
rect 26878 16056 26884 16108
rect 26936 16096 26942 16108
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 26936 16068 27169 16096
rect 26936 16056 26942 16068
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 28994 16056 29000 16108
rect 29052 16056 29058 16108
rect 29362 16056 29368 16108
rect 29420 16056 29426 16108
rect 30116 16105 30144 16136
rect 32309 16133 32321 16136
rect 32355 16164 32367 16167
rect 32600 16164 32628 16192
rect 32677 16167 32735 16173
rect 32677 16164 32689 16167
rect 32355 16136 32689 16164
rect 32355 16133 32367 16136
rect 32309 16127 32367 16133
rect 32677 16133 32689 16136
rect 32723 16133 32735 16167
rect 32677 16127 32735 16133
rect 32858 16124 32864 16176
rect 32916 16124 32922 16176
rect 29636 16099 29694 16105
rect 29636 16096 29648 16099
rect 29564 16068 29648 16096
rect 25648 16000 25728 16028
rect 25869 16031 25927 16037
rect 25648 15988 25654 16000
rect 25869 15997 25881 16031
rect 25915 16028 25927 16031
rect 26145 16031 26203 16037
rect 26145 16028 26157 16031
rect 25915 16000 26157 16028
rect 25915 15997 25927 16000
rect 25869 15991 25927 15997
rect 26145 15997 26157 16000
rect 26191 15997 26203 16031
rect 26145 15991 26203 15997
rect 27430 15988 27436 16040
rect 27488 16028 27494 16040
rect 28166 16028 28172 16040
rect 27488 16000 28172 16028
rect 27488 15988 27494 16000
rect 28166 15988 28172 16000
rect 28224 15988 28230 16040
rect 29012 16028 29040 16056
rect 29564 16028 29592 16068
rect 29636 16065 29648 16068
rect 29682 16065 29694 16099
rect 29636 16059 29694 16065
rect 29825 16099 29883 16105
rect 29825 16065 29837 16099
rect 29871 16065 29883 16099
rect 29825 16059 29883 16065
rect 30008 16099 30066 16105
rect 30008 16065 30020 16099
rect 30054 16065 30066 16099
rect 30008 16059 30066 16065
rect 30101 16099 30159 16105
rect 30101 16065 30113 16099
rect 30147 16065 30159 16099
rect 30101 16059 30159 16065
rect 29012 16000 29592 16028
rect 24029 15963 24087 15969
rect 24029 15929 24041 15963
rect 24075 15929 24087 15963
rect 24029 15923 24087 15929
rect 6420 15864 10916 15892
rect 11057 15895 11115 15901
rect 6420 15852 6426 15864
rect 11057 15861 11069 15895
rect 11103 15892 11115 15895
rect 13078 15892 13084 15904
rect 11103 15864 13084 15892
rect 11103 15861 11115 15864
rect 11057 15855 11115 15861
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15436 15864 15669 15892
rect 15436 15852 15442 15864
rect 15657 15861 15669 15864
rect 15703 15861 15715 15895
rect 15657 15855 15715 15861
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 23290 15892 23296 15904
rect 20312 15864 23296 15892
rect 20312 15852 20318 15864
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 28166 15852 28172 15904
rect 28224 15892 28230 15904
rect 28902 15892 28908 15904
rect 28224 15864 28908 15892
rect 28224 15852 28230 15864
rect 28902 15852 28908 15864
rect 28960 15852 28966 15904
rect 29454 15852 29460 15904
rect 29512 15852 29518 15904
rect 29840 15892 29868 16059
rect 30024 16028 30052 16059
rect 31018 16056 31024 16108
rect 31076 16096 31082 16108
rect 31297 16099 31355 16105
rect 31297 16096 31309 16099
rect 31076 16068 31309 16096
rect 31076 16056 31082 16068
rect 31297 16065 31309 16068
rect 31343 16065 31355 16099
rect 31297 16059 31355 16065
rect 31386 16056 31392 16108
rect 31444 16096 31450 16108
rect 31481 16099 31539 16105
rect 31481 16096 31493 16099
rect 31444 16068 31493 16096
rect 31444 16056 31450 16068
rect 31481 16065 31493 16068
rect 31527 16065 31539 16099
rect 31481 16059 31539 16065
rect 32214 16056 32220 16108
rect 32272 16096 32278 16108
rect 32493 16099 32551 16105
rect 32493 16096 32505 16099
rect 32272 16068 32505 16096
rect 32272 16056 32278 16068
rect 32493 16065 32505 16068
rect 32539 16096 32551 16099
rect 32585 16099 32643 16105
rect 32585 16096 32597 16099
rect 32539 16068 32597 16096
rect 32539 16065 32551 16068
rect 32493 16059 32551 16065
rect 32585 16065 32597 16068
rect 32631 16065 32643 16099
rect 32585 16059 32643 16065
rect 30024 16000 32904 16028
rect 31018 15920 31024 15972
rect 31076 15960 31082 15972
rect 32766 15960 32772 15972
rect 31076 15932 32772 15960
rect 31076 15920 31082 15932
rect 32766 15920 32772 15932
rect 32824 15920 32830 15972
rect 32876 15969 32904 16000
rect 32861 15963 32919 15969
rect 32861 15929 32873 15963
rect 32907 15929 32919 15963
rect 32861 15923 32919 15929
rect 32125 15895 32183 15901
rect 32125 15892 32137 15895
rect 29840 15864 32137 15892
rect 32125 15861 32137 15864
rect 32171 15892 32183 15895
rect 32950 15892 32956 15904
rect 32171 15864 32956 15892
rect 32171 15861 32183 15864
rect 32125 15855 32183 15861
rect 32950 15852 32956 15864
rect 33008 15852 33014 15904
rect 1104 15802 34684 15824
rect 1104 15750 5147 15802
rect 5199 15750 5211 15802
rect 5263 15750 5275 15802
rect 5327 15750 5339 15802
rect 5391 15750 5403 15802
rect 5455 15750 13541 15802
rect 13593 15750 13605 15802
rect 13657 15750 13669 15802
rect 13721 15750 13733 15802
rect 13785 15750 13797 15802
rect 13849 15750 21935 15802
rect 21987 15750 21999 15802
rect 22051 15750 22063 15802
rect 22115 15750 22127 15802
rect 22179 15750 22191 15802
rect 22243 15750 30329 15802
rect 30381 15750 30393 15802
rect 30445 15750 30457 15802
rect 30509 15750 30521 15802
rect 30573 15750 30585 15802
rect 30637 15750 34684 15802
rect 1104 15728 34684 15750
rect 3255 15691 3313 15697
rect 3255 15657 3267 15691
rect 3301 15688 3313 15691
rect 3786 15688 3792 15700
rect 3301 15660 3792 15688
rect 3301 15657 3313 15660
rect 3255 15651 3313 15657
rect 3786 15648 3792 15660
rect 3844 15648 3850 15700
rect 6362 15648 6368 15700
rect 6420 15688 6426 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 6420 15660 7205 15688
rect 6420 15648 6426 15660
rect 7193 15657 7205 15660
rect 7239 15657 7251 15691
rect 7193 15651 7251 15657
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 7558 15688 7564 15700
rect 7423 15660 7564 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 6822 15620 6828 15632
rect 3528 15592 6828 15620
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 3528 15561 3556 15592
rect 6822 15580 6828 15592
rect 6880 15580 6886 15632
rect 7208 15620 7236 15651
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 8018 15648 8024 15700
rect 8076 15648 8082 15700
rect 8570 15648 8576 15700
rect 8628 15648 8634 15700
rect 10042 15688 10048 15700
rect 8956 15660 10048 15688
rect 7208 15592 7512 15620
rect 3513 15555 3571 15561
rect 3513 15552 3525 15555
rect 1452 15524 3525 15552
rect 1452 15512 1458 15524
rect 3513 15521 3525 15524
rect 3559 15521 3571 15555
rect 3513 15515 3571 15521
rect 6270 15512 6276 15564
rect 6328 15512 6334 15564
rect 7374 15512 7380 15564
rect 7432 15512 7438 15564
rect 1486 15444 1492 15496
rect 1544 15444 1550 15496
rect 5626 15444 5632 15496
rect 5684 15444 5690 15496
rect 5997 15487 6055 15493
rect 5997 15453 6009 15487
rect 6043 15453 6055 15487
rect 5997 15447 6055 15453
rect 2958 15416 2964 15428
rect 2806 15388 2964 15416
rect 2958 15376 2964 15388
rect 3016 15376 3022 15428
rect 5644 15348 5672 15444
rect 6012 15416 6040 15447
rect 6086 15444 6092 15496
rect 6144 15444 6150 15496
rect 6288 15416 6316 15512
rect 7009 15487 7067 15493
rect 7009 15484 7021 15487
rect 6012 15388 6316 15416
rect 6380 15456 7021 15484
rect 6086 15348 6092 15360
rect 5644 15320 6092 15348
rect 6086 15308 6092 15320
rect 6144 15348 6150 15360
rect 6380 15348 6408 15456
rect 7009 15453 7021 15456
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 7193 15487 7251 15493
rect 7193 15453 7205 15487
rect 7239 15484 7251 15487
rect 7392 15484 7420 15512
rect 7484 15493 7512 15592
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15552 7619 15555
rect 8036 15552 8064 15648
rect 8956 15632 8984 15660
rect 8386 15580 8392 15632
rect 8444 15580 8450 15632
rect 8938 15580 8944 15632
rect 8996 15580 9002 15632
rect 8404 15552 8432 15580
rect 7607 15524 8248 15552
rect 8404 15524 9260 15552
rect 7607 15521 7619 15524
rect 7561 15515 7619 15521
rect 7239 15456 7420 15484
rect 7239 15453 7251 15456
rect 7193 15447 7251 15453
rect 6917 15419 6975 15425
rect 6917 15385 6929 15419
rect 6963 15385 6975 15419
rect 7392 15416 7420 15456
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15453 7527 15487
rect 7469 15447 7527 15453
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15453 7987 15487
rect 7929 15447 7987 15453
rect 7558 15416 7564 15428
rect 7392 15388 7564 15416
rect 6917 15379 6975 15385
rect 6144 15320 6408 15348
rect 6932 15348 6960 15379
rect 7558 15376 7564 15388
rect 7616 15416 7622 15428
rect 7668 15416 7696 15447
rect 7944 15416 7972 15447
rect 8018 15444 8024 15496
rect 8076 15444 8082 15496
rect 8110 15444 8116 15496
rect 8168 15444 8174 15496
rect 8220 15484 8248 15524
rect 9232 15493 9260 15524
rect 8394 15487 8452 15493
rect 8394 15484 8406 15487
rect 8220 15456 8406 15484
rect 8394 15453 8406 15456
rect 8440 15453 8452 15487
rect 8394 15447 8452 15453
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 9508 15493 9536 15660
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10321 15691 10379 15697
rect 10321 15657 10333 15691
rect 10367 15688 10379 15691
rect 10502 15688 10508 15700
rect 10367 15660 10508 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 10778 15648 10784 15700
rect 10836 15648 10842 15700
rect 13262 15648 13268 15700
rect 13320 15648 13326 15700
rect 14921 15691 14979 15697
rect 14921 15657 14933 15691
rect 14967 15688 14979 15691
rect 15194 15688 15200 15700
rect 14967 15660 15200 15688
rect 14967 15657 14979 15660
rect 14921 15651 14979 15657
rect 15194 15648 15200 15660
rect 15252 15688 15258 15700
rect 15838 15688 15844 15700
rect 15252 15660 15844 15688
rect 15252 15648 15258 15660
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 20898 15688 20904 15700
rect 19904 15660 20904 15688
rect 10686 15512 10692 15564
rect 10744 15512 10750 15564
rect 10796 15552 10824 15648
rect 11514 15580 11520 15632
rect 11572 15580 11578 15632
rect 12066 15620 12072 15632
rect 11808 15592 12072 15620
rect 11532 15552 11560 15580
rect 11808 15564 11836 15592
rect 12066 15580 12072 15592
rect 12124 15620 12130 15632
rect 12124 15592 12940 15620
rect 12124 15580 12130 15592
rect 10796 15524 11468 15552
rect 11532 15524 11652 15552
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9582 15444 9588 15496
rect 9640 15444 9646 15496
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 9916 15456 10609 15484
rect 9916 15444 9922 15456
rect 10597 15453 10609 15456
rect 10643 15484 10655 15487
rect 10778 15484 10784 15496
rect 10643 15456 10784 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 10870 15444 10876 15496
rect 10928 15444 10934 15496
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 11146 15444 11152 15496
rect 11204 15481 11210 15496
rect 11440 15493 11468 15524
rect 11624 15493 11652 15524
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15552 11943 15555
rect 11931 15524 12756 15552
rect 11931 15521 11943 15524
rect 11885 15515 11943 15521
rect 12728 15493 12756 15524
rect 12912 15493 12940 15592
rect 15102 15580 15108 15632
rect 15160 15580 15166 15632
rect 15856 15620 15884 15648
rect 16298 15620 16304 15632
rect 15856 15592 16304 15620
rect 16298 15580 16304 15592
rect 16356 15620 16362 15632
rect 16356 15592 16528 15620
rect 16356 15580 16362 15592
rect 15120 15552 15148 15580
rect 14752 15524 15148 15552
rect 14752 15493 14780 15524
rect 11241 15487 11299 15493
rect 11241 15481 11253 15487
rect 11204 15453 11253 15481
rect 11287 15453 11299 15487
rect 11204 15444 11210 15453
rect 11241 15447 11299 15453
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11517 15487 11575 15493
rect 11517 15453 11529 15487
rect 11563 15453 11575 15487
rect 11517 15447 11575 15453
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15484 11667 15487
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 11655 15456 12357 15484
rect 11655 15453 11667 15456
rect 11609 15447 11667 15453
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 12345 15447 12403 15453
rect 12452 15456 12633 15484
rect 8128 15416 8156 15444
rect 7616 15388 7696 15416
rect 7760 15388 8156 15416
rect 7616 15376 7622 15388
rect 7760 15360 7788 15388
rect 8202 15376 8208 15428
rect 8260 15376 8266 15428
rect 8297 15419 8355 15425
rect 8297 15385 8309 15419
rect 8343 15416 8355 15419
rect 9674 15416 9680 15428
rect 8343 15388 9680 15416
rect 8343 15385 8355 15388
rect 8297 15379 8355 15385
rect 7742 15348 7748 15360
rect 6932 15320 7748 15348
rect 6144 15308 6150 15320
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 7926 15308 7932 15360
rect 7984 15348 7990 15360
rect 8312 15348 8340 15379
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 10686 15376 10692 15428
rect 10744 15416 10750 15428
rect 11532 15416 11560 15447
rect 10744 15388 11560 15416
rect 10744 15376 10750 15388
rect 12158 15376 12164 15428
rect 12216 15376 12222 15428
rect 7984 15320 8340 15348
rect 7984 15308 7990 15320
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9582 15348 9588 15360
rect 8996 15320 9588 15348
rect 8996 15308 9002 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 10042 15308 10048 15360
rect 10100 15348 10106 15360
rect 10870 15348 10876 15360
rect 10100 15320 10876 15348
rect 10100 15308 10106 15320
rect 10870 15308 10876 15320
rect 10928 15308 10934 15360
rect 11882 15308 11888 15360
rect 11940 15348 11946 15360
rect 12452 15348 12480 15456
rect 12621 15453 12633 15456
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 12713 15487 12771 15493
rect 12713 15453 12725 15487
rect 12759 15453 12771 15487
rect 12713 15447 12771 15453
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 14737 15487 14795 15493
rect 13127 15456 13216 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 12986 15376 12992 15428
rect 13044 15376 13050 15428
rect 13188 15360 13216 15456
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14826 15444 14832 15496
rect 14884 15444 14890 15496
rect 15120 15484 15148 15524
rect 16390 15512 16396 15564
rect 16448 15512 16454 15564
rect 16500 15561 16528 15592
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15552 16911 15555
rect 16899 15524 17264 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 16022 15484 16028 15496
rect 15120 15456 16028 15484
rect 16022 15444 16028 15456
rect 16080 15484 16086 15496
rect 16577 15487 16635 15493
rect 16577 15484 16589 15487
rect 16080 15456 16589 15484
rect 16080 15444 16086 15456
rect 16577 15453 16589 15456
rect 16623 15453 16635 15487
rect 16577 15447 16635 15453
rect 16666 15444 16672 15496
rect 16724 15444 16730 15496
rect 17236 15493 17264 15524
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 19904 15552 19932 15660
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 21453 15691 21511 15697
rect 21453 15657 21465 15691
rect 21499 15688 21511 15691
rect 21634 15688 21640 15700
rect 21499 15660 21640 15688
rect 21499 15657 21511 15660
rect 21453 15651 21511 15657
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 22922 15648 22928 15700
rect 22980 15648 22986 15700
rect 26786 15648 26792 15700
rect 26844 15688 26850 15700
rect 27709 15691 27767 15697
rect 26844 15660 27292 15688
rect 26844 15648 26850 15660
rect 21085 15623 21143 15629
rect 21085 15589 21097 15623
rect 21131 15620 21143 15623
rect 22738 15620 22744 15632
rect 21131 15592 22744 15620
rect 21131 15589 21143 15592
rect 21085 15583 21143 15589
rect 22738 15580 22744 15592
rect 22796 15580 22802 15632
rect 23385 15623 23443 15629
rect 23385 15589 23397 15623
rect 23431 15620 23443 15623
rect 23474 15620 23480 15632
rect 23431 15592 23480 15620
rect 23431 15589 23443 15592
rect 23385 15583 23443 15589
rect 23474 15580 23480 15592
rect 23532 15580 23538 15632
rect 22278 15552 22284 15564
rect 19484 15524 19932 15552
rect 19484 15512 19490 15524
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 17589 15487 17647 15493
rect 17589 15484 17601 15487
rect 17451 15456 17601 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 17589 15453 17601 15456
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 19904 15484 19932 15524
rect 21744 15524 22284 15552
rect 21744 15496 21772 15524
rect 22278 15512 22284 15524
rect 22336 15512 22342 15564
rect 23290 15512 23296 15564
rect 23348 15512 23354 15564
rect 19843 15456 19932 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 16960 15416 16988 15447
rect 15120 15388 16988 15416
rect 17865 15419 17923 15425
rect 11940 15320 12480 15348
rect 12529 15351 12587 15357
rect 11940 15308 11946 15320
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 13170 15348 13176 15360
rect 12575 15320 13176 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 15120 15357 15148 15388
rect 17865 15385 17877 15419
rect 17911 15416 17923 15419
rect 19242 15416 19248 15428
rect 17911 15388 19248 15416
rect 17911 15385 17923 15388
rect 17865 15379 17923 15385
rect 19242 15376 19248 15388
rect 19300 15376 19306 15428
rect 19536 15360 19564 15447
rect 19978 15444 19984 15496
rect 20036 15444 20042 15496
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 20622 15484 20628 15496
rect 20220 15456 20628 15484
rect 20220 15444 20226 15456
rect 20622 15444 20628 15456
rect 20680 15484 20686 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 20680 15456 21097 15484
rect 20680 15444 20686 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15453 21235 15487
rect 21177 15447 21235 15453
rect 20438 15376 20444 15428
rect 20496 15416 20502 15428
rect 20990 15416 20996 15428
rect 20496 15388 20996 15416
rect 20496 15376 20502 15388
rect 20990 15376 20996 15388
rect 21048 15416 21054 15428
rect 21192 15416 21220 15447
rect 21634 15444 21640 15496
rect 21692 15444 21698 15496
rect 21726 15444 21732 15496
rect 21784 15444 21790 15496
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15484 22799 15487
rect 23308 15484 23336 15512
rect 23492 15493 23520 15580
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 25777 15555 25835 15561
rect 25777 15552 25789 15555
rect 24176 15524 25789 15552
rect 24176 15512 24182 15524
rect 25777 15521 25789 15524
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 22787 15456 23336 15484
rect 23477 15487 23535 15493
rect 22787 15453 22799 15456
rect 22741 15447 22799 15453
rect 23477 15453 23489 15487
rect 23523 15453 23535 15487
rect 23477 15447 23535 15453
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 21048 15388 21220 15416
rect 21048 15376 21054 15388
rect 22002 15376 22008 15428
rect 22060 15376 22066 15428
rect 22097 15419 22155 15425
rect 22097 15385 22109 15419
rect 22143 15385 22155 15419
rect 22097 15379 22155 15385
rect 15105 15351 15163 15357
rect 15105 15317 15117 15351
rect 15151 15317 15163 15351
rect 15105 15311 15163 15317
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 17037 15351 17095 15357
rect 17037 15348 17049 15351
rect 16540 15320 17049 15348
rect 16540 15308 16546 15320
rect 17037 15317 17049 15320
rect 17083 15348 17095 15351
rect 18138 15348 18144 15360
rect 17083 15320 18144 15348
rect 17083 15317 17095 15320
rect 17037 15311 17095 15317
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 19518 15308 19524 15360
rect 19576 15308 19582 15360
rect 19613 15351 19671 15357
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 19978 15348 19984 15360
rect 19659 15320 19984 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 19978 15308 19984 15320
rect 20036 15348 20042 15360
rect 20346 15348 20352 15360
rect 20036 15320 20352 15348
rect 20036 15308 20042 15320
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 22112 15348 22140 15379
rect 22278 15376 22284 15428
rect 22336 15416 22342 15428
rect 22557 15419 22615 15425
rect 22557 15416 22569 15419
rect 22336 15388 22569 15416
rect 22336 15376 22342 15388
rect 22557 15385 22569 15388
rect 22603 15416 22615 15419
rect 22830 15416 22836 15428
rect 22603 15388 22836 15416
rect 22603 15385 22615 15388
rect 22557 15379 22615 15385
rect 22830 15376 22836 15388
rect 22888 15376 22894 15428
rect 23017 15419 23075 15425
rect 23017 15385 23029 15419
rect 23063 15385 23075 15419
rect 23017 15379 23075 15385
rect 22922 15348 22928 15360
rect 22112 15320 22928 15348
rect 22922 15308 22928 15320
rect 22980 15348 22986 15360
rect 23032 15348 23060 15379
rect 23198 15376 23204 15428
rect 23256 15376 23262 15428
rect 23290 15376 23296 15428
rect 23348 15416 23354 15428
rect 23676 15416 23704 15447
rect 25498 15444 25504 15496
rect 25556 15444 25562 15496
rect 27264 15484 27292 15660
rect 27709 15657 27721 15691
rect 27755 15688 27767 15691
rect 28258 15688 28264 15700
rect 27755 15660 28264 15688
rect 27755 15657 27767 15660
rect 27709 15651 27767 15657
rect 28258 15648 28264 15660
rect 28316 15648 28322 15700
rect 29454 15648 29460 15700
rect 29512 15648 29518 15700
rect 29641 15691 29699 15697
rect 29641 15657 29653 15691
rect 29687 15657 29699 15691
rect 29641 15651 29699 15657
rect 27890 15580 27896 15632
rect 27948 15580 27954 15632
rect 28074 15580 28080 15632
rect 28132 15620 28138 15632
rect 28132 15592 28304 15620
rect 28132 15580 28138 15592
rect 27908 15552 27936 15580
rect 27908 15524 28120 15552
rect 28092 15493 28120 15524
rect 28166 15512 28172 15564
rect 28224 15512 28230 15564
rect 28276 15493 28304 15592
rect 27893 15487 27951 15493
rect 27893 15484 27905 15487
rect 27264 15456 27905 15484
rect 27893 15453 27905 15456
rect 27939 15453 27951 15487
rect 27893 15447 27951 15453
rect 28077 15487 28135 15493
rect 28077 15453 28089 15487
rect 28123 15453 28135 15487
rect 28077 15447 28135 15453
rect 28261 15487 28319 15493
rect 28261 15453 28273 15487
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 28445 15487 28503 15493
rect 28445 15453 28457 15487
rect 28491 15484 28503 15487
rect 29472 15484 29500 15648
rect 28491 15456 29500 15484
rect 28491 15453 28503 15456
rect 28445 15447 28503 15453
rect 29546 15444 29552 15496
rect 29604 15444 29610 15496
rect 29656 15484 29684 15651
rect 29730 15648 29736 15700
rect 29788 15688 29794 15700
rect 30193 15691 30251 15697
rect 30193 15688 30205 15691
rect 29788 15660 30205 15688
rect 29788 15648 29794 15660
rect 30193 15657 30205 15660
rect 30239 15657 30251 15691
rect 30193 15651 30251 15657
rect 30561 15691 30619 15697
rect 30561 15657 30573 15691
rect 30607 15688 30619 15691
rect 31386 15688 31392 15700
rect 30607 15660 31392 15688
rect 30607 15657 30619 15660
rect 30561 15651 30619 15657
rect 31386 15648 31392 15660
rect 31444 15648 31450 15700
rect 30009 15623 30067 15629
rect 30009 15589 30021 15623
rect 30055 15620 30067 15623
rect 31018 15620 31024 15632
rect 30055 15592 31024 15620
rect 30055 15589 30067 15592
rect 30009 15583 30067 15589
rect 31018 15580 31024 15592
rect 31076 15580 31082 15632
rect 30101 15487 30159 15493
rect 30101 15484 30113 15487
rect 29656 15456 30113 15484
rect 26053 15419 26111 15425
rect 26053 15416 26065 15419
rect 23348 15388 23704 15416
rect 25700 15388 26065 15416
rect 23348 15376 23354 15388
rect 22980 15320 23060 15348
rect 23569 15351 23627 15357
rect 22980 15308 22986 15320
rect 23569 15317 23581 15351
rect 23615 15348 23627 15351
rect 24946 15348 24952 15360
rect 23615 15320 24952 15348
rect 23615 15317 23627 15320
rect 23569 15311 23627 15317
rect 24946 15308 24952 15320
rect 25004 15308 25010 15360
rect 25700 15357 25728 15388
rect 26053 15385 26065 15388
rect 26099 15385 26111 15419
rect 27430 15416 27436 15428
rect 27278 15388 27436 15416
rect 26053 15379 26111 15385
rect 27430 15376 27436 15388
rect 27488 15376 27494 15428
rect 29656 15416 29684 15456
rect 30101 15453 30113 15456
rect 30147 15453 30159 15487
rect 30101 15447 30159 15453
rect 27540 15388 29684 15416
rect 27540 15360 27568 15388
rect 25685 15351 25743 15357
rect 25685 15317 25697 15351
rect 25731 15317 25743 15351
rect 25685 15311 25743 15317
rect 27522 15308 27528 15360
rect 27580 15308 27586 15360
rect 28994 15308 29000 15360
rect 29052 15348 29058 15360
rect 31938 15348 31944 15360
rect 29052 15320 31944 15348
rect 29052 15308 29058 15320
rect 31938 15308 31944 15320
rect 31996 15348 32002 15360
rect 33410 15348 33416 15360
rect 31996 15320 33416 15348
rect 31996 15308 32002 15320
rect 33410 15308 33416 15320
rect 33468 15308 33474 15360
rect 1104 15258 34840 15280
rect 1104 15206 9344 15258
rect 9396 15206 9408 15258
rect 9460 15206 9472 15258
rect 9524 15206 9536 15258
rect 9588 15206 9600 15258
rect 9652 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 17930 15258
rect 17982 15206 17994 15258
rect 18046 15206 26132 15258
rect 26184 15206 26196 15258
rect 26248 15206 26260 15258
rect 26312 15206 26324 15258
rect 26376 15206 26388 15258
rect 26440 15206 34526 15258
rect 34578 15206 34590 15258
rect 34642 15206 34654 15258
rect 34706 15206 34718 15258
rect 34770 15206 34782 15258
rect 34834 15206 34840 15258
rect 1104 15184 34840 15206
rect 3145 15147 3203 15153
rect 3145 15113 3157 15147
rect 3191 15144 3203 15147
rect 4798 15144 4804 15156
rect 3191 15116 4804 15144
rect 3191 15113 3203 15116
rect 3145 15107 3203 15113
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 5810 15144 5816 15156
rect 5767 15116 5816 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 5810 15104 5816 15116
rect 5868 15104 5874 15156
rect 6914 15104 6920 15156
rect 6972 15104 6978 15156
rect 7098 15104 7104 15156
rect 7156 15110 7162 15156
rect 7156 15104 7236 15110
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8297 15147 8355 15153
rect 8297 15144 8309 15147
rect 7892 15116 8309 15144
rect 7892 15104 7898 15116
rect 8297 15113 8309 15116
rect 8343 15113 8355 15147
rect 8297 15107 8355 15113
rect 9766 15104 9772 15156
rect 9824 15104 9830 15156
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 10873 15147 10931 15153
rect 10873 15144 10885 15147
rect 10836 15116 10885 15144
rect 10836 15104 10842 15116
rect 10873 15113 10885 15116
rect 10919 15113 10931 15147
rect 10873 15107 10931 15113
rect 12618 15104 12624 15156
rect 12676 15104 12682 15156
rect 13078 15104 13084 15156
rect 13136 15144 13142 15156
rect 17221 15147 17279 15153
rect 13136 15116 14228 15144
rect 13136 15104 13142 15116
rect 3270 15048 4108 15076
rect 3050 14968 3056 15020
rect 3108 14968 3114 15020
rect 3270 15006 3298 15048
rect 4080 15020 4108 15048
rect 4172 15048 4476 15076
rect 3326 15006 3332 15020
rect 3270 14978 3332 15006
rect 3326 14968 3332 14978
rect 3384 14968 3390 15020
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 15008 3663 15011
rect 3970 15008 3976 15020
rect 3651 14980 3976 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 3068 14940 3096 14968
rect 3436 14940 3464 14971
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4062 14968 4068 15020
rect 4120 14968 4126 15020
rect 3988 14940 4016 14968
rect 4172 14940 4200 15048
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 4448 15008 4476 15048
rect 4522 15036 4528 15088
rect 4580 15076 4586 15088
rect 5445 15079 5503 15085
rect 5445 15076 5457 15079
rect 4580 15048 5457 15076
rect 4580 15036 4586 15048
rect 5445 15045 5457 15048
rect 5491 15045 5503 15079
rect 5445 15039 5503 15045
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 7116 15085 7236 15104
rect 7116 15082 7251 15085
rect 7116 15076 7144 15082
rect 6880 15048 7144 15076
rect 7193 15079 7251 15082
rect 6880 15036 6886 15048
rect 7193 15045 7205 15079
rect 7239 15045 7251 15079
rect 7193 15039 7251 15045
rect 7285 15079 7343 15085
rect 7285 15045 7297 15079
rect 7331 15076 7343 15079
rect 12636 15076 12664 15104
rect 13817 15079 13875 15085
rect 13817 15076 13829 15079
rect 7331 15048 7512 15076
rect 7331 15045 7343 15048
rect 7285 15039 7343 15045
rect 7484 15020 7512 15048
rect 7576 15048 12664 15076
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 4448 14980 4629 15008
rect 4249 14971 4307 14977
rect 4617 14977 4629 14980
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 15008 5227 15011
rect 5534 15008 5540 15020
rect 5215 14980 5540 15008
rect 5215 14977 5227 14980
rect 5169 14971 5227 14977
rect 3068 14912 3924 14940
rect 3988 14912 4200 14940
rect 3513 14875 3571 14881
rect 3513 14841 3525 14875
rect 3559 14841 3571 14875
rect 3896 14872 3924 14912
rect 4264 14872 4292 14971
rect 5534 14968 5540 14980
rect 5592 14968 5598 15020
rect 7101 15011 7159 15017
rect 7101 14977 7113 15011
rect 7147 14977 7159 15011
rect 7101 14971 7159 14977
rect 4338 14872 4344 14884
rect 3896 14844 4344 14872
rect 3513 14835 3571 14841
rect 3528 14804 3556 14835
rect 4338 14832 4344 14844
rect 4396 14832 4402 14884
rect 4706 14832 4712 14884
rect 4764 14872 4770 14884
rect 5169 14875 5227 14881
rect 5169 14872 5181 14875
rect 4764 14844 5181 14872
rect 4764 14832 4770 14844
rect 5169 14841 5181 14844
rect 5215 14841 5227 14875
rect 5169 14835 5227 14841
rect 5534 14832 5540 14884
rect 5592 14832 5598 14884
rect 7116 14872 7144 14971
rect 7374 14968 7380 15020
rect 7432 14968 7438 15020
rect 7466 14968 7472 15020
rect 7524 14968 7530 15020
rect 7576 15017 7604 15048
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 14977 7619 15011
rect 7561 14971 7619 14977
rect 8662 14968 8668 15020
rect 8720 15008 8726 15020
rect 8849 15011 8907 15017
rect 8849 15008 8861 15011
rect 8720 14980 8861 15008
rect 8720 14968 8726 14980
rect 8849 14977 8861 14980
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 8938 14968 8944 15020
rect 8996 15008 9002 15020
rect 9309 15011 9367 15017
rect 9309 15008 9321 15011
rect 8996 14980 9321 15008
rect 8996 14968 9002 14980
rect 9309 14977 9321 14980
rect 9355 14977 9367 15011
rect 9309 14971 9367 14977
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 9674 15008 9680 15020
rect 9631 14980 9680 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 10410 14968 10416 15020
rect 10468 15008 10474 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10468 14980 10793 15008
rect 10468 14968 10474 14980
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 15008 11115 15011
rect 11882 15008 11888 15020
rect 11103 14980 11888 15008
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 12032 14980 12265 15008
rect 12032 14968 12038 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 12342 14968 12348 15020
rect 12400 15008 12406 15020
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 12400 14980 12449 15008
rect 12400 14968 12406 14980
rect 12437 14977 12449 14980
rect 12483 14977 12495 15011
rect 12636 15008 12664 15048
rect 13188 15048 13829 15076
rect 13188 15017 13216 15048
rect 13817 15045 13829 15048
rect 13863 15045 13875 15079
rect 13817 15039 13875 15045
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12636 14980 13093 15008
rect 12437 14971 12495 14977
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 14977 13231 15011
rect 13173 14971 13231 14977
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 13446 14968 13452 15020
rect 13504 14968 13510 15020
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 8018 14940 8024 14952
rect 7340 14912 8024 14940
rect 7340 14900 7346 14912
rect 8018 14900 8024 14912
rect 8076 14940 8082 14952
rect 8573 14943 8631 14949
rect 8573 14940 8585 14943
rect 8076 14912 8585 14940
rect 8076 14900 8082 14912
rect 8573 14909 8585 14912
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 9030 14900 9036 14952
rect 9088 14940 9094 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 9088 14912 9413 14940
rect 9088 14900 9094 14912
rect 9401 14909 9413 14912
rect 9447 14940 9459 14943
rect 9766 14940 9772 14952
rect 9447 14912 9772 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 13556 14940 13584 14971
rect 13906 14968 13912 15020
rect 13964 15008 13970 15020
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13964 14980 14013 15008
rect 13964 14968 13970 14980
rect 14001 14977 14013 14980
rect 14047 15008 14059 15011
rect 14090 15008 14096 15020
rect 14047 14980 14096 15008
rect 14047 14977 14059 14980
rect 14001 14971 14059 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14200 15017 14228 15116
rect 17221 15113 17233 15147
rect 17267 15113 17279 15147
rect 17221 15107 17279 15113
rect 16482 15036 16488 15088
rect 16540 15036 16546 15088
rect 17236 15076 17264 15107
rect 19242 15104 19248 15156
rect 19300 15144 19306 15156
rect 20162 15144 20168 15156
rect 19300 15116 20168 15144
rect 19300 15104 19306 15116
rect 17236 15048 18368 15076
rect 18340 15020 18368 15048
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14292 14940 14320 14971
rect 15470 14968 15476 15020
rect 15528 14968 15534 15020
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 16022 14968 16028 15020
rect 16080 15008 16086 15020
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 16080 14980 16129 15008
rect 16080 14968 16086 14980
rect 16117 14977 16129 14980
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 9916 14912 13584 14940
rect 13648 14912 14320 14940
rect 16132 14940 16160 14971
rect 16298 14968 16304 15020
rect 16356 15008 16362 15020
rect 16850 15008 16856 15020
rect 16356 14980 16856 15008
rect 16356 14968 16362 14980
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 17957 15011 18015 15017
rect 17957 14977 17969 15011
rect 18003 15008 18015 15011
rect 18138 15008 18144 15020
rect 18003 14980 18144 15008
rect 18003 14977 18015 14980
rect 17957 14971 18015 14977
rect 16132 14912 16344 14940
rect 9916 14900 9922 14912
rect 9876 14872 9904 14900
rect 11790 14872 11796 14884
rect 7116 14844 9904 14872
rect 10336 14844 11796 14872
rect 3878 14804 3884 14816
rect 3528 14776 3884 14804
rect 3878 14764 3884 14776
rect 3936 14804 3942 14816
rect 5552 14804 5580 14832
rect 10336 14816 10364 14844
rect 11790 14832 11796 14844
rect 11848 14832 11854 14884
rect 13078 14832 13084 14884
rect 13136 14872 13142 14884
rect 13648 14872 13676 14912
rect 16316 14884 16344 14912
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16632 14912 16773 14940
rect 16632 14900 16638 14912
rect 16761 14909 16773 14912
rect 16807 14909 16819 14943
rect 16960 14940 16988 14971
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 18322 14968 18328 15020
rect 18380 14968 18386 15020
rect 19444 15017 19472 15116
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 21726 15144 21732 15156
rect 20404 15116 21732 15144
rect 20404 15104 20410 15116
rect 19518 15036 19524 15088
rect 19576 15076 19582 15088
rect 19613 15079 19671 15085
rect 19613 15076 19625 15079
rect 19576 15048 19625 15076
rect 19576 15036 19582 15048
rect 19613 15045 19625 15048
rect 19659 15076 19671 15079
rect 19659 15048 19840 15076
rect 19659 15045 19671 15048
rect 19613 15039 19671 15045
rect 19245 15011 19303 15017
rect 19245 14977 19257 15011
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 16761 14903 16819 14909
rect 16868 14912 16988 14940
rect 17037 14943 17095 14949
rect 13136 14844 13676 14872
rect 13136 14832 13142 14844
rect 14090 14832 14096 14884
rect 14148 14832 14154 14884
rect 14734 14832 14740 14884
rect 14792 14872 14798 14884
rect 14792 14844 16252 14872
rect 14792 14832 14798 14844
rect 5718 14804 5724 14816
rect 3936 14776 5724 14804
rect 3936 14764 3942 14776
rect 5718 14764 5724 14776
rect 5776 14764 5782 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 8481 14807 8539 14813
rect 8481 14804 8493 14807
rect 7156 14776 8493 14804
rect 7156 14764 7162 14776
rect 8481 14773 8493 14776
rect 8527 14804 8539 14807
rect 8938 14804 8944 14816
rect 8527 14776 8944 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 10318 14764 10324 14816
rect 10376 14764 10382 14816
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11422 14804 11428 14816
rect 11103 14776 11428 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 12437 14807 12495 14813
rect 12437 14773 12449 14807
rect 12483 14804 12495 14807
rect 13446 14804 13452 14816
rect 12483 14776 13452 14804
rect 12483 14773 12495 14776
rect 12437 14767 12495 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 15102 14804 15108 14816
rect 13771 14776 15108 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15562 14764 15568 14816
rect 15620 14764 15626 14816
rect 16224 14804 16252 14844
rect 16298 14832 16304 14884
rect 16356 14872 16362 14884
rect 16868 14872 16896 14912
rect 17037 14909 17049 14943
rect 17083 14940 17095 14943
rect 17126 14940 17132 14952
rect 17083 14912 17132 14940
rect 17083 14909 17095 14912
rect 17037 14903 17095 14909
rect 17126 14900 17132 14912
rect 17184 14900 17190 14952
rect 17681 14943 17739 14949
rect 17681 14909 17693 14943
rect 17727 14909 17739 14943
rect 19260 14940 19288 14971
rect 19702 14968 19708 15020
rect 19760 14968 19766 15020
rect 19812 15017 19840 15048
rect 20456 15017 20484 15116
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 25498 15104 25504 15156
rect 25556 15144 25562 15156
rect 25777 15147 25835 15153
rect 25777 15144 25789 15147
rect 25556 15116 25789 15144
rect 25556 15104 25562 15116
rect 25777 15113 25789 15116
rect 25823 15113 25835 15147
rect 25777 15107 25835 15113
rect 26145 15147 26203 15153
rect 26145 15113 26157 15147
rect 26191 15144 26203 15147
rect 27522 15144 27528 15156
rect 26191 15116 27528 15144
rect 26191 15113 26203 15116
rect 26145 15107 26203 15113
rect 27522 15104 27528 15116
rect 27580 15104 27586 15156
rect 31389 15147 31447 15153
rect 31389 15113 31401 15147
rect 31435 15144 31447 15147
rect 31435 15116 31754 15144
rect 31435 15113 31447 15116
rect 31389 15107 31447 15113
rect 22738 15036 22744 15088
rect 22796 15076 22802 15088
rect 24964 15076 24992 15104
rect 26237 15079 26295 15085
rect 26237 15076 26249 15079
rect 22796 15048 23612 15076
rect 24964 15048 26249 15076
rect 22796 15036 22802 15048
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 14977 19855 15011
rect 19797 14971 19855 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 20530 14968 20536 15020
rect 20588 14968 20594 15020
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 15008 20775 15011
rect 20806 15008 20812 15020
rect 20763 14980 20812 15008
rect 20763 14977 20775 14980
rect 20717 14971 20775 14977
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 21082 14968 21088 15020
rect 21140 14968 21146 15020
rect 22830 14968 22836 15020
rect 22888 15008 22894 15020
rect 23014 15008 23020 15020
rect 22888 14980 23020 15008
rect 22888 14968 22894 14980
rect 23014 14968 23020 14980
rect 23072 14968 23078 15020
rect 23290 14968 23296 15020
rect 23348 15008 23354 15020
rect 23584 15017 23612 15048
rect 26237 15045 26249 15048
rect 26283 15045 26295 15079
rect 26237 15039 26295 15045
rect 28074 15036 28080 15088
rect 28132 15076 28138 15088
rect 28261 15079 28319 15085
rect 28261 15076 28273 15079
rect 28132 15048 28273 15076
rect 28132 15036 28138 15048
rect 28261 15045 28273 15048
rect 28307 15045 28319 15079
rect 28261 15039 28319 15045
rect 30098 15036 30104 15088
rect 30156 15076 30162 15088
rect 30745 15079 30803 15085
rect 30745 15076 30757 15079
rect 30156 15048 30757 15076
rect 30156 15036 30162 15048
rect 30745 15045 30757 15048
rect 30791 15045 30803 15079
rect 30745 15039 30803 15045
rect 30926 15036 30932 15088
rect 30984 15076 30990 15088
rect 31570 15076 31576 15088
rect 30984 15048 31576 15076
rect 30984 15036 30990 15048
rect 31570 15036 31576 15048
rect 31628 15036 31634 15088
rect 31726 15076 31754 15116
rect 31941 15079 31999 15085
rect 31941 15076 31953 15079
rect 31726 15048 31953 15076
rect 31941 15045 31953 15048
rect 31987 15045 31999 15079
rect 31941 15039 31999 15045
rect 33410 15036 33416 15088
rect 33468 15076 33474 15088
rect 33597 15079 33655 15085
rect 33597 15076 33609 15079
rect 33468 15048 33609 15076
rect 33468 15036 33474 15048
rect 33597 15045 33609 15048
rect 33643 15045 33655 15079
rect 33597 15039 33655 15045
rect 23477 15011 23535 15017
rect 23477 15008 23489 15011
rect 23348 14980 23489 15008
rect 23348 14968 23354 14980
rect 23477 14977 23489 14980
rect 23523 14977 23535 15011
rect 23477 14971 23535 14977
rect 23569 15011 23627 15017
rect 23569 14977 23581 15011
rect 23615 14977 23627 15011
rect 23569 14971 23627 14977
rect 28445 15011 28503 15017
rect 28445 14977 28457 15011
rect 28491 15008 28503 15011
rect 29362 15008 29368 15020
rect 28491 14980 29368 15008
rect 28491 14977 28503 14980
rect 28445 14971 28503 14977
rect 29362 14968 29368 14980
rect 29420 14968 29426 15020
rect 31202 14968 31208 15020
rect 31260 14968 31266 15020
rect 31662 14968 31668 15020
rect 31720 14968 31726 15020
rect 32858 14968 32864 15020
rect 32916 15008 32922 15020
rect 33229 15011 33287 15017
rect 33229 15008 33241 15011
rect 32916 14980 33241 15008
rect 32916 14968 32922 14980
rect 33229 14977 33241 14980
rect 33275 14977 33287 15011
rect 33229 14971 33287 14977
rect 34333 15011 34391 15017
rect 34333 14977 34345 15011
rect 34379 14977 34391 15011
rect 34333 14971 34391 14977
rect 19334 14940 19340 14952
rect 19260 14912 19340 14940
rect 17681 14903 17739 14909
rect 16356 14844 16896 14872
rect 16356 14832 16362 14844
rect 17586 14832 17592 14884
rect 17644 14872 17650 14884
rect 17696 14872 17724 14903
rect 19334 14900 19340 14912
rect 19392 14940 19398 14952
rect 20548 14940 20576 14968
rect 19392 14912 20576 14940
rect 21008 14940 21036 14968
rect 21542 14940 21548 14952
rect 21008 14912 21548 14940
rect 19392 14900 19398 14912
rect 21542 14900 21548 14912
rect 21600 14900 21606 14952
rect 22649 14943 22707 14949
rect 22649 14940 22661 14943
rect 21652 14912 22661 14940
rect 17644 14844 17724 14872
rect 17644 14832 17650 14844
rect 18414 14832 18420 14884
rect 18472 14872 18478 14884
rect 19150 14872 19156 14884
rect 18472 14844 19156 14872
rect 18472 14832 18478 14844
rect 19150 14832 19156 14844
rect 19208 14832 19214 14884
rect 20070 14832 20076 14884
rect 20128 14832 20134 14884
rect 20714 14832 20720 14884
rect 20772 14872 20778 14884
rect 21652 14872 21680 14912
rect 22649 14909 22661 14912
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 22922 14900 22928 14952
rect 22980 14940 22986 14952
rect 23201 14943 23259 14949
rect 23201 14940 23213 14943
rect 22980 14912 23213 14940
rect 22980 14900 22986 14912
rect 23201 14909 23213 14912
rect 23247 14909 23259 14943
rect 23201 14903 23259 14909
rect 25958 14900 25964 14952
rect 26016 14940 26022 14952
rect 26329 14943 26387 14949
rect 26329 14940 26341 14943
rect 26016 14912 26341 14940
rect 26016 14900 26022 14912
rect 26329 14909 26341 14912
rect 26375 14940 26387 14943
rect 27338 14940 27344 14952
rect 26375 14912 27344 14940
rect 26375 14909 26387 14912
rect 26329 14903 26387 14909
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 30742 14900 30748 14952
rect 30800 14940 30806 14952
rect 31021 14943 31079 14949
rect 31021 14940 31033 14943
rect 30800 14912 31033 14940
rect 30800 14900 30806 14912
rect 31021 14909 31033 14912
rect 31067 14909 31079 14943
rect 31021 14903 31079 14909
rect 31846 14900 31852 14952
rect 31904 14900 31910 14952
rect 34348 14872 34376 14971
rect 20772 14844 21680 14872
rect 22066 14844 34376 14872
rect 20772 14832 20778 14844
rect 22066 14804 22094 14844
rect 16224 14776 22094 14804
rect 28626 14764 28632 14816
rect 28684 14764 28690 14816
rect 31205 14807 31263 14813
rect 31205 14773 31217 14807
rect 31251 14804 31263 14807
rect 31294 14804 31300 14816
rect 31251 14776 31300 14804
rect 31251 14773 31263 14776
rect 31205 14767 31263 14773
rect 31294 14764 31300 14776
rect 31352 14764 31358 14816
rect 31478 14764 31484 14816
rect 31536 14764 31542 14816
rect 31846 14764 31852 14816
rect 31904 14764 31910 14816
rect 34146 14764 34152 14816
rect 34204 14764 34210 14816
rect 1104 14714 34684 14736
rect 1104 14662 5147 14714
rect 5199 14662 5211 14714
rect 5263 14662 5275 14714
rect 5327 14662 5339 14714
rect 5391 14662 5403 14714
rect 5455 14662 13541 14714
rect 13593 14662 13605 14714
rect 13657 14662 13669 14714
rect 13721 14662 13733 14714
rect 13785 14662 13797 14714
rect 13849 14662 21935 14714
rect 21987 14662 21999 14714
rect 22051 14662 22063 14714
rect 22115 14662 22127 14714
rect 22179 14662 22191 14714
rect 22243 14662 30329 14714
rect 30381 14662 30393 14714
rect 30445 14662 30457 14714
rect 30509 14662 30521 14714
rect 30573 14662 30585 14714
rect 30637 14662 34684 14714
rect 1104 14640 34684 14662
rect 7006 14560 7012 14612
rect 7064 14560 7070 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 10318 14600 10324 14612
rect 8904 14572 10324 14600
rect 8904 14560 8910 14572
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 12526 14600 12532 14612
rect 11020 14572 12532 14600
rect 11020 14560 11026 14572
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13449 14603 13507 14609
rect 13449 14569 13461 14603
rect 13495 14600 13507 14603
rect 14090 14600 14096 14612
rect 13495 14572 14096 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 15102 14560 15108 14612
rect 15160 14560 15166 14612
rect 15194 14560 15200 14612
rect 15252 14560 15258 14612
rect 16850 14560 16856 14612
rect 16908 14600 16914 14612
rect 16945 14603 17003 14609
rect 16945 14600 16957 14603
rect 16908 14572 16957 14600
rect 16908 14560 16914 14572
rect 16945 14569 16957 14572
rect 16991 14569 17003 14603
rect 16945 14563 17003 14569
rect 17126 14560 17132 14612
rect 17184 14560 17190 14612
rect 18322 14560 18328 14612
rect 18380 14560 18386 14612
rect 18509 14603 18567 14609
rect 18509 14569 18521 14603
rect 18555 14600 18567 14603
rect 19334 14600 19340 14612
rect 18555 14572 19340 14600
rect 18555 14569 18567 14572
rect 18509 14563 18567 14569
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 19978 14560 19984 14612
rect 20036 14560 20042 14612
rect 20993 14603 21051 14609
rect 20993 14569 21005 14603
rect 21039 14600 21051 14603
rect 21082 14600 21088 14612
rect 21039 14572 21088 14600
rect 21039 14569 21051 14572
rect 20993 14563 21051 14569
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 21468 14572 23520 14600
rect 3786 14492 3792 14544
rect 3844 14532 3850 14544
rect 4246 14532 4252 14544
rect 3844 14504 4252 14532
rect 3844 14492 3850 14504
rect 4246 14492 4252 14504
rect 4304 14532 4310 14544
rect 6178 14532 6184 14544
rect 4304 14504 6184 14532
rect 4304 14492 4310 14504
rect 6178 14492 6184 14504
rect 6236 14532 6242 14544
rect 7558 14532 7564 14544
rect 6236 14504 7564 14532
rect 6236 14492 6242 14504
rect 5905 14467 5963 14473
rect 5905 14433 5917 14467
rect 5951 14464 5963 14467
rect 5951 14436 6960 14464
rect 5951 14433 5963 14436
rect 5905 14427 5963 14433
rect 4706 14356 4712 14408
rect 4764 14356 4770 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 4856 14368 5181 14396
rect 4856 14356 4862 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 6273 14331 6331 14337
rect 6273 14297 6285 14331
rect 6319 14297 6331 14331
rect 6932 14328 6960 14436
rect 7208 14405 7236 14504
rect 7558 14492 7564 14504
rect 7616 14532 7622 14544
rect 9858 14532 9864 14544
rect 7616 14504 9864 14532
rect 7616 14492 7622 14504
rect 9858 14492 9864 14504
rect 9916 14492 9922 14544
rect 13078 14532 13084 14544
rect 9968 14504 13084 14532
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 7742 14464 7748 14476
rect 7423 14436 7748 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 7576 14408 7604 14436
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 9968 14408 9996 14504
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 13541 14535 13599 14541
rect 13541 14501 13553 14535
rect 13587 14501 13599 14535
rect 15120 14532 15148 14560
rect 16393 14535 16451 14541
rect 15120 14504 16252 14532
rect 13541 14495 13599 14501
rect 11146 14424 11152 14476
rect 11204 14464 11210 14476
rect 11333 14467 11391 14473
rect 11333 14464 11345 14467
rect 11204 14436 11345 14464
rect 11204 14424 11210 14436
rect 11333 14433 11345 14436
rect 11379 14433 11391 14467
rect 11333 14427 11391 14433
rect 11609 14467 11667 14473
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 12989 14467 13047 14473
rect 12989 14464 13001 14467
rect 11655 14436 13001 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 12989 14433 13001 14436
rect 13035 14433 13047 14467
rect 13556 14464 13584 14495
rect 16022 14464 16028 14476
rect 12989 14427 13047 14433
rect 13198 14436 13584 14464
rect 15488 14436 16028 14464
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 7282 14356 7288 14408
rect 7340 14356 7346 14408
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 7484 14328 7512 14359
rect 7558 14356 7564 14408
rect 7616 14356 7622 14408
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14396 7711 14399
rect 9122 14396 9128 14408
rect 7699 14368 9128 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11054 14396 11060 14408
rect 11011 14368 11060 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11238 14396 11244 14408
rect 11164 14368 11244 14396
rect 8110 14328 8116 14340
rect 6932 14300 8116 14328
rect 6273 14291 6331 14297
rect 4522 14220 4528 14272
rect 4580 14220 4586 14272
rect 4890 14220 4896 14272
rect 4948 14260 4954 14272
rect 5442 14260 5448 14272
rect 4948 14232 5448 14260
rect 4948 14220 4954 14232
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5810 14260 5816 14272
rect 5592 14232 5816 14260
rect 5592 14220 5598 14232
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6288 14260 6316 14291
rect 7208 14272 7236 14300
rect 8110 14288 8116 14300
rect 8168 14288 8174 14340
rect 8386 14288 8392 14340
rect 8444 14328 8450 14340
rect 9968 14328 9996 14356
rect 8444 14300 9996 14328
rect 8444 14288 8450 14300
rect 7006 14260 7012 14272
rect 6288 14232 7012 14260
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7190 14220 7196 14272
rect 7248 14220 7254 14272
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 10226 14260 10232 14272
rect 9180 14232 10232 14260
rect 9180 14220 9186 14232
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 11057 14263 11115 14269
rect 11057 14229 11069 14263
rect 11103 14260 11115 14263
rect 11164 14260 11192 14368
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 12434 14396 12440 14408
rect 11480 14368 12440 14396
rect 11480 14356 11486 14368
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 12713 14399 12771 14405
rect 12713 14396 12725 14399
rect 12584 14368 12725 14396
rect 12584 14356 12590 14368
rect 12713 14365 12725 14368
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14365 12955 14399
rect 12897 14359 12955 14365
rect 12912 14328 12940 14359
rect 13078 14356 13084 14408
rect 13136 14356 13142 14408
rect 13198 14328 13226 14436
rect 15488 14408 15516 14436
rect 16022 14424 16028 14436
rect 16080 14464 16086 14476
rect 16224 14464 16252 14504
rect 16393 14501 16405 14535
rect 16439 14532 16451 14535
rect 17144 14532 17172 14560
rect 16439 14504 17172 14532
rect 16439 14501 16451 14504
rect 16393 14495 16451 14501
rect 16850 14464 16856 14476
rect 16080 14436 16160 14464
rect 16224 14436 16856 14464
rect 16080 14424 16086 14436
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 12912 14300 13226 14328
rect 11103 14232 11192 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 11238 14220 11244 14272
rect 11296 14220 11302 14272
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 12066 14260 12072 14272
rect 11388 14232 12072 14260
rect 11388 14220 11394 14232
rect 12066 14220 12072 14232
rect 12124 14260 12130 14272
rect 13280 14260 13308 14359
rect 13446 14356 13452 14408
rect 13504 14396 13510 14408
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 13504 14368 13553 14396
rect 13504 14356 13510 14368
rect 13541 14365 13553 14368
rect 13587 14365 13599 14399
rect 13541 14359 13599 14365
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14396 13783 14399
rect 14274 14396 14280 14408
rect 13771 14368 14280 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 13630 14288 13636 14340
rect 13688 14328 13694 14340
rect 13740 14328 13768 14359
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 15378 14356 15384 14408
rect 15436 14356 15442 14408
rect 15470 14356 15476 14408
rect 15528 14356 15534 14408
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 15620 14368 15669 14396
rect 15620 14356 15626 14368
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 15746 14356 15752 14408
rect 15804 14356 15810 14408
rect 15838 14356 15844 14408
rect 15896 14356 15902 14408
rect 16132 14405 16160 14436
rect 16850 14424 16856 14436
rect 16908 14464 16914 14476
rect 17037 14467 17095 14473
rect 17037 14464 17049 14467
rect 16908 14436 17049 14464
rect 16908 14424 16914 14436
rect 17037 14433 17049 14436
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14365 15991 14399
rect 15933 14359 15991 14365
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 13688 14300 13768 14328
rect 13688 14288 13694 14300
rect 12124 14232 13308 14260
rect 12124 14220 12130 14232
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 14090 14260 14096 14272
rect 13412 14232 14096 14260
rect 13412 14220 13418 14232
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 15396 14260 15424 14356
rect 15764 14328 15792 14356
rect 15948 14328 15976 14359
rect 15764 14300 15976 14328
rect 15930 14260 15936 14272
rect 15396 14232 15936 14260
rect 15930 14220 15936 14232
rect 15988 14260 15994 14272
rect 16224 14260 16252 14359
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16356 14368 16957 14396
rect 16356 14356 16362 14368
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 18138 14356 18144 14408
rect 18196 14356 18202 14408
rect 18340 14405 18368 14560
rect 19429 14535 19487 14541
rect 19429 14532 19441 14535
rect 19260 14504 19441 14532
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 17586 14328 17592 14340
rect 17328 14300 17592 14328
rect 17328 14269 17356 14300
rect 17586 14288 17592 14300
rect 17644 14328 17650 14340
rect 18049 14331 18107 14337
rect 18049 14328 18061 14331
rect 17644 14300 18061 14328
rect 17644 14288 17650 14300
rect 18049 14297 18061 14300
rect 18095 14297 18107 14331
rect 18049 14291 18107 14297
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19260 14328 19288 14504
rect 19429 14501 19441 14504
rect 19475 14501 19487 14535
rect 19429 14495 19487 14501
rect 19517 14535 19575 14541
rect 19517 14501 19529 14535
rect 19563 14532 19575 14535
rect 19563 14504 20392 14532
rect 19563 14501 19575 14504
rect 19517 14495 19575 14501
rect 20364 14464 20392 14504
rect 20622 14464 20628 14476
rect 19352 14436 19748 14464
rect 19352 14405 19380 14436
rect 19720 14408 19748 14436
rect 20364 14436 20628 14464
rect 20364 14408 20392 14436
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 19337 14399 19395 14405
rect 19337 14365 19349 14399
rect 19383 14365 19395 14399
rect 19337 14359 19395 14365
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19484 14368 19625 14396
rect 19484 14356 19490 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20165 14399 20223 14405
rect 20165 14396 20177 14399
rect 19760 14368 20177 14396
rect 19760 14356 19766 14368
rect 20165 14365 20177 14368
rect 20211 14365 20223 14399
rect 20165 14359 20223 14365
rect 20346 14356 20352 14408
rect 20404 14356 20410 14408
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 20809 14399 20867 14405
rect 20809 14396 20821 14399
rect 20487 14368 20821 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 20254 14328 20260 14340
rect 19208 14300 20260 14328
rect 19208 14288 19214 14300
rect 20254 14288 20260 14300
rect 20312 14288 20318 14340
rect 20548 14272 20576 14368
rect 20809 14365 20821 14368
rect 20855 14365 20867 14399
rect 21100 14396 21128 14560
rect 21174 14492 21180 14544
rect 21232 14492 21238 14544
rect 21192 14464 21220 14492
rect 21468 14464 21496 14572
rect 23385 14535 23443 14541
rect 23385 14501 23397 14535
rect 23431 14501 23443 14535
rect 23385 14495 23443 14501
rect 21192 14436 21496 14464
rect 21468 14408 21496 14436
rect 21637 14467 21695 14473
rect 21637 14433 21649 14467
rect 21683 14464 21695 14467
rect 21818 14464 21824 14476
rect 21683 14436 21824 14464
rect 21683 14433 21695 14436
rect 21637 14427 21695 14433
rect 21818 14424 21824 14436
rect 21876 14424 21882 14476
rect 23014 14464 23020 14476
rect 21928 14436 23020 14464
rect 21177 14399 21235 14405
rect 21177 14396 21189 14399
rect 21100 14368 21189 14396
rect 20809 14359 20867 14365
rect 21177 14365 21189 14368
rect 21223 14365 21235 14399
rect 21177 14359 21235 14365
rect 21450 14356 21456 14408
rect 21508 14356 21514 14408
rect 21928 14405 21956 14436
rect 23014 14424 23020 14436
rect 23072 14464 23078 14476
rect 23400 14464 23428 14495
rect 23072 14436 23428 14464
rect 23072 14424 23078 14436
rect 21729 14399 21787 14405
rect 21729 14365 21741 14399
rect 21775 14365 21787 14399
rect 21729 14359 21787 14365
rect 21913 14399 21971 14405
rect 21913 14365 21925 14399
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 21634 14328 21640 14340
rect 20824 14300 21640 14328
rect 20824 14272 20852 14300
rect 21634 14288 21640 14300
rect 21692 14328 21698 14340
rect 21744 14328 21772 14359
rect 22738 14356 22744 14408
rect 22796 14356 22802 14408
rect 22922 14356 22928 14408
rect 22980 14356 22986 14408
rect 23216 14405 23244 14436
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 23290 14356 23296 14408
rect 23348 14356 23354 14408
rect 23492 14405 23520 14572
rect 29362 14560 29368 14612
rect 29420 14560 29426 14612
rect 31205 14603 31263 14609
rect 31205 14569 31217 14603
rect 31251 14600 31263 14603
rect 32214 14600 32220 14612
rect 31251 14572 32220 14600
rect 31251 14569 31263 14572
rect 31205 14563 31263 14569
rect 32214 14560 32220 14572
rect 32272 14560 32278 14612
rect 34241 14603 34299 14609
rect 34241 14569 34253 14603
rect 34287 14600 34299 14603
rect 34287 14572 34744 14600
rect 34287 14569 34299 14572
rect 34241 14563 34299 14569
rect 34716 14544 34744 14572
rect 23952 14504 26188 14532
rect 23477 14399 23535 14405
rect 23477 14365 23489 14399
rect 23523 14365 23535 14399
rect 23477 14359 23535 14365
rect 21692 14300 21772 14328
rect 23109 14331 23167 14337
rect 21692 14288 21698 14300
rect 23109 14297 23121 14331
rect 23155 14328 23167 14331
rect 23952 14328 23980 14504
rect 25958 14424 25964 14476
rect 26016 14424 26022 14476
rect 26160 14473 26188 14504
rect 26878 14492 26884 14544
rect 26936 14492 26942 14544
rect 31938 14492 31944 14544
rect 31996 14492 32002 14544
rect 32493 14535 32551 14541
rect 32493 14501 32505 14535
rect 32539 14501 32551 14535
rect 32493 14495 32551 14501
rect 26145 14467 26203 14473
rect 26145 14433 26157 14467
rect 26191 14433 26203 14467
rect 26896 14464 26924 14492
rect 27614 14464 27620 14476
rect 26896 14436 27620 14464
rect 26145 14427 26203 14433
rect 27614 14424 27620 14436
rect 27672 14424 27678 14476
rect 25682 14356 25688 14408
rect 25740 14396 25746 14408
rect 26881 14399 26939 14405
rect 26881 14396 26893 14399
rect 25740 14368 26893 14396
rect 25740 14356 25746 14368
rect 26881 14365 26893 14368
rect 26927 14365 26939 14399
rect 26881 14359 26939 14365
rect 31205 14399 31263 14405
rect 31205 14365 31217 14399
rect 31251 14396 31263 14399
rect 31386 14396 31392 14408
rect 31251 14368 31392 14396
rect 31251 14365 31263 14368
rect 31205 14359 31263 14365
rect 31386 14356 31392 14368
rect 31444 14356 31450 14408
rect 31481 14399 31539 14405
rect 31481 14365 31493 14399
rect 31527 14365 31539 14399
rect 31481 14359 31539 14365
rect 31757 14399 31815 14405
rect 31757 14365 31769 14399
rect 31803 14396 31815 14399
rect 31956 14396 31984 14492
rect 32508 14464 32536 14495
rect 34698 14492 34704 14544
rect 34756 14492 34762 14544
rect 32140 14436 32536 14464
rect 32140 14405 32168 14436
rect 31803 14368 31984 14396
rect 32125 14399 32183 14405
rect 31803 14365 31815 14368
rect 31757 14359 31815 14365
rect 32125 14365 32137 14399
rect 32171 14365 32183 14399
rect 32125 14359 32183 14365
rect 32217 14399 32275 14405
rect 32217 14365 32229 14399
rect 32263 14365 32275 14399
rect 32217 14359 32275 14365
rect 32493 14399 32551 14405
rect 32493 14365 32505 14399
rect 32539 14396 32551 14399
rect 32858 14396 32864 14408
rect 32539 14368 32864 14396
rect 32539 14365 32551 14368
rect 32493 14359 32551 14365
rect 27522 14328 27528 14340
rect 23155 14300 23980 14328
rect 26068 14300 27528 14328
rect 23155 14297 23167 14300
rect 23109 14291 23167 14297
rect 15988 14232 16252 14260
rect 17313 14263 17371 14269
rect 15988 14220 15994 14232
rect 17313 14229 17325 14263
rect 17359 14229 17371 14263
rect 17313 14223 17371 14229
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 19797 14263 19855 14269
rect 19797 14260 19809 14263
rect 18472 14232 19809 14260
rect 18472 14220 18478 14232
rect 19797 14229 19809 14232
rect 19843 14260 19855 14263
rect 19886 14260 19892 14272
rect 19843 14232 19892 14260
rect 19843 14229 19855 14232
rect 19797 14223 19855 14229
rect 19886 14220 19892 14232
rect 19944 14220 19950 14272
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20806 14220 20812 14272
rect 20864 14220 20870 14272
rect 22554 14220 22560 14272
rect 22612 14260 22618 14272
rect 23124 14260 23152 14291
rect 26068 14272 26096 14300
rect 27522 14288 27528 14300
rect 27580 14288 27586 14340
rect 27890 14288 27896 14340
rect 27948 14288 27954 14340
rect 29362 14328 29368 14340
rect 29118 14300 29368 14328
rect 29362 14288 29368 14300
rect 29420 14288 29426 14340
rect 31110 14288 31116 14340
rect 31168 14328 31174 14340
rect 31496 14328 31524 14359
rect 31168 14300 31432 14328
rect 31496 14300 31754 14328
rect 31168 14288 31174 14300
rect 22612 14232 23152 14260
rect 22612 14220 22618 14232
rect 26050 14220 26056 14272
rect 26108 14220 26114 14272
rect 26237 14263 26295 14269
rect 26237 14229 26249 14263
rect 26283 14260 26295 14263
rect 26510 14260 26516 14272
rect 26283 14232 26516 14260
rect 26283 14229 26295 14232
rect 26237 14223 26295 14229
rect 26510 14220 26516 14232
rect 26568 14220 26574 14272
rect 26602 14220 26608 14272
rect 26660 14220 26666 14272
rect 31404 14269 31432 14300
rect 31389 14263 31447 14269
rect 31389 14229 31401 14263
rect 31435 14229 31447 14263
rect 31389 14223 31447 14229
rect 31570 14220 31576 14272
rect 31628 14220 31634 14272
rect 31726 14260 31754 14300
rect 31846 14288 31852 14340
rect 31904 14288 31910 14340
rect 31938 14288 31944 14340
rect 31996 14288 32002 14340
rect 32232 14272 32260 14359
rect 32858 14356 32864 14368
rect 32916 14356 32922 14408
rect 34057 14399 34115 14405
rect 34057 14365 34069 14399
rect 34103 14396 34115 14399
rect 34146 14396 34152 14408
rect 34103 14368 34152 14396
rect 34103 14365 34115 14368
rect 34057 14359 34115 14365
rect 34146 14356 34152 14368
rect 34204 14356 34210 14408
rect 32214 14260 32220 14272
rect 31726 14232 32220 14260
rect 32214 14220 32220 14232
rect 32272 14220 32278 14272
rect 32306 14220 32312 14272
rect 32364 14220 32370 14272
rect 1104 14170 34840 14192
rect 1104 14118 9344 14170
rect 9396 14118 9408 14170
rect 9460 14118 9472 14170
rect 9524 14118 9536 14170
rect 9588 14118 9600 14170
rect 9652 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 17930 14170
rect 17982 14118 17994 14170
rect 18046 14118 26132 14170
rect 26184 14118 26196 14170
rect 26248 14118 26260 14170
rect 26312 14118 26324 14170
rect 26376 14118 26388 14170
rect 26440 14118 34526 14170
rect 34578 14118 34590 14170
rect 34642 14118 34654 14170
rect 34706 14118 34718 14170
rect 34770 14118 34782 14170
rect 34834 14118 34840 14170
rect 1104 14096 34840 14118
rect 3970 14016 3976 14068
rect 4028 14016 4034 14068
rect 4614 14016 4620 14068
rect 4672 14056 4678 14068
rect 4893 14059 4951 14065
rect 4893 14056 4905 14059
rect 4672 14028 4905 14056
rect 4672 14016 4678 14028
rect 4893 14025 4905 14028
rect 4939 14025 4951 14059
rect 4893 14019 4951 14025
rect 5442 14016 5448 14068
rect 5500 14016 5506 14068
rect 6667 14059 6725 14065
rect 6667 14056 6679 14059
rect 5920 14028 6679 14056
rect 3878 13948 3884 14000
rect 3936 13948 3942 14000
rect 3988 13988 4016 14016
rect 4341 13991 4399 13997
rect 3988 13960 4292 13988
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3421 13923 3479 13929
rect 3421 13920 3433 13923
rect 3384 13892 3433 13920
rect 3384 13880 3390 13892
rect 3421 13889 3433 13892
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 3602 13880 3608 13932
rect 3660 13920 3666 13932
rect 3896 13920 3924 13948
rect 4264 13929 4292 13960
rect 4341 13957 4353 13991
rect 4387 13988 4399 13991
rect 5810 13988 5816 14000
rect 4387 13960 5816 13988
rect 4387 13957 4399 13960
rect 4341 13951 4399 13957
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3660 13892 3985 13920
rect 3660 13880 3666 13892
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 4525 13883 4583 13889
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13852 3755 13855
rect 3786 13852 3792 13864
rect 3743 13824 3792 13852
rect 3743 13821 3755 13824
rect 3697 13815 3755 13821
rect 3786 13812 3792 13824
rect 3844 13812 3850 13864
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13821 4123 13855
rect 4065 13815 4123 13821
rect 4540 13852 4568 13883
rect 4614 13880 4620 13932
rect 4672 13880 4678 13932
rect 4706 13880 4712 13932
rect 4764 13920 4770 13932
rect 5184 13929 5212 13960
rect 5810 13948 5816 13960
rect 5868 13948 5874 14000
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4764 13892 5089 13920
rect 4764 13880 4770 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13920 5595 13923
rect 5718 13920 5724 13932
rect 5583 13892 5724 13920
rect 5583 13889 5595 13892
rect 5537 13883 5595 13889
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 4540 13824 5304 13852
rect 4080 13784 4108 13815
rect 4540 13784 4568 13824
rect 4080 13756 4568 13784
rect 5276 13784 5304 13824
rect 5626 13812 5632 13864
rect 5684 13812 5690 13864
rect 5920 13852 5948 14028
rect 6667 14025 6679 14028
rect 6713 14056 6725 14059
rect 7282 14056 7288 14068
rect 6713 14028 7288 14056
rect 6713 14025 6725 14028
rect 6667 14019 6725 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 7374 14016 7380 14068
rect 7432 14056 7438 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 7432 14028 8217 14056
rect 7432 14016 7438 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 8205 14019 8263 14025
rect 9858 14016 9864 14068
rect 9916 14056 9922 14068
rect 10321 14059 10379 14065
rect 9916 14028 10272 14056
rect 9916 14016 9922 14028
rect 10244 14000 10272 14028
rect 10321 14025 10333 14059
rect 10367 14056 10379 14059
rect 10410 14056 10416 14068
rect 10367 14028 10416 14056
rect 10367 14025 10379 14028
rect 10321 14019 10379 14025
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 10520 14028 10916 14056
rect 6457 13991 6515 13997
rect 6457 13957 6469 13991
rect 6503 13988 6515 13991
rect 6546 13988 6552 14000
rect 6503 13960 6552 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 6546 13948 6552 13960
rect 6604 13948 6610 14000
rect 7006 13988 7012 14000
rect 6840 13960 7012 13988
rect 6840 13920 6868 13960
rect 7006 13948 7012 13960
rect 7064 13988 7070 14000
rect 7064 13960 10088 13988
rect 7064 13948 7070 13960
rect 9646 13932 9674 13960
rect 5736 13824 5948 13852
rect 6012 13892 6868 13920
rect 6917 13923 6975 13929
rect 5736 13784 5764 13824
rect 5276 13756 5764 13784
rect 5905 13787 5963 13793
rect 4338 13676 4344 13728
rect 4396 13716 4402 13728
rect 4525 13719 4583 13725
rect 4525 13716 4537 13719
rect 4396 13688 4537 13716
rect 4396 13676 4402 13688
rect 4525 13685 4537 13688
rect 4571 13716 4583 13719
rect 5074 13716 5080 13728
rect 4571 13688 5080 13716
rect 4571 13685 4583 13688
rect 4525 13679 4583 13685
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 5276 13725 5304 13756
rect 5905 13753 5917 13787
rect 5951 13784 5963 13787
rect 6012 13784 6040 13892
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6932 13852 6960 13883
rect 7098 13880 7104 13932
rect 7156 13880 7162 13932
rect 8386 13880 8392 13932
rect 8444 13880 8450 13932
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13920 8631 13923
rect 8941 13923 8999 13929
rect 8619 13892 8800 13920
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 6144 13824 6960 13852
rect 6144 13812 6150 13824
rect 5951 13756 6040 13784
rect 5951 13753 5963 13756
rect 5905 13747 5963 13753
rect 5261 13719 5319 13725
rect 5261 13685 5273 13719
rect 5307 13685 5319 13719
rect 5261 13679 5319 13685
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 5537 13719 5595 13725
rect 5537 13716 5549 13719
rect 5408 13688 5549 13716
rect 5408 13676 5414 13688
rect 5537 13685 5549 13688
rect 5583 13716 5595 13719
rect 5994 13716 6000 13728
rect 5583 13688 6000 13716
rect 5583 13685 5595 13688
rect 5537 13679 5595 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 6656 13725 6684 13824
rect 7006 13812 7012 13864
rect 7064 13812 7070 13864
rect 8662 13812 8668 13864
rect 8720 13812 8726 13864
rect 8772 13861 8800 13892
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9490 13920 9496 13932
rect 8987 13892 9496 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9646 13890 9680 13932
rect 9674 13880 9680 13890
rect 9732 13880 9738 13932
rect 9766 13880 9772 13932
rect 9824 13880 9830 13932
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 9953 13923 10011 13929
rect 9953 13920 9965 13923
rect 9916 13892 9965 13920
rect 9916 13880 9922 13892
rect 9953 13889 9965 13892
rect 9999 13889 10011 13923
rect 10060 13920 10088 13960
rect 10226 13948 10232 14000
rect 10284 13988 10290 14000
rect 10520 13988 10548 14028
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 10284 13960 10548 13988
rect 10612 13960 10793 13988
rect 10284 13948 10290 13960
rect 10612 13929 10640 13960
rect 10781 13957 10793 13960
rect 10827 13957 10839 13991
rect 10781 13951 10839 13957
rect 10597 13923 10655 13929
rect 10060 13892 10548 13920
rect 9953 13883 10011 13889
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 9030 13812 9036 13864
rect 9088 13812 9094 13864
rect 9122 13812 9128 13864
rect 9180 13812 9186 13864
rect 9214 13812 9220 13864
rect 9272 13812 9278 13864
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 9398 13784 9404 13796
rect 6840 13756 9404 13784
rect 6840 13725 6868 13756
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 9858 13744 9864 13796
rect 9916 13744 9922 13796
rect 10152 13784 10180 13815
rect 10318 13812 10324 13864
rect 10376 13812 10382 13864
rect 10520 13852 10548 13892
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 10704 13852 10732 13883
rect 10520 13824 10732 13852
rect 10888 13852 10916 14028
rect 11606 14016 11612 14068
rect 11664 14016 11670 14068
rect 12897 14059 12955 14065
rect 12897 14025 12909 14059
rect 12943 14056 12955 14059
rect 13078 14056 13084 14068
rect 12943 14028 13084 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13170 14016 13176 14068
rect 13228 14016 13234 14068
rect 15289 14059 15347 14065
rect 15289 14025 15301 14059
rect 15335 14056 15347 14059
rect 16666 14056 16672 14068
rect 15335 14028 16672 14056
rect 15335 14025 15347 14028
rect 15289 14019 15347 14025
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 18877 14059 18935 14065
rect 18064 14028 18644 14056
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13920 11575 13923
rect 11624 13920 11652 14016
rect 13188 13988 13216 14016
rect 13096 13960 13216 13988
rect 11563 13892 11652 13920
rect 11563 13889 11575 13892
rect 11517 13883 11575 13889
rect 12986 13880 12992 13932
rect 13044 13880 13050 13932
rect 13096 13929 13124 13960
rect 13354 13948 13360 14000
rect 13412 13988 13418 14000
rect 13630 13988 13636 14000
rect 13412 13960 13636 13988
rect 13412 13948 13418 13960
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 15378 13948 15384 14000
rect 15436 13948 15442 14000
rect 15657 13991 15715 13997
rect 15657 13957 15669 13991
rect 15703 13988 15715 13991
rect 16117 13991 16175 13997
rect 16117 13988 16129 13991
rect 15703 13960 16129 13988
rect 15703 13957 15715 13960
rect 15657 13951 15715 13957
rect 16117 13957 16129 13960
rect 16163 13957 16175 13991
rect 16117 13951 16175 13957
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 13372 13920 13400 13948
rect 13311 13892 13400 13920
rect 13725 13923 13783 13929
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 11609 13855 11667 13861
rect 11609 13852 11621 13855
rect 10888 13824 11621 13852
rect 11609 13821 11621 13824
rect 11655 13821 11667 13855
rect 13004 13852 13032 13880
rect 13173 13855 13231 13861
rect 13173 13852 13185 13855
rect 11609 13815 11667 13821
rect 12406 13824 13185 13852
rect 11885 13787 11943 13793
rect 10152 13756 10824 13784
rect 10796 13728 10824 13756
rect 11885 13753 11897 13787
rect 11931 13784 11943 13787
rect 12158 13784 12164 13796
rect 11931 13756 12164 13784
rect 11931 13753 11943 13756
rect 11885 13747 11943 13753
rect 12158 13744 12164 13756
rect 12216 13784 12222 13796
rect 12406 13784 12434 13824
rect 13173 13821 13185 13824
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 12216 13756 12434 13784
rect 12216 13744 12222 13756
rect 12710 13744 12716 13796
rect 12768 13784 12774 13796
rect 13740 13784 13768 13883
rect 13814 13880 13820 13932
rect 13872 13880 13878 13932
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13964 13892 14013 13920
rect 13964 13880 13970 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13920 14151 13923
rect 14182 13920 14188 13932
rect 14139 13892 14188 13920
rect 14139 13889 14151 13892
rect 14093 13883 14151 13889
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 15286 13880 15292 13932
rect 15344 13880 15350 13932
rect 15396 13920 15424 13948
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 15396 13892 15485 13920
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 15304 13852 15332 13880
rect 15580 13852 15608 13883
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15804 13892 15853 13920
rect 15804 13880 15810 13892
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 15304 13824 15608 13852
rect 15948 13852 15976 13883
rect 16022 13880 16028 13932
rect 16080 13880 16086 13932
rect 18064 13929 18092 14028
rect 18138 13948 18144 14000
rect 18196 13988 18202 14000
rect 18616 13988 18644 14028
rect 18877 14025 18889 14059
rect 18923 14056 18935 14059
rect 20714 14056 20720 14068
rect 18923 14028 20720 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 24118 14016 24124 14068
rect 24176 14016 24182 14068
rect 25682 14016 25688 14068
rect 25740 14016 25746 14068
rect 26602 14016 26608 14068
rect 26660 14056 26666 14068
rect 26660 14028 27016 14056
rect 26660 14016 26666 14028
rect 24136 13988 24164 14016
rect 25590 13988 25596 14000
rect 18196 13960 18552 13988
rect 18616 13960 19288 13988
rect 18196 13948 18202 13960
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13920 18291 13923
rect 18322 13920 18328 13932
rect 18279 13892 18328 13920
rect 18279 13889 18291 13892
rect 18233 13883 18291 13889
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 18414 13880 18420 13932
rect 18472 13880 18478 13932
rect 16298 13852 16304 13864
rect 15948 13824 16304 13852
rect 12768 13756 13768 13784
rect 15580 13784 15608 13824
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 18524 13861 18552 13960
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13920 18659 13923
rect 18647 13892 18920 13920
rect 18647 13889 18659 13892
rect 18601 13883 18659 13889
rect 18141 13855 18199 13861
rect 18141 13821 18153 13855
rect 18187 13852 18199 13855
rect 18509 13855 18567 13861
rect 18187 13824 18368 13852
rect 18187 13821 18199 13824
rect 18141 13815 18199 13821
rect 16022 13784 16028 13796
rect 15580 13756 16028 13784
rect 12768 13744 12774 13756
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 18340 13784 18368 13824
rect 18509 13821 18521 13855
rect 18555 13821 18567 13855
rect 18693 13855 18751 13861
rect 18693 13852 18705 13855
rect 18509 13815 18567 13821
rect 18616 13824 18705 13852
rect 18616 13784 18644 13824
rect 18693 13821 18705 13824
rect 18739 13821 18751 13855
rect 18693 13815 18751 13821
rect 18340 13756 18644 13784
rect 18892 13784 18920 13892
rect 19150 13880 19156 13932
rect 19208 13880 19214 13932
rect 19260 13929 19288 13960
rect 20548 13960 21772 13988
rect 20548 13932 20576 13960
rect 19245 13923 19303 13929
rect 19245 13889 19257 13923
rect 19291 13920 19303 13923
rect 20346 13920 20352 13932
rect 19291 13892 20352 13920
rect 19291 13889 19303 13892
rect 19245 13883 19303 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 20530 13880 20536 13932
rect 20588 13880 20594 13932
rect 20717 13923 20775 13929
rect 20717 13889 20729 13923
rect 20763 13920 20775 13923
rect 20806 13920 20812 13932
rect 20763 13892 20812 13920
rect 20763 13889 20775 13892
rect 20717 13883 20775 13889
rect 20806 13880 20812 13892
rect 20864 13880 20870 13932
rect 21744 13864 21772 13960
rect 23952 13960 24164 13988
rect 25438 13960 25596 13988
rect 23658 13880 23664 13932
rect 23716 13880 23722 13932
rect 23952 13929 23980 13960
rect 25590 13948 25596 13960
rect 25648 13948 25654 14000
rect 26510 13948 26516 14000
rect 26568 13988 26574 14000
rect 26697 13991 26755 13997
rect 26697 13988 26709 13991
rect 26568 13960 26709 13988
rect 26568 13948 26574 13960
rect 26697 13957 26709 13960
rect 26743 13988 26755 13991
rect 26878 13988 26884 14000
rect 26743 13960 26884 13988
rect 26743 13957 26755 13960
rect 26697 13951 26755 13957
rect 26878 13948 26884 13960
rect 26936 13948 26942 14000
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 25498 13880 25504 13932
rect 25556 13920 25562 13932
rect 26988 13929 27016 14028
rect 27522 14016 27528 14068
rect 27580 14016 27586 14068
rect 27890 14016 27896 14068
rect 27948 14016 27954 14068
rect 30653 14059 30711 14065
rect 30653 14025 30665 14059
rect 30699 14056 30711 14059
rect 31110 14056 31116 14068
rect 30699 14028 31116 14056
rect 30699 14025 30711 14028
rect 30653 14019 30711 14025
rect 31110 14016 31116 14028
rect 31168 14016 31174 14068
rect 31938 14016 31944 14068
rect 31996 14056 32002 14068
rect 32125 14059 32183 14065
rect 32125 14056 32137 14059
rect 31996 14028 32137 14056
rect 31996 14016 32002 14028
rect 32125 14025 32137 14028
rect 32171 14025 32183 14059
rect 32125 14019 32183 14025
rect 25869 13923 25927 13929
rect 25869 13920 25881 13923
rect 25556 13892 25881 13920
rect 25556 13880 25562 13892
rect 25869 13889 25881 13892
rect 25915 13889 25927 13923
rect 25869 13883 25927 13889
rect 26973 13923 27031 13929
rect 26973 13889 26985 13923
rect 27019 13889 27031 13923
rect 27540 13920 27568 14016
rect 31389 13991 31447 13997
rect 28184 13960 30236 13988
rect 28077 13923 28135 13929
rect 28077 13920 28089 13923
rect 27540 13892 28089 13920
rect 26973 13883 27031 13889
rect 28077 13889 28089 13892
rect 28123 13889 28135 13923
rect 28077 13883 28135 13889
rect 18969 13855 19027 13861
rect 18969 13821 18981 13855
rect 19015 13852 19027 13855
rect 19426 13852 19432 13864
rect 19015 13824 19432 13852
rect 19015 13821 19027 13824
rect 18969 13815 19027 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 21726 13812 21732 13864
rect 21784 13812 21790 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23860 13824 24225 13852
rect 19061 13787 19119 13793
rect 19061 13784 19073 13787
rect 18892 13756 19073 13784
rect 19061 13753 19073 13756
rect 19107 13753 19119 13787
rect 19061 13747 19119 13753
rect 21450 13744 21456 13796
rect 21508 13784 21514 13796
rect 22922 13784 22928 13796
rect 21508 13756 22928 13784
rect 21508 13744 21514 13756
rect 22922 13744 22928 13756
rect 22980 13744 22986 13796
rect 23860 13793 23888 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 26694 13812 26700 13864
rect 26752 13852 26758 13864
rect 28184 13852 28212 13960
rect 28350 13880 28356 13932
rect 28408 13880 28414 13932
rect 28445 13923 28503 13929
rect 28445 13889 28457 13923
rect 28491 13889 28503 13923
rect 28445 13883 28503 13889
rect 26752 13824 28212 13852
rect 28261 13855 28319 13861
rect 26752 13812 26758 13824
rect 28261 13821 28273 13855
rect 28307 13821 28319 13855
rect 28460 13852 28488 13883
rect 28626 13880 28632 13932
rect 28684 13880 28690 13932
rect 30208 13929 30236 13960
rect 31389 13957 31401 13991
rect 31435 13988 31447 13991
rect 32306 13988 32312 14000
rect 31435 13960 32312 13988
rect 31435 13957 31447 13960
rect 31389 13951 31447 13957
rect 32306 13948 32312 13960
rect 32364 13948 32370 14000
rect 30193 13923 30251 13929
rect 30193 13889 30205 13923
rect 30239 13920 30251 13923
rect 30650 13920 30656 13932
rect 30239 13892 30656 13920
rect 30239 13889 30251 13892
rect 30193 13883 30251 13889
rect 30650 13880 30656 13892
rect 30708 13880 30714 13932
rect 31110 13880 31116 13932
rect 31168 13920 31174 13932
rect 31297 13923 31355 13929
rect 31297 13920 31309 13923
rect 31168 13892 31309 13920
rect 31168 13880 31174 13892
rect 31297 13889 31309 13892
rect 31343 13889 31355 13923
rect 31297 13883 31355 13889
rect 31478 13880 31484 13932
rect 31536 13880 31542 13932
rect 31570 13880 31576 13932
rect 31628 13880 31634 13932
rect 31938 13880 31944 13932
rect 31996 13920 32002 13932
rect 32214 13920 32220 13932
rect 31996 13892 32220 13920
rect 31996 13880 32002 13892
rect 32214 13880 32220 13892
rect 32272 13920 32278 13932
rect 32493 13923 32551 13929
rect 32493 13920 32505 13923
rect 32272 13892 32505 13920
rect 32272 13880 32278 13892
rect 32493 13889 32505 13892
rect 32539 13889 32551 13923
rect 32493 13883 32551 13889
rect 31588 13852 31616 13880
rect 28460 13824 31616 13852
rect 28261 13815 28319 13821
rect 23845 13787 23903 13793
rect 23845 13753 23857 13787
rect 23891 13753 23903 13787
rect 23845 13747 23903 13753
rect 27982 13744 27988 13796
rect 28040 13784 28046 13796
rect 28276 13784 28304 13815
rect 28810 13784 28816 13796
rect 28040 13756 28816 13784
rect 28040 13744 28046 13756
rect 28810 13744 28816 13756
rect 28868 13744 28874 13796
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13685 6699 13719
rect 6641 13679 6699 13685
rect 6825 13719 6883 13725
rect 6825 13685 6837 13719
rect 6871 13685 6883 13719
rect 6825 13679 6883 13685
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 10505 13719 10563 13725
rect 10505 13716 10517 13719
rect 8904 13688 10517 13716
rect 8904 13676 8910 13688
rect 10505 13685 10517 13688
rect 10551 13685 10563 13719
rect 10505 13679 10563 13685
rect 10778 13676 10784 13728
rect 10836 13676 10842 13728
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 11517 13719 11575 13725
rect 11517 13716 11529 13719
rect 10928 13688 11529 13716
rect 10928 13676 10934 13688
rect 11517 13685 11529 13688
rect 11563 13685 11575 13719
rect 11517 13679 11575 13685
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 12952 13688 13553 13716
rect 12952 13676 12958 13688
rect 13541 13685 13553 13688
rect 13587 13685 13599 13719
rect 13541 13679 13599 13685
rect 27157 13719 27215 13725
rect 27157 13685 27169 13719
rect 27203 13716 27215 13719
rect 27246 13716 27252 13728
rect 27203 13688 27252 13716
rect 27203 13685 27215 13688
rect 27157 13679 27215 13685
rect 27246 13676 27252 13688
rect 27304 13676 27310 13728
rect 30190 13676 30196 13728
rect 30248 13716 30254 13728
rect 30285 13719 30343 13725
rect 30285 13716 30297 13719
rect 30248 13688 30297 13716
rect 30248 13676 30254 13688
rect 30285 13685 30297 13688
rect 30331 13716 30343 13719
rect 31846 13716 31852 13728
rect 30331 13688 31852 13716
rect 30331 13685 30343 13688
rect 30285 13679 30343 13685
rect 31846 13676 31852 13688
rect 31904 13676 31910 13728
rect 1104 13626 34684 13648
rect 1104 13574 5147 13626
rect 5199 13574 5211 13626
rect 5263 13574 5275 13626
rect 5327 13574 5339 13626
rect 5391 13574 5403 13626
rect 5455 13574 13541 13626
rect 13593 13574 13605 13626
rect 13657 13574 13669 13626
rect 13721 13574 13733 13626
rect 13785 13574 13797 13626
rect 13849 13574 21935 13626
rect 21987 13574 21999 13626
rect 22051 13574 22063 13626
rect 22115 13574 22127 13626
rect 22179 13574 22191 13626
rect 22243 13574 30329 13626
rect 30381 13574 30393 13626
rect 30445 13574 30457 13626
rect 30509 13574 30521 13626
rect 30573 13574 30585 13626
rect 30637 13574 34684 13626
rect 1104 13552 34684 13574
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13512 4215 13515
rect 4706 13512 4712 13524
rect 4203 13484 4712 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 7190 13512 7196 13524
rect 6880 13484 7196 13512
rect 6880 13472 6886 13484
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7745 13515 7803 13521
rect 7745 13481 7757 13515
rect 7791 13512 7803 13515
rect 7834 13512 7840 13524
rect 7791 13484 7840 13512
rect 7791 13481 7803 13484
rect 7745 13475 7803 13481
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 7926 13472 7932 13524
rect 7984 13512 7990 13524
rect 8202 13512 8208 13524
rect 7984 13484 8208 13512
rect 7984 13472 7990 13484
rect 8202 13472 8208 13484
rect 8260 13512 8266 13524
rect 8260 13484 9076 13512
rect 8260 13472 8266 13484
rect 4338 13404 4344 13456
rect 4396 13404 4402 13456
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 8168 13416 8984 13444
rect 8168 13404 8174 13416
rect 4356 13376 4384 13404
rect 6178 13376 6184 13388
rect 4080 13348 4384 13376
rect 5736 13348 6184 13376
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 992 13280 1409 13308
rect 992 13268 998 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 3326 13268 3332 13320
rect 3384 13268 3390 13320
rect 3786 13268 3792 13320
rect 3844 13308 3850 13320
rect 4080 13317 4108 13348
rect 5736 13320 5764 13348
rect 6178 13336 6184 13348
rect 6236 13376 6242 13388
rect 6236 13348 6592 13376
rect 6236 13336 6242 13348
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3844 13280 4077 13308
rect 3844 13268 3850 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 3344 13240 3372 13268
rect 3344 13212 4200 13240
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 1670 13172 1676 13184
rect 1627 13144 1676 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 3970 13172 3976 13184
rect 3927 13144 3976 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 4172 13172 4200 13212
rect 5368 13172 5396 13271
rect 5718 13268 5724 13320
rect 5776 13268 5782 13320
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 6454 13308 6460 13320
rect 5868 13280 6460 13308
rect 5868 13268 5874 13280
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 6564 13317 6592 13348
rect 8018 13336 8024 13388
rect 8076 13336 8082 13388
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 7650 13268 7656 13320
rect 7708 13268 7714 13320
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13308 7987 13311
rect 8036 13308 8064 13336
rect 7975 13280 8064 13308
rect 8113 13311 8171 13317
rect 7975 13277 7987 13280
rect 7929 13271 7987 13277
rect 8113 13277 8125 13311
rect 8159 13308 8171 13311
rect 8202 13308 8208 13320
rect 8159 13280 8208 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 5445 13243 5503 13249
rect 5445 13209 5457 13243
rect 5491 13240 5503 13243
rect 5626 13240 5632 13252
rect 5491 13212 5632 13240
rect 5491 13209 5503 13212
rect 5445 13203 5503 13209
rect 5626 13200 5632 13212
rect 5684 13240 5690 13252
rect 6181 13243 6239 13249
rect 6181 13240 6193 13243
rect 5684 13212 6193 13240
rect 5684 13200 5690 13212
rect 6181 13209 6193 13212
rect 6227 13240 6239 13243
rect 6822 13240 6828 13252
rect 6227 13212 6828 13240
rect 6227 13209 6239 13212
rect 6181 13203 6239 13209
rect 6564 13184 6592 13212
rect 6822 13200 6828 13212
rect 6880 13200 6886 13252
rect 7852 13240 7880 13271
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 8956 13317 8984 13416
rect 9048 13376 9076 13484
rect 9490 13472 9496 13524
rect 9548 13512 9554 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 9548 13484 9689 13512
rect 9548 13472 9554 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 11606 13472 11612 13524
rect 11664 13512 11670 13524
rect 12250 13512 12256 13524
rect 11664 13484 12256 13512
rect 11664 13472 11670 13484
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 12710 13472 12716 13524
rect 12768 13472 12774 13524
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 13412 13484 13461 13512
rect 13412 13472 13418 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 15197 13515 15255 13521
rect 15197 13481 15209 13515
rect 15243 13512 15255 13515
rect 15654 13512 15660 13524
rect 15243 13484 15660 13512
rect 15243 13481 15255 13484
rect 15197 13475 15255 13481
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 20530 13512 20536 13524
rect 19996 13484 20536 13512
rect 9214 13404 9220 13456
rect 9272 13444 9278 13456
rect 9309 13447 9367 13453
rect 9309 13444 9321 13447
rect 9272 13416 9321 13444
rect 9272 13404 9278 13416
rect 9309 13413 9321 13416
rect 9355 13413 9367 13447
rect 9309 13407 9367 13413
rect 9401 13447 9459 13453
rect 9401 13413 9413 13447
rect 9447 13444 9459 13447
rect 11422 13444 11428 13456
rect 9447 13416 11428 13444
rect 9447 13413 9459 13416
rect 9401 13407 9459 13413
rect 11422 13404 11428 13416
rect 11480 13444 11486 13456
rect 13078 13444 13084 13456
rect 11480 13416 13084 13444
rect 11480 13404 11486 13416
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 15565 13379 15623 13385
rect 9048 13348 9812 13376
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 8021 13243 8079 13249
rect 8021 13240 8033 13243
rect 7852 13212 8033 13240
rect 8021 13209 8033 13212
rect 8067 13240 8079 13243
rect 9232 13240 9260 13271
rect 9398 13268 9404 13320
rect 9456 13268 9462 13320
rect 9784 13317 9812 13348
rect 9876 13348 13768 13376
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 8067 13212 9260 13240
rect 9416 13240 9444 13268
rect 9876 13240 9904 13348
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10410 13308 10416 13320
rect 10367 13280 10416 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 9416 13212 9904 13240
rect 9968 13240 9996 13271
rect 10410 13268 10416 13280
rect 10468 13308 10474 13320
rect 10870 13308 10876 13320
rect 10468 13280 10876 13308
rect 10468 13268 10474 13280
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 11146 13268 11152 13320
rect 11204 13268 11210 13320
rect 11238 13268 11244 13320
rect 11296 13268 11302 13320
rect 11514 13268 11520 13320
rect 11572 13268 11578 13320
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 12066 13308 12072 13320
rect 11793 13271 11851 13277
rect 11900 13280 12072 13308
rect 11164 13240 11192 13268
rect 9968 13212 11192 13240
rect 11256 13240 11284 13268
rect 11808 13240 11836 13271
rect 11256 13212 11836 13240
rect 8067 13209 8079 13212
rect 8021 13203 8079 13209
rect 4172 13144 5396 13172
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 6270 13172 6276 13184
rect 6052 13144 6276 13172
rect 6052 13132 6058 13144
rect 6270 13132 6276 13144
rect 6328 13172 6334 13184
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6328 13144 6377 13172
rect 6328 13132 6334 13144
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 6546 13132 6552 13184
rect 6604 13132 6610 13184
rect 6733 13175 6791 13181
rect 6733 13141 6745 13175
rect 6779 13172 6791 13175
rect 8846 13172 8852 13184
rect 6779 13144 8852 13172
rect 6779 13141 6791 13144
rect 6733 13135 6791 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8996 13144 9045 13172
rect 8996 13132 9002 13144
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9033 13135 9091 13141
rect 9122 13132 9128 13184
rect 9180 13172 9186 13184
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 9180 13144 9965 13172
rect 9180 13132 9186 13144
rect 9953 13141 9965 13144
rect 9999 13141 10011 13175
rect 9953 13135 10011 13141
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11900 13172 11928 13280
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12575 13311 12633 13317
rect 12216 13280 12261 13308
rect 12216 13268 12222 13280
rect 12575 13277 12587 13311
rect 12621 13308 12633 13311
rect 12710 13308 12716 13320
rect 12621 13280 12716 13308
rect 12621 13277 12633 13280
rect 12575 13271 12633 13277
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 12802 13268 12808 13320
rect 12860 13268 12866 13320
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 13188 13317 13216 13348
rect 13740 13317 13768 13348
rect 15565 13345 15577 13379
rect 15611 13376 15623 13379
rect 16117 13379 16175 13385
rect 16117 13376 16129 13379
rect 15611 13348 16129 13376
rect 15611 13345 15623 13348
rect 15565 13339 15623 13345
rect 16117 13345 16129 13348
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 19797 13379 19855 13385
rect 19797 13345 19809 13379
rect 19843 13376 19855 13379
rect 19996 13376 20024 13484
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 21729 13515 21787 13521
rect 21729 13481 21741 13515
rect 21775 13481 21787 13515
rect 21729 13475 21787 13481
rect 20346 13404 20352 13456
rect 20404 13444 20410 13456
rect 21634 13444 21640 13456
rect 20404 13416 21640 13444
rect 20404 13404 20410 13416
rect 21634 13404 21640 13416
rect 21692 13444 21698 13456
rect 21744 13444 21772 13475
rect 22738 13472 22744 13524
rect 22796 13512 22802 13524
rect 23106 13512 23112 13524
rect 22796 13484 23112 13512
rect 22796 13472 22802 13484
rect 23106 13472 23112 13484
rect 23164 13472 23170 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 23716 13484 24409 13512
rect 23716 13472 23722 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 24397 13475 24455 13481
rect 25869 13515 25927 13521
rect 25869 13481 25881 13515
rect 25915 13512 25927 13515
rect 26694 13512 26700 13524
rect 25915 13484 26700 13512
rect 25915 13481 25927 13484
rect 25869 13475 25927 13481
rect 26694 13472 26700 13484
rect 26752 13472 26758 13524
rect 30650 13512 30656 13524
rect 30484 13484 30656 13512
rect 21692 13416 21772 13444
rect 22097 13447 22155 13453
rect 21692 13404 21698 13416
rect 22097 13413 22109 13447
rect 22143 13413 22155 13447
rect 22097 13407 22155 13413
rect 22373 13447 22431 13453
rect 22373 13413 22385 13447
rect 22419 13444 22431 13447
rect 22646 13444 22652 13456
rect 22419 13416 22652 13444
rect 22419 13413 22431 13416
rect 22373 13407 22431 13413
rect 20364 13376 20392 13404
rect 19843 13348 20024 13376
rect 20272 13348 20392 13376
rect 20441 13379 20499 13385
rect 19843 13345 19855 13348
rect 19797 13339 19855 13345
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12952 13280 13001 13308
rect 12952 13268 12958 13280
rect 12989 13277 13001 13280
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13308 15439 13311
rect 15470 13308 15476 13320
rect 15427 13280 15476 13308
rect 15427 13277 15439 13280
rect 15381 13271 15439 13277
rect 11977 13243 12035 13249
rect 11977 13209 11989 13243
rect 12023 13240 12035 13243
rect 12345 13243 12403 13249
rect 12345 13240 12357 13243
rect 12023 13212 12357 13240
rect 12023 13209 12035 13212
rect 11977 13203 12035 13209
rect 12345 13209 12357 13212
rect 12391 13209 12403 13243
rect 12345 13203 12403 13209
rect 12437 13243 12495 13249
rect 12437 13209 12449 13243
rect 12483 13240 12495 13243
rect 13096 13240 13124 13271
rect 12483 13212 13124 13240
rect 12483 13209 12495 13212
rect 12437 13203 12495 13209
rect 12544 13184 12572 13212
rect 13354 13200 13360 13252
rect 13412 13240 13418 13252
rect 13556 13240 13584 13271
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 15654 13268 15660 13320
rect 15712 13268 15718 13320
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 13412 13212 13584 13240
rect 13412 13200 13418 13212
rect 15764 13184 15792 13271
rect 15930 13268 15936 13320
rect 15988 13268 15994 13320
rect 16022 13268 16028 13320
rect 16080 13268 16086 13320
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13308 19763 13311
rect 20272 13308 20300 13348
rect 20441 13345 20453 13379
rect 20487 13376 20499 13379
rect 21177 13379 21235 13385
rect 21177 13376 21189 13379
rect 20487 13348 21189 13376
rect 20487 13345 20499 13348
rect 20441 13339 20499 13345
rect 21177 13345 21189 13348
rect 21223 13345 21235 13379
rect 21177 13339 21235 13345
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21600 13348 21833 13376
rect 21600 13336 21606 13348
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 19751 13280 20300 13308
rect 20364 13280 20821 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 20364 13184 20392 13280
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13308 20959 13311
rect 21361 13311 21419 13317
rect 21008 13308 21128 13310
rect 20947 13282 21128 13308
rect 20947 13280 21036 13282
rect 20947 13277 20959 13280
rect 20901 13271 20959 13277
rect 20530 13200 20536 13252
rect 20588 13200 20594 13252
rect 21100 13240 21128 13282
rect 21361 13277 21373 13311
rect 21407 13308 21419 13311
rect 21450 13308 21456 13320
rect 21407 13280 21456 13308
rect 21407 13277 21419 13280
rect 21361 13271 21419 13277
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 21634 13268 21640 13320
rect 21692 13268 21698 13320
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 22112 13308 22140 13407
rect 22646 13404 22652 13416
rect 22704 13444 22710 13456
rect 22830 13444 22836 13456
rect 22704 13416 22836 13444
rect 22704 13404 22710 13416
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 30484 13453 30512 13484
rect 30650 13472 30656 13484
rect 30708 13472 30714 13524
rect 31294 13472 31300 13524
rect 31352 13472 31358 13524
rect 31478 13512 31484 13524
rect 31404 13484 31484 13512
rect 30469 13447 30527 13453
rect 30469 13413 30481 13447
rect 30515 13413 30527 13447
rect 31021 13447 31079 13453
rect 31021 13444 31033 13447
rect 30469 13407 30527 13413
rect 30576 13416 31033 13444
rect 24118 13336 24124 13388
rect 24176 13336 24182 13388
rect 24670 13336 24676 13388
rect 24728 13376 24734 13388
rect 24946 13376 24952 13388
rect 24728 13348 24952 13376
rect 24728 13336 24734 13348
rect 24946 13336 24952 13348
rect 25004 13336 25010 13388
rect 27246 13336 27252 13388
rect 27304 13376 27310 13388
rect 27341 13379 27399 13385
rect 27341 13376 27353 13379
rect 27304 13348 27353 13376
rect 27304 13336 27310 13348
rect 27341 13345 27353 13348
rect 27387 13345 27399 13379
rect 27341 13339 27399 13345
rect 27614 13336 27620 13388
rect 27672 13336 27678 13388
rect 30576 13376 30604 13416
rect 31021 13413 31033 13416
rect 31067 13413 31079 13447
rect 31021 13407 31079 13413
rect 31205 13447 31263 13453
rect 31205 13413 31217 13447
rect 31251 13444 31263 13447
rect 31404 13444 31432 13484
rect 31478 13472 31484 13484
rect 31536 13512 31542 13524
rect 31662 13512 31668 13524
rect 31536 13484 31668 13512
rect 31536 13472 31542 13484
rect 31662 13472 31668 13484
rect 31720 13472 31726 13524
rect 31251 13416 31432 13444
rect 31251 13413 31263 13416
rect 31205 13407 31263 13413
rect 30208 13348 30604 13376
rect 30653 13379 30711 13385
rect 22189 13311 22247 13317
rect 22189 13308 22201 13311
rect 22112 13280 22201 13308
rect 22189 13277 22201 13280
rect 22235 13277 22247 13311
rect 22189 13271 22247 13277
rect 22922 13268 22928 13320
rect 22980 13268 22986 13320
rect 23201 13311 23259 13317
rect 23201 13277 23213 13311
rect 23247 13277 23259 13311
rect 23201 13271 23259 13277
rect 23293 13311 23351 13317
rect 23293 13277 23305 13311
rect 23339 13308 23351 13311
rect 23382 13308 23388 13320
rect 23339 13280 23388 13308
rect 23339 13277 23351 13280
rect 23293 13271 23351 13277
rect 21545 13243 21603 13249
rect 21545 13240 21557 13243
rect 21100 13212 21557 13240
rect 21545 13209 21557 13212
rect 21591 13209 21603 13243
rect 21545 13203 21603 13209
rect 11204 13144 11928 13172
rect 11204 13132 11210 13144
rect 12526 13132 12532 13184
rect 12584 13132 12590 13184
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 12952 13144 13553 13172
rect 12952 13132 12958 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 13541 13135 13599 13141
rect 15746 13132 15752 13184
rect 15804 13132 15810 13184
rect 20346 13132 20352 13184
rect 20404 13132 20410 13184
rect 21082 13132 21088 13184
rect 21140 13132 21146 13184
rect 21560 13172 21588 13203
rect 21910 13200 21916 13252
rect 21968 13240 21974 13252
rect 23216 13240 23244 13271
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13308 24823 13311
rect 26050 13308 26056 13320
rect 24811 13280 26056 13308
rect 24811 13277 24823 13280
rect 24765 13271 24823 13277
rect 26050 13268 26056 13280
rect 26108 13268 26114 13320
rect 28166 13268 28172 13320
rect 28224 13308 28230 13320
rect 28445 13311 28503 13317
rect 28445 13308 28457 13311
rect 28224 13280 28457 13308
rect 28224 13268 28230 13280
rect 28445 13277 28457 13280
rect 28491 13277 28503 13311
rect 28445 13271 28503 13277
rect 30208 13252 30236 13348
rect 30653 13345 30665 13379
rect 30699 13376 30711 13379
rect 31110 13376 31116 13388
rect 30699 13348 31116 13376
rect 30699 13345 30711 13348
rect 30653 13339 30711 13345
rect 31110 13336 31116 13348
rect 31168 13376 31174 13388
rect 31573 13379 31631 13385
rect 31573 13376 31585 13379
rect 31168 13348 31585 13376
rect 31168 13336 31174 13348
rect 31573 13345 31585 13348
rect 31619 13345 31631 13379
rect 31573 13339 31631 13345
rect 31665 13311 31723 13317
rect 31665 13277 31677 13311
rect 31711 13277 31723 13311
rect 31665 13271 31723 13277
rect 21968 13212 23612 13240
rect 21968 13200 21974 13212
rect 23584 13184 23612 13212
rect 23658 13200 23664 13252
rect 23716 13240 23722 13252
rect 24857 13243 24915 13249
rect 24857 13240 24869 13243
rect 23716 13212 24869 13240
rect 23716 13200 23722 13212
rect 24857 13209 24869 13212
rect 24903 13209 24915 13243
rect 27430 13240 27436 13252
rect 26910 13212 27436 13240
rect 24857 13203 24915 13209
rect 27430 13200 27436 13212
rect 27488 13200 27494 13252
rect 29546 13200 29552 13252
rect 29604 13240 29610 13252
rect 30190 13240 30196 13252
rect 29604 13212 30196 13240
rect 29604 13200 29610 13212
rect 30190 13200 30196 13212
rect 30248 13200 30254 13252
rect 30650 13200 30656 13252
rect 30708 13240 30714 13252
rect 30745 13243 30803 13249
rect 30745 13240 30757 13243
rect 30708 13212 30757 13240
rect 30708 13200 30714 13212
rect 30745 13209 30757 13212
rect 30791 13209 30803 13243
rect 31680 13240 31708 13271
rect 31680 13212 32720 13240
rect 30745 13203 30803 13209
rect 32692 13184 32720 13212
rect 22278 13172 22284 13184
rect 21560 13144 22284 13172
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 23109 13175 23167 13181
rect 23109 13141 23121 13175
rect 23155 13172 23167 13175
rect 23290 13172 23296 13184
rect 23155 13144 23296 13172
rect 23155 13141 23167 13144
rect 23109 13135 23167 13141
rect 23290 13132 23296 13144
rect 23348 13132 23354 13184
rect 23566 13132 23572 13184
rect 23624 13132 23630 13184
rect 27890 13132 27896 13184
rect 27948 13132 27954 13184
rect 32674 13132 32680 13184
rect 32732 13132 32738 13184
rect 1104 13082 34840 13104
rect 1104 13030 9344 13082
rect 9396 13030 9408 13082
rect 9460 13030 9472 13082
rect 9524 13030 9536 13082
rect 9588 13030 9600 13082
rect 9652 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 17930 13082
rect 17982 13030 17994 13082
rect 18046 13030 26132 13082
rect 26184 13030 26196 13082
rect 26248 13030 26260 13082
rect 26312 13030 26324 13082
rect 26376 13030 26388 13082
rect 26440 13030 34526 13082
rect 34578 13030 34590 13082
rect 34642 13030 34654 13082
rect 34706 13030 34718 13082
rect 34770 13030 34782 13082
rect 34834 13030 34840 13082
rect 1104 13008 34840 13030
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 7466 12968 7472 12980
rect 6328 12940 7472 12968
rect 6328 12928 6334 12940
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 9125 12971 9183 12977
rect 9125 12937 9137 12971
rect 9171 12968 9183 12971
rect 9214 12968 9220 12980
rect 9171 12940 9220 12968
rect 9171 12937 9183 12940
rect 9125 12931 9183 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 12158 12968 12164 12980
rect 12032 12940 12164 12968
rect 12032 12928 12038 12940
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12802 12968 12808 12980
rect 12492 12940 12808 12968
rect 12492 12928 12498 12940
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 15565 12971 15623 12977
rect 15565 12937 15577 12971
rect 15611 12968 15623 12971
rect 16114 12968 16120 12980
rect 15611 12940 16120 12968
rect 15611 12937 15623 12940
rect 15565 12931 15623 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 20346 12928 20352 12980
rect 20404 12968 20410 12980
rect 21910 12968 21916 12980
rect 20404 12940 21916 12968
rect 20404 12928 20410 12940
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 23290 12928 23296 12980
rect 23348 12928 23354 12980
rect 31294 12928 31300 12980
rect 31352 12968 31358 12980
rect 31573 12971 31631 12977
rect 31573 12968 31585 12971
rect 31352 12940 31585 12968
rect 31352 12928 31358 12940
rect 31573 12937 31585 12940
rect 31619 12937 31631 12971
rect 31573 12931 31631 12937
rect 31938 12928 31944 12980
rect 31996 12928 32002 12980
rect 33045 12971 33103 12977
rect 33045 12937 33057 12971
rect 33091 12968 33103 12971
rect 33505 12971 33563 12977
rect 33505 12968 33517 12971
rect 33091 12940 33517 12968
rect 33091 12937 33103 12940
rect 33045 12931 33103 12937
rect 33505 12937 33517 12940
rect 33551 12937 33563 12971
rect 33505 12931 33563 12937
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 9582 12900 9588 12912
rect 8352 12872 9588 12900
rect 8352 12860 8358 12872
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 12452 12900 12480 12928
rect 11940 12872 12480 12900
rect 16025 12903 16083 12909
rect 11940 12860 11946 12872
rect 16025 12869 16037 12903
rect 16071 12900 16083 12903
rect 16206 12900 16212 12912
rect 16071 12872 16212 12900
rect 16071 12869 16083 12872
rect 16025 12863 16083 12869
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 22278 12860 22284 12912
rect 22336 12900 22342 12912
rect 23308 12900 23336 12928
rect 22336 12872 23336 12900
rect 22336 12860 22342 12872
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 8754 12832 8760 12844
rect 6604 12804 8760 12832
rect 6604 12792 6610 12804
rect 8754 12792 8760 12804
rect 8812 12832 8818 12844
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8812 12804 9045 12832
rect 8812 12792 8818 12804
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9048 12764 9076 12795
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 9180 12804 9229 12832
rect 9180 12792 9186 12804
rect 9217 12801 9229 12804
rect 9263 12801 9275 12835
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 9217 12795 9275 12801
rect 15028 12804 15117 12832
rect 11330 12764 11336 12776
rect 9048 12736 11336 12764
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 15028 12708 15056 12804
rect 15105 12801 15117 12804
rect 15151 12832 15163 12835
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15151 12804 15669 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 15746 12764 15752 12776
rect 15488 12736 15752 12764
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 8202 12696 8208 12708
rect 6880 12668 8208 12696
rect 6880 12656 6886 12668
rect 8202 12656 8208 12668
rect 8260 12696 8266 12708
rect 14090 12696 14096 12708
rect 8260 12668 14096 12696
rect 8260 12656 8266 12668
rect 14090 12656 14096 12668
rect 14148 12656 14154 12708
rect 15010 12656 15016 12708
rect 15068 12656 15074 12708
rect 15488 12640 15516 12736
rect 15746 12724 15752 12736
rect 15804 12764 15810 12776
rect 15856 12764 15884 12795
rect 17126 12792 17132 12844
rect 17184 12792 17190 12844
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12832 17371 12835
rect 18322 12832 18328 12844
rect 17359 12804 18328 12832
rect 17359 12801 17371 12804
rect 17313 12795 17371 12801
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 22848 12841 22876 12872
rect 23382 12860 23388 12912
rect 23440 12900 23446 12912
rect 24581 12903 24639 12909
rect 24581 12900 24593 12903
rect 23440 12872 24593 12900
rect 23440 12860 23446 12872
rect 24581 12869 24593 12872
rect 24627 12900 24639 12903
rect 25498 12900 25504 12912
rect 24627 12872 25504 12900
rect 24627 12869 24639 12872
rect 24581 12863 24639 12869
rect 25498 12860 25504 12872
rect 25556 12900 25562 12912
rect 28721 12903 28779 12909
rect 28721 12900 28733 12903
rect 25556 12872 28733 12900
rect 25556 12860 25562 12872
rect 28721 12869 28733 12872
rect 28767 12869 28779 12903
rect 28721 12863 28779 12869
rect 33597 12903 33655 12909
rect 33597 12869 33609 12903
rect 33643 12900 33655 12903
rect 33643 12872 33916 12900
rect 33643 12869 33655 12872
rect 33597 12863 33655 12869
rect 33888 12844 33916 12872
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12801 22891 12835
rect 22833 12795 22891 12801
rect 22922 12792 22928 12844
rect 22980 12792 22986 12844
rect 24854 12792 24860 12844
rect 24912 12792 24918 12844
rect 25038 12792 25044 12844
rect 25096 12832 25102 12844
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 25096 12804 27169 12832
rect 25096 12792 25102 12804
rect 27157 12801 27169 12804
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 27338 12792 27344 12844
rect 27396 12792 27402 12844
rect 27433 12835 27491 12841
rect 27433 12801 27445 12835
rect 27479 12832 27491 12835
rect 27890 12832 27896 12844
rect 27479 12804 27896 12832
rect 27479 12801 27491 12804
rect 27433 12795 27491 12801
rect 27890 12792 27896 12804
rect 27948 12792 27954 12844
rect 31478 12792 31484 12844
rect 31536 12832 31542 12844
rect 31536 12804 31720 12832
rect 31536 12792 31542 12804
rect 15804 12736 15884 12764
rect 22741 12767 22799 12773
rect 15804 12724 15810 12736
rect 22741 12733 22753 12767
rect 22787 12733 22799 12767
rect 22741 12727 22799 12733
rect 23017 12767 23075 12773
rect 23017 12733 23029 12767
rect 23063 12764 23075 12767
rect 23474 12764 23480 12776
rect 23063 12736 23480 12764
rect 23063 12733 23075 12736
rect 23017 12727 23075 12733
rect 22756 12696 22784 12727
rect 23474 12724 23480 12736
rect 23532 12724 23538 12776
rect 23566 12724 23572 12776
rect 23624 12724 23630 12776
rect 23845 12767 23903 12773
rect 23845 12733 23857 12767
rect 23891 12764 23903 12767
rect 24210 12764 24216 12776
rect 23891 12736 24216 12764
rect 23891 12733 23903 12736
rect 23845 12727 23903 12733
rect 24210 12724 24216 12736
rect 24268 12724 24274 12776
rect 27356 12764 27384 12792
rect 27522 12764 27528 12776
rect 27356 12736 27528 12764
rect 27522 12724 27528 12736
rect 27580 12724 27586 12776
rect 27982 12724 27988 12776
rect 28040 12724 28046 12776
rect 31692 12764 31720 12804
rect 31754 12792 31760 12844
rect 31812 12792 31818 12844
rect 32674 12792 32680 12844
rect 32732 12832 32738 12844
rect 32732 12804 33824 12832
rect 32732 12792 32738 12804
rect 32585 12767 32643 12773
rect 32585 12764 32597 12767
rect 31692 12736 32597 12764
rect 32585 12733 32597 12736
rect 32631 12733 32643 12767
rect 32585 12727 32643 12733
rect 33410 12724 33416 12776
rect 33468 12764 33474 12776
rect 33686 12764 33692 12776
rect 33468 12736 33692 12764
rect 33468 12724 33474 12736
rect 33686 12724 33692 12736
rect 33744 12724 33750 12776
rect 33796 12764 33824 12804
rect 33870 12792 33876 12844
rect 33928 12792 33934 12844
rect 33962 12792 33968 12844
rect 34020 12792 34026 12844
rect 34146 12792 34152 12844
rect 34204 12792 34210 12844
rect 34057 12767 34115 12773
rect 34057 12764 34069 12767
rect 33796 12736 34069 12764
rect 34057 12733 34069 12736
rect 34103 12733 34115 12767
rect 34057 12727 34115 12733
rect 23584 12696 23612 12724
rect 22756 12668 23612 12696
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 7650 12628 7656 12640
rect 7340 12600 7656 12628
rect 7340 12588 7346 12600
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 8754 12588 8760 12640
rect 8812 12628 8818 12640
rect 8938 12628 8944 12640
rect 8812 12600 8944 12628
rect 8812 12588 8818 12600
rect 8938 12588 8944 12600
rect 8996 12628 9002 12640
rect 10962 12628 10968 12640
rect 8996 12600 10968 12628
rect 8996 12588 9002 12600
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 15381 12631 15439 12637
rect 15381 12597 15393 12631
rect 15427 12628 15439 12631
rect 15470 12628 15476 12640
rect 15427 12600 15476 12628
rect 15427 12597 15439 12600
rect 15381 12591 15439 12597
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 17494 12588 17500 12640
rect 17552 12588 17558 12640
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 22557 12631 22615 12637
rect 22557 12628 22569 12631
rect 22336 12600 22569 12628
rect 22336 12588 22342 12600
rect 22557 12597 22569 12600
rect 22603 12597 22615 12631
rect 22557 12591 22615 12597
rect 24670 12588 24676 12640
rect 24728 12588 24734 12640
rect 26970 12588 26976 12640
rect 27028 12588 27034 12640
rect 32030 12588 32036 12640
rect 32088 12628 32094 12640
rect 33137 12631 33195 12637
rect 33137 12628 33149 12631
rect 32088 12600 33149 12628
rect 32088 12588 32094 12600
rect 33137 12597 33149 12600
rect 33183 12597 33195 12631
rect 33137 12591 33195 12597
rect 1104 12538 34684 12560
rect 1104 12486 5147 12538
rect 5199 12486 5211 12538
rect 5263 12486 5275 12538
rect 5327 12486 5339 12538
rect 5391 12486 5403 12538
rect 5455 12486 13541 12538
rect 13593 12486 13605 12538
rect 13657 12486 13669 12538
rect 13721 12486 13733 12538
rect 13785 12486 13797 12538
rect 13849 12486 21935 12538
rect 21987 12486 21999 12538
rect 22051 12486 22063 12538
rect 22115 12486 22127 12538
rect 22179 12486 22191 12538
rect 22243 12486 30329 12538
rect 30381 12486 30393 12538
rect 30445 12486 30457 12538
rect 30509 12486 30521 12538
rect 30573 12486 30585 12538
rect 30637 12486 34684 12538
rect 1104 12464 34684 12486
rect 3605 12427 3663 12433
rect 3605 12393 3617 12427
rect 3651 12424 3663 12427
rect 3786 12424 3792 12436
rect 3651 12396 3792 12424
rect 3651 12393 3663 12396
rect 3605 12387 3663 12393
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 4801 12427 4859 12433
rect 4801 12393 4813 12427
rect 4847 12424 4859 12427
rect 7098 12424 7104 12436
rect 4847 12396 7104 12424
rect 4847 12393 4859 12396
rect 4801 12387 4859 12393
rect 7098 12384 7104 12396
rect 7156 12424 7162 12436
rect 8941 12427 8999 12433
rect 7156 12396 7328 12424
rect 7156 12384 7162 12396
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 4157 12359 4215 12365
rect 4157 12356 4169 12359
rect 3476 12328 4169 12356
rect 3476 12316 3482 12328
rect 4157 12325 4169 12328
rect 4203 12356 4215 12359
rect 4203 12328 4660 12356
rect 4203 12325 4215 12328
rect 4157 12319 4215 12325
rect 3326 12248 3332 12300
rect 3384 12288 3390 12300
rect 3513 12291 3571 12297
rect 3513 12288 3525 12291
rect 3384 12260 3525 12288
rect 3384 12248 3390 12260
rect 3513 12257 3525 12260
rect 3559 12257 3571 12291
rect 3513 12251 3571 12257
rect 3896 12260 4200 12288
rect 3528 12152 3556 12251
rect 3896 12232 3924 12260
rect 3602 12180 3608 12232
rect 3660 12220 3666 12232
rect 3789 12223 3847 12229
rect 3789 12220 3801 12223
rect 3660 12192 3801 12220
rect 3660 12180 3666 12192
rect 3789 12189 3801 12192
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 3878 12180 3884 12232
rect 3936 12180 3942 12232
rect 4172 12229 4200 12260
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 3988 12152 4016 12183
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 4632 12229 4660 12328
rect 6104 12328 7052 12356
rect 6104 12232 6132 12328
rect 6270 12248 6276 12300
rect 6328 12288 6334 12300
rect 6328 12260 6408 12288
rect 6328 12248 6334 12260
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12189 5043 12223
rect 4985 12183 5043 12189
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12220 5319 12223
rect 5534 12220 5540 12232
rect 5307 12192 5540 12220
rect 5307 12189 5319 12192
rect 5261 12183 5319 12189
rect 3528 12124 4016 12152
rect 3234 12044 3240 12096
rect 3292 12044 3298 12096
rect 3988 12084 4016 12124
rect 4062 12112 4068 12164
rect 4120 12152 4126 12164
rect 5000 12152 5028 12183
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 6086 12180 6092 12232
rect 6144 12180 6150 12232
rect 6380 12229 6408 12260
rect 6656 12260 6868 12288
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6365 12223 6423 12229
rect 6227 12192 6316 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 4120 12124 5028 12152
rect 4120 12112 4126 12124
rect 5442 12112 5448 12164
rect 5500 12112 5506 12164
rect 4246 12084 4252 12096
rect 3988 12056 4252 12084
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 5074 12044 5080 12096
rect 5132 12084 5138 12096
rect 5810 12084 5816 12096
rect 5132 12056 5816 12084
rect 5132 12044 5138 12056
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 6288 12084 6316 12192
rect 6365 12189 6377 12223
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 6380 12152 6408 12183
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 6656 12220 6684 12260
rect 6840 12229 6868 12260
rect 7024 12229 7052 12328
rect 7300 12288 7328 12396
rect 8941 12393 8953 12427
rect 8987 12424 8999 12427
rect 9030 12424 9036 12436
rect 8987 12396 9036 12424
rect 8987 12393 8999 12396
rect 8941 12387 8999 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11974 12424 11980 12436
rect 11112 12396 11980 12424
rect 11112 12384 11118 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12526 12384 12532 12436
rect 12584 12384 12590 12436
rect 17586 12424 17592 12436
rect 12636 12396 13308 12424
rect 8386 12356 8392 12368
rect 8220 12328 8392 12356
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 7300 12260 7389 12288
rect 7377 12257 7389 12260
rect 7423 12288 7435 12291
rect 7466 12288 7472 12300
rect 7423 12260 7472 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 7650 12248 7656 12300
rect 7708 12288 7714 12300
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 7708 12260 7941 12288
rect 7708 12248 7714 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8220 12232 8248 12328
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 9306 12316 9312 12368
rect 9364 12356 9370 12368
rect 9950 12356 9956 12368
rect 9364 12328 9956 12356
rect 9364 12316 9370 12328
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 8404 12288 8432 12316
rect 8404 12260 9260 12288
rect 6512 12192 6684 12220
rect 6733 12223 6791 12229
rect 6512 12180 6518 12192
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7101 12223 7159 12229
rect 7101 12189 7113 12223
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12220 7619 12223
rect 7742 12220 7748 12232
rect 7607 12192 7748 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 6748 12152 6776 12183
rect 7116 12152 7144 12183
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 8202 12180 8208 12232
rect 8260 12180 8266 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9232 12229 9260 12260
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 12636 12288 12664 12396
rect 9640 12260 12664 12288
rect 12989 12291 13047 12297
rect 9640 12248 9646 12260
rect 12989 12257 13001 12291
rect 13035 12288 13047 12291
rect 13035 12260 13124 12288
rect 13035 12257 13047 12260
rect 12989 12251 13047 12257
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 6380 12124 6776 12152
rect 7024 12124 7144 12152
rect 7285 12155 7343 12161
rect 7024 12096 7052 12124
rect 7285 12121 7297 12155
rect 7331 12152 7343 12155
rect 8294 12152 8300 12164
rect 7331 12124 8300 12152
rect 7331 12121 7343 12124
rect 7285 12115 7343 12121
rect 8294 12112 8300 12124
rect 8352 12112 8358 12164
rect 9232 12152 9260 12183
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 9503 12223 9561 12229
rect 9503 12189 9515 12223
rect 9549 12220 9561 12223
rect 11146 12220 11152 12232
rect 9549 12192 11152 12220
rect 9549 12189 9561 12192
rect 9503 12183 9561 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11238 12180 11244 12232
rect 11296 12180 11302 12232
rect 12526 12180 12532 12232
rect 12584 12180 12590 12232
rect 12710 12180 12716 12232
rect 12768 12180 12774 12232
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12220 12955 12223
rect 12943 12192 13032 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 9858 12152 9864 12164
rect 9232 12124 9864 12152
rect 9858 12112 9864 12124
rect 9916 12152 9922 12164
rect 9916 12124 10272 12152
rect 9916 12112 9922 12124
rect 6236 12056 6316 12084
rect 6236 12044 6242 12056
rect 6638 12044 6644 12096
rect 6696 12044 6702 12096
rect 7006 12044 7012 12096
rect 7064 12044 7070 12096
rect 7834 12044 7840 12096
rect 7892 12044 7898 12096
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 9398 12084 9404 12096
rect 8536 12056 9404 12084
rect 8536 12044 8542 12056
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 10244 12084 10272 12124
rect 10318 12112 10324 12164
rect 10376 12152 10382 12164
rect 11422 12152 11428 12164
rect 10376 12124 11428 12152
rect 10376 12112 10382 12124
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 12544 12152 12572 12180
rect 12820 12152 12848 12183
rect 12544 12124 12848 12152
rect 13004 12096 13032 12192
rect 13096 12152 13124 12260
rect 13280 12254 13308 12396
rect 16776 12396 17592 12424
rect 13446 12316 13452 12368
rect 13504 12316 13510 12368
rect 16776 12297 16804 12396
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 18141 12427 18199 12433
rect 18141 12393 18153 12427
rect 18187 12424 18199 12427
rect 18414 12424 18420 12436
rect 18187 12396 18420 12424
rect 18187 12393 18199 12396
rect 18141 12387 18199 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 18690 12384 18696 12436
rect 18748 12384 18754 12436
rect 20438 12384 20444 12436
rect 20496 12424 20502 12436
rect 21542 12424 21548 12436
rect 20496 12396 21548 12424
rect 20496 12384 20502 12396
rect 21542 12384 21548 12396
rect 21600 12384 21606 12436
rect 21913 12427 21971 12433
rect 21913 12393 21925 12427
rect 21959 12424 21971 12427
rect 22370 12424 22376 12436
rect 21959 12396 22376 12424
rect 21959 12393 21971 12396
rect 21913 12387 21971 12393
rect 22370 12384 22376 12396
rect 22428 12384 22434 12436
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 23937 12427 23995 12433
rect 23937 12424 23949 12427
rect 23532 12396 23949 12424
rect 23532 12384 23538 12396
rect 23937 12393 23949 12396
rect 23983 12393 23995 12427
rect 25038 12424 25044 12436
rect 23937 12387 23995 12393
rect 24412 12396 25044 12424
rect 17957 12359 18015 12365
rect 17957 12356 17969 12359
rect 17236 12328 17969 12356
rect 17236 12297 17264 12328
rect 17957 12325 17969 12328
rect 18003 12356 18015 12359
rect 18708 12356 18736 12384
rect 18003 12328 18736 12356
rect 18003 12325 18015 12328
rect 17957 12319 18015 12325
rect 19702 12316 19708 12368
rect 19760 12356 19766 12368
rect 19760 12328 22784 12356
rect 19760 12316 19766 12328
rect 13198 12236 13308 12254
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 17221 12291 17279 12297
rect 17221 12257 17233 12291
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 17494 12248 17500 12300
rect 17552 12288 17558 12300
rect 17706 12291 17764 12297
rect 17706 12288 17718 12291
rect 17552 12260 17718 12288
rect 17552 12248 17558 12260
rect 17706 12257 17718 12260
rect 17752 12257 17764 12291
rect 17706 12251 17764 12257
rect 18138 12248 18144 12300
rect 18196 12288 18202 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 18196 12260 18828 12288
rect 18196 12248 18202 12260
rect 13188 12229 13308 12236
rect 18800 12232 18828 12260
rect 21560 12260 22017 12288
rect 21560 12232 21588 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22373 12291 22431 12297
rect 22373 12288 22385 12291
rect 22005 12251 22063 12257
rect 22112 12260 22385 12288
rect 13173 12226 13308 12229
rect 13173 12223 13231 12226
rect 13173 12189 13185 12223
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13412 12192 13461 12220
rect 13412 12180 13418 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 17126 12220 17132 12232
rect 16908 12192 17132 12220
rect 16908 12180 16914 12192
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 17880 12192 18613 12220
rect 13372 12152 13400 12180
rect 13096 12124 13400 12152
rect 16644 12155 16702 12161
rect 16644 12121 16656 12155
rect 16690 12152 16702 12155
rect 17034 12152 17040 12164
rect 16690 12124 17040 12152
rect 16690 12121 16702 12124
rect 16644 12115 16702 12121
rect 17034 12112 17040 12124
rect 17092 12112 17098 12164
rect 10686 12084 10692 12096
rect 10244 12056 10692 12084
rect 10686 12044 10692 12056
rect 10744 12084 10750 12096
rect 11882 12084 11888 12096
rect 10744 12056 11888 12084
rect 10744 12044 10750 12056
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13044 12056 13277 12084
rect 13044 12044 13050 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 16482 12044 16488 12096
rect 16540 12044 16546 12096
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 17402 12084 17408 12096
rect 16899 12056 17408 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 17402 12044 17408 12056
rect 17460 12084 17466 12096
rect 17497 12087 17555 12093
rect 17497 12084 17509 12087
rect 17460 12056 17509 12084
rect 17460 12044 17466 12056
rect 17497 12053 17509 12056
rect 17543 12053 17555 12087
rect 17497 12047 17555 12053
rect 17586 12044 17592 12096
rect 17644 12044 17650 12096
rect 17880 12093 17908 12192
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 18840 12192 20085 12220
rect 18840 12180 18846 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20254 12180 20260 12232
rect 20312 12180 20318 12232
rect 21361 12223 21419 12229
rect 21361 12220 21373 12223
rect 21008 12192 21373 12220
rect 18322 12112 18328 12164
rect 18380 12152 18386 12164
rect 19702 12152 19708 12164
rect 18380 12124 19708 12152
rect 18380 12112 18386 12124
rect 19702 12112 19708 12124
rect 19760 12112 19766 12164
rect 21008 12096 21036 12192
rect 21361 12189 21373 12192
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 21542 12180 21548 12232
rect 21600 12180 21606 12232
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 22112 12220 22140 12260
rect 22373 12257 22385 12260
rect 22419 12288 22431 12291
rect 22554 12288 22560 12300
rect 22419 12260 22560 12288
rect 22419 12257 22431 12260
rect 22373 12251 22431 12257
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 21775 12192 22140 12220
rect 22189 12223 22247 12229
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 22189 12189 22201 12223
rect 22235 12220 22247 12223
rect 22278 12220 22284 12232
rect 22235 12192 22284 12220
rect 22235 12189 22247 12192
rect 22189 12183 22247 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 22756 12229 22784 12328
rect 23290 12316 23296 12368
rect 23348 12356 23354 12368
rect 23753 12359 23811 12365
rect 23348 12328 23520 12356
rect 23348 12316 23354 12328
rect 22830 12248 22836 12300
rect 22888 12288 22894 12300
rect 23492 12297 23520 12328
rect 23753 12325 23765 12359
rect 23799 12356 23811 12359
rect 24412 12356 24440 12396
rect 25038 12384 25044 12396
rect 25096 12384 25102 12436
rect 26145 12427 26203 12433
rect 26145 12393 26157 12427
rect 26191 12424 26203 12427
rect 26191 12396 28396 12424
rect 26191 12393 26203 12396
rect 26145 12387 26203 12393
rect 23799 12328 24440 12356
rect 23799 12325 23811 12328
rect 23753 12319 23811 12325
rect 23385 12291 23443 12297
rect 23385 12288 23397 12291
rect 22888 12260 23397 12288
rect 22888 12248 22894 12260
rect 23385 12257 23397 12260
rect 23431 12257 23443 12291
rect 23385 12251 23443 12257
rect 23477 12291 23535 12297
rect 23477 12257 23489 12291
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 23566 12248 23572 12300
rect 23624 12248 23630 12300
rect 24397 12291 24455 12297
rect 24397 12257 24409 12291
rect 24443 12288 24455 12291
rect 26510 12288 26516 12300
rect 24443 12260 26516 12288
rect 24443 12257 24455 12260
rect 24397 12251 24455 12257
rect 26510 12248 26516 12260
rect 26568 12248 26574 12300
rect 26786 12248 26792 12300
rect 26844 12248 26850 12300
rect 27430 12248 27436 12300
rect 27488 12288 27494 12300
rect 28368 12297 28396 12396
rect 29730 12384 29736 12436
rect 29788 12424 29794 12436
rect 29788 12396 30236 12424
rect 29788 12384 29794 12396
rect 30101 12359 30159 12365
rect 30101 12325 30113 12359
rect 30147 12325 30159 12359
rect 30208 12356 30236 12396
rect 30926 12384 30932 12436
rect 30984 12424 30990 12436
rect 31113 12427 31171 12433
rect 31113 12424 31125 12427
rect 30984 12396 31125 12424
rect 30984 12384 30990 12396
rect 31113 12393 31125 12396
rect 31159 12393 31171 12427
rect 31113 12387 31171 12393
rect 31220 12396 31340 12424
rect 31018 12356 31024 12368
rect 30208 12328 31024 12356
rect 30101 12319 30159 12325
rect 28353 12291 28411 12297
rect 27488 12260 27936 12288
rect 27488 12248 27494 12260
rect 22465 12223 22523 12229
rect 22465 12189 22477 12223
rect 22511 12220 22523 12223
rect 22649 12223 22707 12229
rect 22649 12220 22661 12223
rect 22511 12192 22661 12220
rect 22511 12189 22523 12192
rect 22465 12183 22523 12189
rect 22649 12189 22661 12192
rect 22695 12189 22707 12223
rect 22649 12183 22707 12189
rect 22741 12223 22799 12229
rect 22741 12189 22753 12223
rect 22787 12189 22799 12223
rect 22741 12183 22799 12189
rect 23293 12223 23351 12229
rect 23293 12189 23305 12223
rect 23339 12220 23351 12223
rect 23750 12220 23756 12232
rect 23339 12192 23756 12220
rect 23339 12189 23351 12192
rect 23293 12183 23351 12189
rect 21637 12155 21695 12161
rect 21637 12121 21649 12155
rect 21683 12152 21695 12155
rect 22370 12152 22376 12164
rect 21683 12124 22376 12152
rect 21683 12121 21695 12124
rect 21637 12115 21695 12121
rect 22370 12112 22376 12124
rect 22428 12152 22434 12164
rect 22480 12152 22508 12183
rect 22428 12124 22508 12152
rect 22756 12152 22784 12183
rect 23750 12180 23756 12192
rect 23808 12180 23814 12232
rect 24029 12223 24087 12229
rect 24029 12189 24041 12223
rect 24075 12189 24087 12223
rect 24029 12183 24087 12189
rect 23658 12152 23664 12164
rect 22756 12124 23664 12152
rect 22428 12112 22434 12124
rect 23658 12112 23664 12124
rect 23716 12112 23722 12164
rect 24044 12096 24072 12183
rect 25682 12180 25688 12232
rect 25740 12220 25746 12232
rect 27908 12220 27936 12260
rect 28353 12257 28365 12291
rect 28399 12257 28411 12291
rect 28353 12251 28411 12257
rect 28994 12248 29000 12300
rect 29052 12248 29058 12300
rect 29012 12220 29040 12248
rect 25740 12192 25806 12220
rect 27908 12206 29040 12220
rect 27922 12192 29040 12206
rect 25740 12180 25746 12192
rect 29546 12180 29552 12232
rect 29604 12180 29610 12232
rect 29825 12223 29883 12229
rect 29656 12220 29776 12222
rect 29825 12220 29837 12223
rect 29656 12194 29837 12220
rect 24670 12112 24676 12164
rect 24728 12112 24734 12164
rect 28997 12155 29055 12161
rect 28997 12152 29009 12155
rect 28092 12124 29009 12152
rect 18138 12093 18144 12096
rect 17865 12087 17923 12093
rect 17865 12053 17877 12087
rect 17911 12053 17923 12087
rect 17865 12047 17923 12053
rect 18125 12087 18144 12093
rect 18125 12053 18137 12087
rect 18125 12047 18144 12053
rect 18138 12044 18144 12047
rect 18196 12044 18202 12096
rect 18417 12087 18475 12093
rect 18417 12053 18429 12087
rect 18463 12084 18475 12087
rect 18598 12084 18604 12096
rect 18463 12056 18604 12084
rect 18463 12053 18475 12056
rect 18417 12047 18475 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 20162 12044 20168 12096
rect 20220 12044 20226 12096
rect 20990 12044 20996 12096
rect 21048 12044 21054 12096
rect 21082 12044 21088 12096
rect 21140 12084 21146 12096
rect 24026 12084 24032 12096
rect 21140 12056 24032 12084
rect 21140 12044 21146 12056
rect 24026 12044 24032 12056
rect 24084 12044 24090 12096
rect 24946 12044 24952 12096
rect 25004 12084 25010 12096
rect 28092 12084 28120 12124
rect 28997 12121 29009 12124
rect 29043 12152 29055 12155
rect 29656 12152 29684 12194
rect 29748 12192 29837 12194
rect 29825 12189 29837 12192
rect 29871 12189 29883 12223
rect 29825 12183 29883 12189
rect 29917 12223 29975 12229
rect 29917 12189 29929 12223
rect 29963 12220 29975 12223
rect 30006 12220 30012 12232
rect 29963 12192 30012 12220
rect 29963 12189 29975 12192
rect 29917 12183 29975 12189
rect 30006 12180 30012 12192
rect 30064 12180 30070 12232
rect 30116 12220 30144 12319
rect 31018 12316 31024 12328
rect 31076 12316 31082 12368
rect 31220 12288 31248 12396
rect 31312 12356 31340 12396
rect 31386 12384 31392 12436
rect 31444 12424 31450 12436
rect 31570 12424 31576 12436
rect 31444 12396 31576 12424
rect 31444 12384 31450 12396
rect 31570 12384 31576 12396
rect 31628 12384 31634 12436
rect 31754 12384 31760 12436
rect 31812 12424 31818 12436
rect 31849 12427 31907 12433
rect 31849 12424 31861 12427
rect 31812 12396 31861 12424
rect 31812 12384 31818 12396
rect 31849 12393 31861 12396
rect 31895 12393 31907 12427
rect 33045 12427 33103 12433
rect 33045 12424 33057 12427
rect 31849 12387 31907 12393
rect 31956 12396 33057 12424
rect 31312 12328 31754 12356
rect 30484 12260 31248 12288
rect 31726 12288 31754 12328
rect 31956 12288 31984 12396
rect 33045 12393 33057 12396
rect 33091 12393 33103 12427
rect 33781 12427 33839 12433
rect 33781 12424 33793 12427
rect 33045 12387 33103 12393
rect 33152 12396 33793 12424
rect 32033 12359 32091 12365
rect 32033 12325 32045 12359
rect 32079 12356 32091 12359
rect 33152 12356 33180 12396
rect 33781 12393 33793 12396
rect 33827 12424 33839 12427
rect 33870 12424 33876 12436
rect 33827 12396 33876 12424
rect 33827 12393 33839 12396
rect 33781 12387 33839 12393
rect 33870 12384 33876 12396
rect 33928 12384 33934 12436
rect 34146 12384 34152 12436
rect 34204 12384 34210 12436
rect 32079 12328 33180 12356
rect 32079 12325 32091 12328
rect 32033 12319 32091 12325
rect 31726 12260 32352 12288
rect 30377 12223 30435 12229
rect 30377 12220 30389 12223
rect 30116 12192 30389 12220
rect 30377 12189 30389 12192
rect 30423 12189 30435 12223
rect 30377 12183 30435 12189
rect 29043 12124 29684 12152
rect 29043 12121 29055 12124
rect 28997 12115 29055 12121
rect 29730 12112 29736 12164
rect 29788 12112 29794 12164
rect 30484 12152 30512 12260
rect 30653 12223 30711 12229
rect 30653 12189 30665 12223
rect 30699 12189 30711 12223
rect 30653 12183 30711 12189
rect 29840 12124 30512 12152
rect 25004 12056 28120 12084
rect 25004 12044 25010 12056
rect 28166 12044 28172 12096
rect 28224 12084 28230 12096
rect 28261 12087 28319 12093
rect 28261 12084 28273 12087
rect 28224 12056 28273 12084
rect 28224 12044 28230 12056
rect 28261 12053 28273 12056
rect 28307 12084 28319 12087
rect 29840 12084 29868 12124
rect 28307 12056 29868 12084
rect 28307 12053 28319 12056
rect 28261 12047 28319 12053
rect 30190 12044 30196 12096
rect 30248 12044 30254 12096
rect 30558 12044 30564 12096
rect 30616 12044 30622 12096
rect 30668 12084 30696 12183
rect 31202 12180 31208 12232
rect 31260 12180 31266 12232
rect 31294 12180 31300 12232
rect 31352 12180 31358 12232
rect 31389 12223 31447 12229
rect 31389 12189 31401 12223
rect 31435 12220 31447 12223
rect 31435 12192 31616 12220
rect 31435 12189 31447 12192
rect 31389 12183 31447 12189
rect 31220 12152 31248 12180
rect 31404 12152 31432 12183
rect 31220 12124 31432 12152
rect 31478 12112 31484 12164
rect 31536 12112 31542 12164
rect 31588 12152 31616 12192
rect 31662 12180 31668 12232
rect 31720 12180 31726 12232
rect 31754 12180 31760 12232
rect 31812 12180 31818 12232
rect 32324 12229 32352 12260
rect 32309 12223 32367 12229
rect 31956 12192 32260 12220
rect 31956 12152 31984 12192
rect 31588 12124 31984 12152
rect 32030 12112 32036 12164
rect 32088 12112 32094 12164
rect 32048 12084 32076 12112
rect 30668 12056 32076 12084
rect 32232 12084 32260 12192
rect 32309 12189 32321 12223
rect 32355 12189 32367 12223
rect 32309 12183 32367 12189
rect 32953 12223 33011 12229
rect 32953 12189 32965 12223
rect 32999 12220 33011 12223
rect 33152 12220 33180 12328
rect 33413 12359 33471 12365
rect 33413 12325 33425 12359
rect 33459 12356 33471 12359
rect 34164 12356 34192 12384
rect 33459 12328 34192 12356
rect 33459 12325 33471 12328
rect 33413 12319 33471 12325
rect 32999 12192 33180 12220
rect 33505 12223 33563 12229
rect 32999 12189 33011 12192
rect 32953 12183 33011 12189
rect 33505 12189 33517 12223
rect 33551 12189 33563 12223
rect 33505 12183 33563 12189
rect 32324 12152 32352 12183
rect 33520 12152 33548 12183
rect 32324 12124 33548 12152
rect 33962 12084 33968 12096
rect 32232 12056 33968 12084
rect 33962 12044 33968 12056
rect 34020 12044 34026 12096
rect 1104 11994 34840 12016
rect 1104 11942 9344 11994
rect 9396 11942 9408 11994
rect 9460 11942 9472 11994
rect 9524 11942 9536 11994
rect 9588 11942 9600 11994
rect 9652 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 17930 11994
rect 17982 11942 17994 11994
rect 18046 11942 26132 11994
rect 26184 11942 26196 11994
rect 26248 11942 26260 11994
rect 26312 11942 26324 11994
rect 26376 11942 26388 11994
rect 26440 11942 34526 11994
rect 34578 11942 34590 11994
rect 34642 11942 34654 11994
rect 34706 11942 34718 11994
rect 34770 11942 34782 11994
rect 34834 11942 34840 11994
rect 1104 11920 34840 11942
rect 3234 11840 3240 11892
rect 3292 11840 3298 11892
rect 3973 11883 4031 11889
rect 3973 11849 3985 11883
rect 4019 11880 4031 11883
rect 4062 11880 4068 11892
rect 4019 11852 4068 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 4525 11883 4583 11889
rect 4525 11849 4537 11883
rect 4571 11880 4583 11883
rect 5074 11880 5080 11892
rect 4571 11852 5080 11880
rect 4571 11849 4583 11852
rect 4525 11843 4583 11849
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 6454 11840 6460 11892
rect 6512 11840 6518 11892
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 6641 11883 6699 11889
rect 6641 11880 6653 11883
rect 6604 11852 6653 11880
rect 6604 11840 6610 11852
rect 6641 11849 6653 11852
rect 6687 11849 6699 11883
rect 6641 11843 6699 11849
rect 6730 11840 6736 11892
rect 6788 11840 6794 11892
rect 7377 11883 7435 11889
rect 7377 11849 7389 11883
rect 7423 11880 7435 11883
rect 7558 11880 7564 11892
rect 7423 11852 7564 11880
rect 7423 11849 7435 11852
rect 7377 11843 7435 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7653 11883 7711 11889
rect 7653 11849 7665 11883
rect 7699 11880 7711 11883
rect 8478 11880 8484 11892
rect 7699 11852 8484 11880
rect 7699 11849 7711 11852
rect 7653 11843 7711 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 8849 11883 8907 11889
rect 8849 11849 8861 11883
rect 8895 11880 8907 11883
rect 9030 11880 9036 11892
rect 8895 11852 9036 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 10778 11880 10784 11892
rect 9272 11852 9378 11880
rect 9272 11840 9278 11852
rect 3252 11812 3280 11840
rect 3605 11815 3663 11821
rect 3605 11812 3617 11815
rect 3252 11784 3617 11812
rect 3252 11753 3280 11784
rect 3605 11781 3617 11784
rect 3651 11781 3663 11815
rect 4893 11815 4951 11821
rect 3605 11775 3663 11781
rect 3712 11784 4200 11812
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 3476 11716 3525 11744
rect 3476 11704 3482 11716
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3620 11676 3648 11775
rect 3712 11756 3740 11784
rect 3694 11704 3700 11756
rect 3752 11704 3758 11756
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 3878 11744 3884 11756
rect 3835 11716 3884 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 4172 11753 4200 11784
rect 4893 11781 4905 11815
rect 4939 11812 4951 11815
rect 6472 11812 6500 11840
rect 6748 11812 6776 11840
rect 4939 11784 6592 11812
rect 6748 11784 6868 11812
rect 4939 11781 4951 11784
rect 4893 11775 4951 11781
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 4246 11704 4252 11756
rect 4304 11704 4310 11756
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 4430 11676 4436 11688
rect 3620 11648 4436 11676
rect 4430 11636 4436 11648
rect 4488 11676 4494 11688
rect 4724 11676 4752 11707
rect 5074 11704 5080 11756
rect 5132 11704 5138 11756
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 6236 11716 6469 11744
rect 6236 11704 6242 11716
rect 6457 11713 6469 11716
rect 6503 11713 6515 11747
rect 6564 11744 6592 11784
rect 6840 11753 6868 11784
rect 7466 11772 7472 11824
rect 7524 11812 7530 11824
rect 8021 11815 8079 11821
rect 8021 11812 8033 11815
rect 7524 11784 8033 11812
rect 7524 11772 7530 11784
rect 8021 11781 8033 11784
rect 8067 11781 8079 11815
rect 8021 11775 8079 11781
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 9350 11821 9378 11852
rect 10612 11852 10784 11880
rect 8389 11815 8447 11821
rect 8389 11812 8401 11815
rect 8168 11784 8401 11812
rect 8168 11772 8174 11784
rect 8389 11781 8401 11784
rect 8435 11781 8447 11815
rect 8389 11775 8447 11781
rect 9335 11815 9393 11821
rect 9335 11781 9347 11815
rect 9381 11781 9393 11815
rect 9335 11775 9393 11781
rect 9585 11815 9643 11821
rect 9585 11781 9597 11815
rect 9631 11812 9643 11815
rect 9766 11812 9772 11824
rect 9631 11784 9772 11812
rect 9631 11781 9643 11784
rect 9585 11775 9643 11781
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 10410 11812 10416 11824
rect 10152 11784 10416 11812
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 6564 11716 6745 11744
rect 6457 11707 6515 11713
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 4488 11648 4752 11676
rect 4488 11636 4494 11648
rect 6362 11636 6368 11688
rect 6420 11636 6426 11688
rect 6472 11676 6500 11707
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 6972 11716 7205 11744
rect 6972 11704 6978 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 7006 11676 7012 11688
rect 6472 11648 7012 11676
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 6380 11608 6408 11636
rect 4356 11580 6408 11608
rect 7300 11608 7328 11707
rect 7668 11676 7696 11707
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 7837 11747 7895 11753
rect 7837 11744 7849 11747
rect 7800 11716 7849 11744
rect 7800 11704 7806 11716
rect 7837 11713 7849 11716
rect 7883 11744 7895 11747
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 7883 11716 8309 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 8297 11713 8309 11716
rect 8343 11744 8355 11747
rect 8481 11747 8539 11753
rect 8343 11716 8432 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8202 11676 8208 11688
rect 7668 11648 8208 11676
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8110 11608 8116 11620
rect 7300 11580 8116 11608
rect 3326 11500 3332 11552
rect 3384 11500 3390 11552
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 4356 11549 4384 11580
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 8404 11552 8432 11716
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8501 11608 8529 11707
rect 9030 11704 9036 11756
rect 9088 11704 9094 11756
rect 9122 11704 9128 11756
rect 9180 11704 9186 11756
rect 9242 11747 9300 11753
rect 9242 11713 9254 11747
rect 9288 11744 9300 11747
rect 10152 11744 10180 11784
rect 10410 11772 10416 11784
rect 10468 11772 10474 11824
rect 10414 11769 10472 11772
rect 9288 11716 9378 11744
rect 9288 11713 9300 11716
rect 9242 11707 9300 11713
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 9350 11676 9378 11716
rect 9876 11716 10180 11744
rect 9876 11706 9904 11716
rect 9784 11685 9904 11706
rect 10226 11704 10232 11756
rect 10284 11704 10290 11756
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 10414 11735 10426 11769
rect 10460 11735 10472 11769
rect 10414 11729 10472 11735
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 10612 11744 10640 11852
rect 10778 11840 10784 11852
rect 10836 11880 10842 11892
rect 10836 11852 11836 11880
rect 10836 11840 10842 11852
rect 10686 11772 10692 11824
rect 10744 11772 10750 11824
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 11480 11784 11744 11812
rect 11480 11772 11486 11784
rect 10551 11716 10640 11744
rect 10704 11744 10732 11772
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 10704 11716 10793 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 10887 11747 10945 11753
rect 10887 11713 10899 11747
rect 10933 11744 10945 11747
rect 10933 11716 11008 11744
rect 10933 11713 10945 11716
rect 10887 11707 10945 11713
rect 9493 11680 9551 11685
rect 8812 11668 8984 11676
rect 9049 11668 9378 11676
rect 8812 11648 9378 11668
rect 8812 11636 8818 11648
rect 8956 11640 9077 11648
rect 9490 11628 9496 11680
rect 9548 11668 9554 11680
rect 9732 11679 9904 11685
rect 9548 11640 9585 11668
rect 9732 11645 9744 11679
rect 9778 11678 9904 11679
rect 9953 11679 10011 11685
rect 9778 11648 9812 11678
rect 9778 11645 9790 11648
rect 9548 11628 9554 11640
rect 9732 11639 9790 11645
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10244 11676 10272 11704
rect 9999 11648 10272 11676
rect 10336 11676 10364 11704
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10336 11648 10701 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 10689 11645 10701 11648
rect 10735 11645 10747 11679
rect 10980 11676 11008 11716
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11716 11753 11744 11784
rect 11808 11753 11836 11852
rect 11882 11840 11888 11892
rect 11940 11840 11946 11892
rect 12066 11840 12072 11892
rect 12124 11840 12130 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12894 11880 12900 11892
rect 12483 11852 12900 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13357 11883 13415 11889
rect 13357 11880 13369 11883
rect 13320 11852 13369 11880
rect 13320 11840 13326 11852
rect 13357 11849 13369 11852
rect 13403 11849 13415 11883
rect 13357 11843 13415 11849
rect 13446 11840 13452 11892
rect 13504 11840 13510 11892
rect 16482 11840 16488 11892
rect 16540 11840 16546 11892
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 17497 11883 17555 11889
rect 17497 11880 17509 11883
rect 17092 11852 17509 11880
rect 17092 11840 17098 11852
rect 17497 11849 17509 11852
rect 17543 11849 17555 11883
rect 18138 11880 18144 11892
rect 17497 11843 17555 11849
rect 17880 11852 18144 11880
rect 11900 11812 11928 11840
rect 12084 11812 12112 11840
rect 11900 11784 12020 11812
rect 12084 11784 13216 11812
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11296 11716 11529 11744
rect 11296 11704 11302 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 11882 11704 11888 11756
rect 11940 11704 11946 11756
rect 11992 11744 12020 11784
rect 11992 11716 12296 11744
rect 12161 11679 12219 11685
rect 12161 11676 12173 11679
rect 10980 11648 12173 11676
rect 10689 11639 10747 11645
rect 12161 11645 12173 11648
rect 12207 11645 12219 11679
rect 12268 11676 12296 11716
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11713 12679 11747
rect 12621 11707 12679 11713
rect 12636 11676 12664 11707
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 13188 11753 13216 11784
rect 13464 11753 13492 11840
rect 13630 11772 13636 11824
rect 13688 11812 13694 11824
rect 16500 11812 16528 11840
rect 17402 11812 17408 11824
rect 13688 11784 13860 11812
rect 13688 11772 13694 11784
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11713 13507 11747
rect 13449 11707 13507 11713
rect 12268 11648 12664 11676
rect 12912 11676 12940 11707
rect 13538 11704 13544 11756
rect 13596 11704 13602 11756
rect 13722 11704 13728 11756
rect 13780 11704 13786 11756
rect 13832 11753 13860 11784
rect 15580 11784 16528 11812
rect 16684 11784 17408 11812
rect 15580 11753 15608 11784
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16684 11744 16712 11784
rect 17402 11772 17408 11784
rect 17460 11812 17466 11824
rect 17880 11821 17908 11852
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18414 11840 18420 11892
rect 18472 11880 18478 11892
rect 18472 11852 19564 11880
rect 18472 11840 18478 11852
rect 17865 11815 17923 11821
rect 17865 11812 17877 11815
rect 17460 11784 17877 11812
rect 17460 11772 17466 11784
rect 17865 11781 17877 11784
rect 17911 11781 17923 11815
rect 18230 11812 18236 11824
rect 17865 11775 17923 11781
rect 17972 11784 18236 11812
rect 16347 11716 16712 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16758 11704 16764 11756
rect 16816 11744 16822 11756
rect 17218 11744 17224 11756
rect 16816 11716 17224 11744
rect 16816 11704 16822 11716
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17972 11753 18000 11784
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 19536 11812 19564 11852
rect 19702 11840 19708 11892
rect 19760 11840 19766 11892
rect 21082 11880 21088 11892
rect 20548 11852 21088 11880
rect 20548 11812 20576 11852
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 21542 11840 21548 11892
rect 21600 11840 21606 11892
rect 21637 11883 21695 11889
rect 21637 11849 21649 11883
rect 21683 11849 21695 11883
rect 21637 11843 21695 11849
rect 21560 11812 21588 11840
rect 19536 11784 20576 11812
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 17957 11747 18015 11753
rect 17957 11713 17969 11747
rect 18003 11713 18015 11747
rect 19610 11744 19616 11756
rect 19366 11716 19616 11744
rect 17957 11707 18015 11713
rect 14001 11679 14059 11685
rect 14001 11676 14013 11679
rect 12912 11648 14013 11676
rect 12161 11639 12219 11645
rect 14001 11645 14013 11648
rect 14047 11645 14059 11679
rect 14001 11639 14059 11645
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 16485 11679 16543 11685
rect 16485 11645 16497 11679
rect 16531 11676 16543 11679
rect 16850 11676 16856 11688
rect 16531 11648 16856 11676
rect 16531 11645 16543 11648
rect 16485 11639 16543 11645
rect 9968 11608 9996 11639
rect 8501 11580 9168 11608
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4028 11512 4353 11540
rect 4028 11500 4034 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 7101 11543 7159 11549
rect 7101 11509 7113 11543
rect 7147 11540 7159 11543
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 7147 11512 7573 11540
rect 7147 11509 7159 11512
rect 7101 11503 7159 11509
rect 7561 11509 7573 11512
rect 7607 11509 7619 11543
rect 7561 11503 7619 11509
rect 8202 11500 8208 11552
rect 8260 11500 8266 11552
rect 8386 11500 8392 11552
rect 8444 11500 8450 11552
rect 9140 11540 9168 11580
rect 9600 11580 9996 11608
rect 9600 11540 9628 11580
rect 10318 11568 10324 11620
rect 10376 11608 10382 11620
rect 12989 11611 13047 11617
rect 12989 11608 13001 11611
rect 10376 11580 13001 11608
rect 10376 11568 10382 11580
rect 12989 11577 13001 11580
rect 13035 11577 13047 11611
rect 12989 11571 13047 11577
rect 13081 11611 13139 11617
rect 13081 11577 13093 11611
rect 13127 11577 13139 11611
rect 16132 11608 16160 11639
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 17034 11636 17040 11688
rect 17092 11636 17098 11688
rect 17696 11608 17724 11707
rect 19610 11704 19616 11716
rect 19668 11744 19674 11756
rect 19978 11744 19984 11756
rect 19668 11716 19984 11744
rect 19668 11704 19674 11716
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20070 11704 20076 11756
rect 20128 11704 20134 11756
rect 20162 11704 20168 11756
rect 20220 11744 20226 11756
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 20220 11716 20361 11744
rect 20220 11704 20226 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 20438 11704 20444 11756
rect 20496 11704 20502 11756
rect 20548 11753 20576 11784
rect 21100 11784 21588 11812
rect 21100 11753 21128 11784
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11744 21511 11747
rect 21542 11744 21548 11756
rect 21499 11716 21548 11744
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 21652 11744 21680 11843
rect 22370 11840 22376 11892
rect 22428 11840 22434 11892
rect 22462 11840 22468 11892
rect 22520 11840 22526 11892
rect 22664 11852 22876 11880
rect 21726 11772 21732 11824
rect 21784 11812 21790 11824
rect 22097 11815 22155 11821
rect 22097 11812 22109 11815
rect 21784 11784 22109 11812
rect 21784 11772 21790 11784
rect 22097 11781 22109 11784
rect 22143 11781 22155 11815
rect 22388 11812 22416 11840
rect 22664 11824 22692 11852
rect 22097 11775 22155 11781
rect 22204 11784 22416 11812
rect 22204 11753 22232 11784
rect 22646 11772 22652 11824
rect 22704 11772 22710 11824
rect 22848 11821 22876 11852
rect 24026 11840 24032 11892
rect 24084 11840 24090 11892
rect 24581 11883 24639 11889
rect 24581 11849 24593 11883
rect 24627 11880 24639 11883
rect 24854 11880 24860 11892
rect 24627 11852 24860 11880
rect 24627 11849 24639 11852
rect 24581 11843 24639 11849
rect 24854 11840 24860 11852
rect 24912 11840 24918 11892
rect 24946 11840 24952 11892
rect 25004 11840 25010 11892
rect 28000 11852 30420 11880
rect 22833 11815 22891 11821
rect 22833 11781 22845 11815
rect 22879 11781 22891 11815
rect 24044 11812 24072 11840
rect 28000 11824 28028 11852
rect 25041 11815 25099 11821
rect 25041 11812 25053 11815
rect 24044 11784 25053 11812
rect 22833 11775 22891 11781
rect 25041 11781 25053 11784
rect 25087 11781 25099 11815
rect 25041 11775 25099 11781
rect 22742 11769 22800 11775
rect 27982 11772 27988 11824
rect 28040 11772 28046 11824
rect 30101 11815 30159 11821
rect 30101 11781 30113 11815
rect 30147 11812 30159 11815
rect 30190 11812 30196 11824
rect 30147 11784 30196 11812
rect 30147 11781 30159 11784
rect 30101 11775 30159 11781
rect 30190 11772 30196 11784
rect 30248 11772 30254 11824
rect 22742 11756 22754 11769
rect 22788 11756 22800 11769
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21652 11716 21833 11744
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 21914 11747 21972 11753
rect 21914 11713 21926 11747
rect 21960 11713 21972 11747
rect 21914 11707 21972 11713
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 22327 11747 22385 11753
rect 22327 11713 22339 11747
rect 22373 11744 22385 11747
rect 22554 11744 22560 11756
rect 22373 11716 22560 11744
rect 22373 11713 22385 11716
rect 22327 11707 22385 11713
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18598 11676 18604 11688
rect 18279 11648 18604 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 20257 11679 20315 11685
rect 20257 11645 20269 11679
rect 20303 11645 20315 11679
rect 20257 11639 20315 11645
rect 20717 11679 20775 11685
rect 20717 11645 20729 11679
rect 20763 11676 20775 11679
rect 20898 11676 20904 11688
rect 20763 11648 20904 11676
rect 20763 11645 20775 11648
rect 20717 11639 20775 11645
rect 16132 11580 17724 11608
rect 13081 11571 13139 11577
rect 9140 11512 9628 11540
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 9950 11540 9956 11552
rect 9907 11512 9956 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10502 11540 10508 11552
rect 10100 11512 10508 11540
rect 10100 11500 10106 11512
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 10597 11543 10655 11549
rect 10597 11509 10609 11543
rect 10643 11540 10655 11543
rect 11146 11540 11152 11552
rect 10643 11512 11152 11540
rect 10643 11509 10655 11512
rect 10597 11503 10655 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11330 11500 11336 11552
rect 11388 11500 11394 11552
rect 12621 11543 12679 11549
rect 12621 11509 12633 11543
rect 12667 11540 12679 11543
rect 13096 11540 13124 11571
rect 12667 11512 13124 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15252 11512 15393 11540
rect 15252 11500 15258 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 17696 11540 17724 11580
rect 20162 11568 20168 11620
rect 20220 11608 20226 11620
rect 20272 11608 20300 11639
rect 20898 11636 20904 11648
rect 20956 11676 20962 11688
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20956 11648 21005 11676
rect 20956 11636 20962 11648
rect 20993 11645 21005 11648
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 21634 11636 21640 11688
rect 21692 11676 21698 11688
rect 21928 11676 21956 11707
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 22738 11704 22744 11756
rect 22796 11704 22802 11756
rect 22925 11747 22983 11753
rect 22925 11744 22937 11747
rect 22848 11716 22937 11744
rect 21692 11648 21956 11676
rect 22066 11648 22692 11676
rect 21692 11636 21698 11648
rect 22066 11608 22094 11648
rect 20220 11580 22094 11608
rect 22296 11580 22600 11608
rect 20220 11568 20226 11580
rect 17954 11540 17960 11552
rect 17696 11512 17960 11540
rect 15381 11503 15439 11509
rect 17954 11500 17960 11512
rect 18012 11540 18018 11552
rect 18414 11540 18420 11552
rect 18012 11512 18420 11540
rect 18012 11500 18018 11512
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 21450 11500 21456 11552
rect 21508 11540 21514 11552
rect 22296 11540 22324 11580
rect 22572 11549 22600 11580
rect 21508 11512 22324 11540
rect 22557 11543 22615 11549
rect 21508 11500 21514 11512
rect 22557 11509 22569 11543
rect 22603 11509 22615 11543
rect 22664 11540 22692 11648
rect 22848 11620 22876 11716
rect 22925 11713 22937 11716
rect 22971 11713 22983 11747
rect 23043 11747 23101 11753
rect 23043 11744 23055 11747
rect 22925 11707 22983 11713
rect 23032 11713 23055 11744
rect 23089 11713 23101 11747
rect 23032 11707 23101 11713
rect 23032 11676 23060 11707
rect 28994 11704 29000 11756
rect 29052 11704 29058 11756
rect 30392 11753 30420 11852
rect 30558 11840 30564 11892
rect 30616 11880 30622 11892
rect 30616 11852 31754 11880
rect 30616 11840 30622 11852
rect 31294 11812 31300 11824
rect 31220 11784 31300 11812
rect 31220 11753 31248 11784
rect 31294 11772 31300 11784
rect 31352 11772 31358 11824
rect 30377 11747 30435 11753
rect 30377 11713 30389 11747
rect 30423 11713 30435 11747
rect 30377 11707 30435 11713
rect 31205 11747 31263 11753
rect 31205 11713 31217 11747
rect 31251 11713 31263 11747
rect 31205 11707 31263 11713
rect 22940 11648 23060 11676
rect 23201 11679 23259 11685
rect 22940 11620 22968 11648
rect 23201 11645 23213 11679
rect 23247 11676 23259 11679
rect 24302 11676 24308 11688
rect 23247 11648 24308 11676
rect 23247 11645 23259 11648
rect 23201 11639 23259 11645
rect 22830 11568 22836 11620
rect 22888 11568 22894 11620
rect 22922 11568 22928 11620
rect 22980 11568 22986 11620
rect 23216 11540 23244 11639
rect 24302 11636 24308 11648
rect 24360 11636 24366 11688
rect 25038 11636 25044 11688
rect 25096 11676 25102 11688
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 25096 11648 25145 11676
rect 25096 11636 25102 11648
rect 25133 11645 25145 11648
rect 25179 11645 25191 11679
rect 25133 11639 25191 11645
rect 28629 11679 28687 11685
rect 28629 11645 28641 11679
rect 28675 11676 28687 11679
rect 29546 11676 29552 11688
rect 28675 11648 29552 11676
rect 28675 11645 28687 11648
rect 28629 11639 28687 11645
rect 29546 11636 29552 11648
rect 29604 11636 29610 11688
rect 31386 11568 31392 11620
rect 31444 11568 31450 11620
rect 31726 11608 31754 11852
rect 31938 11608 31944 11620
rect 31726 11580 31944 11608
rect 31938 11568 31944 11580
rect 31996 11608 32002 11620
rect 31996 11580 32536 11608
rect 31996 11568 32002 11580
rect 22664 11512 23244 11540
rect 22557 11503 22615 11509
rect 27522 11500 27528 11552
rect 27580 11540 27586 11552
rect 30006 11540 30012 11552
rect 27580 11512 30012 11540
rect 27580 11500 27586 11512
rect 30006 11500 30012 11512
rect 30064 11500 30070 11552
rect 31202 11500 31208 11552
rect 31260 11540 31266 11552
rect 31297 11543 31355 11549
rect 31297 11540 31309 11543
rect 31260 11512 31309 11540
rect 31260 11500 31266 11512
rect 31297 11509 31309 11512
rect 31343 11509 31355 11543
rect 31404 11540 31432 11568
rect 32508 11552 32536 11580
rect 31662 11540 31668 11552
rect 31404 11512 31668 11540
rect 31297 11503 31355 11509
rect 31662 11500 31668 11512
rect 31720 11500 31726 11552
rect 32490 11500 32496 11552
rect 32548 11500 32554 11552
rect 1104 11450 34684 11472
rect 1104 11398 5147 11450
rect 5199 11398 5211 11450
rect 5263 11398 5275 11450
rect 5327 11398 5339 11450
rect 5391 11398 5403 11450
rect 5455 11398 13541 11450
rect 13593 11398 13605 11450
rect 13657 11398 13669 11450
rect 13721 11398 13733 11450
rect 13785 11398 13797 11450
rect 13849 11398 21935 11450
rect 21987 11398 21999 11450
rect 22051 11398 22063 11450
rect 22115 11398 22127 11450
rect 22179 11398 22191 11450
rect 22243 11398 30329 11450
rect 30381 11398 30393 11450
rect 30445 11398 30457 11450
rect 30509 11398 30521 11450
rect 30573 11398 30585 11450
rect 30637 11398 34684 11450
rect 1104 11376 34684 11398
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 4430 11336 4436 11348
rect 4295 11308 4436 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 5534 11296 5540 11348
rect 5592 11296 5598 11348
rect 6362 11296 6368 11348
rect 6420 11296 6426 11348
rect 8110 11296 8116 11348
rect 8168 11296 8174 11348
rect 8665 11339 8723 11345
rect 8665 11305 8677 11339
rect 8711 11336 8723 11339
rect 9030 11336 9036 11348
rect 8711 11308 9036 11336
rect 8711 11305 8723 11308
rect 8665 11299 8723 11305
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 9950 11296 9956 11348
rect 10008 11296 10014 11348
rect 10318 11296 10324 11348
rect 10376 11296 10382 11348
rect 10413 11339 10471 11345
rect 10413 11305 10425 11339
rect 10459 11336 10471 11339
rect 11238 11336 11244 11348
rect 10459 11308 11244 11336
rect 10459 11305 10471 11308
rect 10413 11299 10471 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11330 11296 11336 11348
rect 11388 11296 11394 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 12400 11308 12449 11336
rect 12400 11296 12406 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 12437 11299 12495 11305
rect 12820 11308 13032 11336
rect 1394 11160 1400 11212
rect 1452 11160 1458 11212
rect 1670 11160 1676 11212
rect 1728 11160 1734 11212
rect 2958 11132 2964 11144
rect 2806 11104 2964 11132
rect 2958 11092 2964 11104
rect 3016 11132 3022 11144
rect 3234 11132 3240 11144
rect 3016 11104 3240 11132
rect 3016 11092 3022 11104
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 3436 11132 3464 11296
rect 5552 11268 5580 11296
rect 5552 11240 6776 11268
rect 6178 11160 6184 11212
rect 6236 11200 6242 11212
rect 6236 11172 6408 11200
rect 6236 11160 6242 11172
rect 6380 11141 6408 11172
rect 6454 11160 6460 11212
rect 6512 11160 6518 11212
rect 6748 11200 6776 11240
rect 6822 11228 6828 11280
rect 6880 11228 6886 11280
rect 8128 11268 8156 11296
rect 8128 11240 8294 11268
rect 7466 11200 7472 11212
rect 6748 11172 7472 11200
rect 7466 11160 7472 11172
rect 7524 11200 7530 11212
rect 8266 11200 8294 11240
rect 8938 11228 8944 11280
rect 8996 11268 9002 11280
rect 9677 11271 9735 11277
rect 8996 11240 9444 11268
rect 8996 11228 9002 11240
rect 7524 11172 7788 11200
rect 7524 11160 7530 11172
rect 6365 11135 6423 11141
rect 3436 11104 4200 11132
rect 3970 11024 3976 11076
rect 4028 11064 4034 11076
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 4028 11036 4077 11064
rect 4028 11024 4034 11036
rect 4065 11033 4077 11036
rect 4111 11033 4123 11067
rect 4172 11064 4200 11104
rect 6365 11101 6377 11135
rect 6411 11101 6423 11135
rect 6365 11095 6423 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 6730 11132 6736 11144
rect 6687 11104 6736 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 7282 11092 7288 11144
rect 7340 11092 7346 11144
rect 4265 11067 4323 11073
rect 4265 11064 4277 11067
rect 4172 11036 4277 11064
rect 4065 11027 4123 11033
rect 4265 11033 4277 11036
rect 4311 11033 4323 11067
rect 4706 11064 4712 11076
rect 4265 11027 4323 11033
rect 4448 11036 4712 11064
rect 3142 10956 3148 11008
rect 3200 10956 3206 11008
rect 4448 11005 4476 11036
rect 4706 11024 4712 11036
rect 4764 11064 4770 11076
rect 7300 11064 7328 11092
rect 4764 11036 7328 11064
rect 7760 11064 7788 11172
rect 7944 11172 8156 11200
rect 8266 11172 8529 11200
rect 7944 11144 7972 11172
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 8128 11141 8156 11172
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8114 11135 8172 11141
rect 8114 11101 8126 11135
rect 8160 11101 8172 11135
rect 8114 11095 8172 11101
rect 8036 11064 8064 11095
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8501 11141 8529 11172
rect 8864 11172 9352 11200
rect 8864 11144 8892 11172
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 8260 11104 8309 11132
rect 8260 11092 8266 11104
rect 8297 11101 8309 11104
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8486 11135 8544 11141
rect 8486 11101 8498 11135
rect 8532 11101 8544 11135
rect 8486 11095 8544 11101
rect 8846 11092 8852 11144
rect 8904 11092 8910 11144
rect 9324 11141 9352 11172
rect 9416 11141 9444 11240
rect 9677 11237 9689 11271
rect 9723 11268 9735 11271
rect 10336 11268 10364 11296
rect 9723 11240 10364 11268
rect 11348 11268 11376 11296
rect 12820 11268 12848 11308
rect 11348 11240 12848 11268
rect 9723 11237 9735 11240
rect 9677 11231 9735 11237
rect 12894 11228 12900 11280
rect 12952 11228 12958 11280
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 12805 11203 12863 11209
rect 9824 11172 9996 11200
rect 9824 11160 9830 11172
rect 9968 11141 9996 11172
rect 12805 11169 12817 11203
rect 12851 11200 12863 11203
rect 12912 11200 12940 11228
rect 12851 11172 12940 11200
rect 13004 11200 13032 11308
rect 13078 11296 13084 11348
rect 13136 11296 13142 11348
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 13906 11336 13912 11348
rect 13587 11308 13912 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 16577 11339 16635 11345
rect 16577 11305 16589 11339
rect 16623 11336 16635 11339
rect 17954 11336 17960 11348
rect 16623 11308 17960 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 17954 11296 17960 11308
rect 18012 11296 18018 11348
rect 20898 11296 20904 11348
rect 20956 11296 20962 11348
rect 20990 11296 20996 11348
rect 21048 11296 21054 11348
rect 21450 11296 21456 11348
rect 21508 11296 21514 11348
rect 21542 11296 21548 11348
rect 21600 11336 21606 11348
rect 22557 11339 22615 11345
rect 22557 11336 22569 11339
rect 21600 11308 22569 11336
rect 21600 11296 21606 11308
rect 22557 11305 22569 11308
rect 22603 11305 22615 11339
rect 22557 11299 22615 11305
rect 30561 11339 30619 11345
rect 30561 11305 30573 11339
rect 30607 11336 30619 11339
rect 30650 11336 30656 11348
rect 30607 11308 30656 11336
rect 30607 11305 30619 11308
rect 30561 11299 30619 11305
rect 30650 11296 30656 11308
rect 30708 11296 30714 11348
rect 30745 11339 30803 11345
rect 30745 11305 30757 11339
rect 30791 11336 30803 11339
rect 31294 11336 31300 11348
rect 30791 11308 31300 11336
rect 30791 11305 30803 11308
rect 30745 11299 30803 11305
rect 31294 11296 31300 11308
rect 31352 11296 31358 11348
rect 31570 11296 31576 11348
rect 31628 11336 31634 11348
rect 31665 11339 31723 11345
rect 31665 11336 31677 11339
rect 31628 11308 31677 11336
rect 31628 11296 31634 11308
rect 31665 11305 31677 11308
rect 31711 11305 31723 11339
rect 31665 11299 31723 11305
rect 13096 11268 13124 11296
rect 13096 11240 13400 11268
rect 13004 11172 13124 11200
rect 12851 11169 12863 11172
rect 12805 11163 12863 11169
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 7760 11036 8064 11064
rect 8389 11067 8447 11073
rect 4764 11024 4770 11036
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 8570 11064 8576 11076
rect 8435 11036 8576 11064
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 9048 11064 9076 11095
rect 8812 11036 9076 11064
rect 8812 11024 8818 11036
rect 4433 10999 4491 11005
rect 4433 10965 4445 10999
rect 4479 10965 4491 10999
rect 4433 10959 4491 10965
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 8018 10996 8024 11008
rect 6880 10968 8024 10996
rect 6880 10956 6886 10968
rect 8018 10956 8024 10968
rect 8076 10996 8082 11008
rect 9232 10996 9260 11095
rect 8076 10968 9260 10996
rect 8076 10956 8082 10968
rect 9950 10956 9956 11008
rect 10008 10996 10014 11008
rect 10152 10996 10180 11095
rect 10226 11092 10232 11144
rect 10284 11092 10290 11144
rect 12526 11092 12532 11144
rect 12584 11092 12590 11144
rect 12618 11092 12624 11144
rect 12676 11092 12682 11144
rect 13096 11141 13124 11172
rect 13372 11141 13400 11240
rect 17034 11228 17040 11280
rect 17092 11228 17098 11280
rect 17586 11228 17592 11280
rect 17644 11268 17650 11280
rect 18506 11268 18512 11280
rect 17644 11240 18512 11268
rect 17644 11228 17650 11240
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14550 11200 14556 11212
rect 14056 11172 14556 11200
rect 14056 11160 14062 11172
rect 14550 11160 14556 11172
rect 14608 11200 14614 11212
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 14608 11172 14841 11200
rect 14608 11160 14614 11172
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11200 15163 11203
rect 15194 11200 15200 11212
rect 15151 11172 15200 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11101 12955 11135
rect 12897 11095 12955 11101
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 17052 11132 17080 11228
rect 20916 11141 20944 11296
rect 16238 11118 17080 11132
rect 13357 11095 13415 11101
rect 16224 11104 17080 11118
rect 20901 11135 20959 11141
rect 12544 11064 12572 11092
rect 12728 11064 12756 11095
rect 12544 11036 12756 11064
rect 10008 10968 10180 10996
rect 10008 10956 10014 10968
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 12912 10996 12940 11095
rect 13173 11067 13231 11073
rect 13173 11033 13185 11067
rect 13219 11064 13231 11067
rect 13262 11064 13268 11076
rect 13219 11036 13268 11064
rect 13219 11033 13231 11036
rect 13173 11027 13231 11033
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 13354 10996 13360 11008
rect 12584 10968 13360 10996
rect 12584 10956 12590 10968
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 15930 10956 15936 11008
rect 15988 10996 15994 11008
rect 16224 10996 16252 11104
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 21085 11135 21143 11141
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 21468 11132 21496 11296
rect 23201 11271 23259 11277
rect 23201 11237 23213 11271
rect 23247 11268 23259 11271
rect 26510 11268 26516 11280
rect 23247 11240 26516 11268
rect 23247 11237 23259 11240
rect 23201 11231 23259 11237
rect 26510 11228 26516 11240
rect 26568 11228 26574 11280
rect 30006 11228 30012 11280
rect 30064 11268 30070 11280
rect 31754 11268 31760 11280
rect 30064 11240 31760 11268
rect 30064 11228 30070 11240
rect 31754 11228 31760 11240
rect 31812 11228 31818 11280
rect 22922 11200 22928 11212
rect 21131 11104 21496 11132
rect 22066 11172 22928 11200
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 20070 11024 20076 11076
rect 20128 11064 20134 11076
rect 22066 11064 22094 11172
rect 22922 11160 22928 11172
rect 22980 11200 22986 11212
rect 26973 11203 27031 11209
rect 22980 11172 23704 11200
rect 22980 11160 22986 11172
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 22738 11092 22744 11144
rect 22796 11132 22802 11144
rect 23676 11141 23704 11172
rect 26973 11169 26985 11203
rect 27019 11200 27031 11203
rect 27614 11200 27620 11212
rect 27019 11172 27620 11200
rect 27019 11169 27031 11172
rect 26973 11163 27031 11169
rect 27614 11160 27620 11172
rect 27672 11160 27678 11212
rect 28994 11200 29000 11212
rect 28368 11172 29000 11200
rect 22833 11135 22891 11141
rect 22833 11132 22845 11135
rect 22796 11104 22845 11132
rect 22796 11092 22802 11104
rect 22833 11101 22845 11104
rect 22879 11132 22891 11135
rect 23109 11135 23167 11141
rect 23109 11132 23121 11135
rect 22879 11104 23121 11132
rect 22879 11101 22891 11104
rect 22833 11095 22891 11101
rect 23109 11101 23121 11104
rect 23155 11101 23167 11135
rect 23109 11095 23167 11101
rect 23293 11135 23351 11141
rect 23293 11101 23305 11135
rect 23339 11101 23351 11135
rect 23293 11095 23351 11101
rect 23661 11135 23719 11141
rect 23661 11101 23673 11135
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 20128 11036 22094 11064
rect 20128 11024 20134 11036
rect 22554 11024 22560 11076
rect 22612 11024 22618 11076
rect 22664 11064 22692 11092
rect 23308 11064 23336 11095
rect 26694 11092 26700 11144
rect 26752 11092 26758 11144
rect 28368 11118 28396 11172
rect 28994 11160 29000 11172
rect 29052 11160 29058 11212
rect 30193 11203 30251 11209
rect 30193 11169 30205 11203
rect 30239 11200 30251 11203
rect 30926 11200 30932 11212
rect 30239 11172 30932 11200
rect 30239 11169 30251 11172
rect 30193 11163 30251 11169
rect 30926 11160 30932 11172
rect 30984 11160 30990 11212
rect 32030 11200 32036 11212
rect 31220 11172 32036 11200
rect 28534 11092 28540 11144
rect 28592 11132 28598 11144
rect 29549 11135 29607 11141
rect 29549 11132 29561 11135
rect 28592 11104 29561 11132
rect 28592 11092 28598 11104
rect 29549 11101 29561 11104
rect 29595 11101 29607 11135
rect 30282 11134 30288 11144
rect 30208 11132 30288 11134
rect 29549 11095 29607 11101
rect 29840 11106 30288 11132
rect 29840 11104 30236 11106
rect 22664 11036 23336 11064
rect 23753 11067 23811 11073
rect 15988 10968 16252 10996
rect 22664 10996 22692 11036
rect 23753 11033 23765 11067
rect 23799 11064 23811 11067
rect 25682 11064 25688 11076
rect 23799 11036 25688 11064
rect 23799 11033 23811 11036
rect 23753 11027 23811 11033
rect 25682 11024 25688 11036
rect 25740 11024 25746 11076
rect 27249 11067 27307 11073
rect 27249 11064 27261 11067
rect 26896 11036 27261 11064
rect 26896 11005 26924 11036
rect 27249 11033 27261 11036
rect 27295 11033 27307 11067
rect 29840 11064 29868 11104
rect 30282 11092 30288 11106
rect 30340 11092 30346 11144
rect 31220 11141 31248 11172
rect 32030 11160 32036 11172
rect 32088 11160 32094 11212
rect 31205 11135 31263 11141
rect 31205 11101 31217 11135
rect 31251 11101 31263 11135
rect 31205 11095 31263 11101
rect 31294 11092 31300 11144
rect 31352 11092 31358 11144
rect 31481 11135 31539 11141
rect 31481 11101 31493 11135
rect 31527 11101 31539 11135
rect 31481 11095 31539 11101
rect 31496 11064 31524 11095
rect 31662 11092 31668 11144
rect 31720 11132 31726 11144
rect 31941 11135 31999 11141
rect 31941 11132 31953 11135
rect 31720 11104 31953 11132
rect 31720 11092 31726 11104
rect 31941 11101 31953 11104
rect 31987 11101 31999 11135
rect 31941 11095 31999 11101
rect 27249 11027 27307 11033
rect 28736 11036 29868 11064
rect 31220 11036 31524 11064
rect 28736 11008 28764 11036
rect 31220 11008 31248 11036
rect 22741 10999 22799 11005
rect 22741 10996 22753 10999
rect 22664 10968 22753 10996
rect 15988 10956 15994 10968
rect 22741 10965 22753 10968
rect 22787 10965 22799 10999
rect 22741 10959 22799 10965
rect 26881 10999 26939 11005
rect 26881 10965 26893 10999
rect 26927 10965 26939 10999
rect 26881 10959 26939 10965
rect 28718 10956 28724 11008
rect 28776 10956 28782 11008
rect 31202 10956 31208 11008
rect 31260 10956 31266 11008
rect 32309 10999 32367 11005
rect 32309 10965 32321 10999
rect 32355 10996 32367 10999
rect 33042 10996 33048 11008
rect 32355 10968 33048 10996
rect 32355 10965 32367 10968
rect 32309 10959 32367 10965
rect 33042 10956 33048 10968
rect 33100 10956 33106 11008
rect 1104 10906 34840 10928
rect 1104 10854 9344 10906
rect 9396 10854 9408 10906
rect 9460 10854 9472 10906
rect 9524 10854 9536 10906
rect 9588 10854 9600 10906
rect 9652 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 17930 10906
rect 17982 10854 17994 10906
rect 18046 10854 26132 10906
rect 26184 10854 26196 10906
rect 26248 10854 26260 10906
rect 26312 10854 26324 10906
rect 26376 10854 26388 10906
rect 26440 10854 34526 10906
rect 34578 10854 34590 10906
rect 34642 10854 34654 10906
rect 34706 10854 34718 10906
rect 34770 10854 34782 10906
rect 34834 10854 34840 10906
rect 1104 10832 34840 10854
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 9674 10792 9680 10804
rect 5215 10764 9680 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 17494 10752 17500 10804
rect 17552 10792 17558 10804
rect 17681 10795 17739 10801
rect 17681 10792 17693 10795
rect 17552 10764 17693 10792
rect 17552 10752 17558 10764
rect 17681 10761 17693 10764
rect 17727 10761 17739 10795
rect 17681 10755 17739 10761
rect 18049 10795 18107 10801
rect 18049 10761 18061 10795
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 5445 10727 5503 10733
rect 5445 10724 5457 10727
rect 4908 10696 5457 10724
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3200 10628 3617 10656
rect 3200 10616 3206 10628
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 4908 10665 4936 10696
rect 5445 10693 5457 10696
rect 5491 10693 5503 10727
rect 5445 10687 5503 10693
rect 6270 10684 6276 10736
rect 6328 10684 6334 10736
rect 6362 10684 6368 10736
rect 6420 10684 6426 10736
rect 6840 10696 7604 10724
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4672 10628 4905 10656
rect 4672 10616 4678 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 5040 10628 5273 10656
rect 5040 10616 5046 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 6288 10656 6316 10684
rect 5583 10628 6316 10656
rect 6380 10656 6408 10684
rect 6840 10665 6868 10696
rect 7576 10668 7604 10696
rect 7742 10684 7748 10736
rect 7800 10724 7806 10736
rect 12802 10724 12808 10736
rect 7800 10696 12808 10724
rect 7800 10684 7806 10696
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6380 10628 6561 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6549 10619 6607 10625
rect 6656 10628 6837 10656
rect 4706 10548 4712 10600
rect 4764 10548 4770 10600
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10588 4859 10591
rect 5552 10588 5580 10619
rect 4847 10560 5580 10588
rect 4847 10557 4859 10560
rect 4801 10551 4859 10557
rect 3326 10480 3332 10532
rect 3384 10520 3390 10532
rect 4816 10520 4844 10551
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6656 10588 6684 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 5868 10560 6684 10588
rect 6733 10591 6791 10597
rect 5868 10548 5874 10560
rect 6733 10557 6745 10591
rect 6779 10588 6791 10591
rect 6914 10588 6920 10600
rect 6779 10560 6920 10588
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 6641 10523 6699 10529
rect 3384 10492 4844 10520
rect 5552 10492 6592 10520
rect 3384 10480 3390 10492
rect 5552 10464 5580 10492
rect 3050 10412 3056 10464
rect 3108 10412 3114 10464
rect 5534 10412 5540 10464
rect 5592 10412 5598 10464
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 6564 10452 6592 10492
rect 6641 10489 6653 10523
rect 6687 10520 6699 10523
rect 6822 10520 6828 10532
rect 6687 10492 6828 10520
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 6822 10480 6828 10492
rect 6880 10480 6886 10532
rect 7024 10452 7052 10619
rect 7558 10616 7564 10668
rect 7616 10616 7622 10668
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 12710 10656 12716 10668
rect 11112 10628 12716 10656
rect 11112 10616 11118 10628
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 17402 10616 17408 10668
rect 17460 10616 17466 10668
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17773 10659 17831 10665
rect 17773 10656 17785 10659
rect 17644 10628 17785 10656
rect 17644 10616 17650 10628
rect 17773 10625 17785 10628
rect 17819 10625 17831 10659
rect 18064 10656 18092 10755
rect 18340 10724 18368 10755
rect 20162 10752 20168 10804
rect 20220 10752 20226 10804
rect 24673 10795 24731 10801
rect 24673 10761 24685 10795
rect 24719 10761 24731 10795
rect 24673 10755 24731 10761
rect 18693 10727 18751 10733
rect 18693 10724 18705 10727
rect 18340 10696 18705 10724
rect 18693 10693 18705 10696
rect 18739 10693 18751 10727
rect 24688 10724 24716 10755
rect 25682 10752 25688 10804
rect 25740 10792 25746 10804
rect 25740 10764 26372 10792
rect 25740 10752 25746 10764
rect 25041 10727 25099 10733
rect 25041 10724 25053 10727
rect 24688 10696 25053 10724
rect 18693 10687 18751 10693
rect 25041 10693 25053 10696
rect 25087 10693 25099 10727
rect 25041 10687 25099 10693
rect 25130 10684 25136 10736
rect 25188 10724 25194 10736
rect 26344 10724 26372 10764
rect 26694 10752 26700 10804
rect 26752 10792 26758 10804
rect 26973 10795 27031 10801
rect 26973 10792 26985 10795
rect 26752 10764 26985 10792
rect 26752 10752 26758 10764
rect 26973 10761 26985 10764
rect 27019 10761 27031 10795
rect 26973 10755 27031 10761
rect 31941 10795 31999 10801
rect 31941 10761 31953 10795
rect 31987 10761 31999 10795
rect 31941 10755 31999 10761
rect 32677 10795 32735 10801
rect 32677 10761 32689 10795
rect 32723 10761 32735 10795
rect 32677 10755 32735 10761
rect 27433 10727 27491 10733
rect 27433 10724 27445 10727
rect 25188 10696 25530 10724
rect 26344 10696 27445 10724
rect 25188 10684 25194 10696
rect 27433 10693 27445 10696
rect 27479 10693 27491 10727
rect 27433 10687 27491 10693
rect 30282 10684 30288 10736
rect 30340 10684 30346 10736
rect 30926 10684 30932 10736
rect 30984 10724 30990 10736
rect 31665 10727 31723 10733
rect 31665 10724 31677 10727
rect 30984 10696 31677 10724
rect 30984 10684 30990 10696
rect 31665 10693 31677 10696
rect 31711 10693 31723 10727
rect 31665 10687 31723 10693
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 18064 10628 18153 10656
rect 17773 10619 17831 10625
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 19978 10656 19984 10668
rect 19826 10628 19984 10656
rect 18141 10619 18199 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 23106 10616 23112 10668
rect 23164 10616 23170 10668
rect 24118 10616 24124 10668
rect 24176 10616 24182 10668
rect 24486 10616 24492 10668
rect 24544 10616 24550 10668
rect 27341 10659 27399 10665
rect 27341 10625 27353 10659
rect 27387 10656 27399 10659
rect 28077 10659 28135 10665
rect 28077 10656 28089 10659
rect 27387 10628 28089 10656
rect 27387 10625 27399 10628
rect 27341 10619 27399 10625
rect 28077 10625 28089 10628
rect 28123 10625 28135 10659
rect 28077 10619 28135 10625
rect 28718 10616 28724 10668
rect 28776 10616 28782 10668
rect 31389 10659 31447 10665
rect 31389 10625 31401 10659
rect 31435 10625 31447 10659
rect 31389 10619 31447 10625
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 13078 10588 13084 10600
rect 11296 10560 13084 10588
rect 11296 10548 11302 10560
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 13170 10548 13176 10600
rect 13228 10588 13234 10600
rect 13354 10588 13360 10600
rect 13228 10560 13360 10588
rect 13228 10548 13234 10560
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 17862 10548 17868 10600
rect 17920 10597 17926 10600
rect 17920 10591 17948 10597
rect 17936 10557 17948 10591
rect 17920 10551 17948 10557
rect 17920 10548 17926 10551
rect 18414 10548 18420 10600
rect 18472 10548 18478 10600
rect 24136 10588 24164 10616
rect 24765 10591 24823 10597
rect 24765 10588 24777 10591
rect 24136 10560 24777 10588
rect 24765 10557 24777 10560
rect 24811 10557 24823 10591
rect 24765 10551 24823 10557
rect 27522 10548 27528 10600
rect 27580 10548 27586 10600
rect 31404 10588 31432 10619
rect 31570 10616 31576 10668
rect 31628 10616 31634 10668
rect 31754 10616 31760 10668
rect 31812 10616 31818 10668
rect 31956 10656 31984 10755
rect 32309 10659 32367 10665
rect 32309 10656 32321 10659
rect 31956 10628 32321 10656
rect 32309 10625 32321 10628
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 32490 10616 32496 10668
rect 32548 10616 32554 10668
rect 32585 10659 32643 10665
rect 32585 10625 32597 10659
rect 32631 10656 32643 10659
rect 32692 10656 32720 10755
rect 33042 10752 33048 10804
rect 33100 10752 33106 10804
rect 32631 10628 32720 10656
rect 32631 10625 32643 10628
rect 32585 10619 32643 10625
rect 33042 10616 33048 10668
rect 33100 10656 33106 10668
rect 33100 10628 33272 10656
rect 33100 10616 33106 10628
rect 31404 10560 31708 10588
rect 8570 10480 8576 10532
rect 8628 10520 8634 10532
rect 8628 10492 9674 10520
rect 8628 10480 8634 10492
rect 7098 10452 7104 10464
rect 6564 10424 7104 10452
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 9646 10452 9674 10492
rect 28166 10480 28172 10532
rect 28224 10520 28230 10532
rect 30650 10520 30656 10532
rect 28224 10492 30656 10520
rect 28224 10480 28230 10492
rect 30650 10480 30656 10492
rect 30708 10520 30714 10532
rect 31294 10520 31300 10532
rect 30708 10492 31300 10520
rect 30708 10480 30714 10492
rect 31294 10480 31300 10492
rect 31352 10480 31358 10532
rect 31680 10520 31708 10560
rect 32214 10548 32220 10600
rect 32272 10588 32278 10600
rect 33137 10591 33195 10597
rect 33137 10588 33149 10591
rect 32272 10560 33149 10588
rect 32272 10548 32278 10560
rect 33137 10557 33149 10560
rect 33183 10557 33195 10591
rect 33244 10588 33272 10628
rect 33321 10591 33379 10597
rect 33321 10588 33333 10591
rect 33244 10560 33333 10588
rect 33137 10551 33195 10557
rect 33321 10557 33333 10560
rect 33367 10588 33379 10591
rect 33778 10588 33784 10600
rect 33367 10560 33784 10588
rect 33367 10557 33379 10560
rect 33321 10551 33379 10557
rect 33778 10548 33784 10560
rect 33836 10548 33842 10600
rect 33870 10520 33876 10532
rect 31680 10492 33876 10520
rect 33870 10480 33876 10492
rect 33928 10480 33934 10532
rect 12342 10452 12348 10464
rect 9646 10424 12348 10452
rect 12342 10412 12348 10424
rect 12400 10452 12406 10464
rect 12618 10452 12624 10464
rect 12400 10424 12624 10452
rect 12400 10412 12406 10424
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 22922 10412 22928 10464
rect 22980 10412 22986 10464
rect 26513 10455 26571 10461
rect 26513 10421 26525 10455
rect 26559 10452 26571 10455
rect 26602 10452 26608 10464
rect 26559 10424 26608 10452
rect 26559 10421 26571 10424
rect 26513 10415 26571 10421
rect 26602 10412 26608 10424
rect 26660 10452 26666 10464
rect 28534 10452 28540 10464
rect 26660 10424 28540 10452
rect 26660 10412 26666 10424
rect 28534 10412 28540 10424
rect 28592 10412 28598 10464
rect 30745 10455 30803 10461
rect 30745 10421 30757 10455
rect 30791 10452 30803 10455
rect 31202 10452 31208 10464
rect 30791 10424 31208 10452
rect 30791 10421 30803 10424
rect 30745 10415 30803 10421
rect 31202 10412 31208 10424
rect 31260 10412 31266 10464
rect 31754 10412 31760 10464
rect 31812 10452 31818 10464
rect 31938 10452 31944 10464
rect 31812 10424 31944 10452
rect 31812 10412 31818 10424
rect 31938 10412 31944 10424
rect 31996 10412 32002 10464
rect 32122 10412 32128 10464
rect 32180 10412 32186 10464
rect 1104 10362 34684 10384
rect 1104 10310 5147 10362
rect 5199 10310 5211 10362
rect 5263 10310 5275 10362
rect 5327 10310 5339 10362
rect 5391 10310 5403 10362
rect 5455 10310 13541 10362
rect 13593 10310 13605 10362
rect 13657 10310 13669 10362
rect 13721 10310 13733 10362
rect 13785 10310 13797 10362
rect 13849 10310 21935 10362
rect 21987 10310 21999 10362
rect 22051 10310 22063 10362
rect 22115 10310 22127 10362
rect 22179 10310 22191 10362
rect 22243 10310 30329 10362
rect 30381 10310 30393 10362
rect 30445 10310 30457 10362
rect 30509 10310 30521 10362
rect 30573 10310 30585 10362
rect 30637 10310 34684 10362
rect 1104 10288 34684 10310
rect 6362 10208 6368 10260
rect 6420 10208 6426 10260
rect 6549 10251 6607 10257
rect 6549 10217 6561 10251
rect 6595 10248 6607 10251
rect 6638 10248 6644 10260
rect 6595 10220 6644 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7742 10248 7748 10260
rect 6963 10220 7748 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 5629 10183 5687 10189
rect 5629 10149 5641 10183
rect 5675 10180 5687 10183
rect 5997 10183 6055 10189
rect 5997 10180 6009 10183
rect 5675 10152 6009 10180
rect 5675 10149 5687 10152
rect 5629 10143 5687 10149
rect 5997 10149 6009 10152
rect 6043 10149 6055 10183
rect 5997 10143 6055 10149
rect 6089 10183 6147 10189
rect 6089 10149 6101 10183
rect 6135 10180 6147 10183
rect 6380 10180 6408 10208
rect 6135 10152 6408 10180
rect 6135 10149 6147 10152
rect 6089 10143 6147 10149
rect 5810 10112 5816 10124
rect 5384 10084 5816 10112
rect 5384 10053 5412 10084
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 6932 10112 6960 10211
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8570 10248 8576 10260
rect 7975 10220 8576 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8720 10220 8953 10248
rect 8720 10208 8726 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 11054 10248 11060 10260
rect 8941 10211 8999 10217
rect 9324 10220 11060 10248
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8297 10183 8355 10189
rect 8297 10180 8309 10183
rect 8260 10152 8309 10180
rect 8260 10140 8266 10152
rect 8297 10149 8309 10152
rect 8343 10149 8355 10183
rect 8297 10143 8355 10149
rect 8478 10140 8484 10192
rect 8536 10140 8542 10192
rect 5920 10084 6960 10112
rect 7469 10115 7527 10121
rect 5356 10047 5414 10053
rect 5356 10013 5368 10047
rect 5402 10013 5414 10047
rect 5356 10007 5414 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5534 10044 5540 10056
rect 5491 10016 5540 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5920 10053 5948 10084
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 8496 10112 8524 10140
rect 9324 10112 9352 10220
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 11287 10220 12909 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 12897 10217 12909 10220
rect 12943 10248 12955 10251
rect 13446 10248 13452 10260
rect 12943 10220 13452 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 17402 10208 17408 10260
rect 17460 10208 17466 10260
rect 17862 10208 17868 10260
rect 17920 10208 17926 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 19058 10248 19064 10260
rect 18196 10220 19064 10248
rect 18196 10208 18202 10220
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 22728 10251 22786 10257
rect 22728 10217 22740 10251
rect 22774 10248 22786 10251
rect 22922 10248 22928 10260
rect 22774 10220 22928 10248
rect 22774 10217 22786 10220
rect 22728 10211 22786 10217
rect 22922 10208 22928 10220
rect 22980 10208 22986 10260
rect 24486 10208 24492 10260
rect 24544 10248 24550 10260
rect 24949 10251 25007 10257
rect 24949 10248 24961 10251
rect 24544 10220 24961 10248
rect 24544 10208 24550 10220
rect 24949 10217 24961 10220
rect 24995 10217 25007 10251
rect 24949 10211 25007 10217
rect 27614 10208 27620 10260
rect 27672 10248 27678 10260
rect 27672 10220 29592 10248
rect 27672 10208 27678 10220
rect 11146 10180 11152 10192
rect 10980 10152 11152 10180
rect 10980 10121 11008 10152
rect 11146 10140 11152 10152
rect 11204 10180 11210 10192
rect 12345 10183 12403 10189
rect 11204 10152 11744 10180
rect 11204 10140 11210 10152
rect 11716 10124 11744 10152
rect 12345 10149 12357 10183
rect 12391 10180 12403 10183
rect 13170 10180 13176 10192
rect 12391 10152 13176 10180
rect 12391 10149 12403 10152
rect 12345 10143 12403 10149
rect 13170 10140 13176 10152
rect 13228 10180 13234 10192
rect 17420 10180 17448 10208
rect 17957 10183 18015 10189
rect 17957 10180 17969 10183
rect 13228 10152 13308 10180
rect 17420 10152 17969 10180
rect 13228 10140 13234 10152
rect 7515 10084 8524 10112
rect 9140 10084 9352 10112
rect 10965 10115 11023 10121
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6178 10004 6184 10056
rect 6236 10004 6242 10056
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6307 10016 6469 10044
rect 4522 9936 4528 9988
rect 4580 9976 4586 9988
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 4580 9948 5641 9976
rect 4580 9936 4586 9948
rect 5629 9945 5641 9948
rect 5675 9945 5687 9979
rect 5629 9939 5687 9945
rect 6307 9908 6335 10016
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10044 6791 10047
rect 7190 10044 7196 10056
rect 6779 10016 7196 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7558 10004 7564 10056
rect 7616 10004 7622 10056
rect 7926 10004 7932 10056
rect 7984 10004 7990 10056
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8386 10044 8392 10056
rect 8067 10016 8392 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 9140 10053 9168 10084
rect 10965 10081 10977 10115
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 11238 10112 11244 10124
rect 11103 10084 11244 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10112 11391 10115
rect 11422 10112 11428 10124
rect 11379 10084 11428 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 11698 10072 11704 10124
rect 11756 10072 11762 10124
rect 12526 10112 12532 10124
rect 11808 10084 12532 10112
rect 11808 10056 11836 10084
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 9272 10016 9321 10044
rect 9272 10004 9278 10016
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 6365 9979 6423 9985
rect 6365 9945 6377 9979
rect 6411 9976 6423 9979
rect 7006 9976 7012 9988
rect 6411 9948 7012 9976
rect 6411 9945 6423 9948
rect 6365 9939 6423 9945
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 7098 9936 7104 9988
rect 7156 9936 7162 9988
rect 7285 9979 7343 9985
rect 7285 9945 7297 9979
rect 7331 9976 7343 9979
rect 7466 9976 7472 9988
rect 7331 9948 7472 9976
rect 7331 9945 7343 9948
rect 7285 9939 7343 9945
rect 7466 9936 7472 9948
rect 7524 9976 7530 9988
rect 7745 9979 7803 9985
rect 7745 9976 7757 9979
rect 7524 9948 7757 9976
rect 7524 9936 7530 9948
rect 7745 9945 7757 9948
rect 7791 9945 7803 9979
rect 7944 9976 7972 10004
rect 8113 9979 8171 9985
rect 8113 9976 8125 9979
rect 7944 9948 8125 9976
rect 7745 9939 7803 9945
rect 8113 9945 8125 9948
rect 8159 9945 8171 9979
rect 8113 9939 8171 9945
rect 8297 9979 8355 9985
rect 8297 9945 8309 9979
rect 8343 9945 8355 9979
rect 9416 9976 9444 10007
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 9732 10016 10609 10044
rect 9732 10004 9738 10016
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 10870 10044 10876 10056
rect 10735 10016 10876 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 11606 10004 11612 10056
rect 11664 10004 11670 10056
rect 11790 10004 11796 10056
rect 11848 10004 11854 10056
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 12124 10016 12173 10044
rect 12124 10004 12130 10016
rect 12161 10013 12173 10016
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12250 10004 12256 10056
rect 12308 10044 12314 10056
rect 12452 10053 12480 10084
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10112 12863 10115
rect 12851 10084 13032 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 12345 10047 12403 10053
rect 12345 10044 12357 10047
rect 12308 10016 12357 10044
rect 12308 10004 12314 10016
rect 12345 10013 12357 10016
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 12894 10044 12900 10056
rect 12676 10016 12900 10044
rect 12676 10004 12682 10016
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 12713 9979 12771 9985
rect 12713 9976 12725 9979
rect 9416 9948 12725 9976
rect 8297 9939 8355 9945
rect 12713 9945 12725 9948
rect 12759 9945 12771 9979
rect 12713 9939 12771 9945
rect 7650 9908 7656 9920
rect 6307 9880 7656 9908
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 7760 9908 7788 9939
rect 8312 9908 8340 9939
rect 13004 9920 13032 10084
rect 13280 10053 13308 10152
rect 17957 10149 17969 10152
rect 18003 10149 18015 10183
rect 17957 10143 18015 10149
rect 24213 10183 24271 10189
rect 24213 10149 24225 10183
rect 24259 10180 24271 10183
rect 24394 10180 24400 10192
rect 24259 10152 24400 10180
rect 24259 10149 24271 10152
rect 24213 10143 24271 10149
rect 24394 10140 24400 10152
rect 24452 10180 24458 10192
rect 27341 10183 27399 10189
rect 24452 10152 26740 10180
rect 24452 10140 24458 10152
rect 22465 10115 22523 10121
rect 22465 10081 22477 10115
rect 22511 10112 22523 10115
rect 23474 10112 23480 10124
rect 22511 10084 23480 10112
rect 22511 10081 22523 10084
rect 22465 10075 22523 10081
rect 23474 10072 23480 10084
rect 23532 10112 23538 10124
rect 24118 10112 24124 10124
rect 23532 10084 24124 10112
rect 23532 10072 23538 10084
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 24302 10072 24308 10124
rect 24360 10112 24366 10124
rect 25409 10115 25467 10121
rect 25409 10112 25421 10115
rect 24360 10084 25421 10112
rect 24360 10072 24366 10084
rect 25409 10081 25421 10084
rect 25455 10081 25467 10115
rect 25409 10075 25467 10081
rect 25501 10115 25559 10121
rect 25501 10081 25513 10115
rect 25547 10081 25559 10115
rect 25501 10075 25559 10081
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 17681 10047 17739 10053
rect 17681 10013 17693 10047
rect 17727 10044 17739 10047
rect 25130 10044 25136 10056
rect 17727 10016 18368 10044
rect 23874 10030 25136 10044
rect 17727 10013 17739 10016
rect 17681 10007 17739 10013
rect 13173 9979 13231 9985
rect 13173 9945 13185 9979
rect 13219 9976 13231 9979
rect 13725 9979 13783 9985
rect 13725 9976 13737 9979
rect 13219 9948 13737 9976
rect 13219 9945 13231 9948
rect 13173 9939 13231 9945
rect 13725 9945 13737 9948
rect 13771 9945 13783 9979
rect 13725 9939 13783 9945
rect 17402 9936 17408 9988
rect 17460 9976 17466 9988
rect 18340 9985 18368 10016
rect 23860 10016 25136 10030
rect 17497 9979 17555 9985
rect 17497 9976 17509 9979
rect 17460 9948 17509 9976
rect 17460 9936 17466 9948
rect 17497 9945 17509 9948
rect 17543 9945 17555 9979
rect 18109 9979 18167 9985
rect 18109 9976 18121 9979
rect 17497 9939 17555 9945
rect 17788 9948 18121 9976
rect 10318 9908 10324 9920
rect 7760 9880 10324 9908
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 10410 9868 10416 9920
rect 10468 9908 10474 9920
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10468 9880 10793 9908
rect 10468 9868 10474 9880
rect 10781 9877 10793 9880
rect 10827 9877 10839 9911
rect 10781 9871 10839 9877
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11333 9911 11391 9917
rect 11333 9908 11345 9911
rect 11112 9880 11345 9908
rect 11112 9868 11118 9880
rect 11333 9877 11345 9880
rect 11379 9877 11391 9911
rect 11333 9871 11391 9877
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12986 9908 12992 9920
rect 12575 9880 12992 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 13078 9868 13084 9920
rect 13136 9868 13142 9920
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 14090 9908 14096 9920
rect 13403 9880 14096 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 17788 9908 17816 9948
rect 18109 9945 18121 9948
rect 18155 9945 18167 9979
rect 18109 9939 18167 9945
rect 18325 9979 18383 9985
rect 18325 9945 18337 9979
rect 18371 9976 18383 9979
rect 20162 9976 20168 9988
rect 18371 9948 20168 9976
rect 18371 9945 18383 9948
rect 18325 9939 18383 9945
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 17368 9880 17816 9908
rect 17368 9868 17374 9880
rect 19978 9868 19984 9920
rect 20036 9908 20042 9920
rect 23860 9908 23888 10016
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25516 10044 25544 10075
rect 26602 10072 26608 10124
rect 26660 10072 26666 10124
rect 26712 10121 26740 10152
rect 27341 10149 27353 10183
rect 27387 10180 27399 10183
rect 27387 10152 29040 10180
rect 27387 10149 27399 10152
rect 27341 10143 27399 10149
rect 26697 10115 26755 10121
rect 26697 10081 26709 10115
rect 26743 10081 26755 10115
rect 26697 10075 26755 10081
rect 28644 10084 28948 10112
rect 25240 10016 25544 10044
rect 27985 10047 28043 10053
rect 25038 9936 25044 9988
rect 25096 9976 25102 9988
rect 25240 9976 25268 10016
rect 27985 10013 27997 10047
rect 28031 10044 28043 10047
rect 28258 10044 28264 10056
rect 28031 10016 28264 10044
rect 28031 10013 28043 10016
rect 27985 10007 28043 10013
rect 28258 10004 28264 10016
rect 28316 10004 28322 10056
rect 28644 10053 28672 10084
rect 28353 10047 28411 10053
rect 28353 10013 28365 10047
rect 28399 10044 28411 10047
rect 28445 10047 28503 10053
rect 28445 10044 28457 10047
rect 28399 10016 28457 10044
rect 28399 10013 28411 10016
rect 28353 10007 28411 10013
rect 28445 10013 28457 10016
rect 28491 10013 28503 10047
rect 28445 10007 28503 10013
rect 28629 10047 28687 10053
rect 28629 10013 28641 10047
rect 28675 10013 28687 10047
rect 28629 10007 28687 10013
rect 28721 10047 28779 10053
rect 28721 10013 28733 10047
rect 28767 10013 28779 10047
rect 28721 10007 28779 10013
rect 25096 9948 25268 9976
rect 25317 9979 25375 9985
rect 25096 9936 25102 9948
rect 25317 9945 25329 9979
rect 25363 9976 25375 9979
rect 25961 9979 26019 9985
rect 25961 9976 25973 9979
rect 25363 9948 25973 9976
rect 25363 9945 25375 9948
rect 25317 9939 25375 9945
rect 25961 9945 25973 9948
rect 26007 9945 26019 9979
rect 25961 9939 26019 9945
rect 28166 9936 28172 9988
rect 28224 9936 28230 9988
rect 28736 9976 28764 10007
rect 28810 10004 28816 10056
rect 28868 10004 28874 10056
rect 28368 9948 28764 9976
rect 28368 9920 28396 9948
rect 20036 9880 23888 9908
rect 20036 9868 20042 9880
rect 28350 9868 28356 9920
rect 28408 9868 28414 9920
rect 28920 9908 28948 10084
rect 29012 10053 29040 10152
rect 29564 10121 29592 10220
rect 31294 10208 31300 10260
rect 31352 10248 31358 10260
rect 31352 10220 31708 10248
rect 31352 10208 31358 10220
rect 31018 10140 31024 10192
rect 31076 10180 31082 10192
rect 31570 10180 31576 10192
rect 31076 10152 31576 10180
rect 31076 10140 31082 10152
rect 31570 10140 31576 10152
rect 31628 10140 31634 10192
rect 31680 10180 31708 10220
rect 32122 10208 32128 10260
rect 32180 10248 32186 10260
rect 32842 10251 32900 10257
rect 32842 10248 32854 10251
rect 32180 10220 32854 10248
rect 32180 10208 32186 10220
rect 32842 10217 32854 10220
rect 32888 10217 32900 10251
rect 32842 10211 32900 10217
rect 33870 10208 33876 10260
rect 33928 10248 33934 10260
rect 34333 10251 34391 10257
rect 34333 10248 34345 10251
rect 33928 10220 34345 10248
rect 33928 10208 33934 10220
rect 34333 10217 34345 10220
rect 34379 10217 34391 10251
rect 34333 10211 34391 10217
rect 32214 10180 32220 10192
rect 31680 10152 32220 10180
rect 32214 10140 32220 10152
rect 32272 10140 32278 10192
rect 29549 10115 29607 10121
rect 29549 10081 29561 10115
rect 29595 10112 29607 10115
rect 32585 10115 32643 10121
rect 32585 10112 32597 10115
rect 29595 10084 32597 10112
rect 29595 10081 29607 10084
rect 29549 10075 29607 10081
rect 32585 10081 32597 10084
rect 32631 10112 32643 10115
rect 32631 10084 34376 10112
rect 32631 10081 32643 10084
rect 32585 10075 32643 10081
rect 34348 10056 34376 10084
rect 28997 10047 29055 10053
rect 28997 10013 29009 10047
rect 29043 10013 29055 10047
rect 30958 10016 32352 10044
rect 28997 10007 29055 10013
rect 29181 9979 29239 9985
rect 29181 9945 29193 9979
rect 29227 9976 29239 9979
rect 29825 9979 29883 9985
rect 29825 9976 29837 9979
rect 29227 9948 29837 9976
rect 29227 9945 29239 9948
rect 29181 9939 29239 9945
rect 29825 9945 29837 9948
rect 29871 9945 29883 9979
rect 32214 9976 32220 9988
rect 29825 9939 29883 9945
rect 31726 9948 32220 9976
rect 31726 9908 31754 9948
rect 32214 9936 32220 9948
rect 32272 9936 32278 9988
rect 32324 9976 32352 10016
rect 34330 10004 34336 10056
rect 34388 10004 34394 10056
rect 32324 9948 33350 9976
rect 32968 9920 32996 9948
rect 28920 9880 31754 9908
rect 32950 9868 32956 9920
rect 33008 9868 33014 9920
rect 1104 9818 34840 9840
rect 1104 9766 9344 9818
rect 9396 9766 9408 9818
rect 9460 9766 9472 9818
rect 9524 9766 9536 9818
rect 9588 9766 9600 9818
rect 9652 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 17930 9818
rect 17982 9766 17994 9818
rect 18046 9766 26132 9818
rect 26184 9766 26196 9818
rect 26248 9766 26260 9818
rect 26312 9766 26324 9818
rect 26376 9766 26388 9818
rect 26440 9766 34526 9818
rect 34578 9766 34590 9818
rect 34642 9766 34654 9818
rect 34706 9766 34718 9818
rect 34770 9766 34782 9818
rect 34834 9766 34840 9818
rect 1104 9744 34840 9766
rect 6178 9664 6184 9716
rect 6236 9704 6242 9716
rect 8754 9704 8760 9716
rect 6236 9676 8760 9704
rect 6236 9664 6242 9676
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 9125 9707 9183 9713
rect 9125 9673 9137 9707
rect 9171 9704 9183 9707
rect 9214 9704 9220 9716
rect 9171 9676 9220 9704
rect 9171 9673 9183 9676
rect 9125 9667 9183 9673
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 9490 9664 9496 9716
rect 9548 9664 9554 9716
rect 9582 9664 9588 9716
rect 9640 9664 9646 9716
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 9732 9676 9996 9704
rect 9732 9664 9738 9676
rect 2961 9639 3019 9645
rect 2961 9605 2973 9639
rect 3007 9636 3019 9639
rect 3050 9636 3056 9648
rect 3007 9608 3056 9636
rect 3007 9605 3019 9608
rect 2961 9599 3019 9605
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 3234 9596 3240 9648
rect 3292 9636 3298 9648
rect 8573 9639 8631 9645
rect 3292 9608 3450 9636
rect 8128 9608 8524 9636
rect 3292 9596 3298 9608
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 2682 9568 2688 9580
rect 1452 9540 2688 9568
rect 1452 9528 1458 9540
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 8018 9528 8024 9580
rect 8076 9528 8082 9580
rect 8128 9577 8156 9608
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8202 9528 8208 9580
rect 8260 9528 8266 9580
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8496 9568 8524 9608
rect 8573 9605 8585 9639
rect 8619 9636 8631 9639
rect 9306 9636 9312 9648
rect 8619 9608 9312 9636
rect 8619 9605 8631 9608
rect 8573 9599 8631 9605
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 9508 9636 9536 9664
rect 9416 9608 9536 9636
rect 9600 9636 9628 9664
rect 9600 9608 9775 9636
rect 8941 9571 8999 9577
rect 8496 9540 8616 9568
rect 8389 9531 8447 9537
rect 8036 9500 8064 9528
rect 8404 9500 8432 9531
rect 8036 9472 8432 9500
rect 8588 9432 8616 9540
rect 8941 9537 8953 9571
rect 8987 9568 8999 9571
rect 9416 9568 9444 9608
rect 9747 9577 9775 9608
rect 9473 9571 9531 9577
rect 9473 9568 9485 9571
rect 8987 9540 9352 9568
rect 9416 9540 9485 9568
rect 8987 9537 8999 9540
rect 8941 9531 8999 9537
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 8711 9472 9229 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9217 9463 9275 9469
rect 8938 9432 8944 9444
rect 8588 9404 8944 9432
rect 8938 9392 8944 9404
rect 8996 9392 9002 9444
rect 4430 9324 4436 9376
rect 4488 9324 4494 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 7064 9336 8769 9364
rect 7064 9324 7070 9336
rect 8757 9333 8769 9336
rect 8803 9333 8815 9367
rect 9324 9364 9352 9540
rect 9473 9537 9485 9540
rect 9519 9537 9531 9571
rect 9473 9531 9531 9537
rect 9585 9571 9643 9577
rect 9585 9537 9597 9571
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 9698 9571 9775 9577
rect 9698 9537 9710 9571
rect 9744 9540 9775 9571
rect 9744 9537 9756 9540
rect 9698 9531 9756 9537
rect 9600 9500 9628 9531
rect 9858 9528 9864 9580
rect 9916 9528 9922 9580
rect 9968 9577 9996 9676
rect 10042 9664 10048 9716
rect 10100 9664 10106 9716
rect 10318 9664 10324 9716
rect 10376 9704 10382 9716
rect 10376 9676 11376 9704
rect 10376 9664 10382 9676
rect 10502 9596 10508 9648
rect 10560 9596 10566 9648
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 10689 9639 10747 9645
rect 10689 9636 10701 9639
rect 10652 9608 10701 9636
rect 10652 9596 10658 9608
rect 10689 9605 10701 9608
rect 10735 9605 10747 9639
rect 10689 9599 10747 9605
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11348 9636 11376 9676
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 11517 9707 11575 9713
rect 11517 9704 11529 9707
rect 11480 9676 11529 9704
rect 11480 9664 11486 9676
rect 11517 9673 11529 9676
rect 11563 9673 11575 9707
rect 11517 9667 11575 9673
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 11664 9676 12756 9704
rect 11664 9664 11670 9676
rect 11698 9636 11704 9648
rect 11112 9608 11192 9636
rect 11348 9608 11704 9636
rect 11112 9596 11118 9608
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10520 9568 10548 9596
rect 10459 9540 10548 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10226 9500 10232 9512
rect 9600 9472 10232 9500
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 10520 9500 10548 9540
rect 10870 9528 10876 9580
rect 10928 9528 10934 9580
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 11164 9577 11192 9608
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 12618 9636 12624 9648
rect 11900 9608 12624 9636
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 11333 9571 11391 9577
rect 11333 9568 11345 9571
rect 11296 9540 11345 9568
rect 11296 9528 11302 9540
rect 11333 9537 11345 9540
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11790 9568 11796 9580
rect 11480 9540 11796 9568
rect 11480 9528 11486 9540
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 11900 9577 11928 9608
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 12728 9645 12756 9676
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13541 9707 13599 9713
rect 13541 9704 13553 9707
rect 13136 9676 13553 9704
rect 13136 9664 13142 9676
rect 13541 9673 13553 9676
rect 13587 9673 13599 9707
rect 13541 9667 13599 9673
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17586 9704 17592 9716
rect 17276 9676 17592 9704
rect 17276 9664 17282 9676
rect 17586 9664 17592 9676
rect 17644 9704 17650 9716
rect 17865 9707 17923 9713
rect 17865 9704 17877 9707
rect 17644 9676 17877 9704
rect 17644 9664 17650 9676
rect 17865 9673 17877 9676
rect 17911 9673 17923 9707
rect 22925 9707 22983 9713
rect 17865 9667 17923 9673
rect 21560 9676 21772 9704
rect 12713 9639 12771 9645
rect 12713 9605 12725 9639
rect 12759 9605 12771 9639
rect 12713 9599 12771 9605
rect 13170 9596 13176 9648
rect 13228 9596 13234 9648
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 13320 9608 13461 9636
rect 13320 9596 13326 9608
rect 13449 9605 13461 9608
rect 13495 9605 13507 9639
rect 13449 9599 13507 9605
rect 14553 9639 14611 9645
rect 14553 9605 14565 9639
rect 14599 9636 14611 9639
rect 14642 9636 14648 9648
rect 14599 9608 14648 9636
rect 14599 9605 14611 9608
rect 14553 9599 14611 9605
rect 14642 9596 14648 9608
rect 14700 9596 14706 9648
rect 14844 9608 15424 9636
rect 13174 9593 13232 9596
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 11900 9500 11928 9531
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 12137 9571 12195 9577
rect 12137 9537 12149 9571
rect 12183 9568 12195 9571
rect 12434 9568 12440 9580
rect 12183 9566 12204 9568
rect 12360 9566 12440 9568
rect 12183 9540 12440 9566
rect 12183 9538 12388 9540
rect 12183 9537 12195 9538
rect 12137 9531 12195 9537
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 12526 9528 12532 9580
rect 12584 9528 12590 9580
rect 13174 9559 13186 9593
rect 13220 9559 13232 9593
rect 13174 9553 13232 9559
rect 13354 9528 13360 9580
rect 13412 9528 13418 9580
rect 13538 9528 13544 9580
rect 13596 9528 13602 9580
rect 13722 9528 13728 9580
rect 13780 9528 13786 9580
rect 14844 9577 14872 9608
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 10520 9472 11928 9500
rect 12253 9503 12311 9509
rect 12253 9492 12265 9503
rect 12084 9469 12265 9492
rect 12299 9469 12311 9503
rect 13372 9500 13400 9528
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 13372 9472 13461 9500
rect 12084 9464 12311 9469
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 11057 9435 11115 9441
rect 11057 9432 11069 9435
rect 9456 9404 11069 9432
rect 9456 9392 9462 9404
rect 11057 9401 11069 9404
rect 11103 9401 11115 9435
rect 11057 9395 11115 9401
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 12084 9432 12112 9464
rect 12253 9463 12311 9464
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 13449 9463 13507 9469
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 15120 9500 15148 9531
rect 15396 9509 15424 9608
rect 15470 9596 15476 9648
rect 15528 9596 15534 9648
rect 15749 9639 15807 9645
rect 15749 9605 15761 9639
rect 15795 9636 15807 9639
rect 15838 9636 15844 9648
rect 15795 9608 15844 9636
rect 15795 9605 15807 9608
rect 15749 9599 15807 9605
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17310 9636 17316 9648
rect 17083 9608 17316 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 17405 9639 17463 9645
rect 17405 9605 17417 9639
rect 17451 9636 17463 9639
rect 17982 9639 18040 9645
rect 17982 9636 17994 9639
rect 17451 9608 17994 9636
rect 17451 9605 17463 9608
rect 17405 9599 17463 9605
rect 17982 9605 17994 9608
rect 18028 9605 18040 9639
rect 17982 9599 18040 9605
rect 18138 9596 18144 9648
rect 18196 9596 18202 9648
rect 20993 9639 21051 9645
rect 20993 9605 21005 9639
rect 21039 9636 21051 9639
rect 21560 9636 21588 9676
rect 21744 9648 21772 9676
rect 21039 9608 21588 9636
rect 21039 9605 21051 9608
rect 20993 9599 21051 9605
rect 21634 9596 21640 9648
rect 21692 9596 21698 9648
rect 21726 9596 21732 9648
rect 21784 9596 21790 9648
rect 21818 9634 21824 9686
rect 21876 9634 21882 9686
rect 22925 9673 22937 9707
rect 22971 9704 22983 9707
rect 23106 9704 23112 9716
rect 22971 9676 23112 9704
rect 22971 9673 22983 9676
rect 22925 9667 22983 9673
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 27890 9664 27896 9716
rect 27948 9704 27954 9716
rect 28810 9704 28816 9716
rect 27948 9676 28816 9704
rect 27948 9664 27954 9676
rect 28810 9664 28816 9676
rect 28868 9664 28874 9716
rect 15488 9568 15516 9596
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15488 9540 16037 9568
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 17221 9571 17279 9577
rect 17221 9537 17233 9571
rect 17267 9568 17279 9571
rect 18156 9568 18184 9596
rect 17267 9540 18184 9568
rect 17267 9537 17279 9540
rect 17221 9531 17279 9537
rect 14792 9472 15148 9500
rect 15381 9503 15439 9509
rect 14792 9460 14798 9472
rect 15381 9469 15393 9503
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 11756 9404 12112 9432
rect 11756 9392 11762 9404
rect 15010 9392 15016 9444
rect 15068 9392 15074 9444
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 15396 9432 15424 9463
rect 15746 9460 15752 9512
rect 15804 9460 15810 9512
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 16132 9500 16160 9531
rect 18414 9528 18420 9580
rect 18472 9528 18478 9580
rect 19978 9568 19984 9580
rect 19826 9540 19984 9568
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 20548 9540 20729 9568
rect 20548 9512 20576 9540
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 21075 9571 21133 9577
rect 21075 9568 21087 9571
rect 20717 9531 20775 9537
rect 21008 9540 21087 9568
rect 15896 9472 16160 9500
rect 15896 9460 15902 9472
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 17497 9503 17555 9509
rect 17497 9500 17509 9503
rect 17460 9472 17509 9500
rect 17460 9460 17466 9472
rect 17497 9469 17509 9472
rect 17543 9469 17555 9503
rect 17497 9463 17555 9469
rect 17773 9503 17831 9509
rect 17773 9469 17785 9503
rect 17819 9469 17831 9503
rect 17773 9463 17831 9469
rect 15160 9404 15424 9432
rect 15160 9392 15166 9404
rect 11238 9364 11244 9376
rect 9324 9336 11244 9364
rect 8757 9327 8815 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 12345 9367 12403 9373
rect 12345 9333 12357 9367
rect 12391 9364 12403 9367
rect 12434 9364 12440 9376
rect 12391 9336 12440 9364
rect 12391 9333 12403 9336
rect 12345 9327 12403 9333
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 13044 9336 13277 9364
rect 13044 9324 13050 9336
rect 13265 9333 13277 9336
rect 13311 9333 13323 9367
rect 13265 9327 13323 9333
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 14553 9367 14611 9373
rect 14553 9364 14565 9367
rect 14516 9336 14565 9364
rect 14516 9324 14522 9336
rect 14553 9333 14565 9336
rect 14599 9364 14611 9367
rect 15194 9364 15200 9376
rect 14599 9336 15200 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 15654 9324 15660 9376
rect 15712 9324 15718 9376
rect 15933 9367 15991 9373
rect 15933 9333 15945 9367
rect 15979 9364 15991 9367
rect 16114 9364 16120 9376
rect 15979 9336 16120 9364
rect 15979 9333 15991 9336
rect 15933 9327 15991 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16206 9324 16212 9376
rect 16264 9324 16270 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 17788 9364 17816 9463
rect 18690 9460 18696 9512
rect 18748 9460 18754 9512
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 20162 9500 20168 9512
rect 19116 9472 20168 9500
rect 19116 9460 19122 9472
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 20530 9460 20536 9512
rect 20588 9460 20594 9512
rect 21008 9509 21036 9540
rect 21075 9537 21087 9540
rect 21121 9537 21133 9571
rect 21075 9531 21133 9537
rect 21174 9528 21180 9580
rect 21232 9528 21238 9580
rect 21358 9528 21364 9580
rect 21416 9528 21422 9580
rect 21836 9577 21864 9634
rect 22554 9596 22560 9648
rect 22612 9636 22618 9648
rect 23385 9639 23443 9645
rect 23385 9636 23397 9639
rect 22612 9608 23397 9636
rect 22612 9596 22618 9608
rect 23385 9605 23397 9608
rect 23431 9605 23443 9639
rect 23385 9599 23443 9605
rect 26510 9596 26516 9648
rect 26568 9636 26574 9648
rect 27433 9639 27491 9645
rect 27433 9636 27445 9639
rect 26568 9608 27445 9636
rect 26568 9596 26574 9608
rect 27433 9605 27445 9608
rect 27479 9605 27491 9639
rect 27433 9599 27491 9605
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9568 21511 9571
rect 21821 9571 21879 9577
rect 21499 9540 21588 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 20993 9503 21051 9509
rect 20993 9500 21005 9503
rect 20916 9472 21005 9500
rect 19886 9392 19892 9444
rect 19944 9392 19950 9444
rect 17552 9336 17816 9364
rect 17552 9324 17558 9336
rect 18138 9324 18144 9376
rect 18196 9324 18202 9376
rect 19904 9364 19932 9392
rect 20916 9376 20944 9472
rect 20993 9469 21005 9472
rect 21039 9469 21051 9503
rect 21560 9500 21588 9540
rect 21821 9537 21833 9571
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9568 23351 9571
rect 23845 9571 23903 9577
rect 23845 9568 23857 9571
rect 23339 9540 23857 9568
rect 23339 9537 23351 9540
rect 23293 9531 23351 9537
rect 23845 9537 23857 9540
rect 23891 9537 23903 9571
rect 23845 9531 23903 9537
rect 21560 9472 21934 9500
rect 20993 9463 21051 9469
rect 21906 9441 21934 9472
rect 22002 9460 22008 9512
rect 22060 9460 22066 9512
rect 21891 9435 21949 9441
rect 21891 9401 21903 9435
rect 21937 9401 21949 9435
rect 22204 9432 22232 9531
rect 24394 9528 24400 9580
rect 24452 9528 24458 9580
rect 26421 9571 26479 9577
rect 26421 9537 26433 9571
rect 26467 9568 26479 9571
rect 27341 9571 27399 9577
rect 26467 9540 27016 9568
rect 26467 9537 26479 9540
rect 26421 9531 26479 9537
rect 22278 9460 22284 9512
rect 22336 9500 22342 9512
rect 23569 9503 23627 9509
rect 23569 9500 23581 9503
rect 22336 9472 23581 9500
rect 22336 9460 22342 9472
rect 23569 9469 23581 9472
rect 23615 9500 23627 9503
rect 25038 9500 25044 9512
rect 23615 9472 25044 9500
rect 23615 9469 23627 9472
rect 23569 9463 23627 9469
rect 25038 9460 25044 9472
rect 25096 9460 25102 9512
rect 22554 9432 22560 9444
rect 22204 9404 22560 9432
rect 21891 9395 21949 9401
rect 22554 9392 22560 9404
rect 22612 9392 22618 9444
rect 26988 9441 27016 9540
rect 27341 9537 27353 9571
rect 27387 9568 27399 9571
rect 27798 9568 27804 9580
rect 27387 9540 27804 9568
rect 27387 9537 27399 9540
rect 27341 9531 27399 9537
rect 27798 9528 27804 9540
rect 27856 9528 27862 9580
rect 29546 9528 29552 9580
rect 29604 9568 29610 9580
rect 29641 9571 29699 9577
rect 29641 9568 29653 9571
rect 29604 9540 29653 9568
rect 29604 9528 29610 9540
rect 29641 9537 29653 9540
rect 29687 9537 29699 9571
rect 29641 9531 29699 9537
rect 30834 9528 30840 9580
rect 30892 9568 30898 9580
rect 31113 9571 31171 9577
rect 31113 9568 31125 9571
rect 30892 9540 31125 9568
rect 30892 9528 30898 9540
rect 31113 9537 31125 9540
rect 31159 9568 31171 9571
rect 31662 9568 31668 9580
rect 31159 9540 31668 9568
rect 31159 9537 31171 9540
rect 31113 9531 31171 9537
rect 31662 9528 31668 9540
rect 31720 9528 31726 9580
rect 27154 9460 27160 9512
rect 27212 9500 27218 9512
rect 27522 9500 27528 9512
rect 27212 9472 27528 9500
rect 27212 9460 27218 9472
rect 27522 9460 27528 9472
rect 27580 9460 27586 9512
rect 29914 9460 29920 9512
rect 29972 9460 29978 9512
rect 31294 9460 31300 9512
rect 31352 9500 31358 9512
rect 31389 9503 31447 9509
rect 31389 9500 31401 9503
rect 31352 9472 31401 9500
rect 31352 9460 31358 9472
rect 31389 9469 31401 9472
rect 31435 9469 31447 9503
rect 31389 9463 31447 9469
rect 26973 9435 27031 9441
rect 23676 9404 26556 9432
rect 20622 9364 20628 9376
rect 19904 9336 20628 9364
rect 20622 9324 20628 9336
rect 20680 9364 20686 9376
rect 20809 9367 20867 9373
rect 20809 9364 20821 9367
rect 20680 9336 20821 9364
rect 20680 9324 20686 9336
rect 20809 9333 20821 9336
rect 20855 9333 20867 9367
rect 20809 9327 20867 9333
rect 20898 9324 20904 9376
rect 20956 9324 20962 9376
rect 20990 9324 20996 9376
rect 21048 9364 21054 9376
rect 22097 9367 22155 9373
rect 22097 9364 22109 9367
rect 21048 9336 22109 9364
rect 21048 9324 21054 9336
rect 22097 9333 22109 9336
rect 22143 9364 22155 9367
rect 23676 9364 23704 9404
rect 26528 9376 26556 9404
rect 26973 9401 26985 9435
rect 27019 9401 27031 9435
rect 26973 9395 27031 9401
rect 30193 9435 30251 9441
rect 30193 9401 30205 9435
rect 30239 9432 30251 9435
rect 31110 9432 31116 9444
rect 30239 9404 31116 9432
rect 30239 9401 30251 9404
rect 30193 9395 30251 9401
rect 31110 9392 31116 9404
rect 31168 9392 31174 9444
rect 31478 9392 31484 9444
rect 31536 9432 31542 9444
rect 31665 9435 31723 9441
rect 31665 9432 31677 9435
rect 31536 9404 31677 9432
rect 31536 9392 31542 9404
rect 31665 9401 31677 9404
rect 31711 9401 31723 9435
rect 31665 9395 31723 9401
rect 22143 9336 23704 9364
rect 26237 9367 26295 9373
rect 22143 9333 22155 9336
rect 22097 9327 22155 9333
rect 26237 9333 26249 9367
rect 26283 9364 26295 9367
rect 26326 9364 26332 9376
rect 26283 9336 26332 9364
rect 26283 9333 26295 9336
rect 26237 9327 26295 9333
rect 26326 9324 26332 9336
rect 26384 9324 26390 9376
rect 26510 9324 26516 9376
rect 26568 9324 26574 9376
rect 29822 9324 29828 9376
rect 29880 9324 29886 9376
rect 31202 9324 31208 9376
rect 31260 9324 31266 9376
rect 1104 9274 34684 9296
rect 1104 9222 5147 9274
rect 5199 9222 5211 9274
rect 5263 9222 5275 9274
rect 5327 9222 5339 9274
rect 5391 9222 5403 9274
rect 5455 9222 13541 9274
rect 13593 9222 13605 9274
rect 13657 9222 13669 9274
rect 13721 9222 13733 9274
rect 13785 9222 13797 9274
rect 13849 9222 21935 9274
rect 21987 9222 21999 9274
rect 22051 9222 22063 9274
rect 22115 9222 22127 9274
rect 22179 9222 22191 9274
rect 22243 9222 30329 9274
rect 30381 9222 30393 9274
rect 30445 9222 30457 9274
rect 30509 9222 30521 9274
rect 30573 9222 30585 9274
rect 30637 9222 34684 9274
rect 1104 9200 34684 9222
rect 4430 9120 4436 9172
rect 4488 9120 4494 9172
rect 8018 9120 8024 9172
rect 8076 9120 8082 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8904 9132 9045 9160
rect 8904 9120 8910 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9582 9160 9588 9172
rect 9171 9132 9588 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 10229 9163 10287 9169
rect 10229 9129 10241 9163
rect 10275 9160 10287 9163
rect 10962 9160 10968 9172
rect 10275 9132 10968 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 11572 9132 11621 9160
rect 11572 9120 11578 9132
rect 11609 9129 11621 9132
rect 11655 9129 11667 9163
rect 11609 9123 11667 9129
rect 12342 9120 12348 9172
rect 12400 9120 12406 9172
rect 14458 9160 14464 9172
rect 14016 9132 14464 9160
rect 4448 8888 4476 9120
rect 8036 9024 8064 9120
rect 11241 9095 11299 9101
rect 11241 9061 11253 9095
rect 11287 9092 11299 9095
rect 12360 9092 12388 9120
rect 11287 9064 12388 9092
rect 11287 9061 11299 9064
rect 11241 9055 11299 9061
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8036 8996 9229 9024
rect 9217 8993 9229 8996
rect 9263 9024 9275 9027
rect 9490 9024 9496 9036
rect 9263 8996 9496 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9490 8984 9496 8996
rect 9548 9024 9554 9036
rect 9950 9024 9956 9036
rect 9548 8996 9956 9024
rect 9548 8984 9554 8996
rect 9950 8984 9956 8996
rect 10008 9024 10014 9036
rect 10008 8996 10364 9024
rect 10008 8984 10014 8996
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 10060 8965 10088 8996
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 10226 8916 10232 8968
rect 10284 8916 10290 8968
rect 10336 8956 10364 8996
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11204 8996 12296 9024
rect 11204 8984 11210 8996
rect 12268 8968 12296 8996
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 10336 8928 11437 8956
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 12250 8916 12256 8968
rect 12308 8916 12314 8968
rect 14016 8888 14044 9132
rect 14458 9120 14464 9132
rect 14516 9160 14522 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 14516 9132 14657 9160
rect 14516 9120 14522 9132
rect 14645 9129 14657 9132
rect 14691 9129 14703 9163
rect 14645 9123 14703 9129
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 15746 9160 15752 9172
rect 15335 9132 15752 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 16206 9120 16212 9172
rect 16264 9120 16270 9172
rect 16298 9120 16304 9172
rect 16356 9120 16362 9172
rect 16390 9120 16396 9172
rect 16448 9120 16454 9172
rect 17402 9120 17408 9172
rect 17460 9120 17466 9172
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 17635 9132 17724 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 15197 9095 15255 9101
rect 15197 9061 15209 9095
rect 15243 9061 15255 9095
rect 15197 9055 15255 9061
rect 15565 9095 15623 9101
rect 15565 9061 15577 9095
rect 15611 9092 15623 9095
rect 16224 9092 16252 9120
rect 15611 9064 16252 9092
rect 16316 9092 16344 9120
rect 16485 9095 16543 9101
rect 16485 9092 16497 9095
rect 16316 9064 16497 9092
rect 15611 9061 15623 9064
rect 15565 9055 15623 9061
rect 16485 9061 16497 9064
rect 16531 9061 16543 9095
rect 16485 9055 16543 9061
rect 15212 9024 15240 9055
rect 16114 9024 16120 9036
rect 15212 8996 16120 9024
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 14829 8959 14887 8965
rect 14829 8956 14841 8959
rect 14792 8928 14841 8956
rect 14792 8916 14798 8928
rect 14829 8925 14841 8928
rect 14875 8925 14887 8959
rect 14829 8919 14887 8925
rect 15013 8959 15071 8965
rect 15013 8925 15025 8959
rect 15059 8956 15071 8959
rect 15102 8956 15108 8968
rect 15059 8928 15108 8956
rect 15059 8925 15071 8928
rect 15013 8919 15071 8925
rect 4448 8860 14044 8888
rect 14553 8891 14611 8897
rect 14553 8857 14565 8891
rect 14599 8888 14611 8891
rect 14642 8888 14648 8900
rect 14599 8860 14648 8888
rect 14599 8857 14611 8860
rect 14553 8851 14611 8857
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 15028 8820 15056 8919
rect 15102 8916 15108 8928
rect 15160 8956 15166 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15160 8928 15485 8956
rect 15160 8916 15166 8928
rect 15473 8925 15485 8928
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 15562 8916 15568 8968
rect 15620 8956 15626 8968
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 15620 8928 15669 8956
rect 15620 8916 15626 8928
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 15657 8919 15715 8925
rect 15746 8916 15752 8968
rect 15804 8916 15810 8968
rect 16040 8965 16068 8996
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 15856 8928 15945 8956
rect 15856 8900 15884 8928
rect 15933 8925 15945 8928
rect 15979 8925 15991 8959
rect 15933 8919 15991 8925
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8925 16083 8959
rect 16025 8919 16083 8925
rect 16482 8916 16488 8968
rect 16540 8916 16546 8968
rect 15838 8848 15844 8900
rect 15896 8848 15902 8900
rect 16666 8888 16672 8900
rect 16224 8860 16672 8888
rect 13964 8792 15056 8820
rect 13964 8780 13970 8792
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 16224 8829 16252 8860
rect 16666 8848 16672 8860
rect 16724 8848 16730 8900
rect 17586 8829 17592 8832
rect 16117 8823 16175 8829
rect 16117 8820 16129 8823
rect 15712 8792 16129 8820
rect 15712 8780 15718 8792
rect 16117 8789 16129 8792
rect 16163 8789 16175 8823
rect 16117 8783 16175 8789
rect 16209 8823 16267 8829
rect 16209 8789 16221 8823
rect 16255 8789 16267 8823
rect 16209 8783 16267 8789
rect 17573 8823 17592 8829
rect 17573 8789 17585 8823
rect 17573 8783 17592 8789
rect 17586 8780 17592 8783
rect 17644 8780 17650 8832
rect 17696 8820 17724 9132
rect 18138 9120 18144 9172
rect 18196 9120 18202 9172
rect 18417 9163 18475 9169
rect 18417 9129 18429 9163
rect 18463 9160 18475 9163
rect 18690 9160 18696 9172
rect 18463 9132 18696 9160
rect 18463 9129 18475 9132
rect 18417 9123 18475 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 20898 9120 20904 9172
rect 20956 9120 20962 9172
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 21821 9163 21879 9169
rect 21821 9160 21833 9163
rect 21232 9132 21833 9160
rect 21232 9120 21238 9132
rect 21821 9129 21833 9132
rect 21867 9129 21879 9163
rect 21821 9123 21879 9129
rect 23569 9163 23627 9169
rect 23569 9129 23581 9163
rect 23615 9160 23627 9163
rect 23750 9160 23756 9172
rect 23615 9132 23756 9160
rect 23615 9129 23627 9132
rect 23569 9123 23627 9129
rect 18156 8956 18184 9120
rect 21100 9064 21956 9092
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 18156 8928 18245 8956
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21100 8965 21128 9064
rect 21928 9036 21956 9064
rect 21634 8984 21640 9036
rect 21692 9024 21698 9036
rect 21821 9027 21879 9033
rect 21821 9024 21833 9027
rect 21692 8996 21833 9024
rect 21692 8984 21698 8996
rect 21821 8993 21833 8996
rect 21867 8993 21879 9027
rect 21821 8987 21879 8993
rect 21910 8984 21916 9036
rect 21968 8984 21974 9036
rect 22370 8984 22376 9036
rect 22428 9024 22434 9036
rect 22428 8996 23520 9024
rect 22428 8984 22434 8996
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 20680 8928 21097 8956
rect 20680 8916 20686 8928
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21085 8919 21143 8925
rect 21266 8916 21272 8968
rect 21324 8916 21330 8968
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8956 21511 8959
rect 21652 8956 21680 8984
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21499 8928 21680 8956
rect 21963 8928 22017 8956
rect 21499 8925 21511 8928
rect 21453 8919 21511 8925
rect 22005 8925 22017 8928
rect 22051 8956 22063 8959
rect 22462 8956 22468 8968
rect 22051 8928 22468 8956
rect 22051 8925 22063 8928
rect 22005 8919 22063 8925
rect 17773 8891 17831 8897
rect 17773 8857 17785 8891
rect 17819 8888 17831 8891
rect 18046 8888 18052 8900
rect 17819 8860 18052 8888
rect 17819 8857 17831 8860
rect 17773 8851 17831 8857
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 20530 8888 20536 8900
rect 18156 8860 20536 8888
rect 18156 8832 18184 8860
rect 20530 8848 20536 8860
rect 20588 8888 20594 8900
rect 21177 8891 21235 8897
rect 21177 8888 21189 8891
rect 20588 8860 21189 8888
rect 20588 8848 20594 8860
rect 21177 8857 21189 8860
rect 21223 8857 21235 8891
rect 21284 8888 21312 8916
rect 21637 8891 21695 8897
rect 21637 8888 21649 8891
rect 21284 8860 21649 8888
rect 21177 8851 21235 8857
rect 21637 8857 21649 8860
rect 21683 8888 21695 8891
rect 21726 8888 21732 8900
rect 21683 8860 21732 8888
rect 21683 8857 21695 8860
rect 21637 8851 21695 8857
rect 18138 8820 18144 8832
rect 17696 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 21192 8820 21220 8851
rect 21726 8848 21732 8860
rect 21784 8848 21790 8900
rect 22020 8820 22048 8919
rect 22462 8916 22468 8928
rect 22520 8916 22526 8968
rect 23492 8965 23520 8996
rect 23477 8959 23535 8965
rect 23477 8925 23489 8959
rect 23523 8925 23535 8959
rect 23676 8956 23704 9132
rect 23750 9120 23756 9132
rect 23808 9160 23814 9172
rect 23808 9132 27568 9160
rect 23808 9120 23814 9132
rect 23753 9027 23811 9033
rect 23753 8993 23765 9027
rect 23799 9024 23811 9027
rect 24489 9027 24547 9033
rect 24489 9024 24501 9027
rect 23799 8996 24501 9024
rect 23799 8993 23811 8996
rect 23753 8987 23811 8993
rect 24489 8993 24501 8996
rect 24535 8993 24547 9027
rect 24489 8987 24547 8993
rect 26326 8984 26332 9036
rect 26384 8984 26390 9036
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 23676 8928 24409 8956
rect 23477 8919 23535 8925
rect 24397 8925 24409 8928
rect 24443 8925 24455 8959
rect 24397 8919 24455 8925
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 24949 8959 25007 8965
rect 24949 8956 24961 8959
rect 24627 8928 24961 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 24949 8925 24961 8928
rect 24995 8925 25007 8959
rect 24949 8919 25007 8925
rect 25593 8959 25651 8965
rect 25593 8925 25605 8959
rect 25639 8925 25651 8959
rect 25593 8919 25651 8925
rect 25608 8832 25636 8919
rect 26050 8916 26056 8968
rect 26108 8916 26114 8968
rect 27540 8956 27568 9132
rect 27798 9120 27804 9172
rect 27856 9120 27862 9172
rect 30834 9120 30840 9172
rect 30892 9120 30898 9172
rect 31021 9163 31079 9169
rect 31021 9129 31033 9163
rect 31067 9129 31079 9163
rect 31754 9160 31760 9172
rect 31021 9123 31079 9129
rect 31312 9132 31760 9160
rect 27816 9092 27844 9120
rect 31036 9092 31064 9123
rect 27816 9064 31064 9092
rect 28258 8984 28264 9036
rect 28316 8984 28322 9036
rect 27890 8956 27896 8968
rect 27540 8928 27896 8956
rect 27890 8916 27896 8928
rect 27948 8916 27954 8968
rect 28169 8959 28227 8965
rect 28169 8925 28181 8959
rect 28215 8925 28227 8959
rect 28276 8956 28304 8984
rect 28353 8959 28411 8965
rect 28353 8956 28365 8959
rect 28276 8928 28365 8956
rect 28169 8919 28227 8925
rect 28353 8925 28365 8928
rect 28399 8925 28411 8959
rect 28353 8919 28411 8925
rect 26602 8848 26608 8900
rect 26660 8888 26666 8900
rect 28184 8888 28212 8919
rect 28537 8891 28595 8897
rect 26660 8860 26818 8888
rect 28184 8860 28396 8888
rect 26660 8848 26666 8860
rect 28368 8832 28396 8860
rect 28537 8857 28549 8891
rect 28583 8888 28595 8891
rect 29822 8888 29828 8900
rect 28583 8860 29828 8888
rect 28583 8857 28595 8860
rect 28537 8851 28595 8857
rect 29822 8848 29828 8860
rect 29880 8848 29886 8900
rect 31036 8888 31064 9064
rect 31312 8965 31340 9132
rect 31754 9120 31760 9132
rect 31812 9120 31818 9172
rect 32030 9120 32036 9172
rect 32088 9120 32094 9172
rect 32214 9120 32220 9172
rect 32272 9160 32278 9172
rect 32677 9163 32735 9169
rect 32677 9160 32689 9163
rect 32272 9132 32689 9160
rect 32272 9120 32278 9132
rect 32677 9129 32689 9132
rect 32723 9129 32735 9163
rect 32677 9123 32735 9129
rect 31570 9052 31576 9104
rect 31628 9092 31634 9104
rect 32125 9095 32183 9101
rect 32125 9092 32137 9095
rect 31628 9064 32137 9092
rect 31628 9052 31634 9064
rect 32125 9061 32137 9064
rect 32171 9061 32183 9095
rect 32125 9055 32183 9061
rect 31662 8984 31668 9036
rect 31720 9024 31726 9036
rect 31941 9027 31999 9033
rect 31941 9024 31953 9027
rect 31720 8996 31953 9024
rect 31720 8984 31726 8996
rect 31941 8993 31953 8996
rect 31987 8993 31999 9027
rect 31941 8987 31999 8993
rect 32398 8984 32404 9036
rect 32456 9024 32462 9036
rect 33042 9024 33048 9036
rect 32456 8996 33048 9024
rect 32456 8984 32462 8996
rect 33042 8984 33048 8996
rect 33100 9024 33106 9036
rect 33229 9027 33287 9033
rect 33229 9024 33241 9027
rect 33100 8996 33241 9024
rect 33100 8984 33106 8996
rect 33229 8993 33241 8996
rect 33275 8993 33287 9027
rect 33229 8987 33287 8993
rect 31297 8959 31355 8965
rect 31297 8925 31309 8959
rect 31343 8925 31355 8959
rect 31849 8959 31907 8965
rect 31849 8956 31861 8959
rect 31297 8919 31355 8925
rect 31404 8928 31861 8956
rect 31404 8888 31432 8928
rect 31849 8925 31861 8928
rect 31895 8925 31907 8959
rect 31849 8919 31907 8925
rect 32217 8959 32275 8965
rect 32217 8925 32229 8959
rect 32263 8925 32275 8959
rect 32217 8919 32275 8925
rect 31036 8860 31432 8888
rect 31478 8848 31484 8900
rect 31536 8888 31542 8900
rect 32232 8888 32260 8919
rect 33137 8891 33195 8897
rect 33137 8888 33149 8891
rect 31536 8860 32260 8888
rect 32324 8860 33149 8888
rect 31536 8848 31542 8860
rect 21192 8792 22048 8820
rect 23750 8780 23756 8832
rect 23808 8780 23814 8832
rect 25590 8780 25596 8832
rect 25648 8820 25654 8832
rect 27338 8820 27344 8832
rect 25648 8792 27344 8820
rect 25648 8780 25654 8792
rect 27338 8780 27344 8792
rect 27396 8780 27402 8832
rect 28350 8780 28356 8832
rect 28408 8780 28414 8832
rect 28718 8780 28724 8832
rect 28776 8780 28782 8832
rect 31386 8780 31392 8832
rect 31444 8780 31450 8832
rect 31754 8780 31760 8832
rect 31812 8820 31818 8832
rect 32324 8820 32352 8860
rect 33137 8857 33149 8860
rect 33183 8857 33195 8891
rect 33137 8851 33195 8857
rect 31812 8792 32352 8820
rect 31812 8780 31818 8792
rect 33042 8780 33048 8832
rect 33100 8780 33106 8832
rect 1104 8730 34840 8752
rect 1104 8678 9344 8730
rect 9396 8678 9408 8730
rect 9460 8678 9472 8730
rect 9524 8678 9536 8730
rect 9588 8678 9600 8730
rect 9652 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 17930 8730
rect 17982 8678 17994 8730
rect 18046 8678 26132 8730
rect 26184 8678 26196 8730
rect 26248 8678 26260 8730
rect 26312 8678 26324 8730
rect 26376 8678 26388 8730
rect 26440 8678 34526 8730
rect 34578 8678 34590 8730
rect 34642 8678 34654 8730
rect 34706 8678 34718 8730
rect 34770 8678 34782 8730
rect 34834 8678 34840 8730
rect 1104 8656 34840 8678
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 16482 8616 16488 8628
rect 15804 8588 16488 8616
rect 15804 8576 15810 8588
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17368 8588 17509 8616
rect 17368 8576 17374 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 18984 8588 19748 8616
rect 17604 8480 17632 8576
rect 18984 8560 19012 8588
rect 18966 8508 18972 8560
rect 19024 8508 19030 8560
rect 19720 8557 19748 8588
rect 21358 8576 21364 8628
rect 21416 8576 21422 8628
rect 21910 8576 21916 8628
rect 21968 8616 21974 8628
rect 25225 8619 25283 8625
rect 21968 8588 23244 8616
rect 21968 8576 21974 8588
rect 19705 8551 19763 8557
rect 19475 8517 19533 8523
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 17604 8452 17693 8480
rect 17681 8449 17693 8452
rect 17727 8480 17739 8483
rect 18230 8480 18236 8492
rect 17727 8452 18236 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 19475 8483 19487 8517
rect 19521 8514 19533 8517
rect 19705 8517 19717 8551
rect 19751 8548 19763 8551
rect 21818 8548 21824 8560
rect 19751 8520 21824 8548
rect 19751 8517 19763 8520
rect 19521 8483 19548 8514
rect 19705 8511 19763 8517
rect 21818 8508 21824 8520
rect 21876 8508 21882 8560
rect 19475 8477 19548 8483
rect 17865 8415 17923 8421
rect 17865 8381 17877 8415
rect 17911 8412 17923 8415
rect 18046 8412 18052 8424
rect 17911 8384 18052 8412
rect 17911 8381 17923 8384
rect 17865 8375 17923 8381
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18248 8344 18276 8440
rect 19337 8347 19395 8353
rect 19337 8344 19349 8347
rect 18248 8316 19349 8344
rect 19337 8313 19349 8316
rect 19383 8313 19395 8347
rect 19520 8344 19548 8477
rect 20990 8440 20996 8492
rect 21048 8480 21054 8492
rect 21177 8483 21235 8489
rect 21177 8480 21189 8483
rect 21048 8452 21189 8480
rect 21048 8440 21054 8452
rect 21177 8449 21189 8452
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 21450 8480 21456 8492
rect 21407 8452 21456 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 21376 8344 21404 8443
rect 21450 8440 21456 8452
rect 21508 8480 21514 8492
rect 22554 8480 22560 8492
rect 21508 8452 22560 8480
rect 21508 8440 21514 8452
rect 22554 8440 22560 8452
rect 22612 8440 22618 8492
rect 23106 8440 23112 8492
rect 23164 8440 23170 8492
rect 23216 8489 23244 8588
rect 25225 8585 25237 8619
rect 25271 8616 25283 8619
rect 25590 8616 25596 8628
rect 25271 8588 25596 8616
rect 25271 8585 25283 8588
rect 25225 8579 25283 8585
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 28994 8616 29000 8628
rect 28736 8588 29000 8616
rect 26602 8508 26608 8560
rect 26660 8548 26666 8560
rect 28736 8548 28764 8588
rect 28994 8576 29000 8588
rect 29052 8616 29058 8628
rect 29052 8588 29776 8616
rect 29052 8576 29058 8588
rect 29748 8548 29776 8588
rect 29822 8576 29828 8628
rect 29880 8576 29886 8628
rect 29932 8588 32996 8616
rect 29932 8548 29960 8588
rect 32968 8560 32996 8588
rect 33042 8576 33048 8628
rect 33100 8576 33106 8628
rect 26660 8520 28842 8548
rect 29748 8520 29960 8548
rect 26660 8508 26666 8520
rect 31478 8508 31484 8560
rect 31536 8548 31542 8560
rect 31536 8520 31754 8548
rect 31536 8508 31542 8520
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 23474 8440 23480 8492
rect 23532 8440 23538 8492
rect 24854 8440 24860 8492
rect 24912 8440 24918 8492
rect 26050 8440 26056 8492
rect 26108 8440 26114 8492
rect 26510 8440 26516 8492
rect 26568 8480 26574 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26568 8452 26985 8480
rect 26568 8440 26574 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 30834 8440 30840 8492
rect 30892 8480 30898 8492
rect 31205 8483 31263 8489
rect 31205 8480 31217 8483
rect 30892 8452 31217 8480
rect 30892 8440 30898 8452
rect 31205 8449 31217 8452
rect 31251 8449 31263 8483
rect 31205 8443 31263 8449
rect 31386 8440 31392 8492
rect 31444 8440 31450 8492
rect 31726 8480 31754 8520
rect 32950 8508 32956 8560
rect 33008 8508 33014 8560
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 31726 8452 32321 8480
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 23750 8372 23756 8424
rect 23808 8372 23814 8424
rect 24946 8372 24952 8424
rect 25004 8412 25010 8424
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 25004 8384 25973 8412
rect 25004 8372 25010 8384
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 26068 8412 26096 8440
rect 27614 8412 27620 8424
rect 26068 8384 27620 8412
rect 25961 8375 26019 8381
rect 27614 8372 27620 8384
rect 27672 8412 27678 8424
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27672 8384 28089 8412
rect 27672 8372 27678 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 28350 8372 28356 8424
rect 28408 8372 28414 8424
rect 31018 8372 31024 8424
rect 31076 8412 31082 8424
rect 31570 8412 31576 8424
rect 31076 8384 31576 8412
rect 31076 8372 31082 8384
rect 31570 8372 31576 8384
rect 31628 8412 31634 8424
rect 32217 8415 32275 8421
rect 32217 8412 32229 8415
rect 31628 8384 32229 8412
rect 31628 8372 31634 8384
rect 32217 8381 32229 8384
rect 32263 8381 32275 8415
rect 32217 8375 32275 8381
rect 32677 8415 32735 8421
rect 32677 8381 32689 8415
rect 32723 8412 32735 8415
rect 33060 8412 33088 8576
rect 34333 8483 34391 8489
rect 34333 8449 34345 8483
rect 34379 8480 34391 8483
rect 34379 8452 34836 8480
rect 34379 8449 34391 8452
rect 34333 8443 34391 8449
rect 32723 8384 33088 8412
rect 32723 8381 32735 8384
rect 32677 8375 32735 8381
rect 34808 8356 34836 8452
rect 19337 8307 19395 8313
rect 19444 8316 21404 8344
rect 19242 8236 19248 8288
rect 19300 8276 19306 8288
rect 19444 8276 19472 8316
rect 21726 8304 21732 8356
rect 21784 8344 21790 8356
rect 22370 8344 22376 8356
rect 21784 8316 22376 8344
rect 21784 8304 21790 8316
rect 22370 8304 22376 8316
rect 22428 8304 22434 8356
rect 23293 8347 23351 8353
rect 23293 8313 23305 8347
rect 23339 8344 23351 8347
rect 23474 8344 23480 8356
rect 23339 8316 23480 8344
rect 23339 8313 23351 8316
rect 23293 8307 23351 8313
rect 23474 8304 23480 8316
rect 23532 8304 23538 8356
rect 26605 8347 26663 8353
rect 26605 8313 26617 8347
rect 26651 8344 26663 8347
rect 27706 8344 27712 8356
rect 26651 8316 27712 8344
rect 26651 8313 26663 8316
rect 26605 8307 26663 8313
rect 27706 8304 27712 8316
rect 27764 8304 27770 8356
rect 34790 8304 34796 8356
rect 34848 8304 34854 8356
rect 19300 8248 19472 8276
rect 19521 8279 19579 8285
rect 19300 8236 19306 8248
rect 19521 8245 19533 8279
rect 19567 8276 19579 8279
rect 20438 8276 20444 8288
rect 19567 8248 20444 8276
rect 19567 8245 19579 8248
rect 19521 8239 19579 8245
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 22922 8236 22928 8288
rect 22980 8236 22986 8288
rect 27062 8236 27068 8288
rect 27120 8236 27126 8288
rect 31297 8279 31355 8285
rect 31297 8245 31309 8279
rect 31343 8276 31355 8279
rect 31478 8276 31484 8288
rect 31343 8248 31484 8276
rect 31343 8245 31355 8248
rect 31297 8239 31355 8245
rect 31478 8236 31484 8248
rect 31536 8236 31542 8288
rect 34054 8236 34060 8288
rect 34112 8276 34118 8288
rect 34149 8279 34207 8285
rect 34149 8276 34161 8279
rect 34112 8248 34161 8276
rect 34112 8236 34118 8248
rect 34149 8245 34161 8248
rect 34195 8245 34207 8279
rect 34149 8239 34207 8245
rect 1104 8186 34684 8208
rect 1104 8134 5147 8186
rect 5199 8134 5211 8186
rect 5263 8134 5275 8186
rect 5327 8134 5339 8186
rect 5391 8134 5403 8186
rect 5455 8134 13541 8186
rect 13593 8134 13605 8186
rect 13657 8134 13669 8186
rect 13721 8134 13733 8186
rect 13785 8134 13797 8186
rect 13849 8134 21935 8186
rect 21987 8134 21999 8186
rect 22051 8134 22063 8186
rect 22115 8134 22127 8186
rect 22179 8134 22191 8186
rect 22243 8134 30329 8186
rect 30381 8134 30393 8186
rect 30445 8134 30457 8186
rect 30509 8134 30521 8186
rect 30573 8134 30585 8186
rect 30637 8134 34684 8186
rect 1104 8112 34684 8134
rect 13906 8032 13912 8084
rect 13964 8032 13970 8084
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 17218 8032 17224 8084
rect 17276 8072 17282 8084
rect 17586 8072 17592 8084
rect 17276 8044 17592 8072
rect 17276 8032 17282 8044
rect 17586 8032 17592 8044
rect 17644 8072 17650 8084
rect 19886 8072 19892 8084
rect 17644 8044 19892 8072
rect 17644 8032 17650 8044
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 22833 8075 22891 8081
rect 22833 8041 22845 8075
rect 22879 8072 22891 8075
rect 23106 8072 23112 8084
rect 22879 8044 23112 8072
rect 22879 8041 22891 8044
rect 22833 8035 22891 8041
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 27985 8075 28043 8081
rect 27172 8044 27384 8072
rect 17402 7964 17408 8016
rect 17460 8004 17466 8016
rect 17773 8007 17831 8013
rect 17773 8004 17785 8007
rect 17460 7976 17785 8004
rect 17460 7964 17466 7976
rect 17773 7973 17785 7976
rect 17819 7973 17831 8007
rect 17773 7967 17831 7973
rect 18230 7964 18236 8016
rect 18288 7964 18294 8016
rect 19702 7964 19708 8016
rect 19760 8004 19766 8016
rect 20165 8007 20223 8013
rect 20165 8004 20177 8007
rect 19760 7976 20177 8004
rect 19760 7964 19766 7976
rect 20165 7973 20177 7976
rect 20211 7973 20223 8007
rect 27172 8004 27200 8044
rect 20165 7967 20223 7973
rect 22066 7976 25268 8004
rect 12158 7896 12164 7948
rect 12216 7896 12222 7948
rect 17129 7939 17187 7945
rect 15580 7908 16252 7936
rect 15580 7877 15608 7908
rect 16224 7880 16252 7908
rect 17129 7905 17141 7939
rect 17175 7936 17187 7939
rect 17310 7936 17316 7948
rect 17175 7908 17316 7936
rect 17175 7905 17187 7908
rect 17129 7899 17187 7905
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 18248 7936 18276 7964
rect 19521 7939 19579 7945
rect 19521 7936 19533 7939
rect 18248 7908 19533 7936
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 16114 7828 16120 7880
rect 16172 7828 16178 7880
rect 16206 7828 16212 7880
rect 16264 7828 16270 7880
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7868 17463 7871
rect 17494 7868 17500 7880
rect 17451 7840 17500 7868
rect 17451 7837 17463 7840
rect 17405 7831 17463 7837
rect 17494 7828 17500 7840
rect 17552 7868 17558 7880
rect 18248 7877 18276 7908
rect 19521 7905 19533 7908
rect 19567 7905 19579 7939
rect 19521 7899 19579 7905
rect 19610 7896 19616 7948
rect 19668 7936 19674 7948
rect 22066 7936 22094 7976
rect 19668 7908 22094 7936
rect 19668 7896 19674 7908
rect 22278 7896 22284 7948
rect 22336 7936 22342 7948
rect 22646 7936 22652 7948
rect 22336 7908 22652 7936
rect 22336 7896 22342 7908
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 23474 7896 23480 7948
rect 23532 7936 23538 7948
rect 24857 7939 24915 7945
rect 24857 7936 24869 7939
rect 23532 7908 24869 7936
rect 23532 7896 23538 7908
rect 24857 7905 24869 7908
rect 24903 7905 24915 7939
rect 24857 7899 24915 7905
rect 24946 7896 24952 7948
rect 25004 7896 25010 7948
rect 25240 7945 25268 7976
rect 25884 7976 27200 8004
rect 27356 8004 27384 8044
rect 27985 8041 27997 8075
rect 28031 8072 28043 8075
rect 28350 8072 28356 8084
rect 28031 8044 28356 8072
rect 28031 8041 28043 8044
rect 27985 8035 28043 8041
rect 28350 8032 28356 8044
rect 28408 8032 28414 8084
rect 30837 8075 30895 8081
rect 30837 8041 30849 8075
rect 30883 8072 30895 8075
rect 31386 8072 31392 8084
rect 30883 8044 31392 8072
rect 30883 8041 30895 8044
rect 30837 8035 30895 8041
rect 31386 8032 31392 8044
rect 31444 8032 31450 8084
rect 32585 8007 32643 8013
rect 27356 7976 31754 8004
rect 25884 7945 25912 7976
rect 25041 7939 25099 7945
rect 25041 7905 25053 7939
rect 25087 7905 25099 7939
rect 25041 7899 25099 7905
rect 25225 7939 25283 7945
rect 25225 7905 25237 7939
rect 25271 7905 25283 7939
rect 25225 7899 25283 7905
rect 25869 7939 25927 7945
rect 25869 7905 25881 7939
rect 25915 7905 25927 7939
rect 25869 7899 25927 7905
rect 26421 7939 26479 7945
rect 26421 7905 26433 7939
rect 26467 7905 26479 7939
rect 26421 7899 26479 7905
rect 26513 7939 26571 7945
rect 26513 7905 26525 7939
rect 26559 7936 26571 7939
rect 27062 7936 27068 7948
rect 26559 7908 27068 7936
rect 26559 7905 26571 7908
rect 26513 7899 26571 7905
rect 18233 7871 18291 7877
rect 17552 7840 18000 7868
rect 17552 7828 17558 7840
rect 12434 7760 12440 7812
rect 12492 7760 12498 7812
rect 13906 7800 13912 7812
rect 13662 7772 13912 7800
rect 13906 7760 13912 7772
rect 13964 7760 13970 7812
rect 15841 7803 15899 7809
rect 15841 7769 15853 7803
rect 15887 7800 15899 7803
rect 16390 7800 16396 7812
rect 15887 7772 16396 7800
rect 15887 7769 15899 7772
rect 15841 7763 15899 7769
rect 16390 7760 16396 7772
rect 16448 7760 16454 7812
rect 17614 7803 17672 7809
rect 17614 7769 17626 7803
rect 17660 7800 17672 7803
rect 17865 7803 17923 7809
rect 17865 7800 17877 7803
rect 17660 7772 17877 7800
rect 17660 7769 17672 7772
rect 17614 7763 17672 7769
rect 17865 7769 17877 7772
rect 17911 7769 17923 7803
rect 17865 7763 17923 7769
rect 15657 7735 15715 7741
rect 15657 7701 15669 7735
rect 15703 7732 15715 7735
rect 16025 7735 16083 7741
rect 16025 7732 16037 7735
rect 15703 7704 16037 7732
rect 15703 7701 15715 7704
rect 15657 7695 15715 7701
rect 16025 7701 16037 7704
rect 16071 7701 16083 7735
rect 16025 7695 16083 7701
rect 17494 7692 17500 7744
rect 17552 7692 17558 7744
rect 17972 7732 18000 7840
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 19024 7840 20392 7868
rect 19024 7828 19030 7840
rect 18046 7760 18052 7812
rect 18104 7800 18110 7812
rect 18782 7800 18788 7812
rect 18104 7772 18788 7800
rect 18104 7760 18110 7772
rect 18782 7760 18788 7772
rect 18840 7760 18846 7812
rect 20006 7803 20064 7809
rect 20006 7769 20018 7803
rect 20052 7800 20064 7803
rect 20257 7803 20315 7809
rect 20257 7800 20269 7803
rect 20052 7772 20269 7800
rect 20052 7769 20064 7772
rect 20006 7763 20064 7769
rect 20257 7769 20269 7772
rect 20303 7769 20315 7803
rect 20364 7800 20392 7840
rect 20438 7828 20444 7880
rect 20496 7828 20502 7880
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 20763 7840 21496 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 20625 7803 20683 7809
rect 20625 7800 20637 7803
rect 20364 7772 20637 7800
rect 20257 7763 20315 7769
rect 20625 7769 20637 7772
rect 20671 7769 20683 7803
rect 20625 7763 20683 7769
rect 21468 7744 21496 7840
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 24964 7868 24992 7896
rect 23808 7840 24992 7868
rect 25056 7868 25084 7899
rect 26436 7868 26464 7899
rect 27062 7896 27068 7908
rect 27120 7896 27126 7948
rect 27154 7896 27160 7948
rect 27212 7896 27218 7948
rect 27890 7896 27896 7948
rect 27948 7936 27954 7948
rect 28353 7939 28411 7945
rect 28353 7936 28365 7939
rect 27948 7908 28365 7936
rect 27948 7896 27954 7908
rect 28353 7905 28365 7908
rect 28399 7905 28411 7939
rect 28353 7899 28411 7905
rect 28442 7896 28448 7948
rect 28500 7896 28506 7948
rect 31726 7936 31754 7976
rect 32585 7973 32597 8007
rect 32631 7973 32643 8007
rect 32585 7967 32643 7973
rect 32600 7936 32628 7967
rect 31726 7908 32628 7936
rect 34054 7896 34060 7948
rect 34112 7896 34118 7948
rect 27172 7868 27200 7896
rect 27246 7877 27252 7880
rect 25056 7840 27200 7868
rect 23808 7828 23814 7840
rect 27241 7831 27252 7877
rect 27304 7868 27310 7880
rect 27304 7840 27341 7868
rect 27246 7828 27252 7831
rect 27304 7828 27310 7840
rect 27706 7828 27712 7880
rect 27764 7868 27770 7880
rect 28169 7871 28227 7877
rect 28169 7868 28181 7871
rect 27764 7840 28181 7868
rect 27764 7828 27770 7840
rect 28169 7837 28181 7840
rect 28215 7837 28227 7871
rect 28169 7831 28227 7837
rect 28534 7828 28540 7880
rect 28592 7828 28598 7880
rect 28718 7828 28724 7880
rect 28776 7828 28782 7880
rect 32950 7828 32956 7880
rect 33008 7828 33014 7880
rect 34330 7828 34336 7880
rect 34388 7828 34394 7880
rect 22465 7803 22523 7809
rect 22465 7769 22477 7803
rect 22511 7800 22523 7803
rect 23109 7803 23167 7809
rect 23109 7800 23121 7803
rect 22511 7772 23121 7800
rect 22511 7769 22523 7772
rect 22465 7763 22523 7769
rect 23109 7769 23121 7772
rect 23155 7769 23167 7803
rect 23109 7763 23167 7769
rect 26605 7803 26663 7809
rect 26605 7769 26617 7803
rect 26651 7800 26663 7803
rect 27798 7800 27804 7812
rect 26651 7772 27804 7800
rect 26651 7769 26663 7772
rect 26605 7763 26663 7769
rect 27798 7760 27804 7772
rect 27856 7760 27862 7812
rect 29730 7760 29736 7812
rect 29788 7800 29794 7812
rect 30653 7803 30711 7809
rect 30653 7800 30665 7803
rect 29788 7772 30665 7800
rect 29788 7760 29794 7772
rect 30653 7769 30665 7772
rect 30699 7769 30711 7803
rect 30653 7763 30711 7769
rect 31294 7760 31300 7812
rect 31352 7760 31358 7812
rect 19794 7732 19800 7744
rect 17972 7704 19800 7732
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 19886 7692 19892 7744
rect 19944 7692 19950 7744
rect 21450 7692 21456 7744
rect 21508 7692 21514 7744
rect 21634 7692 21640 7744
rect 21692 7732 21698 7744
rect 22373 7735 22431 7741
rect 22373 7732 22385 7735
rect 21692 7704 22385 7732
rect 21692 7692 21698 7704
rect 22373 7701 22385 7704
rect 22419 7701 22431 7735
rect 22373 7695 22431 7701
rect 24394 7692 24400 7744
rect 24452 7692 24458 7744
rect 24762 7692 24768 7744
rect 24820 7692 24826 7744
rect 26970 7692 26976 7744
rect 27028 7692 27034 7744
rect 27062 7692 27068 7744
rect 27120 7692 27126 7744
rect 30834 7692 30840 7744
rect 30892 7741 30898 7744
rect 30892 7735 30911 7741
rect 30899 7701 30911 7735
rect 30892 7695 30911 7701
rect 31021 7735 31079 7741
rect 31021 7701 31033 7735
rect 31067 7732 31079 7735
rect 31312 7732 31340 7760
rect 31067 7704 31340 7732
rect 31067 7701 31079 7704
rect 31021 7695 31079 7701
rect 30892 7692 30898 7695
rect 1104 7642 34840 7664
rect 1104 7590 9344 7642
rect 9396 7590 9408 7642
rect 9460 7590 9472 7642
rect 9524 7590 9536 7642
rect 9588 7590 9600 7642
rect 9652 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 17930 7642
rect 17982 7590 17994 7642
rect 18046 7590 26132 7642
rect 26184 7590 26196 7642
rect 26248 7590 26260 7642
rect 26312 7590 26324 7642
rect 26376 7590 26388 7642
rect 26440 7590 34526 7642
rect 34578 7590 34590 7642
rect 34642 7590 34654 7642
rect 34706 7590 34718 7642
rect 34770 7590 34782 7642
rect 34834 7590 34840 7642
rect 1104 7568 34840 7590
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 12434 7528 12440 7540
rect 11379 7500 12440 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 15838 7528 15844 7540
rect 15212 7500 15844 7528
rect 8573 7463 8631 7469
rect 8573 7429 8585 7463
rect 8619 7460 8631 7463
rect 12621 7463 12679 7469
rect 12621 7460 12633 7463
rect 8619 7432 12633 7460
rect 8619 7429 8631 7432
rect 8573 7423 8631 7429
rect 12621 7429 12633 7432
rect 12667 7429 12679 7463
rect 13906 7460 13912 7472
rect 13846 7432 13912 7460
rect 12621 7423 12679 7429
rect 13906 7420 13912 7432
rect 13964 7460 13970 7472
rect 14826 7460 14832 7472
rect 13964 7432 14832 7460
rect 13964 7420 13970 7432
rect 14826 7420 14832 7432
rect 14884 7460 14890 7472
rect 15212 7460 15240 7500
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 16390 7528 16396 7540
rect 16347 7500 16396 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 16666 7488 16672 7540
rect 16724 7528 16730 7540
rect 16761 7531 16819 7537
rect 16761 7528 16773 7531
rect 16724 7500 16773 7528
rect 16724 7488 16730 7500
rect 16761 7497 16773 7500
rect 16807 7497 16819 7531
rect 16761 7491 16819 7497
rect 17402 7488 17408 7540
rect 17460 7488 17466 7540
rect 18966 7488 18972 7540
rect 19024 7488 19030 7540
rect 19702 7488 19708 7540
rect 19760 7488 19766 7540
rect 19797 7531 19855 7537
rect 19797 7497 19809 7531
rect 19843 7497 19855 7531
rect 19797 7491 19855 7497
rect 14884 7432 15318 7460
rect 14884 7420 14890 7432
rect 7926 7284 7932 7336
rect 7984 7284 7990 7336
rect 10686 7284 10692 7336
rect 10744 7284 10750 7336
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 12216 7296 12357 7324
rect 12216 7284 12222 7296
rect 12345 7293 12357 7296
rect 12391 7324 12403 7327
rect 13262 7324 13268 7336
rect 12391 7296 13268 7324
rect 12391 7293 12403 7296
rect 12345 7287 12403 7293
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 13924 7324 13952 7420
rect 14550 7352 14556 7404
rect 14608 7352 14614 7404
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 16669 7395 16727 7401
rect 16669 7392 16681 7395
rect 16264 7364 16681 7392
rect 16264 7352 16270 7364
rect 16669 7361 16681 7364
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7361 16911 7395
rect 17420 7392 17448 7488
rect 18984 7460 19012 7488
rect 18800 7432 19012 7460
rect 17589 7395 17647 7401
rect 17589 7392 17601 7395
rect 17420 7364 17601 7392
rect 16853 7355 16911 7361
rect 17589 7361 17601 7364
rect 17635 7361 17647 7395
rect 17589 7355 17647 7361
rect 13412 7296 13952 7324
rect 14829 7327 14887 7333
rect 13412 7284 13418 7296
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 14875 7296 16068 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 16040 7256 16068 7296
rect 16114 7284 16120 7336
rect 16172 7324 16178 7336
rect 16868 7324 16896 7355
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 18414 7352 18420 7404
rect 18472 7352 18478 7404
rect 18800 7401 18828 7432
rect 19242 7420 19248 7472
rect 19300 7420 19306 7472
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 18966 7352 18972 7404
rect 19024 7392 19030 7404
rect 19260 7392 19288 7420
rect 19024 7364 19288 7392
rect 19613 7395 19671 7401
rect 19024 7352 19030 7364
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 19720 7392 19748 7488
rect 19812 7460 19840 7491
rect 20438 7488 20444 7540
rect 20496 7528 20502 7540
rect 21634 7528 21640 7540
rect 20496 7500 21640 7528
rect 20496 7488 20502 7500
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 22922 7528 22928 7540
rect 22204 7500 22928 7528
rect 20165 7463 20223 7469
rect 20165 7460 20177 7463
rect 19812 7432 20177 7460
rect 20165 7429 20177 7432
rect 20211 7429 20223 7463
rect 22094 7460 22100 7472
rect 21390 7432 22100 7460
rect 20165 7423 20223 7429
rect 22094 7420 22100 7432
rect 22152 7420 22158 7472
rect 22204 7469 22232 7500
rect 22922 7488 22928 7500
rect 22980 7488 22986 7540
rect 23661 7531 23719 7537
rect 23661 7497 23673 7531
rect 23707 7528 23719 7531
rect 23750 7528 23756 7540
rect 23707 7500 23756 7528
rect 23707 7497 23719 7500
rect 23661 7491 23719 7497
rect 23750 7488 23756 7500
rect 23808 7488 23814 7540
rect 24394 7488 24400 7540
rect 24452 7488 24458 7540
rect 24762 7488 24768 7540
rect 24820 7528 24826 7540
rect 26145 7531 26203 7537
rect 26145 7528 26157 7531
rect 24820 7500 26157 7528
rect 24820 7488 24826 7500
rect 26145 7497 26157 7500
rect 26191 7497 26203 7531
rect 26145 7491 26203 7497
rect 22189 7463 22247 7469
rect 22189 7429 22201 7463
rect 22235 7429 22247 7463
rect 24412 7460 24440 7488
rect 22189 7423 22247 7429
rect 24136 7432 24440 7460
rect 23750 7392 23756 7404
rect 19659 7364 19748 7392
rect 23322 7378 23756 7392
rect 23308 7364 23756 7378
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 18248 7324 18276 7352
rect 16172 7296 18276 7324
rect 18432 7324 18460 7352
rect 19242 7324 19248 7336
rect 18432 7296 19248 7324
rect 16172 7284 16178 7296
rect 19242 7284 19248 7296
rect 19300 7324 19306 7336
rect 19889 7327 19947 7333
rect 19889 7324 19901 7327
rect 19300 7296 19901 7324
rect 19300 7284 19306 7296
rect 19889 7293 19901 7296
rect 19935 7324 19947 7327
rect 21913 7327 21971 7333
rect 21913 7324 21925 7327
rect 19935 7296 21925 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 21913 7293 21925 7296
rect 21959 7293 21971 7327
rect 21913 7287 21971 7293
rect 19610 7256 19616 7268
rect 16040 7228 19616 7256
rect 19610 7216 19616 7228
rect 19668 7216 19674 7268
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 16022 7188 16028 7200
rect 14139 7160 16028 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 17402 7148 17408 7200
rect 17460 7148 17466 7200
rect 18877 7191 18935 7197
rect 18877 7157 18889 7191
rect 18923 7188 18935 7191
rect 19518 7188 19524 7200
rect 18923 7160 19524 7188
rect 18923 7157 18935 7160
rect 18877 7151 18935 7157
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 21928 7188 21956 7287
rect 22186 7284 22192 7336
rect 22244 7324 22250 7336
rect 23308 7324 23336 7364
rect 23750 7352 23756 7364
rect 23808 7352 23814 7404
rect 24136 7401 24164 7432
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7361 24179 7395
rect 24121 7355 24179 7361
rect 24210 7352 24216 7404
rect 24268 7392 24274 7404
rect 24397 7395 24455 7401
rect 24397 7392 24409 7395
rect 24268 7364 24409 7392
rect 24268 7352 24274 7364
rect 24397 7361 24409 7364
rect 24443 7361 24455 7395
rect 26160 7392 26188 7491
rect 26970 7488 26976 7540
rect 27028 7528 27034 7540
rect 27246 7528 27252 7540
rect 27028 7500 27252 7528
rect 27028 7488 27034 7500
rect 27246 7488 27252 7500
rect 27304 7488 27310 7540
rect 31846 7488 31852 7540
rect 31904 7488 31910 7540
rect 30377 7463 30435 7469
rect 30377 7460 30389 7463
rect 29840 7432 30389 7460
rect 29840 7401 29868 7432
rect 30377 7429 30389 7432
rect 30423 7429 30435 7463
rect 30377 7423 30435 7429
rect 30834 7420 30840 7472
rect 30892 7420 30898 7472
rect 29825 7395 29883 7401
rect 29825 7392 29837 7395
rect 24397 7355 24455 7361
rect 25700 7364 25806 7392
rect 26160 7364 29837 7392
rect 22244 7296 23336 7324
rect 22244 7284 22250 7296
rect 22278 7188 22284 7200
rect 21928 7160 22284 7188
rect 22278 7148 22284 7160
rect 22336 7148 22342 7200
rect 23768 7188 23796 7352
rect 24673 7327 24731 7333
rect 24673 7324 24685 7327
rect 24320 7296 24685 7324
rect 24320 7265 24348 7296
rect 24673 7293 24685 7296
rect 24719 7293 24731 7327
rect 24673 7287 24731 7293
rect 24305 7259 24363 7265
rect 24305 7225 24317 7259
rect 24351 7225 24363 7259
rect 24305 7219 24363 7225
rect 24854 7188 24860 7200
rect 23768 7160 24860 7188
rect 24854 7148 24860 7160
rect 24912 7188 24918 7200
rect 25700 7188 25728 7364
rect 29825 7361 29837 7364
rect 29871 7361 29883 7395
rect 30852 7392 30880 7420
rect 30929 7395 30987 7401
rect 30929 7392 30941 7395
rect 29825 7355 29883 7361
rect 30300 7364 30941 7392
rect 30300 7333 30328 7364
rect 30929 7361 30941 7364
rect 30975 7361 30987 7395
rect 30929 7355 30987 7361
rect 31478 7352 31484 7404
rect 31536 7352 31542 7404
rect 30285 7327 30343 7333
rect 30285 7293 30297 7327
rect 30331 7293 30343 7327
rect 30285 7287 30343 7293
rect 31389 7327 31447 7333
rect 31389 7293 31401 7327
rect 31435 7324 31447 7327
rect 31570 7324 31576 7336
rect 31435 7296 31576 7324
rect 31435 7293 31447 7296
rect 31389 7287 31447 7293
rect 31570 7284 31576 7296
rect 31628 7284 31634 7336
rect 30653 7259 30711 7265
rect 30653 7256 30665 7259
rect 29932 7228 30665 7256
rect 24912 7160 25728 7188
rect 24912 7148 24918 7160
rect 29822 7148 29828 7200
rect 29880 7188 29886 7200
rect 29932 7197 29960 7228
rect 30653 7225 30665 7228
rect 30699 7256 30711 7259
rect 32582 7256 32588 7268
rect 30699 7228 32588 7256
rect 30699 7225 30711 7228
rect 30653 7219 30711 7225
rect 32582 7216 32588 7228
rect 32640 7216 32646 7268
rect 29917 7191 29975 7197
rect 29917 7188 29929 7191
rect 29880 7160 29929 7188
rect 29880 7148 29886 7160
rect 29917 7157 29929 7160
rect 29963 7157 29975 7191
rect 29917 7151 29975 7157
rect 30837 7191 30895 7197
rect 30837 7157 30849 7191
rect 30883 7188 30895 7191
rect 30926 7188 30932 7200
rect 30883 7160 30932 7188
rect 30883 7157 30895 7160
rect 30837 7151 30895 7157
rect 30926 7148 30932 7160
rect 30984 7188 30990 7200
rect 31021 7191 31079 7197
rect 31021 7188 31033 7191
rect 30984 7160 31033 7188
rect 30984 7148 30990 7160
rect 31021 7157 31033 7160
rect 31067 7157 31079 7191
rect 31021 7151 31079 7157
rect 31478 7148 31484 7200
rect 31536 7148 31542 7200
rect 1104 7098 34684 7120
rect 1104 7046 5147 7098
rect 5199 7046 5211 7098
rect 5263 7046 5275 7098
rect 5327 7046 5339 7098
rect 5391 7046 5403 7098
rect 5455 7046 13541 7098
rect 13593 7046 13605 7098
rect 13657 7046 13669 7098
rect 13721 7046 13733 7098
rect 13785 7046 13797 7098
rect 13849 7046 21935 7098
rect 21987 7046 21999 7098
rect 22051 7046 22063 7098
rect 22115 7046 22127 7098
rect 22179 7046 22191 7098
rect 22243 7046 30329 7098
rect 30381 7046 30393 7098
rect 30445 7046 30457 7098
rect 30509 7046 30521 7098
rect 30573 7046 30585 7098
rect 30637 7046 34684 7098
rect 1104 7024 34684 7046
rect 7926 6944 7932 6996
rect 7984 6944 7990 6996
rect 16209 6987 16267 6993
rect 16209 6953 16221 6987
rect 16255 6984 16267 6987
rect 16390 6984 16396 6996
rect 16255 6956 16396 6984
rect 16255 6953 16267 6956
rect 16209 6947 16267 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 17300 6987 17358 6993
rect 17300 6953 17312 6987
rect 17346 6984 17358 6987
rect 17402 6984 17408 6996
rect 17346 6956 17408 6984
rect 17346 6953 17358 6956
rect 17300 6947 17358 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 18414 6944 18420 6996
rect 18472 6944 18478 6996
rect 18782 6944 18788 6996
rect 18840 6944 18846 6996
rect 26316 6987 26374 6993
rect 26316 6953 26328 6987
rect 26362 6984 26374 6987
rect 27062 6984 27068 6996
rect 26362 6956 27068 6984
rect 26362 6953 26374 6956
rect 26316 6947 26374 6953
rect 27062 6944 27068 6956
rect 27120 6944 27126 6996
rect 27798 6944 27804 6996
rect 27856 6944 27862 6996
rect 31018 6944 31024 6996
rect 31076 6944 31082 6996
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 3145 6851 3203 6857
rect 1443 6820 2728 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2700 6792 2728 6820
rect 3145 6817 3157 6851
rect 3191 6848 3203 6851
rect 7944 6848 7972 6944
rect 3191 6820 7972 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 16114 6808 16120 6860
rect 16172 6808 16178 6860
rect 17037 6851 17095 6857
rect 17037 6817 17049 6851
rect 17083 6848 17095 6851
rect 18432 6848 18460 6944
rect 19794 6876 19800 6928
rect 19852 6876 19858 6928
rect 17083 6820 18460 6848
rect 19444 6820 20024 6848
rect 17083 6817 17095 6820
rect 17037 6811 17095 6817
rect 2682 6740 2688 6792
rect 2740 6740 2746 6792
rect 3234 6780 3240 6792
rect 2806 6752 3240 6780
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 15930 6740 15936 6792
rect 15988 6740 15994 6792
rect 19444 6780 19472 6820
rect 18446 6752 19472 6780
rect 19518 6740 19524 6792
rect 19576 6740 19582 6792
rect 19613 6783 19671 6789
rect 19613 6749 19625 6783
rect 19659 6780 19671 6783
rect 19886 6780 19892 6792
rect 19659 6752 19892 6780
rect 19659 6749 19671 6752
rect 19613 6743 19671 6749
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 19996 6724 20024 6820
rect 26050 6808 26056 6860
rect 26108 6848 26114 6860
rect 26970 6848 26976 6860
rect 26108 6820 26976 6848
rect 26108 6808 26114 6820
rect 26970 6808 26976 6820
rect 27028 6808 27034 6860
rect 27522 6808 27528 6860
rect 27580 6848 27586 6860
rect 27580 6820 29592 6848
rect 27580 6808 27586 6820
rect 23566 6740 23572 6792
rect 23624 6740 23630 6792
rect 29564 6789 29592 6820
rect 29914 6808 29920 6860
rect 29972 6808 29978 6860
rect 31757 6851 31815 6857
rect 31757 6848 31769 6851
rect 30760 6820 31769 6848
rect 29549 6783 29607 6789
rect 29549 6749 29561 6783
rect 29595 6780 29607 6783
rect 29932 6780 29960 6808
rect 30760 6792 30788 6820
rect 31757 6817 31769 6820
rect 31803 6817 31815 6851
rect 31757 6811 31815 6817
rect 32398 6808 32404 6860
rect 32456 6808 32462 6860
rect 32582 6808 32588 6860
rect 32640 6808 32646 6860
rect 29595 6752 29960 6780
rect 29595 6749 29607 6752
rect 29549 6743 29607 6749
rect 30742 6740 30748 6792
rect 30800 6740 30806 6792
rect 30834 6740 30840 6792
rect 30892 6740 30898 6792
rect 31570 6740 31576 6792
rect 31628 6780 31634 6792
rect 31665 6783 31723 6789
rect 31665 6780 31677 6783
rect 31628 6752 31677 6780
rect 31628 6740 31634 6752
rect 31665 6749 31677 6752
rect 31711 6749 31723 6783
rect 31665 6743 31723 6749
rect 1670 6672 1676 6724
rect 1728 6672 1734 6724
rect 15194 6672 15200 6724
rect 15252 6712 15258 6724
rect 16206 6712 16212 6724
rect 15252 6684 16212 6712
rect 15252 6672 15258 6684
rect 16206 6672 16212 6684
rect 16264 6672 16270 6724
rect 19150 6672 19156 6724
rect 19208 6712 19214 6724
rect 19429 6715 19487 6721
rect 19429 6712 19441 6715
rect 19208 6684 19441 6712
rect 19208 6672 19214 6684
rect 19429 6681 19441 6684
rect 19475 6681 19487 6715
rect 19429 6675 19487 6681
rect 19978 6672 19984 6724
rect 20036 6672 20042 6724
rect 26602 6672 26608 6724
rect 26660 6712 26666 6724
rect 26660 6684 26818 6712
rect 26660 6672 26666 6684
rect 28810 6672 28816 6724
rect 28868 6712 28874 6724
rect 28868 6684 29776 6712
rect 28868 6672 28874 6684
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15749 6647 15807 6653
rect 15749 6644 15761 6647
rect 15620 6616 15761 6644
rect 15620 6604 15626 6616
rect 15749 6613 15761 6616
rect 15795 6613 15807 6647
rect 15749 6607 15807 6613
rect 19245 6647 19303 6653
rect 19245 6613 19257 6647
rect 19291 6644 19303 6647
rect 19334 6644 19340 6656
rect 19291 6616 19340 6644
rect 19291 6613 19303 6616
rect 19245 6607 19303 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 23382 6604 23388 6656
rect 23440 6604 23446 6656
rect 29638 6604 29644 6656
rect 29696 6604 29702 6656
rect 29748 6644 29776 6684
rect 30190 6672 30196 6724
rect 30248 6712 30254 6724
rect 30926 6712 30932 6724
rect 30248 6684 30932 6712
rect 30248 6672 30254 6684
rect 30926 6672 30932 6684
rect 30984 6712 30990 6724
rect 31021 6715 31079 6721
rect 31021 6712 31033 6715
rect 30984 6684 31033 6712
rect 30984 6672 30990 6684
rect 31021 6681 31033 6684
rect 31067 6681 31079 6715
rect 32416 6712 32444 6808
rect 31021 6675 31079 6681
rect 31726 6684 32444 6712
rect 31726 6644 31754 6684
rect 29748 6616 31754 6644
rect 32033 6647 32091 6653
rect 32033 6613 32045 6647
rect 32079 6644 32091 6647
rect 32677 6647 32735 6653
rect 32677 6644 32689 6647
rect 32079 6616 32689 6644
rect 32079 6613 32091 6616
rect 32033 6607 32091 6613
rect 32677 6613 32689 6616
rect 32723 6613 32735 6647
rect 32677 6607 32735 6613
rect 33042 6604 33048 6656
rect 33100 6604 33106 6656
rect 1104 6554 34840 6576
rect 1104 6502 9344 6554
rect 9396 6502 9408 6554
rect 9460 6502 9472 6554
rect 9524 6502 9536 6554
rect 9588 6502 9600 6554
rect 9652 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 17930 6554
rect 17982 6502 17994 6554
rect 18046 6502 26132 6554
rect 26184 6502 26196 6554
rect 26248 6502 26260 6554
rect 26312 6502 26324 6554
rect 26376 6502 26388 6554
rect 26440 6502 34526 6554
rect 34578 6502 34590 6554
rect 34642 6502 34654 6554
rect 34706 6502 34718 6554
rect 34770 6502 34782 6554
rect 34834 6502 34840 6554
rect 1104 6480 34840 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 8941 6443 8999 6449
rect 7852 6412 8800 6440
rect 3234 6332 3240 6384
rect 3292 6372 3298 6384
rect 7852 6372 7880 6412
rect 8772 6372 8800 6412
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 10686 6440 10692 6452
rect 8987 6412 10692 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 11716 6412 13124 6440
rect 11716 6372 11744 6412
rect 3292 6344 7958 6372
rect 8772 6344 11744 6372
rect 3292 6332 3298 6344
rect 11790 6332 11796 6384
rect 11848 6332 11854 6384
rect 13096 6372 13124 6412
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 14550 6440 14556 6452
rect 13320 6412 14556 6440
rect 13320 6400 13326 6412
rect 13354 6372 13360 6384
rect 13018 6344 13360 6372
rect 13354 6332 13360 6344
rect 13412 6332 13418 6384
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 13464 6313 13492 6412
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 15194 6400 15200 6452
rect 15252 6400 15258 6452
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 19245 6443 19303 6449
rect 19245 6440 19257 6443
rect 19208 6412 19257 6440
rect 19208 6400 19214 6412
rect 19245 6409 19257 6412
rect 19291 6409 19303 6443
rect 19245 6403 19303 6409
rect 19334 6400 19340 6452
rect 19392 6400 19398 6452
rect 22462 6400 22468 6452
rect 22520 6440 22526 6452
rect 22833 6443 22891 6449
rect 22833 6440 22845 6443
rect 22520 6412 22845 6440
rect 22520 6400 22526 6412
rect 22833 6409 22845 6412
rect 22879 6409 22891 6443
rect 22833 6403 22891 6409
rect 23293 6443 23351 6449
rect 23293 6409 23305 6443
rect 23339 6440 23351 6443
rect 23566 6440 23572 6452
rect 23339 6412 23572 6440
rect 23339 6409 23351 6412
rect 23293 6403 23351 6409
rect 23566 6400 23572 6412
rect 23624 6400 23630 6452
rect 24673 6443 24731 6449
rect 24673 6409 24685 6443
rect 24719 6440 24731 6443
rect 27338 6440 27344 6452
rect 24719 6412 27344 6440
rect 24719 6409 24731 6412
rect 24673 6403 24731 6409
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 29546 6440 29552 6452
rect 27724 6412 29552 6440
rect 18877 6375 18935 6381
rect 18877 6341 18889 6375
rect 18923 6372 18935 6375
rect 18966 6372 18972 6384
rect 18923 6344 18972 6372
rect 18923 6341 18935 6344
rect 18877 6335 18935 6341
rect 18966 6332 18972 6344
rect 19024 6332 19030 6384
rect 19058 6332 19064 6384
rect 19116 6332 19122 6384
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 2740 6276 7205 6304
rect 2740 6264 2746 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 7466 6196 7472 6248
rect 7524 6196 7530 6248
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 12802 6236 12808 6248
rect 11563 6208 12808 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 12802 6196 12808 6208
rect 12860 6236 12866 6248
rect 13464 6236 13492 6267
rect 14826 6264 14832 6316
rect 14884 6264 14890 6316
rect 19352 6313 19380 6400
rect 27724 6372 27752 6412
rect 29546 6400 29552 6412
rect 29604 6400 29610 6452
rect 29730 6400 29736 6452
rect 29788 6400 29794 6452
rect 30469 6443 30527 6449
rect 30469 6440 30481 6443
rect 30300 6412 30481 6440
rect 27448 6344 27752 6372
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 20530 6264 20536 6316
rect 20588 6264 20594 6316
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6304 22431 6307
rect 22462 6304 22468 6316
rect 22419 6276 22468 6304
rect 22419 6273 22431 6276
rect 22373 6267 22431 6273
rect 22462 6264 22468 6276
rect 22520 6304 22526 6316
rect 22925 6307 22983 6313
rect 22520 6276 22784 6304
rect 22520 6264 22526 6276
rect 12860 6208 13492 6236
rect 13725 6239 13783 6245
rect 12860 6196 12866 6208
rect 13725 6205 13737 6239
rect 13771 6236 13783 6239
rect 14090 6236 14096 6248
rect 13771 6208 14096 6236
rect 13771 6205 13783 6208
rect 13725 6199 13783 6205
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 22646 6196 22652 6248
rect 22704 6196 22710 6248
rect 22756 6236 22784 6276
rect 22925 6273 22937 6307
rect 22971 6304 22983 6307
rect 24305 6307 24363 6313
rect 22971 6276 24072 6304
rect 22971 6273 22983 6276
rect 22925 6267 22983 6273
rect 23477 6239 23535 6245
rect 23477 6236 23489 6239
rect 22756 6208 23489 6236
rect 23477 6205 23489 6208
rect 23523 6205 23535 6239
rect 23477 6199 23535 6205
rect 24044 6168 24072 6276
rect 24305 6273 24317 6307
rect 24351 6304 24363 6307
rect 24351 6276 27384 6304
rect 24351 6273 24363 6276
rect 24305 6267 24363 6273
rect 27356 6248 27384 6276
rect 24121 6239 24179 6245
rect 24121 6205 24133 6239
rect 24167 6236 24179 6239
rect 24946 6236 24952 6248
rect 24167 6208 24952 6236
rect 24167 6205 24179 6208
rect 24121 6199 24179 6205
rect 24946 6196 24952 6208
rect 25004 6196 25010 6248
rect 25866 6196 25872 6248
rect 25924 6196 25930 6248
rect 27338 6196 27344 6248
rect 27396 6196 27402 6248
rect 27448 6245 27476 6344
rect 27798 6332 27804 6384
rect 27856 6372 27862 6384
rect 27985 6375 28043 6381
rect 27985 6372 27997 6375
rect 27856 6344 27997 6372
rect 27856 6332 27862 6344
rect 27985 6341 27997 6344
rect 28031 6341 28043 6375
rect 30300 6372 30328 6412
rect 30469 6409 30481 6412
rect 30515 6409 30527 6443
rect 30469 6403 30527 6409
rect 30742 6400 30748 6452
rect 30800 6440 30806 6452
rect 30837 6443 30895 6449
rect 30837 6440 30849 6443
rect 30800 6412 30849 6440
rect 30800 6400 30806 6412
rect 30837 6409 30849 6412
rect 30883 6409 30895 6443
rect 30837 6403 30895 6409
rect 31754 6400 31760 6452
rect 31812 6440 31818 6452
rect 32585 6443 32643 6449
rect 32585 6440 32597 6443
rect 31812 6412 32597 6440
rect 31812 6400 31818 6412
rect 32585 6409 32597 6412
rect 32631 6409 32643 6443
rect 32585 6403 32643 6409
rect 32490 6372 32496 6384
rect 27985 6335 28043 6341
rect 29932 6344 30328 6372
rect 31726 6344 32496 6372
rect 27522 6264 27528 6316
rect 27580 6264 27586 6316
rect 28000 6304 28028 6335
rect 29932 6316 29960 6344
rect 28537 6307 28595 6313
rect 28537 6304 28549 6307
rect 28000 6276 28549 6304
rect 28537 6273 28549 6276
rect 28583 6273 28595 6307
rect 28537 6267 28595 6273
rect 29914 6264 29920 6316
rect 29972 6264 29978 6316
rect 30009 6307 30067 6313
rect 30009 6273 30021 6307
rect 30055 6273 30067 6307
rect 30009 6267 30067 6273
rect 27433 6239 27491 6245
rect 27433 6205 27445 6239
rect 27479 6205 27491 6239
rect 28445 6239 28503 6245
rect 27433 6199 27491 6205
rect 27540 6208 28396 6236
rect 26786 6168 26792 6180
rect 24044 6140 24164 6168
rect 24136 6112 24164 6140
rect 24688 6140 26792 6168
rect 13262 6060 13268 6112
rect 13320 6060 13326 6112
rect 19518 6060 19524 6112
rect 19576 6060 19582 6112
rect 20254 6060 20260 6112
rect 20312 6100 20318 6112
rect 20349 6103 20407 6109
rect 20349 6100 20361 6103
rect 20312 6072 20361 6100
rect 20312 6060 20318 6072
rect 20349 6069 20361 6072
rect 20395 6069 20407 6103
rect 20349 6063 20407 6069
rect 21818 6060 21824 6112
rect 21876 6060 21882 6112
rect 24118 6060 24124 6112
rect 24176 6060 24182 6112
rect 24688 6109 24716 6140
rect 26786 6128 26792 6140
rect 26844 6168 26850 6180
rect 27540 6168 27568 6208
rect 26844 6140 27568 6168
rect 26844 6128 26850 6140
rect 27890 6128 27896 6180
rect 27948 6168 27954 6180
rect 28261 6171 28319 6177
rect 28261 6168 28273 6171
rect 27948 6140 28273 6168
rect 27948 6128 27954 6140
rect 28261 6137 28273 6140
rect 28307 6137 28319 6171
rect 28368 6168 28396 6208
rect 28445 6205 28457 6239
rect 28491 6236 28503 6239
rect 29089 6239 29147 6245
rect 29089 6236 29101 6239
rect 28491 6208 29101 6236
rect 28491 6205 28503 6208
rect 28445 6199 28503 6205
rect 29089 6205 29101 6208
rect 29135 6236 29147 6239
rect 29822 6236 29828 6248
rect 29135 6208 29828 6236
rect 29135 6205 29147 6208
rect 29089 6199 29147 6205
rect 29822 6196 29828 6208
rect 29880 6236 29886 6248
rect 30024 6236 30052 6267
rect 30190 6264 30196 6316
rect 30248 6264 30254 6316
rect 30285 6307 30343 6313
rect 30285 6273 30297 6307
rect 30331 6273 30343 6307
rect 30285 6267 30343 6273
rect 29880 6208 30052 6236
rect 29880 6196 29886 6208
rect 30098 6196 30104 6248
rect 30156 6236 30162 6248
rect 30300 6236 30328 6267
rect 30374 6264 30380 6316
rect 30432 6264 30438 6316
rect 30653 6307 30711 6313
rect 30653 6304 30665 6307
rect 30576 6276 30665 6304
rect 30576 6236 30604 6276
rect 30653 6273 30665 6276
rect 30699 6273 30711 6307
rect 30653 6267 30711 6273
rect 30156 6208 30604 6236
rect 30156 6196 30162 6208
rect 28997 6171 29055 6177
rect 28368 6140 28764 6168
rect 28261 6131 28319 6137
rect 24673 6103 24731 6109
rect 24673 6069 24685 6103
rect 24719 6069 24731 6103
rect 24673 6063 24731 6069
rect 24854 6060 24860 6112
rect 24912 6060 24918 6112
rect 25314 6060 25320 6112
rect 25372 6060 25378 6112
rect 27798 6060 27804 6112
rect 27856 6060 27862 6112
rect 28276 6100 28304 6131
rect 28629 6103 28687 6109
rect 28629 6100 28641 6103
rect 28276 6072 28641 6100
rect 28629 6069 28641 6072
rect 28675 6069 28687 6103
rect 28736 6100 28764 6140
rect 28997 6137 29009 6171
rect 29043 6168 29055 6171
rect 29362 6168 29368 6180
rect 29043 6140 29368 6168
rect 29043 6137 29055 6140
rect 28997 6131 29055 6137
rect 29362 6128 29368 6140
rect 29420 6128 29426 6180
rect 31726 6100 31754 6344
rect 32490 6332 32496 6344
rect 32548 6332 32554 6384
rect 32122 6264 32128 6316
rect 32180 6304 32186 6316
rect 32950 6304 32956 6316
rect 32180 6276 32956 6304
rect 32180 6264 32186 6276
rect 32950 6264 32956 6276
rect 33008 6264 33014 6316
rect 34330 6264 34336 6316
rect 34388 6264 34394 6316
rect 34054 6196 34060 6248
rect 34112 6196 34118 6248
rect 28736 6072 31754 6100
rect 28629 6063 28687 6069
rect 1104 6010 34684 6032
rect 1104 5958 5147 6010
rect 5199 5958 5211 6010
rect 5263 5958 5275 6010
rect 5327 5958 5339 6010
rect 5391 5958 5403 6010
rect 5455 5958 13541 6010
rect 13593 5958 13605 6010
rect 13657 5958 13669 6010
rect 13721 5958 13733 6010
rect 13785 5958 13797 6010
rect 13849 5958 21935 6010
rect 21987 5958 21999 6010
rect 22051 5958 22063 6010
rect 22115 5958 22127 6010
rect 22179 5958 22191 6010
rect 22243 5958 30329 6010
rect 30381 5958 30393 6010
rect 30445 5958 30457 6010
rect 30509 5958 30521 6010
rect 30573 5958 30585 6010
rect 30637 5958 34684 6010
rect 1104 5936 34684 5958
rect 13262 5856 13268 5908
rect 13320 5856 13326 5908
rect 14090 5856 14096 5908
rect 14148 5856 14154 5908
rect 15930 5856 15936 5908
rect 15988 5856 15994 5908
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 21361 5899 21419 5905
rect 21361 5896 21373 5899
rect 20588 5868 21373 5896
rect 20588 5856 20594 5868
rect 21361 5865 21373 5868
rect 21407 5865 21419 5899
rect 21361 5859 21419 5865
rect 21818 5856 21824 5908
rect 21876 5856 21882 5908
rect 22554 5856 22560 5908
rect 22612 5856 22618 5908
rect 22728 5899 22786 5905
rect 22728 5865 22740 5899
rect 22774 5896 22786 5899
rect 23382 5896 23388 5908
rect 22774 5868 23388 5896
rect 22774 5865 22786 5868
rect 22728 5859 22786 5865
rect 23382 5856 23388 5868
rect 23440 5856 23446 5908
rect 26694 5896 26700 5908
rect 24780 5868 26700 5896
rect 13280 5760 13308 5856
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 13280 5732 14657 5760
rect 14645 5729 14657 5732
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 17681 5763 17739 5769
rect 17681 5729 17693 5763
rect 17727 5760 17739 5763
rect 19242 5760 19248 5772
rect 17727 5732 19248 5760
rect 17727 5729 17739 5732
rect 17681 5723 17739 5729
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 19518 5720 19524 5772
rect 19576 5720 19582 5772
rect 21729 5695 21787 5701
rect 21729 5661 21741 5695
rect 21775 5692 21787 5695
rect 21836 5692 21864 5856
rect 22572 5828 22600 5856
rect 24780 5840 24808 5868
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 29362 5856 29368 5908
rect 29420 5856 29426 5908
rect 29638 5856 29644 5908
rect 29696 5856 29702 5908
rect 29822 5856 29828 5908
rect 29880 5856 29886 5908
rect 30009 5899 30067 5905
rect 30009 5865 30021 5899
rect 30055 5896 30067 5899
rect 30190 5896 30196 5908
rect 30055 5868 30196 5896
rect 30055 5865 30067 5868
rect 30009 5859 30067 5865
rect 30190 5856 30196 5868
rect 30248 5856 30254 5908
rect 31754 5896 31760 5908
rect 31726 5856 31760 5896
rect 31812 5856 31818 5908
rect 32217 5899 32275 5905
rect 32217 5865 32229 5899
rect 32263 5896 32275 5899
rect 34054 5896 34060 5908
rect 32263 5868 34060 5896
rect 32263 5865 32275 5868
rect 32217 5859 32275 5865
rect 34054 5856 34060 5868
rect 34112 5856 34118 5908
rect 21928 5800 22600 5828
rect 21928 5769 21956 5800
rect 24762 5788 24768 5840
rect 24820 5788 24826 5840
rect 21913 5763 21971 5769
rect 21913 5729 21925 5763
rect 21959 5729 21971 5763
rect 21913 5723 21971 5729
rect 22278 5720 22284 5772
rect 22336 5760 22342 5772
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 22336 5732 22477 5760
rect 22336 5720 22342 5732
rect 22465 5729 22477 5732
rect 22511 5760 22523 5763
rect 24210 5760 24216 5772
rect 22511 5732 24216 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 24210 5720 24216 5732
rect 24268 5760 24274 5772
rect 24949 5763 25007 5769
rect 24949 5760 24961 5763
rect 24268 5732 24961 5760
rect 24268 5720 24274 5732
rect 24949 5729 24961 5732
rect 24995 5729 25007 5763
rect 24949 5723 25007 5729
rect 25225 5763 25283 5769
rect 25225 5729 25237 5763
rect 25271 5760 25283 5763
rect 25314 5760 25320 5772
rect 25271 5732 25320 5760
rect 25271 5729 25283 5732
rect 25225 5723 25283 5729
rect 25314 5720 25320 5732
rect 25372 5720 25378 5772
rect 26602 5760 26608 5772
rect 26344 5732 26608 5760
rect 21775 5664 21864 5692
rect 26344 5678 26372 5732
rect 26602 5720 26608 5732
rect 26660 5720 26666 5772
rect 27614 5720 27620 5772
rect 27672 5760 27678 5772
rect 28077 5763 28135 5769
rect 28077 5760 28089 5763
rect 27672 5732 28089 5760
rect 27672 5720 27678 5732
rect 28077 5729 28089 5732
rect 28123 5760 28135 5763
rect 28810 5760 28816 5772
rect 28123 5732 28816 5760
rect 28123 5729 28135 5732
rect 28077 5723 28135 5729
rect 28810 5720 28816 5732
rect 28868 5720 28874 5772
rect 29380 5692 29408 5856
rect 29656 5701 29684 5856
rect 29840 5701 29868 5856
rect 31726 5760 31754 5856
rect 31496 5732 31754 5760
rect 31496 5701 31524 5732
rect 29549 5695 29607 5701
rect 29549 5692 29561 5695
rect 26528 5664 28028 5692
rect 29380 5664 29561 5692
rect 21775 5661 21787 5664
rect 21729 5655 21787 5661
rect 17126 5624 17132 5636
rect 16974 5596 17132 5624
rect 17126 5584 17132 5596
rect 17184 5584 17190 5636
rect 17405 5627 17463 5633
rect 17405 5593 17417 5627
rect 17451 5593 17463 5627
rect 17405 5587 17463 5593
rect 17420 5556 17448 5587
rect 19978 5584 19984 5636
rect 20036 5584 20042 5636
rect 21269 5627 21327 5633
rect 21269 5593 21281 5627
rect 21315 5624 21327 5627
rect 21450 5624 21456 5636
rect 21315 5596 21456 5624
rect 21315 5593 21327 5596
rect 21269 5587 21327 5593
rect 21450 5584 21456 5596
rect 21508 5584 21514 5636
rect 21744 5596 22094 5624
rect 21744 5556 21772 5596
rect 17420 5528 21772 5556
rect 21818 5516 21824 5568
rect 21876 5516 21882 5568
rect 22066 5556 22094 5596
rect 23750 5584 23756 5636
rect 23808 5584 23814 5636
rect 23474 5556 23480 5568
rect 22066 5528 23480 5556
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 24118 5516 24124 5568
rect 24176 5556 24182 5568
rect 24213 5559 24271 5565
rect 24213 5556 24225 5559
rect 24176 5528 24225 5556
rect 24176 5516 24182 5528
rect 24213 5525 24225 5528
rect 24259 5556 24271 5559
rect 26528 5556 26556 5664
rect 26694 5584 26700 5636
rect 26752 5624 26758 5636
rect 27890 5624 27896 5636
rect 26752 5596 27896 5624
rect 26752 5584 26758 5596
rect 27890 5584 27896 5596
rect 27948 5584 27954 5636
rect 28000 5624 28028 5664
rect 29549 5661 29561 5664
rect 29595 5661 29607 5695
rect 29549 5655 29607 5661
rect 29641 5695 29699 5701
rect 29641 5661 29653 5695
rect 29687 5661 29699 5695
rect 29641 5655 29699 5661
rect 29825 5695 29883 5701
rect 29825 5661 29837 5695
rect 29871 5661 29883 5695
rect 29825 5655 29883 5661
rect 31481 5695 31539 5701
rect 31481 5661 31493 5695
rect 31527 5661 31539 5695
rect 31757 5695 31815 5701
rect 31757 5692 31769 5695
rect 31481 5655 31539 5661
rect 31588 5664 31769 5692
rect 31588 5624 31616 5664
rect 31757 5661 31769 5664
rect 31803 5661 31815 5695
rect 31757 5655 31815 5661
rect 31846 5652 31852 5704
rect 31904 5652 31910 5704
rect 32401 5695 32459 5701
rect 32401 5692 32413 5695
rect 32048 5664 32413 5692
rect 28000 5596 31616 5624
rect 31665 5627 31723 5633
rect 31665 5593 31677 5627
rect 31711 5593 31723 5627
rect 31665 5587 31723 5593
rect 24259 5528 26556 5556
rect 24259 5525 24271 5528
rect 24213 5519 24271 5525
rect 26878 5516 26884 5568
rect 26936 5556 26942 5568
rect 27433 5559 27491 5565
rect 27433 5556 27445 5559
rect 26936 5528 27445 5556
rect 26936 5516 26942 5528
rect 27433 5525 27445 5528
rect 27479 5525 27491 5559
rect 27433 5519 27491 5525
rect 27798 5516 27804 5568
rect 27856 5516 27862 5568
rect 30374 5516 30380 5568
rect 30432 5556 30438 5568
rect 31110 5556 31116 5568
rect 30432 5528 31116 5556
rect 30432 5516 30438 5528
rect 31110 5516 31116 5528
rect 31168 5556 31174 5568
rect 31680 5556 31708 5587
rect 32048 5565 32076 5664
rect 32401 5661 32413 5664
rect 32447 5661 32459 5695
rect 32401 5655 32459 5661
rect 32490 5652 32496 5704
rect 32548 5692 32554 5704
rect 32585 5695 32643 5701
rect 32585 5692 32597 5695
rect 32548 5664 32597 5692
rect 32548 5652 32554 5664
rect 32585 5661 32597 5664
rect 32631 5661 32643 5695
rect 32585 5655 32643 5661
rect 32677 5695 32735 5701
rect 32677 5661 32689 5695
rect 32723 5692 32735 5695
rect 33042 5692 33048 5704
rect 32723 5664 33048 5692
rect 32723 5661 32735 5664
rect 32677 5655 32735 5661
rect 33042 5652 33048 5664
rect 33100 5652 33106 5704
rect 31168 5528 31708 5556
rect 32033 5559 32091 5565
rect 31168 5516 31174 5528
rect 32033 5525 32045 5559
rect 32079 5525 32091 5559
rect 32033 5519 32091 5525
rect 1104 5466 34840 5488
rect 1104 5414 9344 5466
rect 9396 5414 9408 5466
rect 9460 5414 9472 5466
rect 9524 5414 9536 5466
rect 9588 5414 9600 5466
rect 9652 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 17930 5466
rect 17982 5414 17994 5466
rect 18046 5414 26132 5466
rect 26184 5414 26196 5466
rect 26248 5414 26260 5466
rect 26312 5414 26324 5466
rect 26376 5414 26388 5466
rect 26440 5414 34526 5466
rect 34578 5414 34590 5466
rect 34642 5414 34654 5466
rect 34706 5414 34718 5466
rect 34770 5414 34782 5466
rect 34834 5414 34840 5466
rect 1104 5392 34840 5414
rect 19978 5312 19984 5364
rect 20036 5352 20042 5364
rect 21637 5355 21695 5361
rect 20036 5324 21312 5352
rect 20036 5312 20042 5324
rect 15746 5244 15752 5296
rect 15804 5284 15810 5296
rect 17126 5284 17132 5296
rect 15804 5256 17132 5284
rect 15804 5244 15810 5256
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 20165 5287 20223 5293
rect 20165 5253 20177 5287
rect 20211 5284 20223 5287
rect 20254 5284 20260 5296
rect 20211 5256 20260 5284
rect 20211 5253 20223 5256
rect 20165 5247 20223 5253
rect 20254 5244 20260 5256
rect 20312 5244 20318 5296
rect 20456 5284 20484 5324
rect 20456 5256 20654 5284
rect 12802 5176 12808 5228
rect 12860 5216 12866 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12860 5188 12909 5216
rect 12860 5176 12866 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 14826 5216 14832 5228
rect 14306 5188 14832 5216
rect 12897 5179 12955 5185
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 16482 5176 16488 5228
rect 16540 5176 16546 5228
rect 13170 5108 13176 5160
rect 13228 5108 13234 5160
rect 14642 5108 14648 5160
rect 14700 5108 14706 5160
rect 14734 5108 14740 5160
rect 14792 5108 14798 5160
rect 14844 5148 14872 5176
rect 15746 5148 15752 5160
rect 14844 5120 15752 5148
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 16206 5108 16212 5160
rect 16264 5108 16270 5160
rect 19886 5108 19892 5160
rect 19944 5148 19950 5160
rect 21174 5148 21180 5160
rect 19944 5120 21180 5148
rect 19944 5108 19950 5120
rect 21174 5108 21180 5120
rect 21232 5108 21238 5160
rect 21284 5080 21312 5324
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 22462 5352 22468 5364
rect 21683 5324 22468 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 23845 5355 23903 5361
rect 23845 5352 23857 5355
rect 23532 5324 23857 5352
rect 23532 5312 23538 5324
rect 23845 5321 23857 5324
rect 23891 5321 23903 5355
rect 23845 5315 23903 5321
rect 24854 5312 24860 5364
rect 24912 5312 24918 5364
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 25409 5355 25467 5361
rect 25004 5324 25176 5352
rect 25004 5312 25010 5324
rect 21450 5244 21456 5296
rect 21508 5284 21514 5296
rect 22281 5287 22339 5293
rect 22281 5284 22293 5287
rect 21508 5256 22293 5284
rect 21508 5244 21514 5256
rect 22281 5253 22293 5256
rect 22327 5253 22339 5287
rect 24872 5284 24900 5312
rect 25148 5293 25176 5324
rect 25409 5321 25421 5355
rect 25455 5352 25467 5355
rect 25866 5352 25872 5364
rect 25455 5324 25872 5352
rect 25455 5321 25467 5324
rect 25409 5315 25467 5321
rect 25866 5312 25872 5324
rect 25924 5312 25930 5364
rect 26421 5355 26479 5361
rect 26421 5321 26433 5355
rect 26467 5352 26479 5355
rect 26786 5352 26792 5364
rect 26467 5324 26792 5352
rect 26467 5321 26479 5324
rect 26421 5315 26479 5321
rect 26786 5312 26792 5324
rect 26844 5312 26850 5364
rect 26878 5312 26884 5364
rect 26936 5312 26942 5364
rect 26973 5355 27031 5361
rect 26973 5321 26985 5355
rect 27019 5321 27031 5355
rect 26973 5315 27031 5321
rect 28445 5355 28503 5361
rect 28445 5321 28457 5355
rect 28491 5352 28503 5355
rect 28534 5352 28540 5364
rect 28491 5324 28540 5352
rect 28491 5321 28503 5324
rect 28445 5315 28503 5321
rect 22281 5247 22339 5253
rect 24780 5256 24900 5284
rect 25133 5287 25191 5293
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5216 22247 5219
rect 23017 5219 23075 5225
rect 23017 5216 23029 5219
rect 22235 5188 23029 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 23017 5185 23029 5188
rect 23063 5185 23075 5219
rect 23017 5179 23075 5185
rect 23658 5176 23664 5228
rect 23716 5216 23722 5228
rect 24780 5225 24808 5256
rect 25133 5253 25145 5287
rect 25179 5253 25191 5287
rect 26896 5284 26924 5312
rect 25133 5247 25191 5253
rect 26344 5256 26924 5284
rect 24765 5219 24823 5225
rect 23716 5188 24532 5216
rect 23716 5176 23722 5188
rect 22465 5151 22523 5157
rect 22465 5117 22477 5151
rect 22511 5148 22523 5151
rect 22554 5148 22560 5160
rect 22511 5120 22560 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 22554 5108 22560 5120
rect 22612 5108 22618 5160
rect 24397 5151 24455 5157
rect 24397 5117 24409 5151
rect 24443 5117 24455 5151
rect 24397 5111 24455 5117
rect 23750 5080 23756 5092
rect 21284 5052 23756 5080
rect 23750 5040 23756 5052
rect 23808 5040 23814 5092
rect 21818 4972 21824 5024
rect 21876 4972 21882 5024
rect 24412 5012 24440 5111
rect 24504 5080 24532 5188
rect 24765 5185 24777 5219
rect 24811 5185 24823 5219
rect 24765 5179 24823 5185
rect 24854 5176 24860 5228
rect 24912 5176 24918 5228
rect 25038 5176 25044 5228
rect 25096 5176 25102 5228
rect 25222 5176 25228 5228
rect 25280 5225 25286 5228
rect 26344 5225 26372 5256
rect 25280 5216 25288 5225
rect 26329 5219 26387 5225
rect 25280 5188 25325 5216
rect 25280 5179 25288 5188
rect 26329 5185 26341 5219
rect 26375 5185 26387 5219
rect 26329 5179 26387 5185
rect 26605 5219 26663 5225
rect 26605 5185 26617 5219
rect 26651 5216 26663 5219
rect 26988 5216 27016 5315
rect 28534 5312 28540 5324
rect 28592 5312 28598 5364
rect 28813 5355 28871 5361
rect 28813 5321 28825 5355
rect 28859 5352 28871 5355
rect 30009 5355 30067 5361
rect 30009 5352 30021 5355
rect 28859 5324 30021 5352
rect 28859 5321 28871 5324
rect 28813 5315 28871 5321
rect 30009 5321 30021 5324
rect 30055 5321 30067 5355
rect 30374 5352 30380 5364
rect 30009 5315 30067 5321
rect 30300 5324 30380 5352
rect 30300 5284 30328 5324
rect 30374 5312 30380 5324
rect 30432 5312 30438 5364
rect 30837 5355 30895 5361
rect 30837 5321 30849 5355
rect 30883 5352 30895 5355
rect 31478 5352 31484 5364
rect 30883 5324 31484 5352
rect 30883 5321 30895 5324
rect 30837 5315 30895 5321
rect 30852 5284 30880 5315
rect 31478 5312 31484 5324
rect 31536 5312 31542 5364
rect 27356 5256 30328 5284
rect 30392 5256 30880 5284
rect 26651 5188 27016 5216
rect 26651 5185 26663 5188
rect 26605 5179 26663 5185
rect 25280 5176 25286 5179
rect 27154 5176 27160 5228
rect 27212 5176 27218 5228
rect 27356 5225 27384 5256
rect 27249 5219 27307 5225
rect 27249 5185 27261 5219
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5185 27399 5219
rect 27341 5179 27399 5185
rect 27525 5219 27583 5225
rect 27525 5185 27537 5219
rect 27571 5216 27583 5219
rect 28902 5216 28908 5228
rect 27571 5188 28908 5216
rect 27571 5185 27583 5188
rect 27525 5179 27583 5185
rect 25501 5151 25559 5157
rect 25501 5117 25513 5151
rect 25547 5117 25559 5151
rect 25501 5111 25559 5117
rect 26145 5151 26203 5157
rect 26145 5117 26157 5151
rect 26191 5148 26203 5151
rect 27264 5148 27292 5179
rect 26191 5120 27292 5148
rect 26191 5117 26203 5120
rect 26145 5111 26203 5117
rect 25516 5080 25544 5111
rect 27356 5092 27384 5179
rect 28902 5176 28908 5188
rect 28960 5176 28966 5228
rect 30392 5225 30420 5256
rect 30377 5219 30435 5225
rect 30377 5185 30389 5219
rect 30423 5185 30435 5219
rect 30377 5179 30435 5185
rect 30650 5176 30656 5228
rect 30708 5176 30714 5228
rect 30837 5219 30895 5225
rect 30837 5216 30849 5219
rect 30760 5188 30849 5216
rect 28810 5108 28816 5160
rect 28868 5148 28874 5160
rect 28997 5151 29055 5157
rect 28997 5148 29009 5151
rect 28868 5120 29009 5148
rect 28868 5108 28874 5120
rect 28997 5117 29009 5120
rect 29043 5117 29055 5151
rect 28997 5111 29055 5117
rect 29362 5108 29368 5160
rect 29420 5108 29426 5160
rect 30190 5108 30196 5160
rect 30248 5148 30254 5160
rect 30285 5151 30343 5157
rect 30285 5148 30297 5151
rect 30248 5120 30297 5148
rect 30248 5108 30254 5120
rect 30285 5117 30297 5120
rect 30331 5117 30343 5151
rect 30285 5111 30343 5117
rect 24504 5052 25544 5080
rect 26786 5040 26792 5092
rect 26844 5040 26850 5092
rect 27338 5040 27344 5092
rect 27396 5040 27402 5092
rect 29380 5080 29408 5108
rect 29914 5080 29920 5092
rect 29380 5052 29920 5080
rect 29914 5040 29920 5052
rect 29972 5080 29978 5092
rect 30760 5080 30788 5188
rect 30837 5185 30849 5188
rect 30883 5185 30895 5219
rect 30837 5179 30895 5185
rect 29972 5052 30788 5080
rect 29972 5040 29978 5052
rect 30190 5012 30196 5024
rect 24412 4984 30196 5012
rect 30190 4972 30196 4984
rect 30248 4972 30254 5024
rect 1104 4922 34684 4944
rect 1104 4870 5147 4922
rect 5199 4870 5211 4922
rect 5263 4870 5275 4922
rect 5327 4870 5339 4922
rect 5391 4870 5403 4922
rect 5455 4870 13541 4922
rect 13593 4870 13605 4922
rect 13657 4870 13669 4922
rect 13721 4870 13733 4922
rect 13785 4870 13797 4922
rect 13849 4870 21935 4922
rect 21987 4870 21999 4922
rect 22051 4870 22063 4922
rect 22115 4870 22127 4922
rect 22179 4870 22191 4922
rect 22243 4870 30329 4922
rect 30381 4870 30393 4922
rect 30445 4870 30457 4922
rect 30509 4870 30521 4922
rect 30573 4870 30585 4922
rect 30637 4870 34684 4922
rect 1104 4848 34684 4870
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 13228 4780 13277 4808
rect 13228 4768 13234 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 16206 4808 16212 4820
rect 15335 4780 16212 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 23658 4768 23664 4820
rect 23716 4768 23722 4820
rect 25038 4768 25044 4820
rect 25096 4808 25102 4820
rect 27338 4808 27344 4820
rect 25096 4780 27344 4808
rect 25096 4768 25102 4780
rect 27338 4768 27344 4780
rect 27396 4768 27402 4820
rect 28902 4768 28908 4820
rect 28960 4808 28966 4820
rect 28997 4811 29055 4817
rect 28997 4808 29009 4811
rect 28960 4780 29009 4808
rect 28960 4768 28966 4780
rect 28997 4777 29009 4780
rect 29043 4808 29055 4811
rect 30009 4811 30067 4817
rect 29043 4780 29868 4808
rect 29043 4777 29055 4780
rect 28997 4771 29055 4777
rect 25222 4740 25228 4752
rect 25056 4712 25228 4740
rect 21174 4632 21180 4684
rect 21232 4672 21238 4684
rect 21913 4675 21971 4681
rect 21913 4672 21925 4675
rect 21232 4644 21925 4672
rect 21232 4632 21238 4644
rect 21913 4641 21925 4644
rect 21959 4672 21971 4675
rect 22278 4672 22284 4684
rect 21959 4644 22284 4672
rect 21959 4641 21971 4644
rect 21913 4635 21971 4641
rect 22278 4632 22284 4644
rect 22336 4632 22342 4684
rect 25056 4681 25084 4712
rect 25222 4700 25228 4712
rect 25280 4740 25286 4752
rect 27154 4740 27160 4752
rect 25280 4712 27160 4740
rect 25280 4700 25286 4712
rect 27154 4700 27160 4712
rect 27212 4700 27218 4752
rect 29362 4700 29368 4752
rect 29420 4700 29426 4752
rect 29840 4749 29868 4780
rect 30009 4777 30021 4811
rect 30055 4808 30067 4811
rect 30098 4808 30104 4820
rect 30055 4780 30104 4808
rect 30055 4777 30067 4780
rect 30009 4771 30067 4777
rect 30098 4768 30104 4780
rect 30156 4768 30162 4820
rect 30193 4811 30251 4817
rect 30193 4777 30205 4811
rect 30239 4808 30251 4811
rect 30650 4808 30656 4820
rect 30239 4780 30656 4808
rect 30239 4777 30251 4780
rect 30193 4771 30251 4777
rect 30650 4768 30656 4780
rect 30708 4768 30714 4820
rect 29825 4743 29883 4749
rect 29825 4709 29837 4743
rect 29871 4709 29883 4743
rect 29825 4703 29883 4709
rect 25041 4675 25099 4681
rect 25041 4641 25053 4675
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 13814 4564 13820 4616
rect 13872 4564 13878 4616
rect 14642 4564 14648 4616
rect 14700 4564 14706 4616
rect 18138 4564 18144 4616
rect 18196 4564 18202 4616
rect 21637 4607 21695 4613
rect 21637 4573 21649 4607
rect 21683 4604 21695 4607
rect 21818 4604 21824 4616
rect 21683 4576 21824 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 21818 4564 21824 4576
rect 21876 4564 21882 4616
rect 23750 4604 23756 4616
rect 23322 4576 23756 4604
rect 23750 4564 23756 4576
rect 23808 4604 23814 4616
rect 24486 4604 24492 4616
rect 23808 4576 24492 4604
rect 23808 4564 23814 4576
rect 24486 4564 24492 4576
rect 24544 4564 24550 4616
rect 30116 4613 30144 4768
rect 28905 4607 28963 4613
rect 28905 4604 28917 4607
rect 25976 4576 28917 4604
rect 22189 4539 22247 4545
rect 22189 4536 22201 4539
rect 22066 4508 22201 4536
rect 14366 4428 14372 4480
rect 14424 4468 14430 4480
rect 16758 4468 16764 4480
rect 14424 4440 16764 4468
rect 14424 4428 14430 4440
rect 16758 4428 16764 4440
rect 16816 4428 16822 4480
rect 18785 4471 18843 4477
rect 18785 4437 18797 4471
rect 18831 4468 18843 4471
rect 19426 4468 19432 4480
rect 18831 4440 19432 4468
rect 18831 4437 18843 4440
rect 18785 4431 18843 4437
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 21821 4471 21879 4477
rect 21821 4437 21833 4471
rect 21867 4468 21879 4471
rect 22066 4468 22094 4508
rect 22189 4505 22201 4508
rect 22235 4505 22247 4539
rect 22189 4499 22247 4505
rect 23474 4496 23480 4548
rect 23532 4536 23538 4548
rect 24857 4539 24915 4545
rect 24857 4536 24869 4539
rect 23532 4508 24869 4536
rect 23532 4496 23538 4508
rect 24857 4505 24869 4508
rect 24903 4505 24915 4539
rect 24857 4499 24915 4505
rect 25976 4480 26004 4576
rect 28905 4573 28917 4576
rect 28951 4604 28963 4607
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 28951 4576 29561 4604
rect 28951 4573 28963 4576
rect 28905 4567 28963 4573
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29549 4567 29607 4573
rect 30101 4607 30159 4613
rect 30101 4573 30113 4607
rect 30147 4573 30159 4607
rect 30101 4567 30159 4573
rect 21867 4440 22094 4468
rect 21867 4437 21879 4440
rect 21821 4431 21879 4437
rect 24394 4428 24400 4480
rect 24452 4428 24458 4480
rect 24765 4471 24823 4477
rect 24765 4437 24777 4471
rect 24811 4468 24823 4471
rect 25958 4468 25964 4480
rect 24811 4440 25964 4468
rect 24811 4437 24823 4440
rect 24765 4431 24823 4437
rect 25958 4428 25964 4440
rect 26016 4428 26022 4480
rect 1104 4378 34840 4400
rect 1104 4326 9344 4378
rect 9396 4326 9408 4378
rect 9460 4326 9472 4378
rect 9524 4326 9536 4378
rect 9588 4326 9600 4378
rect 9652 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 17930 4378
rect 17982 4326 17994 4378
rect 18046 4326 26132 4378
rect 26184 4326 26196 4378
rect 26248 4326 26260 4378
rect 26312 4326 26324 4378
rect 26376 4326 26388 4378
rect 26440 4326 34526 4378
rect 34578 4326 34590 4378
rect 34642 4326 34654 4378
rect 34706 4326 34718 4378
rect 34770 4326 34782 4378
rect 34834 4326 34840 4378
rect 1104 4304 34840 4326
rect 12802 4264 12808 4276
rect 11900 4236 12808 4264
rect 11900 4137 11928 4236
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 14185 4267 14243 4273
rect 14185 4233 14197 4267
rect 14231 4264 14243 4267
rect 14642 4264 14648 4276
rect 14231 4236 14648 4264
rect 14231 4233 14243 4236
rect 14185 4227 14243 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 23474 4224 23480 4276
rect 23532 4224 23538 4276
rect 24394 4224 24400 4276
rect 24452 4224 24458 4276
rect 25958 4224 25964 4276
rect 26016 4224 26022 4276
rect 28721 4267 28779 4273
rect 26620 4236 27660 4264
rect 14366 4196 14372 4208
rect 13386 4168 14372 4196
rect 14366 4156 14372 4168
rect 14424 4156 14430 4208
rect 17126 4196 17132 4208
rect 15226 4168 17132 4196
rect 17126 4156 17132 4168
rect 17184 4156 17190 4208
rect 19978 4196 19984 4208
rect 18998 4168 19984 4196
rect 19978 4156 19984 4168
rect 20036 4156 20042 4208
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 19705 4131 19763 4137
rect 19705 4097 19717 4131
rect 19751 4128 19763 4131
rect 19886 4128 19892 4140
rect 19751 4100 19892 4128
rect 19751 4097 19763 4100
rect 19705 4091 19763 4097
rect 19886 4088 19892 4100
rect 19944 4088 19950 4140
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 22189 4131 22247 4137
rect 22189 4097 22201 4131
rect 22235 4128 22247 4131
rect 23492 4128 23520 4224
rect 24412 4196 24440 4224
rect 26620 4208 26648 4236
rect 23952 4168 24440 4196
rect 23952 4137 23980 4168
rect 24486 4156 24492 4208
rect 24544 4196 24550 4208
rect 24544 4168 24978 4196
rect 24544 4156 24550 4168
rect 26602 4156 26608 4208
rect 26660 4156 26666 4208
rect 26786 4156 26792 4208
rect 26844 4196 26850 4208
rect 27249 4199 27307 4205
rect 27249 4196 27261 4199
rect 26844 4168 27261 4196
rect 26844 4156 26850 4168
rect 27249 4165 27261 4168
rect 27295 4165 27307 4199
rect 27632 4196 27660 4236
rect 28721 4233 28733 4267
rect 28767 4264 28779 4267
rect 28902 4264 28908 4276
rect 28767 4236 28908 4264
rect 28767 4233 28779 4236
rect 28721 4227 28779 4233
rect 28902 4224 28908 4236
rect 28960 4224 28966 4276
rect 30190 4224 30196 4276
rect 30248 4224 30254 4276
rect 32122 4196 32128 4208
rect 27632 4168 27738 4196
rect 31234 4168 32128 4196
rect 27249 4159 27307 4165
rect 32122 4156 32128 4168
rect 32180 4156 32186 4208
rect 22235 4100 23520 4128
rect 23937 4131 23995 4137
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 23937 4097 23949 4131
rect 23983 4097 23995 4131
rect 23937 4091 23995 4097
rect 12158 4020 12164 4072
rect 12216 4020 12222 4072
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 13633 4063 13691 4069
rect 12860 4032 13584 4060
rect 12860 4020 12866 4032
rect 13556 3924 13584 4032
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 13814 4060 13820 4072
rect 13679 4032 13820 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 15654 4020 15660 4072
rect 15712 4020 15718 4072
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15856 4032 15945 4060
rect 15856 3924 15884 4032
rect 15933 4029 15945 4032
rect 15979 4060 15991 4063
rect 16482 4060 16488 4072
rect 15979 4032 16488 4060
rect 15979 4029 15991 4032
rect 15933 4023 15991 4029
rect 16482 4020 16488 4032
rect 16540 4020 16546 4072
rect 17957 4063 18015 4069
rect 17957 4029 17969 4063
rect 18003 4060 18015 4063
rect 18230 4060 18236 4072
rect 18003 4032 18236 4060
rect 18003 4029 18015 4032
rect 17957 4023 18015 4029
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 19426 4020 19432 4072
rect 19484 4020 19490 4072
rect 22112 4060 22140 4091
rect 24210 4088 24216 4140
rect 24268 4088 24274 4140
rect 26970 4088 26976 4140
rect 27028 4088 27034 4140
rect 31941 4131 31999 4137
rect 31941 4097 31953 4131
rect 31987 4128 31999 4131
rect 34330 4128 34336 4140
rect 31987 4100 34336 4128
rect 31987 4097 31999 4100
rect 31941 4091 31999 4097
rect 34330 4088 34336 4100
rect 34388 4088 34394 4140
rect 22370 4060 22376 4072
rect 22112 4032 22376 4060
rect 22370 4020 22376 4032
rect 22428 4020 22434 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 24136 4032 24501 4060
rect 24136 4001 24164 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 31662 4020 31668 4072
rect 31720 4020 31726 4072
rect 24121 3995 24179 4001
rect 24121 3961 24133 3995
rect 24167 3961 24179 3995
rect 24121 3955 24179 3961
rect 13556 3896 15884 3924
rect 1104 3834 34684 3856
rect 1104 3782 5147 3834
rect 5199 3782 5211 3834
rect 5263 3782 5275 3834
rect 5327 3782 5339 3834
rect 5391 3782 5403 3834
rect 5455 3782 13541 3834
rect 13593 3782 13605 3834
rect 13657 3782 13669 3834
rect 13721 3782 13733 3834
rect 13785 3782 13797 3834
rect 13849 3782 21935 3834
rect 21987 3782 21999 3834
rect 22051 3782 22063 3834
rect 22115 3782 22127 3834
rect 22179 3782 22191 3834
rect 22243 3782 30329 3834
rect 30381 3782 30393 3834
rect 30445 3782 30457 3834
rect 30509 3782 30521 3834
rect 30573 3782 30585 3834
rect 30637 3782 34684 3834
rect 1104 3760 34684 3782
rect 16761 3723 16819 3729
rect 16761 3689 16773 3723
rect 16807 3720 16819 3723
rect 18138 3720 18144 3732
rect 16807 3692 18144 3720
rect 16807 3689 16819 3692
rect 16761 3683 16819 3689
rect 18138 3680 18144 3692
rect 18196 3680 18202 3732
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3584 18567 3587
rect 19334 3584 19340 3596
rect 18555 3556 19340 3584
rect 18555 3553 18567 3556
rect 18509 3547 18567 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 17126 3476 17132 3528
rect 17184 3476 17190 3528
rect 18233 3451 18291 3457
rect 18233 3417 18245 3451
rect 18279 3448 18291 3451
rect 24578 3448 24584 3460
rect 18279 3420 24584 3448
rect 18279 3417 18291 3420
rect 18233 3411 18291 3417
rect 24578 3408 24584 3420
rect 24636 3408 24642 3460
rect 1104 3290 34840 3312
rect 1104 3238 9344 3290
rect 9396 3238 9408 3290
rect 9460 3238 9472 3290
rect 9524 3238 9536 3290
rect 9588 3238 9600 3290
rect 9652 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 17930 3290
rect 17982 3238 17994 3290
rect 18046 3238 26132 3290
rect 26184 3238 26196 3290
rect 26248 3238 26260 3290
rect 26312 3238 26324 3290
rect 26376 3238 26388 3290
rect 26440 3238 34526 3290
rect 34578 3238 34590 3290
rect 34642 3238 34654 3290
rect 34706 3238 34718 3290
rect 34770 3238 34782 3290
rect 34834 3238 34840 3290
rect 1104 3216 34840 3238
rect 1104 2746 34684 2768
rect 1104 2694 5147 2746
rect 5199 2694 5211 2746
rect 5263 2694 5275 2746
rect 5327 2694 5339 2746
rect 5391 2694 5403 2746
rect 5455 2694 13541 2746
rect 13593 2694 13605 2746
rect 13657 2694 13669 2746
rect 13721 2694 13733 2746
rect 13785 2694 13797 2746
rect 13849 2694 21935 2746
rect 21987 2694 21999 2746
rect 22051 2694 22063 2746
rect 22115 2694 22127 2746
rect 22179 2694 22191 2746
rect 22243 2694 30329 2746
rect 30381 2694 30393 2746
rect 30445 2694 30457 2746
rect 30509 2694 30521 2746
rect 30573 2694 30585 2746
rect 30637 2694 34684 2746
rect 1104 2672 34684 2694
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 7466 2632 7472 2644
rect 6135 2604 7472 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 12216 2604 12357 2632
rect 12216 2592 12222 2604
rect 12345 2601 12357 2604
rect 12391 2601 12403 2635
rect 12345 2595 12403 2601
rect 24578 2592 24584 2644
rect 24636 2592 24642 2644
rect 31205 2635 31263 2641
rect 31205 2601 31217 2635
rect 31251 2632 31263 2635
rect 31662 2632 31668 2644
rect 31251 2604 31668 2632
rect 31251 2601 31263 2604
rect 31205 2595 31263 2601
rect 31662 2592 31668 2604
rect 31720 2592 31726 2644
rect 34149 2567 34207 2573
rect 34149 2564 34161 2567
rect 26206 2536 34161 2564
rect 15654 2456 15660 2508
rect 15712 2496 15718 2508
rect 26206 2496 26234 2536
rect 34149 2533 34161 2536
rect 34195 2533 34207 2567
rect 34149 2527 34207 2533
rect 15712 2468 26234 2496
rect 15712 2456 15718 2468
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 5902 2388 5908 2440
rect 5960 2388 5966 2440
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12308 2400 12541 2428
rect 12308 2388 12314 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 17000 2400 19349 2428
rect 17000 2388 17006 2400
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 19337 2391 19395 2397
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24544 2400 24777 2428
rect 24544 2388 24550 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 31018 2388 31024 2440
rect 31076 2388 31082 2440
rect 34333 2431 34391 2437
rect 34333 2397 34345 2431
rect 34379 2428 34391 2431
rect 34379 2400 34468 2428
rect 34379 2397 34391 2400
rect 34333 2391 34391 2397
rect 34440 2304 34468 2400
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 11790 2292 11796 2304
rect 1627 2264 11796 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 11790 2252 11796 2264
rect 11848 2252 11854 2304
rect 19058 2252 19064 2304
rect 19116 2292 19122 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 19116 2264 19441 2292
rect 19116 2252 19122 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 34422 2252 34428 2304
rect 34480 2252 34486 2304
rect 1104 2202 34840 2224
rect 1104 2150 9344 2202
rect 9396 2150 9408 2202
rect 9460 2150 9472 2202
rect 9524 2150 9536 2202
rect 9588 2150 9600 2202
rect 9652 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 17930 2202
rect 17982 2150 17994 2202
rect 18046 2150 26132 2202
rect 26184 2150 26196 2202
rect 26248 2150 26260 2202
rect 26312 2150 26324 2202
rect 26376 2150 26388 2202
rect 26440 2150 34526 2202
rect 34578 2150 34590 2202
rect 34642 2150 34654 2202
rect 34706 2150 34718 2202
rect 34770 2150 34782 2202
rect 34834 2150 34840 2202
rect 1104 2128 34840 2150
<< via1 >>
rect 5147 35334 5199 35386
rect 5211 35334 5263 35386
rect 5275 35334 5327 35386
rect 5339 35334 5391 35386
rect 5403 35334 5455 35386
rect 13541 35334 13593 35386
rect 13605 35334 13657 35386
rect 13669 35334 13721 35386
rect 13733 35334 13785 35386
rect 13797 35334 13849 35386
rect 21935 35334 21987 35386
rect 21999 35334 22051 35386
rect 22063 35334 22115 35386
rect 22127 35334 22179 35386
rect 22191 35334 22243 35386
rect 30329 35334 30381 35386
rect 30393 35334 30445 35386
rect 30457 35334 30509 35386
rect 30521 35334 30573 35386
rect 30585 35334 30637 35386
rect 1308 35232 1360 35284
rect 26424 35232 26476 35284
rect 9220 35164 9272 35216
rect 15752 35164 15804 35216
rect 13912 35096 13964 35148
rect 7748 35028 7800 35080
rect 8116 35071 8168 35080
rect 8116 35037 8125 35071
rect 8125 35037 8159 35071
rect 8159 35037 8168 35071
rect 8116 35028 8168 35037
rect 1768 35003 1820 35012
rect 1768 34969 1777 35003
rect 1777 34969 1811 35003
rect 1811 34969 1820 35003
rect 1768 34960 1820 34969
rect 16580 35028 16632 35080
rect 17132 35071 17184 35080
rect 17132 35037 17141 35071
rect 17141 35037 17175 35071
rect 17175 35037 17184 35071
rect 17132 35028 17184 35037
rect 19984 35028 20036 35080
rect 12532 34960 12584 35012
rect 7932 34935 7984 34944
rect 7932 34901 7941 34935
rect 7941 34901 7975 34935
rect 7975 34901 7984 34935
rect 7932 34892 7984 34901
rect 9772 34892 9824 34944
rect 13636 34935 13688 34944
rect 13636 34901 13645 34935
rect 13645 34901 13679 34935
rect 13679 34901 13688 34935
rect 13636 34892 13688 34901
rect 13912 34892 13964 34944
rect 15660 34892 15712 34944
rect 32864 35028 32916 35080
rect 22284 34960 22336 35012
rect 24216 34960 24268 35012
rect 27068 35003 27120 35012
rect 27068 34969 27077 35003
rect 27077 34969 27111 35003
rect 27111 34969 27120 35003
rect 27068 34960 27120 34969
rect 32680 34892 32732 34944
rect 9344 34790 9396 34842
rect 9408 34790 9460 34842
rect 9472 34790 9524 34842
rect 9536 34790 9588 34842
rect 9600 34790 9652 34842
rect 17738 34790 17790 34842
rect 17802 34790 17854 34842
rect 17866 34790 17918 34842
rect 17930 34790 17982 34842
rect 17994 34790 18046 34842
rect 26132 34790 26184 34842
rect 26196 34790 26248 34842
rect 26260 34790 26312 34842
rect 26324 34790 26376 34842
rect 26388 34790 26440 34842
rect 34526 34790 34578 34842
rect 34590 34790 34642 34842
rect 34654 34790 34706 34842
rect 34718 34790 34770 34842
rect 34782 34790 34834 34842
rect 7932 34663 7984 34672
rect 7932 34629 7941 34663
rect 7941 34629 7975 34663
rect 7975 34629 7984 34663
rect 7932 34620 7984 34629
rect 9220 34620 9272 34672
rect 9588 34620 9640 34672
rect 9772 34620 9824 34672
rect 12532 34688 12584 34740
rect 13636 34688 13688 34740
rect 5724 34552 5776 34604
rect 3608 34527 3660 34536
rect 3608 34493 3617 34527
rect 3617 34493 3651 34527
rect 3651 34493 3660 34527
rect 3608 34484 3660 34493
rect 5908 34484 5960 34536
rect 10600 34484 10652 34536
rect 13912 34620 13964 34672
rect 14188 34595 14240 34604
rect 14188 34561 14197 34595
rect 14197 34561 14231 34595
rect 14231 34561 14240 34595
rect 14188 34552 14240 34561
rect 11336 34527 11388 34536
rect 11336 34493 11345 34527
rect 11345 34493 11379 34527
rect 11379 34493 11388 34527
rect 11336 34484 11388 34493
rect 14464 34527 14516 34536
rect 14464 34493 14473 34527
rect 14473 34493 14507 34527
rect 14507 34493 14516 34527
rect 14464 34484 14516 34493
rect 19340 34688 19392 34740
rect 22560 34688 22612 34740
rect 24308 34688 24360 34740
rect 27068 34688 27120 34740
rect 23112 34620 23164 34672
rect 15752 34552 15804 34604
rect 16580 34552 16632 34604
rect 16488 34484 16540 34536
rect 16764 34527 16816 34536
rect 16764 34493 16773 34527
rect 16773 34493 16807 34527
rect 16807 34493 16816 34527
rect 16764 34484 16816 34493
rect 17316 34595 17368 34604
rect 17316 34561 17325 34595
rect 17325 34561 17359 34595
rect 17359 34561 17368 34595
rect 17316 34552 17368 34561
rect 19616 34595 19668 34604
rect 19616 34561 19625 34595
rect 19625 34561 19659 34595
rect 19659 34561 19668 34595
rect 19616 34552 19668 34561
rect 17592 34527 17644 34536
rect 17592 34493 17601 34527
rect 17601 34493 17635 34527
rect 17635 34493 17644 34527
rect 17592 34484 17644 34493
rect 19340 34484 19392 34536
rect 22284 34552 22336 34604
rect 22376 34527 22428 34536
rect 22376 34493 22385 34527
rect 22385 34493 22419 34527
rect 22419 34493 22428 34527
rect 22376 34484 22428 34493
rect 22652 34527 22704 34536
rect 22652 34493 22661 34527
rect 22661 34493 22695 34527
rect 22695 34493 22704 34527
rect 22652 34484 22704 34493
rect 23112 34484 23164 34536
rect 32680 34620 32732 34672
rect 24308 34595 24360 34604
rect 24308 34561 24317 34595
rect 24317 34561 24351 34595
rect 24351 34561 24360 34595
rect 24308 34552 24360 34561
rect 4620 34348 4672 34400
rect 5632 34348 5684 34400
rect 7012 34391 7064 34400
rect 7012 34357 7021 34391
rect 7021 34357 7055 34391
rect 7055 34357 7064 34391
rect 7012 34348 7064 34357
rect 7656 34348 7708 34400
rect 8944 34348 8996 34400
rect 9404 34391 9456 34400
rect 9404 34357 9413 34391
rect 9413 34357 9447 34391
rect 9447 34357 9456 34391
rect 9404 34348 9456 34357
rect 14096 34391 14148 34400
rect 14096 34357 14105 34391
rect 14105 34357 14139 34391
rect 14139 34357 14148 34391
rect 14096 34348 14148 34357
rect 18788 34348 18840 34400
rect 19340 34348 19392 34400
rect 19984 34348 20036 34400
rect 21640 34391 21692 34400
rect 21640 34357 21649 34391
rect 21649 34357 21683 34391
rect 21683 34357 21692 34391
rect 21640 34348 21692 34357
rect 21824 34416 21876 34468
rect 32404 34484 32456 34536
rect 24124 34391 24176 34400
rect 24124 34357 24133 34391
rect 24133 34357 24167 34391
rect 24167 34357 24176 34391
rect 24124 34348 24176 34357
rect 32956 34348 33008 34400
rect 33876 34391 33928 34400
rect 33876 34357 33885 34391
rect 33885 34357 33919 34391
rect 33919 34357 33928 34391
rect 33876 34348 33928 34357
rect 5147 34246 5199 34298
rect 5211 34246 5263 34298
rect 5275 34246 5327 34298
rect 5339 34246 5391 34298
rect 5403 34246 5455 34298
rect 13541 34246 13593 34298
rect 13605 34246 13657 34298
rect 13669 34246 13721 34298
rect 13733 34246 13785 34298
rect 13797 34246 13849 34298
rect 21935 34246 21987 34298
rect 21999 34246 22051 34298
rect 22063 34246 22115 34298
rect 22127 34246 22179 34298
rect 22191 34246 22243 34298
rect 30329 34246 30381 34298
rect 30393 34246 30445 34298
rect 30457 34246 30509 34298
rect 30521 34246 30573 34298
rect 30585 34246 30637 34298
rect 4160 34076 4212 34128
rect 4620 34187 4672 34196
rect 4620 34153 4629 34187
rect 4629 34153 4663 34187
rect 4663 34153 4672 34187
rect 4620 34144 4672 34153
rect 7932 34144 7984 34196
rect 8116 34144 8168 34196
rect 14464 34144 14516 34196
rect 16764 34144 16816 34196
rect 17592 34144 17644 34196
rect 19616 34144 19668 34196
rect 22652 34144 22704 34196
rect 9588 34076 9640 34128
rect 7656 34008 7708 34060
rect 14096 34008 14148 34060
rect 14188 34008 14240 34060
rect 15108 34008 15160 34060
rect 17316 34008 17368 34060
rect 18788 34051 18840 34060
rect 18788 34017 18797 34051
rect 18797 34017 18831 34051
rect 18831 34017 18840 34051
rect 18788 34008 18840 34017
rect 23388 34008 23440 34060
rect 3976 33983 4028 33992
rect 3976 33949 3985 33983
rect 3985 33949 4019 33983
rect 4019 33949 4028 33983
rect 3976 33940 4028 33949
rect 4344 33847 4396 33856
rect 4344 33813 4353 33847
rect 4353 33813 4387 33847
rect 4387 33813 4396 33847
rect 4344 33804 4396 33813
rect 5724 33940 5776 33992
rect 6828 33915 6880 33924
rect 6828 33881 6837 33915
rect 6837 33881 6871 33915
rect 6871 33881 6880 33915
rect 6828 33872 6880 33881
rect 9404 33940 9456 33992
rect 8024 33872 8076 33924
rect 8300 33915 8352 33924
rect 8300 33881 8309 33915
rect 8309 33881 8343 33915
rect 8343 33881 8352 33915
rect 8300 33872 8352 33881
rect 15660 33872 15712 33924
rect 5908 33804 5960 33856
rect 7104 33804 7156 33856
rect 16488 33804 16540 33856
rect 19340 33940 19392 33992
rect 24216 34008 24268 34060
rect 19340 33804 19392 33856
rect 20168 33847 20220 33856
rect 20168 33813 20177 33847
rect 20177 33813 20211 33847
rect 20211 33813 20220 33847
rect 20168 33804 20220 33813
rect 20720 33804 20772 33856
rect 24124 33940 24176 33992
rect 26792 33983 26844 33992
rect 26792 33949 26801 33983
rect 26801 33949 26835 33983
rect 26835 33949 26844 33983
rect 26792 33940 26844 33949
rect 23756 33847 23808 33856
rect 23756 33813 23765 33847
rect 23765 33813 23799 33847
rect 23799 33813 23808 33847
rect 23756 33804 23808 33813
rect 23940 33804 23992 33856
rect 25044 33847 25096 33856
rect 25044 33813 25053 33847
rect 25053 33813 25087 33847
rect 25087 33813 25096 33847
rect 25044 33804 25096 33813
rect 26516 33915 26568 33924
rect 26516 33881 26525 33915
rect 26525 33881 26559 33915
rect 26559 33881 26568 33915
rect 26516 33872 26568 33881
rect 33876 34008 33928 34060
rect 32956 33872 33008 33924
rect 27160 33804 27212 33856
rect 34336 33847 34388 33856
rect 34336 33813 34345 33847
rect 34345 33813 34379 33847
rect 34379 33813 34388 33847
rect 34336 33804 34388 33813
rect 9344 33702 9396 33754
rect 9408 33702 9460 33754
rect 9472 33702 9524 33754
rect 9536 33702 9588 33754
rect 9600 33702 9652 33754
rect 17738 33702 17790 33754
rect 17802 33702 17854 33754
rect 17866 33702 17918 33754
rect 17930 33702 17982 33754
rect 17994 33702 18046 33754
rect 26132 33702 26184 33754
rect 26196 33702 26248 33754
rect 26260 33702 26312 33754
rect 26324 33702 26376 33754
rect 26388 33702 26440 33754
rect 34526 33702 34578 33754
rect 34590 33702 34642 33754
rect 34654 33702 34706 33754
rect 34718 33702 34770 33754
rect 34782 33702 34834 33754
rect 4344 33600 4396 33652
rect 5908 33600 5960 33652
rect 6828 33600 6880 33652
rect 5816 33532 5868 33584
rect 17500 33600 17552 33652
rect 5816 33439 5868 33448
rect 5816 33405 5825 33439
rect 5825 33405 5859 33439
rect 5859 33405 5868 33439
rect 5816 33396 5868 33405
rect 5908 33439 5960 33448
rect 5908 33405 5917 33439
rect 5917 33405 5951 33439
rect 5951 33405 5960 33439
rect 5908 33396 5960 33405
rect 6000 33439 6052 33448
rect 6000 33405 6009 33439
rect 6009 33405 6043 33439
rect 6043 33405 6052 33439
rect 6000 33396 6052 33405
rect 6552 33507 6604 33516
rect 6552 33473 6561 33507
rect 6561 33473 6595 33507
rect 6595 33473 6604 33507
rect 6552 33464 6604 33473
rect 7012 33507 7064 33516
rect 7012 33473 7021 33507
rect 7021 33473 7055 33507
rect 7055 33473 7064 33507
rect 7012 33464 7064 33473
rect 19984 33600 20036 33652
rect 20168 33600 20220 33652
rect 21088 33600 21140 33652
rect 21640 33600 21692 33652
rect 23756 33600 23808 33652
rect 24768 33600 24820 33652
rect 25044 33600 25096 33652
rect 26516 33600 26568 33652
rect 19708 33532 19760 33584
rect 7104 33439 7156 33448
rect 7104 33405 7113 33439
rect 7113 33405 7147 33439
rect 7147 33405 7156 33439
rect 7104 33396 7156 33405
rect 6184 33328 6236 33380
rect 8300 33464 8352 33516
rect 8852 33507 8904 33516
rect 8852 33473 8861 33507
rect 8861 33473 8895 33507
rect 8895 33473 8904 33507
rect 8852 33464 8904 33473
rect 16672 33507 16724 33516
rect 16672 33473 16681 33507
rect 16681 33473 16715 33507
rect 16715 33473 16724 33507
rect 16672 33464 16724 33473
rect 19248 33464 19300 33516
rect 17224 33439 17276 33448
rect 17224 33405 17233 33439
rect 17233 33405 17267 33439
rect 17267 33405 17276 33439
rect 17224 33396 17276 33405
rect 13452 33328 13504 33380
rect 3976 33260 4028 33312
rect 5632 33260 5684 33312
rect 5908 33260 5960 33312
rect 6368 33260 6420 33312
rect 9128 33260 9180 33312
rect 17040 33260 17092 33312
rect 20536 33464 20588 33516
rect 23112 33532 23164 33584
rect 20720 33396 20772 33448
rect 21824 33439 21876 33448
rect 21824 33405 21833 33439
rect 21833 33405 21867 33439
rect 21867 33405 21876 33439
rect 21824 33396 21876 33405
rect 22192 33396 22244 33448
rect 25964 33439 26016 33448
rect 25964 33405 25973 33439
rect 25973 33405 26007 33439
rect 26007 33405 26016 33439
rect 25964 33396 26016 33405
rect 19340 33328 19392 33380
rect 19524 33303 19576 33312
rect 19524 33269 19533 33303
rect 19533 33269 19567 33303
rect 19567 33269 19576 33303
rect 19524 33260 19576 33269
rect 20536 33260 20588 33312
rect 20996 33260 21048 33312
rect 23572 33303 23624 33312
rect 23572 33269 23581 33303
rect 23581 33269 23615 33303
rect 23615 33269 23624 33303
rect 23572 33260 23624 33269
rect 5147 33158 5199 33210
rect 5211 33158 5263 33210
rect 5275 33158 5327 33210
rect 5339 33158 5391 33210
rect 5403 33158 5455 33210
rect 13541 33158 13593 33210
rect 13605 33158 13657 33210
rect 13669 33158 13721 33210
rect 13733 33158 13785 33210
rect 13797 33158 13849 33210
rect 21935 33158 21987 33210
rect 21999 33158 22051 33210
rect 22063 33158 22115 33210
rect 22127 33158 22179 33210
rect 22191 33158 22243 33210
rect 30329 33158 30381 33210
rect 30393 33158 30445 33210
rect 30457 33158 30509 33210
rect 30521 33158 30573 33210
rect 30585 33158 30637 33210
rect 6552 33056 6604 33108
rect 7932 33056 7984 33108
rect 8300 33056 8352 33108
rect 8852 33056 8904 33108
rect 6184 32988 6236 33040
rect 940 32852 992 32904
rect 3976 32852 4028 32904
rect 5816 32852 5868 32904
rect 6184 32895 6236 32904
rect 6184 32861 6193 32895
rect 6193 32861 6227 32895
rect 6227 32861 6236 32895
rect 6184 32852 6236 32861
rect 6276 32895 6328 32904
rect 6276 32861 6285 32895
rect 6285 32861 6319 32895
rect 6319 32861 6328 32895
rect 6276 32852 6328 32861
rect 6368 32895 6420 32904
rect 6368 32861 6377 32895
rect 6377 32861 6411 32895
rect 6411 32861 6420 32895
rect 6368 32852 6420 32861
rect 8024 32852 8076 32904
rect 8944 32895 8996 32904
rect 8944 32861 8953 32895
rect 8953 32861 8987 32895
rect 8987 32861 8996 32895
rect 8944 32852 8996 32861
rect 12808 32895 12860 32904
rect 12808 32861 12817 32895
rect 12817 32861 12851 32895
rect 12851 32861 12860 32895
rect 12808 32852 12860 32861
rect 13452 32920 13504 32972
rect 14740 32895 14792 32904
rect 14740 32861 14749 32895
rect 14749 32861 14783 32895
rect 14783 32861 14792 32895
rect 14740 32852 14792 32861
rect 19708 33056 19760 33108
rect 22284 33056 22336 33108
rect 23020 33056 23072 33108
rect 24584 33056 24636 33108
rect 25964 33056 26016 33108
rect 15108 32963 15160 32972
rect 15108 32929 15117 32963
rect 15117 32929 15151 32963
rect 15151 32929 15160 32963
rect 15108 32920 15160 32929
rect 16672 32988 16724 33040
rect 16580 32920 16632 32972
rect 17224 32963 17276 32972
rect 17224 32929 17233 32963
rect 17233 32929 17267 32963
rect 17267 32929 17276 32963
rect 17224 32920 17276 32929
rect 19248 32895 19300 32904
rect 19248 32861 19257 32895
rect 19257 32861 19291 32895
rect 19291 32861 19300 32895
rect 19248 32852 19300 32861
rect 3516 32716 3568 32768
rect 3884 32759 3936 32768
rect 3884 32725 3893 32759
rect 3893 32725 3927 32759
rect 3927 32725 3936 32759
rect 3884 32716 3936 32725
rect 4896 32716 4948 32768
rect 8484 32759 8536 32768
rect 8484 32725 8493 32759
rect 8493 32725 8527 32759
rect 8527 32725 8536 32759
rect 8484 32716 8536 32725
rect 9128 32784 9180 32836
rect 9680 32784 9732 32836
rect 15384 32784 15436 32836
rect 19340 32784 19392 32836
rect 20996 32852 21048 32904
rect 23388 32920 23440 32972
rect 23572 32920 23624 32972
rect 24308 32920 24360 32972
rect 9864 32716 9916 32768
rect 10692 32759 10744 32768
rect 10692 32725 10701 32759
rect 10701 32725 10735 32759
rect 10735 32725 10744 32759
rect 10692 32716 10744 32725
rect 17592 32716 17644 32768
rect 19524 32716 19576 32768
rect 19616 32759 19668 32768
rect 19616 32725 19625 32759
rect 19625 32725 19659 32759
rect 19659 32725 19668 32759
rect 19616 32716 19668 32725
rect 24768 32895 24820 32904
rect 24768 32861 24777 32895
rect 24777 32861 24811 32895
rect 24811 32861 24820 32895
rect 24768 32852 24820 32861
rect 24400 32784 24452 32836
rect 24952 32827 25004 32836
rect 24952 32793 24961 32827
rect 24961 32793 24995 32827
rect 24995 32793 25004 32827
rect 24952 32784 25004 32793
rect 25044 32827 25096 32836
rect 25044 32793 25053 32827
rect 25053 32793 25087 32827
rect 25087 32793 25096 32827
rect 25044 32784 25096 32793
rect 32404 32920 32456 32972
rect 26976 32895 27028 32904
rect 26976 32861 26985 32895
rect 26985 32861 27019 32895
rect 27019 32861 27028 32895
rect 26976 32852 27028 32861
rect 32956 32852 33008 32904
rect 34336 32784 34388 32836
rect 28356 32716 28408 32768
rect 32588 32759 32640 32768
rect 32588 32725 32597 32759
rect 32597 32725 32631 32759
rect 32631 32725 32640 32759
rect 32588 32716 32640 32725
rect 9344 32614 9396 32666
rect 9408 32614 9460 32666
rect 9472 32614 9524 32666
rect 9536 32614 9588 32666
rect 9600 32614 9652 32666
rect 17738 32614 17790 32666
rect 17802 32614 17854 32666
rect 17866 32614 17918 32666
rect 17930 32614 17982 32666
rect 17994 32614 18046 32666
rect 26132 32614 26184 32666
rect 26196 32614 26248 32666
rect 26260 32614 26312 32666
rect 26324 32614 26376 32666
rect 26388 32614 26440 32666
rect 34526 32614 34578 32666
rect 34590 32614 34642 32666
rect 34654 32614 34706 32666
rect 34718 32614 34770 32666
rect 34782 32614 34834 32666
rect 3884 32555 3936 32564
rect 3884 32521 3893 32555
rect 3893 32521 3927 32555
rect 3927 32521 3936 32555
rect 3884 32512 3936 32521
rect 8024 32555 8076 32564
rect 8024 32521 8033 32555
rect 8033 32521 8067 32555
rect 8067 32521 8076 32555
rect 8024 32512 8076 32521
rect 8484 32512 8536 32564
rect 9680 32512 9732 32564
rect 10324 32512 10376 32564
rect 10692 32512 10744 32564
rect 4344 32444 4396 32496
rect 6276 32444 6328 32496
rect 8208 32487 8260 32496
rect 8208 32453 8235 32487
rect 8235 32453 8260 32487
rect 8208 32444 8260 32453
rect 9036 32444 9088 32496
rect 2136 32351 2188 32360
rect 2136 32317 2145 32351
rect 2145 32317 2179 32351
rect 2179 32317 2188 32351
rect 2136 32308 2188 32317
rect 2780 32172 2832 32224
rect 3608 32308 3660 32360
rect 4620 32419 4672 32428
rect 4620 32385 4629 32419
rect 4629 32385 4663 32419
rect 4663 32385 4672 32419
rect 4620 32376 4672 32385
rect 6920 32351 6972 32360
rect 6920 32317 6929 32351
rect 6929 32317 6963 32351
rect 6963 32317 6972 32351
rect 6920 32308 6972 32317
rect 6368 32240 6420 32292
rect 3608 32215 3660 32224
rect 3608 32181 3617 32215
rect 3617 32181 3651 32215
rect 3651 32181 3660 32215
rect 3608 32172 3660 32181
rect 3700 32215 3752 32224
rect 3700 32181 3709 32215
rect 3709 32181 3743 32215
rect 3743 32181 3752 32215
rect 3700 32172 3752 32181
rect 4160 32172 4212 32224
rect 4252 32172 4304 32224
rect 4988 32172 5040 32224
rect 6552 32215 6604 32224
rect 6552 32181 6561 32215
rect 6561 32181 6595 32215
rect 6595 32181 6604 32215
rect 6552 32172 6604 32181
rect 15108 32512 15160 32564
rect 15384 32555 15436 32564
rect 15384 32521 15393 32555
rect 15393 32521 15427 32555
rect 15427 32521 15436 32555
rect 15384 32512 15436 32521
rect 16672 32512 16724 32564
rect 17040 32555 17092 32564
rect 17040 32521 17049 32555
rect 17049 32521 17083 32555
rect 17083 32521 17092 32555
rect 17040 32512 17092 32521
rect 17592 32512 17644 32564
rect 14096 32444 14148 32496
rect 14740 32444 14792 32496
rect 12348 32376 12400 32428
rect 13820 32376 13872 32428
rect 15016 32376 15068 32428
rect 9128 32351 9180 32360
rect 9128 32317 9137 32351
rect 9137 32317 9171 32351
rect 9171 32317 9180 32351
rect 9128 32308 9180 32317
rect 9680 32308 9732 32360
rect 12716 32351 12768 32360
rect 12716 32317 12725 32351
rect 12725 32317 12759 32351
rect 12759 32317 12768 32351
rect 12716 32308 12768 32317
rect 9128 32172 9180 32224
rect 19616 32512 19668 32564
rect 17592 32419 17644 32428
rect 17592 32385 17601 32419
rect 17601 32385 17635 32419
rect 17635 32385 17644 32419
rect 17592 32376 17644 32385
rect 17776 32419 17828 32428
rect 17776 32385 17785 32419
rect 17785 32385 17819 32419
rect 17819 32385 17828 32419
rect 17776 32376 17828 32385
rect 20352 32419 20404 32428
rect 20352 32385 20361 32419
rect 20361 32385 20395 32419
rect 20395 32385 20404 32419
rect 20352 32376 20404 32385
rect 20536 32419 20588 32428
rect 20536 32385 20545 32419
rect 20545 32385 20579 32419
rect 20579 32385 20588 32419
rect 20536 32376 20588 32385
rect 20720 32376 20772 32428
rect 25044 32512 25096 32564
rect 23848 32487 23900 32496
rect 23848 32453 23857 32487
rect 23857 32453 23891 32487
rect 23891 32453 23900 32487
rect 23848 32444 23900 32453
rect 24308 32444 24360 32496
rect 26976 32444 27028 32496
rect 27160 32444 27212 32496
rect 28540 32444 28592 32496
rect 14004 32240 14056 32292
rect 14188 32215 14240 32224
rect 14188 32181 14197 32215
rect 14197 32181 14231 32215
rect 14231 32181 14240 32215
rect 14188 32172 14240 32181
rect 14280 32215 14332 32224
rect 14280 32181 14289 32215
rect 14289 32181 14323 32215
rect 14323 32181 14332 32215
rect 14280 32172 14332 32181
rect 17408 32351 17460 32360
rect 17408 32317 17417 32351
rect 17417 32317 17451 32351
rect 17451 32317 17460 32351
rect 17408 32308 17460 32317
rect 20996 32351 21048 32360
rect 20996 32317 21005 32351
rect 21005 32317 21039 32351
rect 21039 32317 21048 32351
rect 20996 32308 21048 32317
rect 21088 32351 21140 32360
rect 21088 32317 21097 32351
rect 21097 32317 21131 32351
rect 21131 32317 21140 32351
rect 21088 32308 21140 32317
rect 17592 32240 17644 32292
rect 19984 32240 20036 32292
rect 20720 32240 20772 32292
rect 23756 32419 23808 32428
rect 23756 32385 23765 32419
rect 23765 32385 23799 32419
rect 23799 32385 23808 32419
rect 23756 32376 23808 32385
rect 24400 32376 24452 32428
rect 24584 32376 24636 32428
rect 26516 32419 26568 32428
rect 26516 32385 26525 32419
rect 26525 32385 26559 32419
rect 26559 32385 26568 32419
rect 26516 32376 26568 32385
rect 26792 32376 26844 32428
rect 20168 32172 20220 32224
rect 20628 32215 20680 32224
rect 20628 32181 20637 32215
rect 20637 32181 20671 32215
rect 20671 32181 20680 32215
rect 20628 32172 20680 32181
rect 23940 32172 23992 32224
rect 24124 32215 24176 32224
rect 24124 32181 24133 32215
rect 24133 32181 24167 32215
rect 24167 32181 24176 32215
rect 24124 32172 24176 32181
rect 25136 32308 25188 32360
rect 25688 32351 25740 32360
rect 25688 32317 25697 32351
rect 25697 32317 25731 32351
rect 25731 32317 25740 32351
rect 25688 32308 25740 32317
rect 28816 32444 28868 32496
rect 32404 32376 32456 32428
rect 28908 32308 28960 32360
rect 26976 32215 27028 32224
rect 26976 32181 26985 32215
rect 26985 32181 27019 32215
rect 27019 32181 27028 32215
rect 26976 32172 27028 32181
rect 27160 32172 27212 32224
rect 27988 32172 28040 32224
rect 28816 32172 28868 32224
rect 5147 32070 5199 32122
rect 5211 32070 5263 32122
rect 5275 32070 5327 32122
rect 5339 32070 5391 32122
rect 5403 32070 5455 32122
rect 13541 32070 13593 32122
rect 13605 32070 13657 32122
rect 13669 32070 13721 32122
rect 13733 32070 13785 32122
rect 13797 32070 13849 32122
rect 21935 32070 21987 32122
rect 21999 32070 22051 32122
rect 22063 32070 22115 32122
rect 22127 32070 22179 32122
rect 22191 32070 22243 32122
rect 30329 32070 30381 32122
rect 30393 32070 30445 32122
rect 30457 32070 30509 32122
rect 30521 32070 30573 32122
rect 30585 32070 30637 32122
rect 2136 31968 2188 32020
rect 3700 31968 3752 32020
rect 4252 31968 4304 32020
rect 3608 31832 3660 31884
rect 3976 31764 4028 31816
rect 4896 31968 4948 32020
rect 8208 31968 8260 32020
rect 6276 31900 6328 31952
rect 5816 31832 5868 31884
rect 4436 31696 4488 31748
rect 4804 31671 4856 31680
rect 4804 31637 4813 31671
rect 4813 31637 4847 31671
rect 4847 31637 4856 31671
rect 4804 31628 4856 31637
rect 4988 31739 5040 31748
rect 4988 31705 4997 31739
rect 4997 31705 5031 31739
rect 5031 31705 5040 31739
rect 4988 31696 5040 31705
rect 5540 31764 5592 31816
rect 6368 31807 6420 31816
rect 6368 31773 6377 31807
rect 6377 31773 6411 31807
rect 6411 31773 6420 31807
rect 6368 31764 6420 31773
rect 5632 31696 5684 31748
rect 8576 31832 8628 31884
rect 8300 31807 8352 31816
rect 8300 31773 8309 31807
rect 8309 31773 8343 31807
rect 8343 31773 8352 31807
rect 8300 31764 8352 31773
rect 9220 31900 9272 31952
rect 9864 31968 9916 32020
rect 12716 31968 12768 32020
rect 14096 32011 14148 32020
rect 14096 31977 14105 32011
rect 14105 31977 14139 32011
rect 14139 31977 14148 32011
rect 14096 31968 14148 31977
rect 14280 31968 14332 32020
rect 17408 31968 17460 32020
rect 17776 32011 17828 32020
rect 17776 31977 17785 32011
rect 17785 31977 17819 32011
rect 17819 31977 17828 32011
rect 17776 31968 17828 31977
rect 9680 31764 9732 31816
rect 10600 31764 10652 31816
rect 12348 31832 12400 31884
rect 14004 31900 14056 31952
rect 11704 31739 11756 31748
rect 11704 31705 11713 31739
rect 11713 31705 11747 31739
rect 11747 31705 11756 31739
rect 11704 31696 11756 31705
rect 5724 31628 5776 31680
rect 5908 31628 5960 31680
rect 6092 31671 6144 31680
rect 6092 31637 6101 31671
rect 6101 31637 6135 31671
rect 6135 31637 6144 31671
rect 6092 31628 6144 31637
rect 8116 31628 8168 31680
rect 9128 31628 9180 31680
rect 9956 31671 10008 31680
rect 9956 31637 9965 31671
rect 9965 31637 9999 31671
rect 9999 31637 10008 31671
rect 9956 31628 10008 31637
rect 10416 31628 10468 31680
rect 14188 31764 14240 31816
rect 15016 31764 15068 31816
rect 17132 31807 17184 31816
rect 17132 31773 17141 31807
rect 17141 31773 17175 31807
rect 17175 31773 17184 31807
rect 17132 31764 17184 31773
rect 19524 31968 19576 32020
rect 20628 31968 20680 32020
rect 19984 31943 20036 31952
rect 19984 31909 19993 31943
rect 19993 31909 20027 31943
rect 20027 31909 20036 31943
rect 19984 31900 20036 31909
rect 20168 31900 20220 31952
rect 17592 31807 17644 31816
rect 17592 31773 17606 31807
rect 17606 31773 17640 31807
rect 17640 31773 17644 31807
rect 17592 31764 17644 31773
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 19708 31807 19760 31816
rect 19708 31773 19717 31807
rect 19717 31773 19751 31807
rect 19751 31773 19760 31807
rect 19708 31764 19760 31773
rect 23388 31968 23440 32020
rect 25688 31968 25740 32020
rect 26516 31968 26568 32020
rect 28080 31968 28132 32020
rect 24124 31832 24176 31884
rect 26976 31832 27028 31884
rect 27160 31875 27212 31884
rect 27160 31841 27169 31875
rect 27169 31841 27203 31875
rect 27203 31841 27212 31875
rect 27160 31832 27212 31841
rect 17500 31739 17552 31748
rect 17500 31705 17509 31739
rect 17509 31705 17543 31739
rect 17543 31705 17552 31739
rect 17500 31696 17552 31705
rect 18880 31739 18932 31748
rect 18880 31705 18889 31739
rect 18889 31705 18923 31739
rect 18923 31705 18932 31739
rect 18880 31696 18932 31705
rect 21824 31764 21876 31816
rect 20536 31696 20588 31748
rect 22284 31739 22336 31748
rect 22284 31705 22293 31739
rect 22293 31705 22327 31739
rect 22327 31705 22336 31739
rect 22284 31696 22336 31705
rect 23020 31696 23072 31748
rect 12808 31628 12860 31680
rect 19616 31671 19668 31680
rect 19616 31637 19625 31671
rect 19625 31637 19659 31671
rect 19659 31637 19668 31671
rect 19616 31628 19668 31637
rect 23756 31628 23808 31680
rect 24860 31628 24912 31680
rect 26976 31671 27028 31680
rect 26976 31637 26985 31671
rect 26985 31637 27019 31671
rect 27019 31637 27028 31671
rect 26976 31628 27028 31637
rect 28080 31807 28132 31816
rect 28080 31773 28089 31807
rect 28089 31773 28123 31807
rect 28123 31773 28132 31807
rect 28080 31764 28132 31773
rect 28356 31807 28408 31816
rect 28356 31773 28365 31807
rect 28365 31773 28399 31807
rect 28399 31773 28408 31807
rect 28356 31764 28408 31773
rect 28908 32011 28960 32020
rect 28908 31977 28917 32011
rect 28917 31977 28951 32011
rect 28951 31977 28960 32011
rect 28908 31968 28960 31977
rect 27804 31696 27856 31748
rect 28448 31696 28500 31748
rect 28356 31628 28408 31680
rect 9344 31526 9396 31578
rect 9408 31526 9460 31578
rect 9472 31526 9524 31578
rect 9536 31526 9588 31578
rect 9600 31526 9652 31578
rect 17738 31526 17790 31578
rect 17802 31526 17854 31578
rect 17866 31526 17918 31578
rect 17930 31526 17982 31578
rect 17994 31526 18046 31578
rect 26132 31526 26184 31578
rect 26196 31526 26248 31578
rect 26260 31526 26312 31578
rect 26324 31526 26376 31578
rect 26388 31526 26440 31578
rect 34526 31526 34578 31578
rect 34590 31526 34642 31578
rect 34654 31526 34706 31578
rect 34718 31526 34770 31578
rect 34782 31526 34834 31578
rect 4436 31424 4488 31476
rect 6368 31424 6420 31476
rect 8576 31467 8628 31476
rect 8576 31433 8585 31467
rect 8585 31433 8619 31467
rect 8619 31433 8628 31467
rect 8576 31424 8628 31433
rect 9956 31424 10008 31476
rect 11704 31424 11756 31476
rect 17132 31467 17184 31476
rect 17132 31433 17141 31467
rect 17141 31433 17175 31467
rect 17175 31433 17184 31467
rect 17132 31424 17184 31433
rect 19432 31467 19484 31476
rect 19432 31433 19441 31467
rect 19441 31433 19475 31467
rect 19475 31433 19484 31467
rect 19432 31424 19484 31433
rect 20352 31424 20404 31476
rect 22284 31424 22336 31476
rect 4344 31356 4396 31408
rect 5908 31356 5960 31408
rect 6092 31356 6144 31408
rect 9220 31356 9272 31408
rect 15200 31356 15252 31408
rect 17500 31356 17552 31408
rect 2780 31331 2832 31340
rect 2780 31297 2789 31331
rect 2789 31297 2823 31331
rect 2823 31297 2832 31331
rect 2780 31288 2832 31297
rect 5724 31331 5776 31340
rect 5724 31297 5733 31331
rect 5733 31297 5767 31331
rect 5767 31297 5776 31331
rect 5724 31288 5776 31297
rect 6920 31288 6972 31340
rect 8116 31331 8168 31340
rect 8116 31297 8125 31331
rect 8125 31297 8159 31331
rect 8159 31297 8168 31331
rect 8116 31288 8168 31297
rect 9680 31288 9732 31340
rect 10416 31331 10468 31340
rect 10416 31297 10425 31331
rect 10425 31297 10459 31331
rect 10459 31297 10468 31331
rect 10416 31288 10468 31297
rect 14832 31288 14884 31340
rect 15016 31288 15068 31340
rect 3056 31263 3108 31272
rect 3056 31229 3065 31263
rect 3065 31229 3099 31263
rect 3099 31229 3108 31263
rect 3056 31220 3108 31229
rect 8760 31220 8812 31272
rect 9128 31263 9180 31272
rect 9128 31229 9137 31263
rect 9137 31229 9171 31263
rect 9171 31229 9180 31263
rect 9128 31220 9180 31229
rect 6000 31127 6052 31136
rect 6000 31093 6009 31127
rect 6009 31093 6043 31127
rect 6043 31093 6052 31127
rect 6000 31084 6052 31093
rect 7380 31084 7432 31136
rect 14004 31084 14056 31136
rect 14372 31084 14424 31136
rect 15568 31127 15620 31136
rect 15568 31093 15577 31127
rect 15577 31093 15611 31127
rect 15611 31093 15620 31127
rect 15568 31084 15620 31093
rect 17684 31331 17736 31340
rect 17684 31297 17693 31331
rect 17693 31297 17727 31331
rect 17727 31297 17736 31331
rect 17684 31288 17736 31297
rect 17868 31331 17920 31340
rect 17868 31297 17877 31331
rect 17877 31297 17911 31331
rect 17911 31297 17920 31331
rect 17868 31288 17920 31297
rect 19616 31356 19668 31408
rect 19708 31288 19760 31340
rect 20996 31356 21048 31408
rect 21088 31356 21140 31408
rect 23388 31467 23440 31476
rect 23388 31433 23397 31467
rect 23397 31433 23431 31467
rect 23431 31433 23440 31467
rect 23388 31424 23440 31433
rect 23848 31424 23900 31476
rect 26976 31424 27028 31476
rect 28448 31467 28500 31476
rect 28448 31433 28457 31467
rect 28457 31433 28491 31467
rect 28491 31433 28500 31467
rect 28448 31424 28500 31433
rect 24952 31331 25004 31340
rect 24952 31297 24961 31331
rect 24961 31297 24995 31331
rect 24995 31297 25004 31331
rect 24952 31288 25004 31297
rect 17684 31152 17736 31204
rect 21088 31263 21140 31272
rect 21088 31229 21097 31263
rect 21097 31229 21131 31263
rect 21131 31229 21140 31263
rect 21088 31220 21140 31229
rect 23388 31220 23440 31272
rect 27620 31263 27672 31272
rect 27620 31229 27629 31263
rect 27629 31229 27663 31263
rect 27663 31229 27672 31263
rect 27620 31220 27672 31229
rect 29736 31220 29788 31272
rect 21364 31152 21416 31204
rect 17776 31084 17828 31136
rect 20168 31084 20220 31136
rect 24768 31127 24820 31136
rect 24768 31093 24777 31127
rect 24777 31093 24811 31127
rect 24811 31093 24820 31127
rect 24768 31084 24820 31093
rect 25872 31084 25924 31136
rect 5147 30982 5199 31034
rect 5211 30982 5263 31034
rect 5275 30982 5327 31034
rect 5339 30982 5391 31034
rect 5403 30982 5455 31034
rect 13541 30982 13593 31034
rect 13605 30982 13657 31034
rect 13669 30982 13721 31034
rect 13733 30982 13785 31034
rect 13797 30982 13849 31034
rect 21935 30982 21987 31034
rect 21999 30982 22051 31034
rect 22063 30982 22115 31034
rect 22127 30982 22179 31034
rect 22191 30982 22243 31034
rect 30329 30982 30381 31034
rect 30393 30982 30445 31034
rect 30457 30982 30509 31034
rect 30521 30982 30573 31034
rect 30585 30982 30637 31034
rect 3056 30880 3108 30932
rect 6000 30880 6052 30932
rect 6920 30923 6972 30932
rect 6920 30889 6929 30923
rect 6929 30889 6963 30923
rect 6963 30889 6972 30923
rect 6920 30880 6972 30889
rect 7380 30880 7432 30932
rect 14832 30923 14884 30932
rect 14832 30889 14841 30923
rect 14841 30889 14875 30923
rect 14875 30889 14884 30923
rect 14832 30880 14884 30889
rect 8944 30744 8996 30796
rect 12348 30744 12400 30796
rect 2780 30676 2832 30728
rect 4804 30676 4856 30728
rect 10324 30676 10376 30728
rect 5908 30608 5960 30660
rect 8760 30583 8812 30592
rect 8760 30549 8769 30583
rect 8769 30549 8803 30583
rect 8803 30549 8812 30583
rect 8760 30540 8812 30549
rect 9772 30540 9824 30592
rect 10600 30540 10652 30592
rect 13912 30676 13964 30728
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 14556 30719 14608 30728
rect 14556 30685 14565 30719
rect 14565 30685 14599 30719
rect 14599 30685 14608 30719
rect 14556 30676 14608 30685
rect 17868 30880 17920 30932
rect 18880 30880 18932 30932
rect 21088 30880 21140 30932
rect 21364 30880 21416 30932
rect 24768 30880 24820 30932
rect 27620 30880 27672 30932
rect 17040 30855 17092 30864
rect 17040 30821 17049 30855
rect 17049 30821 17083 30855
rect 17083 30821 17092 30855
rect 17040 30812 17092 30821
rect 17500 30812 17552 30864
rect 17684 30812 17736 30864
rect 17776 30812 17828 30864
rect 15292 30787 15344 30796
rect 15292 30753 15301 30787
rect 15301 30753 15335 30787
rect 15335 30753 15344 30787
rect 15292 30744 15344 30753
rect 15568 30787 15620 30796
rect 15568 30753 15577 30787
rect 15577 30753 15611 30787
rect 15611 30753 15620 30787
rect 15568 30744 15620 30753
rect 17592 30744 17644 30796
rect 13820 30583 13872 30592
rect 13820 30549 13829 30583
rect 13829 30549 13863 30583
rect 13863 30549 13872 30583
rect 16672 30676 16724 30728
rect 15660 30608 15712 30660
rect 17408 30608 17460 30660
rect 13820 30540 13872 30549
rect 15568 30540 15620 30592
rect 18144 30676 18196 30728
rect 21180 30812 21232 30864
rect 20536 30744 20588 30796
rect 21824 30744 21876 30796
rect 21364 30719 21416 30728
rect 21364 30685 21373 30719
rect 21373 30685 21407 30719
rect 21407 30685 21416 30719
rect 21364 30676 21416 30685
rect 21272 30651 21324 30660
rect 21272 30617 21281 30651
rect 21281 30617 21315 30651
rect 21315 30617 21324 30651
rect 21272 30608 21324 30617
rect 25136 30608 25188 30660
rect 26516 30651 26568 30660
rect 26516 30617 26525 30651
rect 26525 30617 26559 30651
rect 26559 30617 26568 30651
rect 26516 30608 26568 30617
rect 27988 30608 28040 30660
rect 28908 30608 28960 30660
rect 25596 30540 25648 30592
rect 27804 30540 27856 30592
rect 28080 30583 28132 30592
rect 28080 30549 28089 30583
rect 28089 30549 28123 30583
rect 28123 30549 28132 30583
rect 28080 30540 28132 30549
rect 9344 30438 9396 30490
rect 9408 30438 9460 30490
rect 9472 30438 9524 30490
rect 9536 30438 9588 30490
rect 9600 30438 9652 30490
rect 17738 30438 17790 30490
rect 17802 30438 17854 30490
rect 17866 30438 17918 30490
rect 17930 30438 17982 30490
rect 17994 30438 18046 30490
rect 26132 30438 26184 30490
rect 26196 30438 26248 30490
rect 26260 30438 26312 30490
rect 26324 30438 26376 30490
rect 26388 30438 26440 30490
rect 34526 30438 34578 30490
rect 34590 30438 34642 30490
rect 34654 30438 34706 30490
rect 34718 30438 34770 30490
rect 34782 30438 34834 30490
rect 14280 30336 14332 30388
rect 15200 30379 15252 30388
rect 15200 30345 15209 30379
rect 15209 30345 15243 30379
rect 15243 30345 15252 30379
rect 15200 30336 15252 30345
rect 15568 30336 15620 30388
rect 15660 30336 15712 30388
rect 17040 30336 17092 30388
rect 21364 30336 21416 30388
rect 24952 30336 25004 30388
rect 25596 30379 25648 30388
rect 25596 30345 25605 30379
rect 25605 30345 25639 30379
rect 25639 30345 25648 30379
rect 25596 30336 25648 30345
rect 6552 30268 6604 30320
rect 8760 30268 8812 30320
rect 6276 30132 6328 30184
rect 6736 30175 6788 30184
rect 6736 30141 6745 30175
rect 6745 30141 6779 30175
rect 6779 30141 6788 30175
rect 6736 30132 6788 30141
rect 6920 29996 6972 30048
rect 9220 30200 9272 30252
rect 9680 30132 9732 30184
rect 9036 30064 9088 30116
rect 13452 30200 13504 30252
rect 13820 30243 13872 30252
rect 13820 30209 13829 30243
rect 13829 30209 13863 30243
rect 13863 30209 13872 30243
rect 13820 30200 13872 30209
rect 13912 30243 13964 30252
rect 13912 30209 13921 30243
rect 13921 30209 13955 30243
rect 13955 30209 13964 30243
rect 13912 30200 13964 30209
rect 14004 30175 14056 30184
rect 14004 30141 14013 30175
rect 14013 30141 14047 30175
rect 14047 30141 14056 30175
rect 21272 30200 21324 30252
rect 23112 30268 23164 30320
rect 24676 30268 24728 30320
rect 26056 30268 26108 30320
rect 26516 30336 26568 30388
rect 28172 30336 28224 30388
rect 29736 30379 29788 30388
rect 29736 30345 29745 30379
rect 29745 30345 29779 30379
rect 29779 30345 29788 30379
rect 29736 30336 29788 30345
rect 14004 30132 14056 30141
rect 15752 30132 15804 30184
rect 16580 30132 16632 30184
rect 17408 30132 17460 30184
rect 20996 30175 21048 30184
rect 20996 30141 21005 30175
rect 21005 30141 21039 30175
rect 21039 30141 21048 30175
rect 20996 30132 21048 30141
rect 21088 30175 21140 30184
rect 21088 30141 21097 30175
rect 21097 30141 21131 30175
rect 21131 30141 21140 30175
rect 21088 30132 21140 30141
rect 21180 30175 21232 30184
rect 21180 30141 21189 30175
rect 21189 30141 21223 30175
rect 21223 30141 21232 30175
rect 21180 30132 21232 30141
rect 9128 29996 9180 30048
rect 9680 29996 9732 30048
rect 9864 30039 9916 30048
rect 9864 30005 9873 30039
rect 9873 30005 9907 30039
rect 9907 30005 9916 30039
rect 9864 29996 9916 30005
rect 10048 30039 10100 30048
rect 10048 30005 10057 30039
rect 10057 30005 10091 30039
rect 10091 30005 10100 30039
rect 10048 29996 10100 30005
rect 17592 29996 17644 30048
rect 20168 30039 20220 30048
rect 20168 30005 20177 30039
rect 20177 30005 20211 30039
rect 20211 30005 20220 30039
rect 20168 29996 20220 30005
rect 24216 30200 24268 30252
rect 24768 30200 24820 30252
rect 25872 30200 25924 30252
rect 21824 30132 21876 30184
rect 22376 30175 22428 30184
rect 22376 30141 22385 30175
rect 22385 30141 22419 30175
rect 22419 30141 22428 30175
rect 22376 30132 22428 30141
rect 23112 30132 23164 30184
rect 23848 30039 23900 30048
rect 23848 30005 23857 30039
rect 23857 30005 23891 30039
rect 23891 30005 23900 30039
rect 23848 29996 23900 30005
rect 25872 29996 25924 30048
rect 26240 30243 26292 30252
rect 26240 30209 26249 30243
rect 26249 30209 26283 30243
rect 26283 30209 26292 30243
rect 26240 30200 26292 30209
rect 28264 30268 28316 30320
rect 28540 30268 28592 30320
rect 29276 30200 29328 30252
rect 28356 30132 28408 30184
rect 28080 29996 28132 30048
rect 5147 29894 5199 29946
rect 5211 29894 5263 29946
rect 5275 29894 5327 29946
rect 5339 29894 5391 29946
rect 5403 29894 5455 29946
rect 13541 29894 13593 29946
rect 13605 29894 13657 29946
rect 13669 29894 13721 29946
rect 13733 29894 13785 29946
rect 13797 29894 13849 29946
rect 21935 29894 21987 29946
rect 21999 29894 22051 29946
rect 22063 29894 22115 29946
rect 22127 29894 22179 29946
rect 22191 29894 22243 29946
rect 30329 29894 30381 29946
rect 30393 29894 30445 29946
rect 30457 29894 30509 29946
rect 30521 29894 30573 29946
rect 30585 29894 30637 29946
rect 9036 29792 9088 29844
rect 9680 29792 9732 29844
rect 2780 29656 2832 29708
rect 4068 29563 4120 29572
rect 4068 29529 4077 29563
rect 4077 29529 4111 29563
rect 4111 29529 4120 29563
rect 4068 29520 4120 29529
rect 4988 29452 5040 29504
rect 5540 29495 5592 29504
rect 5540 29461 5549 29495
rect 5549 29461 5583 29495
rect 5583 29461 5592 29495
rect 5540 29452 5592 29461
rect 7656 29452 7708 29504
rect 9312 29724 9364 29776
rect 8576 29699 8628 29708
rect 8576 29665 8585 29699
rect 8585 29665 8619 29699
rect 8619 29665 8628 29699
rect 8576 29656 8628 29665
rect 9588 29699 9640 29708
rect 9588 29665 9597 29699
rect 9597 29665 9631 29699
rect 9631 29665 9640 29699
rect 9588 29656 9640 29665
rect 14556 29792 14608 29844
rect 18144 29835 18196 29844
rect 18144 29801 18153 29835
rect 18153 29801 18187 29835
rect 18187 29801 18196 29835
rect 18144 29792 18196 29801
rect 20996 29792 21048 29844
rect 22376 29792 22428 29844
rect 10692 29724 10744 29776
rect 11244 29656 11296 29708
rect 11704 29656 11756 29708
rect 12348 29656 12400 29708
rect 14096 29656 14148 29708
rect 9128 29520 9180 29572
rect 9220 29563 9272 29572
rect 9220 29529 9245 29563
rect 9245 29529 9272 29563
rect 9220 29520 9272 29529
rect 10600 29588 10652 29640
rect 11428 29520 11480 29572
rect 14004 29588 14056 29640
rect 13912 29520 13964 29572
rect 15476 29588 15528 29640
rect 10232 29495 10284 29504
rect 10232 29461 10241 29495
rect 10241 29461 10275 29495
rect 10275 29461 10284 29495
rect 10232 29452 10284 29461
rect 11520 29452 11572 29504
rect 12256 29452 12308 29504
rect 12992 29452 13044 29504
rect 15016 29452 15068 29504
rect 16672 29452 16724 29504
rect 17132 29452 17184 29504
rect 17408 29631 17460 29640
rect 17408 29597 17417 29631
rect 17417 29597 17451 29631
rect 17451 29597 17460 29631
rect 17408 29588 17460 29597
rect 17500 29588 17552 29640
rect 17592 29631 17644 29640
rect 17592 29597 17601 29631
rect 17601 29597 17635 29631
rect 17635 29597 17644 29631
rect 17592 29588 17644 29597
rect 19248 29656 19300 29708
rect 19892 29699 19944 29708
rect 19892 29665 19901 29699
rect 19901 29665 19935 29699
rect 19935 29665 19944 29699
rect 19892 29656 19944 29665
rect 19340 29588 19392 29640
rect 20076 29631 20128 29640
rect 20076 29597 20085 29631
rect 20085 29597 20119 29631
rect 20119 29597 20128 29631
rect 20076 29588 20128 29597
rect 18144 29520 18196 29572
rect 20812 29520 20864 29572
rect 21364 29520 21416 29572
rect 23848 29792 23900 29844
rect 23572 29656 23624 29708
rect 25872 29792 25924 29844
rect 27344 29792 27396 29844
rect 31116 29724 31168 29776
rect 24860 29656 24912 29708
rect 26056 29656 26108 29708
rect 26792 29656 26844 29708
rect 24492 29588 24544 29640
rect 25044 29588 25096 29640
rect 26056 29563 26108 29572
rect 26056 29529 26065 29563
rect 26065 29529 26099 29563
rect 26099 29529 26108 29563
rect 26056 29520 26108 29529
rect 26516 29520 26568 29572
rect 18604 29452 18656 29504
rect 20352 29452 20404 29504
rect 21180 29452 21232 29504
rect 29460 29588 29512 29640
rect 30840 29631 30892 29640
rect 30840 29597 30849 29631
rect 30849 29597 30883 29631
rect 30883 29597 30892 29631
rect 30840 29588 30892 29597
rect 29368 29452 29420 29504
rect 29552 29495 29604 29504
rect 29552 29461 29561 29495
rect 29561 29461 29595 29495
rect 29595 29461 29604 29495
rect 29552 29452 29604 29461
rect 9344 29350 9396 29402
rect 9408 29350 9460 29402
rect 9472 29350 9524 29402
rect 9536 29350 9588 29402
rect 9600 29350 9652 29402
rect 17738 29350 17790 29402
rect 17802 29350 17854 29402
rect 17866 29350 17918 29402
rect 17930 29350 17982 29402
rect 17994 29350 18046 29402
rect 26132 29350 26184 29402
rect 26196 29350 26248 29402
rect 26260 29350 26312 29402
rect 26324 29350 26376 29402
rect 26388 29350 26440 29402
rect 34526 29350 34578 29402
rect 34590 29350 34642 29402
rect 34654 29350 34706 29402
rect 34718 29350 34770 29402
rect 34782 29350 34834 29402
rect 4068 29291 4120 29300
rect 4068 29257 4077 29291
rect 4077 29257 4111 29291
rect 4111 29257 4120 29291
rect 4068 29248 4120 29257
rect 6736 29248 6788 29300
rect 3240 29112 3292 29164
rect 7656 29180 7708 29232
rect 3884 29155 3936 29164
rect 3884 29121 3893 29155
rect 3893 29121 3927 29155
rect 3927 29121 3936 29155
rect 3884 29112 3936 29121
rect 4436 29112 4488 29164
rect 5540 29112 5592 29164
rect 7012 29155 7064 29164
rect 7012 29121 7021 29155
rect 7021 29121 7055 29155
rect 7055 29121 7064 29155
rect 7012 29112 7064 29121
rect 8484 29180 8536 29232
rect 15016 29248 15068 29300
rect 8944 29180 8996 29232
rect 5632 29087 5684 29096
rect 5632 29053 5641 29087
rect 5641 29053 5675 29087
rect 5675 29053 5684 29087
rect 5632 29044 5684 29053
rect 6000 29044 6052 29096
rect 4896 28976 4948 29028
rect 8852 29112 8904 29164
rect 9680 29180 9732 29232
rect 10048 29180 10100 29232
rect 9220 29112 9272 29164
rect 4160 28908 4212 28960
rect 5724 28908 5776 28960
rect 7196 28908 7248 28960
rect 10692 29044 10744 29096
rect 11428 29180 11480 29232
rect 11244 29112 11296 29164
rect 11704 29180 11756 29232
rect 13820 29180 13872 29232
rect 15476 29291 15528 29300
rect 15476 29257 15485 29291
rect 15485 29257 15519 29291
rect 15519 29257 15528 29291
rect 15476 29248 15528 29257
rect 17408 29248 17460 29300
rect 18144 29248 18196 29300
rect 19892 29248 19944 29300
rect 26056 29248 26108 29300
rect 26516 29248 26568 29300
rect 28264 29248 28316 29300
rect 12900 29112 12952 29164
rect 14004 29112 14056 29164
rect 11520 28976 11572 29028
rect 7380 28951 7432 28960
rect 7380 28917 7389 28951
rect 7389 28917 7423 28951
rect 7423 28917 7432 28951
rect 7380 28908 7432 28917
rect 9128 28908 9180 28960
rect 12348 29044 12400 29096
rect 12992 29044 13044 29096
rect 14556 29044 14608 29096
rect 14648 29087 14700 29096
rect 14648 29053 14657 29087
rect 14657 29053 14691 29087
rect 14691 29053 14700 29087
rect 14648 29044 14700 29053
rect 14372 28976 14424 29028
rect 16948 29112 17000 29164
rect 17500 29044 17552 29096
rect 17776 29044 17828 29096
rect 16580 28976 16632 29028
rect 17040 28976 17092 29028
rect 18512 29112 18564 29164
rect 18604 29155 18656 29164
rect 18604 29121 18613 29155
rect 18613 29121 18647 29155
rect 18647 29121 18656 29155
rect 18604 29112 18656 29121
rect 18788 29112 18840 29164
rect 19708 29180 19760 29232
rect 23112 29223 23164 29232
rect 20444 29112 20496 29164
rect 19524 29087 19576 29096
rect 19524 29053 19533 29087
rect 19533 29053 19567 29087
rect 19567 29053 19576 29087
rect 19524 29044 19576 29053
rect 19616 29087 19668 29096
rect 19616 29053 19625 29087
rect 19625 29053 19659 29087
rect 19659 29053 19668 29087
rect 19616 29044 19668 29053
rect 19708 29087 19760 29096
rect 19708 29053 19717 29087
rect 19717 29053 19751 29087
rect 19751 29053 19760 29087
rect 19708 29044 19760 29053
rect 20352 29044 20404 29096
rect 20076 28976 20128 29028
rect 14280 28908 14332 28960
rect 18880 28908 18932 28960
rect 20996 29112 21048 29164
rect 21180 29112 21232 29164
rect 20720 29087 20772 29096
rect 20720 29053 20729 29087
rect 20729 29053 20763 29087
rect 20763 29053 20772 29087
rect 20720 29044 20772 29053
rect 21088 28976 21140 29028
rect 23112 29189 23121 29223
rect 23121 29189 23155 29223
rect 23155 29189 23164 29223
rect 23112 29180 23164 29189
rect 23572 29112 23624 29164
rect 23388 29044 23440 29096
rect 24492 29155 24544 29164
rect 24492 29121 24501 29155
rect 24501 29121 24535 29155
rect 24535 29121 24544 29155
rect 24492 29112 24544 29121
rect 24676 29155 24728 29164
rect 24676 29121 24685 29155
rect 24685 29121 24719 29155
rect 24719 29121 24728 29155
rect 24676 29112 24728 29121
rect 24768 29112 24820 29164
rect 29184 29180 29236 29232
rect 26792 29112 26844 29164
rect 29460 29180 29512 29232
rect 31116 29223 31168 29232
rect 31116 29189 31125 29223
rect 31125 29189 31159 29223
rect 31159 29189 31168 29223
rect 31116 29180 31168 29189
rect 27160 28976 27212 29028
rect 29552 29112 29604 29164
rect 29368 28976 29420 29028
rect 22284 28951 22336 28960
rect 22284 28917 22293 28951
rect 22293 28917 22327 28951
rect 22327 28917 22336 28951
rect 22284 28908 22336 28917
rect 29184 28908 29236 28960
rect 29644 28951 29696 28960
rect 29644 28917 29653 28951
rect 29653 28917 29687 28951
rect 29687 28917 29696 28951
rect 29644 28908 29696 28917
rect 5147 28806 5199 28858
rect 5211 28806 5263 28858
rect 5275 28806 5327 28858
rect 5339 28806 5391 28858
rect 5403 28806 5455 28858
rect 13541 28806 13593 28858
rect 13605 28806 13657 28858
rect 13669 28806 13721 28858
rect 13733 28806 13785 28858
rect 13797 28806 13849 28858
rect 21935 28806 21987 28858
rect 21999 28806 22051 28858
rect 22063 28806 22115 28858
rect 22127 28806 22179 28858
rect 22191 28806 22243 28858
rect 30329 28806 30381 28858
rect 30393 28806 30445 28858
rect 30457 28806 30509 28858
rect 30521 28806 30573 28858
rect 30585 28806 30637 28858
rect 3884 28704 3936 28756
rect 3608 28611 3660 28620
rect 3608 28577 3617 28611
rect 3617 28577 3651 28611
rect 3651 28577 3660 28611
rect 3608 28568 3660 28577
rect 3240 28500 3292 28552
rect 3976 28543 4028 28552
rect 3976 28509 3985 28543
rect 3985 28509 4019 28543
rect 4019 28509 4028 28543
rect 3976 28500 4028 28509
rect 4344 28500 4396 28552
rect 3700 28432 3752 28484
rect 4436 28475 4488 28484
rect 4436 28441 4445 28475
rect 4445 28441 4479 28475
rect 4479 28441 4488 28475
rect 4436 28432 4488 28441
rect 5816 28704 5868 28756
rect 7288 28747 7340 28756
rect 7288 28713 7297 28747
rect 7297 28713 7331 28747
rect 7331 28713 7340 28747
rect 7288 28704 7340 28713
rect 10692 28747 10744 28756
rect 10692 28713 10701 28747
rect 10701 28713 10735 28747
rect 10735 28713 10744 28747
rect 10692 28704 10744 28713
rect 15752 28704 15804 28756
rect 16580 28704 16632 28756
rect 4896 28636 4948 28688
rect 5540 28568 5592 28620
rect 7196 28636 7248 28688
rect 17960 28704 18012 28756
rect 18880 28704 18932 28756
rect 19524 28704 19576 28756
rect 19616 28704 19668 28756
rect 20720 28704 20772 28756
rect 20996 28747 21048 28756
rect 20996 28713 21005 28747
rect 21005 28713 21039 28747
rect 21039 28713 21048 28747
rect 20996 28704 21048 28713
rect 21824 28704 21876 28756
rect 23112 28704 23164 28756
rect 28448 28704 28500 28756
rect 28540 28704 28592 28756
rect 4896 28543 4948 28552
rect 4896 28509 4905 28543
rect 4905 28509 4939 28543
rect 4939 28509 4948 28543
rect 4896 28500 4948 28509
rect 5632 28500 5684 28552
rect 5724 28543 5776 28552
rect 5724 28509 5733 28543
rect 5733 28509 5767 28543
rect 5767 28509 5776 28543
rect 5724 28500 5776 28509
rect 6000 28543 6052 28552
rect 6000 28509 6009 28543
rect 6009 28509 6043 28543
rect 6043 28509 6052 28543
rect 6000 28500 6052 28509
rect 6460 28500 6512 28552
rect 16948 28636 17000 28688
rect 8944 28611 8996 28620
rect 8944 28577 8953 28611
rect 8953 28577 8987 28611
rect 8987 28577 8996 28611
rect 8944 28568 8996 28577
rect 11336 28568 11388 28620
rect 14096 28611 14148 28620
rect 14096 28577 14105 28611
rect 14105 28577 14139 28611
rect 14139 28577 14148 28611
rect 14096 28568 14148 28577
rect 18604 28611 18656 28620
rect 18604 28577 18613 28611
rect 18613 28577 18647 28611
rect 18647 28577 18656 28611
rect 18604 28568 18656 28577
rect 18512 28543 18564 28552
rect 18512 28509 18521 28543
rect 18521 28509 18555 28543
rect 18555 28509 18564 28543
rect 18512 28500 18564 28509
rect 18788 28543 18840 28552
rect 18788 28509 18797 28543
rect 18797 28509 18831 28543
rect 18831 28509 18840 28543
rect 18788 28500 18840 28509
rect 18880 28500 18932 28552
rect 19340 28543 19392 28552
rect 19340 28509 19349 28543
rect 19349 28509 19383 28543
rect 19383 28509 19392 28543
rect 19340 28500 19392 28509
rect 2504 28364 2556 28416
rect 3240 28407 3292 28416
rect 3240 28373 3249 28407
rect 3249 28373 3283 28407
rect 3283 28373 3292 28407
rect 3240 28364 3292 28373
rect 5448 28407 5500 28416
rect 5448 28373 5457 28407
rect 5457 28373 5491 28407
rect 5491 28373 5500 28407
rect 5448 28364 5500 28373
rect 7380 28432 7432 28484
rect 7656 28475 7708 28484
rect 7656 28441 7665 28475
rect 7665 28441 7699 28475
rect 7699 28441 7708 28475
rect 7656 28432 7708 28441
rect 8852 28432 8904 28484
rect 9128 28432 9180 28484
rect 9772 28432 9824 28484
rect 14280 28432 14332 28484
rect 16580 28432 16632 28484
rect 17040 28475 17092 28484
rect 17040 28441 17049 28475
rect 17049 28441 17083 28475
rect 17083 28441 17092 28475
rect 17040 28432 17092 28441
rect 8576 28407 8628 28416
rect 8576 28373 8585 28407
rect 8585 28373 8619 28407
rect 8619 28373 8628 28407
rect 8576 28364 8628 28373
rect 13176 28364 13228 28416
rect 17500 28364 17552 28416
rect 20076 28432 20128 28484
rect 20444 28543 20496 28552
rect 20444 28509 20453 28543
rect 20453 28509 20487 28543
rect 20487 28509 20496 28543
rect 20444 28500 20496 28509
rect 20812 28500 20864 28552
rect 23572 28543 23624 28552
rect 23572 28509 23581 28543
rect 23581 28509 23615 28543
rect 23615 28509 23624 28543
rect 23572 28500 23624 28509
rect 24492 28568 24544 28620
rect 24676 28500 24728 28552
rect 25136 28500 25188 28552
rect 28816 28636 28868 28688
rect 29368 28747 29420 28756
rect 29368 28713 29377 28747
rect 29377 28713 29411 28747
rect 29411 28713 29420 28747
rect 29368 28704 29420 28713
rect 30840 28704 30892 28756
rect 28954 28568 29006 28620
rect 29552 28568 29604 28620
rect 29644 28611 29696 28620
rect 29644 28577 29653 28611
rect 29653 28577 29687 28611
rect 29687 28577 29696 28611
rect 29644 28568 29696 28577
rect 26700 28543 26752 28552
rect 26700 28509 26709 28543
rect 26709 28509 26743 28543
rect 26743 28509 26752 28543
rect 26700 28500 26752 28509
rect 27712 28500 27764 28552
rect 28632 28543 28684 28552
rect 28632 28509 28642 28543
rect 28642 28509 28676 28543
rect 28676 28509 28684 28543
rect 28632 28500 28684 28509
rect 30564 28543 30616 28552
rect 22284 28432 22336 28484
rect 23296 28432 23348 28484
rect 23848 28475 23900 28484
rect 23848 28441 23857 28475
rect 23857 28441 23891 28475
rect 23891 28441 23900 28475
rect 23848 28432 23900 28441
rect 25780 28432 25832 28484
rect 24308 28364 24360 28416
rect 26976 28364 27028 28416
rect 28356 28364 28408 28416
rect 30564 28509 30573 28543
rect 30573 28509 30607 28543
rect 30607 28509 30616 28543
rect 30564 28500 30616 28509
rect 28954 28432 29006 28484
rect 29092 28364 29144 28416
rect 30656 28364 30708 28416
rect 9344 28262 9396 28314
rect 9408 28262 9460 28314
rect 9472 28262 9524 28314
rect 9536 28262 9588 28314
rect 9600 28262 9652 28314
rect 17738 28262 17790 28314
rect 17802 28262 17854 28314
rect 17866 28262 17918 28314
rect 17930 28262 17982 28314
rect 17994 28262 18046 28314
rect 26132 28262 26184 28314
rect 26196 28262 26248 28314
rect 26260 28262 26312 28314
rect 26324 28262 26376 28314
rect 26388 28262 26440 28314
rect 34526 28262 34578 28314
rect 34590 28262 34642 28314
rect 34654 28262 34706 28314
rect 34718 28262 34770 28314
rect 34782 28262 34834 28314
rect 2504 28160 2556 28212
rect 3608 28160 3660 28212
rect 3700 28160 3752 28212
rect 5448 28160 5500 28212
rect 7012 28160 7064 28212
rect 7656 28160 7708 28212
rect 4160 28024 4212 28076
rect 8576 28135 8628 28144
rect 8576 28101 8585 28135
rect 8585 28101 8619 28135
rect 8619 28101 8628 28135
rect 8576 28092 8628 28101
rect 5816 28024 5868 28076
rect 5908 28024 5960 28076
rect 12348 28160 12400 28212
rect 21824 28160 21876 28212
rect 9772 28092 9824 28144
rect 3976 27956 4028 28008
rect 6184 27956 6236 28008
rect 11980 28024 12032 28076
rect 12348 28067 12400 28076
rect 12348 28033 12357 28067
rect 12357 28033 12391 28067
rect 12391 28033 12400 28067
rect 12348 28024 12400 28033
rect 11244 27956 11296 28008
rect 12164 27956 12216 28008
rect 13452 28092 13504 28144
rect 17040 28092 17092 28144
rect 20076 28092 20128 28144
rect 22376 28092 22428 28144
rect 23388 28092 23440 28144
rect 26976 28160 27028 28212
rect 27712 28203 27764 28212
rect 27712 28169 27721 28203
rect 27721 28169 27755 28203
rect 27755 28169 27764 28203
rect 27712 28160 27764 28169
rect 30564 28160 30616 28212
rect 3240 27820 3292 27872
rect 4344 27888 4396 27940
rect 18972 27888 19024 27940
rect 23480 27999 23532 28008
rect 23480 27965 23489 27999
rect 23489 27965 23523 27999
rect 23523 27965 23532 27999
rect 23480 27956 23532 27965
rect 25596 28067 25648 28076
rect 25596 28033 25605 28067
rect 25605 28033 25639 28067
rect 25639 28033 25648 28067
rect 25596 28024 25648 28033
rect 26792 28024 26844 28076
rect 30748 28092 30800 28144
rect 24952 27956 25004 28008
rect 25780 27956 25832 28008
rect 27896 27956 27948 28008
rect 28356 27956 28408 28008
rect 32588 28160 32640 28212
rect 23572 27888 23624 27940
rect 34796 27956 34848 28008
rect 4988 27820 5040 27872
rect 5540 27820 5592 27872
rect 12532 27863 12584 27872
rect 12532 27829 12541 27863
rect 12541 27829 12575 27863
rect 12575 27829 12584 27863
rect 12532 27820 12584 27829
rect 22284 27820 22336 27872
rect 25136 27820 25188 27872
rect 30932 27888 30984 27940
rect 27620 27863 27672 27872
rect 27620 27829 27629 27863
rect 27629 27829 27663 27863
rect 27663 27829 27672 27863
rect 27620 27820 27672 27829
rect 5147 27718 5199 27770
rect 5211 27718 5263 27770
rect 5275 27718 5327 27770
rect 5339 27718 5391 27770
rect 5403 27718 5455 27770
rect 13541 27718 13593 27770
rect 13605 27718 13657 27770
rect 13669 27718 13721 27770
rect 13733 27718 13785 27770
rect 13797 27718 13849 27770
rect 21935 27718 21987 27770
rect 21999 27718 22051 27770
rect 22063 27718 22115 27770
rect 22127 27718 22179 27770
rect 22191 27718 22243 27770
rect 30329 27718 30381 27770
rect 30393 27718 30445 27770
rect 30457 27718 30509 27770
rect 30521 27718 30573 27770
rect 30585 27718 30637 27770
rect 5540 27616 5592 27668
rect 22376 27616 22428 27668
rect 23848 27616 23900 27668
rect 27620 27659 27672 27668
rect 27620 27625 27641 27659
rect 27641 27625 27672 27659
rect 27620 27616 27672 27625
rect 30748 27659 30800 27668
rect 30748 27625 30757 27659
rect 30757 27625 30791 27659
rect 30791 27625 30800 27659
rect 30748 27616 30800 27625
rect 30932 27616 30984 27668
rect 6460 27548 6512 27600
rect 16028 27591 16080 27600
rect 16028 27557 16037 27591
rect 16037 27557 16071 27591
rect 16071 27557 16080 27591
rect 16028 27548 16080 27557
rect 14648 27480 14700 27532
rect 3240 27412 3292 27464
rect 10324 27455 10376 27464
rect 10324 27421 10333 27455
rect 10333 27421 10367 27455
rect 10367 27421 10376 27455
rect 10324 27412 10376 27421
rect 11244 27455 11296 27464
rect 11244 27421 11253 27455
rect 11253 27421 11287 27455
rect 11287 27421 11296 27455
rect 11244 27412 11296 27421
rect 11980 27412 12032 27464
rect 13912 27412 13964 27464
rect 14096 27412 14148 27464
rect 15384 27455 15436 27464
rect 15384 27421 15393 27455
rect 15393 27421 15427 27455
rect 15427 27421 15436 27455
rect 15384 27412 15436 27421
rect 15844 27455 15896 27464
rect 15844 27421 15853 27455
rect 15853 27421 15887 27455
rect 15887 27421 15896 27455
rect 15844 27412 15896 27421
rect 16856 27412 16908 27464
rect 17500 27412 17552 27464
rect 23480 27480 23532 27532
rect 26884 27480 26936 27532
rect 28080 27480 28132 27532
rect 4988 27344 5040 27396
rect 5908 27344 5960 27396
rect 12900 27344 12952 27396
rect 13360 27387 13412 27396
rect 13360 27353 13369 27387
rect 13369 27353 13403 27387
rect 13403 27353 13412 27387
rect 13360 27344 13412 27353
rect 16672 27344 16724 27396
rect 18880 27412 18932 27464
rect 19064 27412 19116 27464
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 22928 27412 22980 27464
rect 20812 27387 20864 27396
rect 20812 27353 20821 27387
rect 20821 27353 20855 27387
rect 20855 27353 20864 27387
rect 20812 27344 20864 27353
rect 23296 27344 23348 27396
rect 25872 27387 25924 27396
rect 25872 27353 25881 27387
rect 25881 27353 25915 27387
rect 25915 27353 25924 27387
rect 25872 27344 25924 27353
rect 27160 27344 27212 27396
rect 27528 27344 27580 27396
rect 27712 27344 27764 27396
rect 28908 27548 28960 27600
rect 28264 27480 28316 27532
rect 33600 27480 33652 27532
rect 28172 27455 28224 27464
rect 28172 27421 28181 27455
rect 28181 27421 28215 27455
rect 28215 27421 28224 27455
rect 28172 27412 28224 27421
rect 32956 27412 33008 27464
rect 29092 27344 29144 27396
rect 30656 27344 30708 27396
rect 31760 27344 31812 27396
rect 32772 27344 32824 27396
rect 10140 27319 10192 27328
rect 10140 27285 10149 27319
rect 10149 27285 10183 27319
rect 10183 27285 10192 27319
rect 10140 27276 10192 27285
rect 11060 27319 11112 27328
rect 11060 27285 11069 27319
rect 11069 27285 11103 27319
rect 11103 27285 11112 27319
rect 11060 27276 11112 27285
rect 11888 27319 11940 27328
rect 11888 27285 11897 27319
rect 11897 27285 11931 27319
rect 11931 27285 11940 27319
rect 11888 27276 11940 27285
rect 14280 27319 14332 27328
rect 14280 27285 14289 27319
rect 14289 27285 14323 27319
rect 14323 27285 14332 27319
rect 14280 27276 14332 27285
rect 17040 27276 17092 27328
rect 17592 27276 17644 27328
rect 19248 27319 19300 27328
rect 19248 27285 19257 27319
rect 19257 27285 19291 27319
rect 19291 27285 19300 27319
rect 19248 27276 19300 27285
rect 28448 27276 28500 27328
rect 32588 27319 32640 27328
rect 32588 27285 32597 27319
rect 32597 27285 32631 27319
rect 32631 27285 32640 27319
rect 32588 27276 32640 27285
rect 9344 27174 9396 27226
rect 9408 27174 9460 27226
rect 9472 27174 9524 27226
rect 9536 27174 9588 27226
rect 9600 27174 9652 27226
rect 17738 27174 17790 27226
rect 17802 27174 17854 27226
rect 17866 27174 17918 27226
rect 17930 27174 17982 27226
rect 17994 27174 18046 27226
rect 26132 27174 26184 27226
rect 26196 27174 26248 27226
rect 26260 27174 26312 27226
rect 26324 27174 26376 27226
rect 26388 27174 26440 27226
rect 34526 27174 34578 27226
rect 34590 27174 34642 27226
rect 34654 27174 34706 27226
rect 34718 27174 34770 27226
rect 34782 27174 34834 27226
rect 10140 27072 10192 27124
rect 11244 27072 11296 27124
rect 12348 27072 12400 27124
rect 13360 27072 13412 27124
rect 11888 27047 11940 27056
rect 11888 27013 11897 27047
rect 11897 27013 11931 27047
rect 11931 27013 11940 27047
rect 14280 27072 14332 27124
rect 16028 27072 16080 27124
rect 16672 27115 16724 27124
rect 16672 27081 16681 27115
rect 16681 27081 16715 27115
rect 16715 27081 16724 27115
rect 16672 27072 16724 27081
rect 16856 27072 16908 27124
rect 16948 27072 17000 27124
rect 11888 27004 11940 27013
rect 15384 27004 15436 27056
rect 7012 26911 7064 26920
rect 7012 26877 7021 26911
rect 7021 26877 7055 26911
rect 7055 26877 7064 26911
rect 7012 26868 7064 26877
rect 7656 26868 7708 26920
rect 9220 26868 9272 26920
rect 10876 26868 10928 26920
rect 17592 27072 17644 27124
rect 18880 27115 18932 27124
rect 18880 27081 18889 27115
rect 18889 27081 18923 27115
rect 18923 27081 18932 27115
rect 18880 27072 18932 27081
rect 19248 27072 19300 27124
rect 18972 27004 19024 27056
rect 20812 27072 20864 27124
rect 20076 27004 20128 27056
rect 22928 27072 22980 27124
rect 23480 27072 23532 27124
rect 25872 27072 25924 27124
rect 26700 27072 26752 27124
rect 12900 26868 12952 26920
rect 13084 26911 13136 26920
rect 13084 26877 13093 26911
rect 13093 26877 13127 26911
rect 13127 26877 13136 26911
rect 13084 26868 13136 26877
rect 7288 26843 7340 26852
rect 7288 26809 7297 26843
rect 7297 26809 7331 26843
rect 7331 26809 7340 26843
rect 7288 26800 7340 26809
rect 14464 26868 14516 26920
rect 16212 26868 16264 26920
rect 16764 26868 16816 26920
rect 19064 26911 19116 26920
rect 19064 26877 19073 26911
rect 19073 26877 19107 26911
rect 19107 26877 19116 26911
rect 19064 26868 19116 26877
rect 22284 26936 22336 26988
rect 25228 26979 25280 26988
rect 25228 26945 25237 26979
rect 25237 26945 25271 26979
rect 25271 26945 25280 26979
rect 25228 26936 25280 26945
rect 25320 26979 25372 26988
rect 25320 26945 25329 26979
rect 25329 26945 25363 26979
rect 25363 26945 25372 26979
rect 25320 26936 25372 26945
rect 25596 26936 25648 26988
rect 23848 26868 23900 26920
rect 24860 26911 24912 26920
rect 24860 26877 24869 26911
rect 24869 26877 24903 26911
rect 24903 26877 24912 26911
rect 24860 26868 24912 26877
rect 27344 26979 27396 26988
rect 27344 26945 27353 26979
rect 27353 26945 27387 26979
rect 27387 26945 27396 26979
rect 27344 26936 27396 26945
rect 27896 27004 27948 27056
rect 29184 27072 29236 27124
rect 31760 27004 31812 27056
rect 26516 26868 26568 26920
rect 27252 26868 27304 26920
rect 27988 26936 28040 26988
rect 28264 26979 28316 26988
rect 28264 26945 28273 26979
rect 28273 26945 28307 26979
rect 28307 26945 28316 26979
rect 28264 26936 28316 26945
rect 30656 26936 30708 26988
rect 32496 26936 32548 26988
rect 28540 26911 28592 26920
rect 28540 26877 28549 26911
rect 28549 26877 28583 26911
rect 28583 26877 28592 26911
rect 28540 26868 28592 26877
rect 28632 26868 28684 26920
rect 25688 26800 25740 26852
rect 27160 26800 27212 26852
rect 7472 26775 7524 26784
rect 7472 26741 7481 26775
rect 7481 26741 7515 26775
rect 7515 26741 7524 26775
rect 7472 26732 7524 26741
rect 11520 26775 11572 26784
rect 11520 26741 11529 26775
rect 11529 26741 11563 26775
rect 11563 26741 11572 26775
rect 11520 26732 11572 26741
rect 11980 26732 12032 26784
rect 13912 26732 13964 26784
rect 14832 26732 14884 26784
rect 16488 26775 16540 26784
rect 16488 26741 16497 26775
rect 16497 26741 16531 26775
rect 16531 26741 16540 26775
rect 16488 26732 16540 26741
rect 20904 26775 20956 26784
rect 20904 26741 20913 26775
rect 20913 26741 20947 26775
rect 20947 26741 20956 26775
rect 20904 26732 20956 26741
rect 23296 26732 23348 26784
rect 28080 26732 28132 26784
rect 29920 26732 29972 26784
rect 31576 26732 31628 26784
rect 5147 26630 5199 26682
rect 5211 26630 5263 26682
rect 5275 26630 5327 26682
rect 5339 26630 5391 26682
rect 5403 26630 5455 26682
rect 13541 26630 13593 26682
rect 13605 26630 13657 26682
rect 13669 26630 13721 26682
rect 13733 26630 13785 26682
rect 13797 26630 13849 26682
rect 21935 26630 21987 26682
rect 21999 26630 22051 26682
rect 22063 26630 22115 26682
rect 22127 26630 22179 26682
rect 22191 26630 22243 26682
rect 30329 26630 30381 26682
rect 30393 26630 30445 26682
rect 30457 26630 30509 26682
rect 30521 26630 30573 26682
rect 30585 26630 30637 26682
rect 7288 26528 7340 26580
rect 9956 26528 10008 26580
rect 10324 26571 10376 26580
rect 10324 26537 10333 26571
rect 10333 26537 10367 26571
rect 10367 26537 10376 26571
rect 10324 26528 10376 26537
rect 12256 26571 12308 26580
rect 12256 26537 12265 26571
rect 12265 26537 12299 26571
rect 12299 26537 12308 26571
rect 12256 26528 12308 26537
rect 13084 26528 13136 26580
rect 14096 26571 14148 26580
rect 14096 26537 14105 26571
rect 14105 26537 14139 26571
rect 14139 26537 14148 26571
rect 14096 26528 14148 26537
rect 14372 26528 14424 26580
rect 16488 26528 16540 26580
rect 17500 26528 17552 26580
rect 19432 26528 19484 26580
rect 11520 26460 11572 26512
rect 3240 26392 3292 26444
rect 7656 26392 7708 26444
rect 11060 26392 11112 26444
rect 12348 26392 12400 26444
rect 3424 26367 3476 26376
rect 3424 26333 3433 26367
rect 3433 26333 3467 26367
rect 3467 26333 3476 26367
rect 3424 26324 3476 26333
rect 5080 26324 5132 26376
rect 5632 26324 5684 26376
rect 1400 26299 1452 26308
rect 1400 26265 1409 26299
rect 1409 26265 1443 26299
rect 1443 26265 1452 26299
rect 1400 26256 1452 26265
rect 1860 26256 1912 26308
rect 9772 26324 9824 26376
rect 7196 26299 7248 26308
rect 7196 26265 7205 26299
rect 7205 26265 7239 26299
rect 7239 26265 7248 26299
rect 7196 26256 7248 26265
rect 16764 26392 16816 26444
rect 19064 26392 19116 26444
rect 19984 26435 20036 26444
rect 19984 26401 19993 26435
rect 19993 26401 20027 26435
rect 20027 26401 20036 26435
rect 19984 26392 20036 26401
rect 20904 26392 20956 26444
rect 25228 26528 25280 26580
rect 27896 26528 27948 26580
rect 28540 26528 28592 26580
rect 28908 26460 28960 26512
rect 33600 26528 33652 26580
rect 12532 26324 12584 26376
rect 13912 26324 13964 26376
rect 14556 26324 14608 26376
rect 14832 26324 14884 26376
rect 20996 26367 21048 26376
rect 20996 26333 21005 26367
rect 21005 26333 21039 26367
rect 21039 26333 21048 26367
rect 20996 26324 21048 26333
rect 25044 26367 25096 26376
rect 25044 26333 25053 26367
rect 25053 26333 25087 26367
rect 25087 26333 25096 26367
rect 25044 26324 25096 26333
rect 5540 26231 5592 26240
rect 5540 26197 5549 26231
rect 5549 26197 5583 26231
rect 5583 26197 5592 26231
rect 5540 26188 5592 26197
rect 5908 26188 5960 26240
rect 8668 26231 8720 26240
rect 8668 26197 8677 26231
rect 8677 26197 8711 26231
rect 8711 26197 8720 26231
rect 8668 26188 8720 26197
rect 14740 26299 14792 26308
rect 14740 26265 14749 26299
rect 14749 26265 14783 26299
rect 14783 26265 14792 26299
rect 14740 26256 14792 26265
rect 16580 26256 16632 26308
rect 20720 26256 20772 26308
rect 23296 26256 23348 26308
rect 23572 26256 23624 26308
rect 28080 26324 28132 26376
rect 28448 26367 28500 26376
rect 28448 26333 28457 26367
rect 28457 26333 28491 26367
rect 28491 26333 28500 26367
rect 28448 26324 28500 26333
rect 28540 26367 28592 26376
rect 28540 26333 28549 26367
rect 28549 26333 28583 26367
rect 28583 26333 28592 26367
rect 28540 26324 28592 26333
rect 25504 26299 25556 26308
rect 25504 26265 25513 26299
rect 25513 26265 25547 26299
rect 25547 26265 25556 26299
rect 25504 26256 25556 26265
rect 27988 26256 28040 26308
rect 28632 26256 28684 26308
rect 23112 26231 23164 26240
rect 23112 26197 23121 26231
rect 23121 26197 23155 26231
rect 23155 26197 23164 26231
rect 23112 26188 23164 26197
rect 25412 26188 25464 26240
rect 29092 26324 29144 26376
rect 29828 26324 29880 26376
rect 31576 26367 31628 26376
rect 31576 26333 31585 26367
rect 31585 26333 31619 26367
rect 31619 26333 31628 26367
rect 31576 26324 31628 26333
rect 31392 26299 31444 26308
rect 31392 26265 31401 26299
rect 31401 26265 31435 26299
rect 31435 26265 31444 26299
rect 31392 26256 31444 26265
rect 32864 26256 32916 26308
rect 33048 26256 33100 26308
rect 30472 26231 30524 26240
rect 30472 26197 30481 26231
rect 30481 26197 30515 26231
rect 30515 26197 30524 26231
rect 30472 26188 30524 26197
rect 32312 26188 32364 26240
rect 9344 26086 9396 26138
rect 9408 26086 9460 26138
rect 9472 26086 9524 26138
rect 9536 26086 9588 26138
rect 9600 26086 9652 26138
rect 17738 26086 17790 26138
rect 17802 26086 17854 26138
rect 17866 26086 17918 26138
rect 17930 26086 17982 26138
rect 17994 26086 18046 26138
rect 26132 26086 26184 26138
rect 26196 26086 26248 26138
rect 26260 26086 26312 26138
rect 26324 26086 26376 26138
rect 26388 26086 26440 26138
rect 34526 26086 34578 26138
rect 34590 26086 34642 26138
rect 34654 26086 34706 26138
rect 34718 26086 34770 26138
rect 34782 26086 34834 26138
rect 3424 25984 3476 26036
rect 3976 26027 4028 26036
rect 3976 25993 3985 26027
rect 3985 25993 4019 26027
rect 4019 25993 4028 26027
rect 3976 25984 4028 25993
rect 7196 25984 7248 26036
rect 7472 25984 7524 26036
rect 20996 25984 21048 26036
rect 23112 25984 23164 26036
rect 4160 25848 4212 25900
rect 5540 25916 5592 25968
rect 6920 25916 6972 25968
rect 4712 25823 4764 25832
rect 4712 25789 4721 25823
rect 4721 25789 4755 25823
rect 4755 25789 4764 25823
rect 4712 25780 4764 25789
rect 5724 25848 5776 25900
rect 12072 25916 12124 25968
rect 23296 25916 23348 25968
rect 23664 25916 23716 25968
rect 25504 25984 25556 26036
rect 30472 25984 30524 26036
rect 33048 25984 33100 26036
rect 29000 25916 29052 25968
rect 4988 25712 5040 25764
rect 6920 25780 6972 25832
rect 14740 25848 14792 25900
rect 14832 25848 14884 25900
rect 19984 25848 20036 25900
rect 20996 25848 21048 25900
rect 21640 25780 21692 25832
rect 23112 25891 23164 25900
rect 23112 25857 23121 25891
rect 23121 25857 23155 25891
rect 23155 25857 23164 25891
rect 23112 25848 23164 25857
rect 24676 25848 24728 25900
rect 22928 25780 22980 25832
rect 12532 25712 12584 25764
rect 12716 25755 12768 25764
rect 12716 25721 12725 25755
rect 12725 25721 12759 25755
rect 12759 25721 12768 25755
rect 12716 25712 12768 25721
rect 25044 25823 25096 25832
rect 25044 25789 25053 25823
rect 25053 25789 25087 25823
rect 25087 25789 25096 25823
rect 25044 25780 25096 25789
rect 25596 25891 25648 25900
rect 25596 25857 25605 25891
rect 25605 25857 25639 25891
rect 25639 25857 25648 25891
rect 25596 25848 25648 25857
rect 26516 25848 26568 25900
rect 26608 25891 26660 25900
rect 26608 25857 26617 25891
rect 26617 25857 26651 25891
rect 26651 25857 26660 25891
rect 26608 25848 26660 25857
rect 27160 25848 27212 25900
rect 27252 25891 27304 25900
rect 27252 25857 27261 25891
rect 27261 25857 27295 25891
rect 27295 25857 27304 25891
rect 27252 25848 27304 25857
rect 28172 25848 28224 25900
rect 30012 25891 30064 25900
rect 30012 25857 30021 25891
rect 30021 25857 30055 25891
rect 30055 25857 30064 25891
rect 30012 25848 30064 25857
rect 32312 25891 32364 25900
rect 32312 25857 32321 25891
rect 32321 25857 32355 25891
rect 32355 25857 32364 25891
rect 32312 25848 32364 25857
rect 32496 25891 32548 25900
rect 32496 25857 32505 25891
rect 32505 25857 32539 25891
rect 32539 25857 32548 25891
rect 32496 25848 32548 25857
rect 32588 25891 32640 25900
rect 32588 25857 32597 25891
rect 32597 25857 32631 25891
rect 32631 25857 32640 25891
rect 32588 25848 32640 25857
rect 25688 25712 25740 25764
rect 27160 25712 27212 25764
rect 30656 25780 30708 25832
rect 5816 25687 5868 25696
rect 5816 25653 5825 25687
rect 5825 25653 5859 25687
rect 5859 25653 5868 25687
rect 5816 25644 5868 25653
rect 5908 25644 5960 25696
rect 7012 25644 7064 25696
rect 7196 25644 7248 25696
rect 7840 25644 7892 25696
rect 9128 25644 9180 25696
rect 9956 25644 10008 25696
rect 14556 25687 14608 25696
rect 14556 25653 14565 25687
rect 14565 25653 14599 25687
rect 14599 25653 14608 25687
rect 14556 25644 14608 25653
rect 24860 25687 24912 25696
rect 24860 25653 24869 25687
rect 24869 25653 24903 25687
rect 24903 25653 24912 25687
rect 24860 25644 24912 25653
rect 25320 25644 25372 25696
rect 28448 25644 28500 25696
rect 5147 25542 5199 25594
rect 5211 25542 5263 25594
rect 5275 25542 5327 25594
rect 5339 25542 5391 25594
rect 5403 25542 5455 25594
rect 13541 25542 13593 25594
rect 13605 25542 13657 25594
rect 13669 25542 13721 25594
rect 13733 25542 13785 25594
rect 13797 25542 13849 25594
rect 21935 25542 21987 25594
rect 21999 25542 22051 25594
rect 22063 25542 22115 25594
rect 22127 25542 22179 25594
rect 22191 25542 22243 25594
rect 30329 25542 30381 25594
rect 30393 25542 30445 25594
rect 30457 25542 30509 25594
rect 30521 25542 30573 25594
rect 30585 25542 30637 25594
rect 4160 25440 4212 25492
rect 5540 25440 5592 25492
rect 7196 25483 7248 25492
rect 7196 25449 7205 25483
rect 7205 25449 7239 25483
rect 7239 25449 7248 25483
rect 7196 25440 7248 25449
rect 4436 25347 4488 25356
rect 4436 25313 4445 25347
rect 4445 25313 4479 25347
rect 4479 25313 4488 25347
rect 4436 25304 4488 25313
rect 3332 25236 3384 25288
rect 3424 25279 3476 25288
rect 3424 25245 3433 25279
rect 3433 25245 3467 25279
rect 3467 25245 3476 25279
rect 3424 25236 3476 25245
rect 5816 25304 5868 25356
rect 7196 25304 7248 25356
rect 7840 25483 7892 25492
rect 7840 25449 7849 25483
rect 7849 25449 7883 25483
rect 7883 25449 7892 25483
rect 7840 25440 7892 25449
rect 8668 25440 8720 25492
rect 9220 25440 9272 25492
rect 20720 25440 20772 25492
rect 26516 25440 26568 25492
rect 28816 25483 28868 25492
rect 28816 25449 28825 25483
rect 28825 25449 28859 25483
rect 28859 25449 28868 25483
rect 28816 25440 28868 25449
rect 4988 25211 5040 25220
rect 4988 25177 4997 25211
rect 4997 25177 5031 25211
rect 5031 25177 5040 25211
rect 4988 25168 5040 25177
rect 7748 25236 7800 25288
rect 2872 25100 2924 25152
rect 4804 25143 4856 25152
rect 4804 25109 4831 25143
rect 4831 25109 4856 25143
rect 4804 25100 4856 25109
rect 6460 25143 6512 25152
rect 6460 25109 6469 25143
rect 6469 25109 6503 25143
rect 6503 25109 6512 25143
rect 6460 25100 6512 25109
rect 6920 25100 6972 25152
rect 7012 25143 7064 25152
rect 7012 25109 7021 25143
rect 7021 25109 7055 25143
rect 7055 25109 7064 25143
rect 7012 25100 7064 25109
rect 7196 25143 7248 25152
rect 7196 25109 7223 25143
rect 7223 25109 7248 25143
rect 7196 25100 7248 25109
rect 9036 25100 9088 25152
rect 10876 25236 10928 25288
rect 11336 25236 11388 25288
rect 11704 25279 11756 25288
rect 11704 25245 11713 25279
rect 11713 25245 11747 25279
rect 11747 25245 11756 25279
rect 11704 25236 11756 25245
rect 9864 25168 9916 25220
rect 11980 25236 12032 25288
rect 12164 25236 12216 25288
rect 13912 25279 13964 25288
rect 13912 25245 13921 25279
rect 13921 25245 13955 25279
rect 13955 25245 13964 25279
rect 13912 25236 13964 25245
rect 16764 25304 16816 25356
rect 27804 25372 27856 25424
rect 12256 25168 12308 25220
rect 13636 25211 13688 25220
rect 13636 25177 13645 25211
rect 13645 25177 13679 25211
rect 13679 25177 13688 25211
rect 13636 25168 13688 25177
rect 14556 25168 14608 25220
rect 16488 25279 16540 25288
rect 16488 25245 16497 25279
rect 16497 25245 16531 25279
rect 16531 25245 16540 25279
rect 16488 25236 16540 25245
rect 26608 25279 26660 25288
rect 16212 25211 16264 25220
rect 16212 25177 16221 25211
rect 16221 25177 16255 25211
rect 16255 25177 16264 25211
rect 16212 25168 16264 25177
rect 16580 25168 16632 25220
rect 9956 25100 10008 25152
rect 11152 25143 11204 25152
rect 11152 25109 11161 25143
rect 11161 25109 11195 25143
rect 11195 25109 11204 25143
rect 11152 25100 11204 25109
rect 11244 25100 11296 25152
rect 12164 25143 12216 25152
rect 12164 25109 12173 25143
rect 12173 25109 12207 25143
rect 12207 25109 12216 25143
rect 12164 25100 12216 25109
rect 15844 25143 15896 25152
rect 15844 25109 15853 25143
rect 15853 25109 15887 25143
rect 15887 25109 15896 25143
rect 15844 25100 15896 25109
rect 16948 25168 17000 25220
rect 18236 25100 18288 25152
rect 19064 25143 19116 25152
rect 19064 25109 19073 25143
rect 19073 25109 19107 25143
rect 19107 25109 19116 25143
rect 19064 25100 19116 25109
rect 19524 25211 19576 25220
rect 19524 25177 19533 25211
rect 19533 25177 19567 25211
rect 19567 25177 19576 25211
rect 19524 25168 19576 25177
rect 19984 25168 20036 25220
rect 20076 25168 20128 25220
rect 23480 25168 23532 25220
rect 24676 25211 24728 25220
rect 24676 25177 24685 25211
rect 24685 25177 24719 25211
rect 24719 25177 24728 25211
rect 24676 25168 24728 25177
rect 25412 25211 25464 25220
rect 25412 25177 25421 25211
rect 25421 25177 25455 25211
rect 25455 25177 25464 25211
rect 25412 25168 25464 25177
rect 26608 25245 26617 25279
rect 26617 25245 26651 25279
rect 26651 25245 26660 25279
rect 26608 25236 26660 25245
rect 29828 25483 29880 25492
rect 29828 25449 29837 25483
rect 29837 25449 29871 25483
rect 29871 25449 29880 25483
rect 29828 25440 29880 25449
rect 30012 25440 30064 25492
rect 32588 25440 32640 25492
rect 31392 25304 31444 25356
rect 33416 25347 33468 25356
rect 33416 25313 33425 25347
rect 33425 25313 33459 25347
rect 33459 25313 33468 25347
rect 33416 25304 33468 25313
rect 29184 25168 29236 25220
rect 29828 25168 29880 25220
rect 31852 25236 31904 25288
rect 32588 25168 32640 25220
rect 26976 25100 27028 25152
rect 30196 25100 30248 25152
rect 30840 25143 30892 25152
rect 30840 25109 30849 25143
rect 30849 25109 30883 25143
rect 30883 25109 30892 25143
rect 30840 25100 30892 25109
rect 9344 24998 9396 25050
rect 9408 24998 9460 25050
rect 9472 24998 9524 25050
rect 9536 24998 9588 25050
rect 9600 24998 9652 25050
rect 17738 24998 17790 25050
rect 17802 24998 17854 25050
rect 17866 24998 17918 25050
rect 17930 24998 17982 25050
rect 17994 24998 18046 25050
rect 26132 24998 26184 25050
rect 26196 24998 26248 25050
rect 26260 24998 26312 25050
rect 26324 24998 26376 25050
rect 26388 24998 26440 25050
rect 34526 24998 34578 25050
rect 34590 24998 34642 25050
rect 34654 24998 34706 25050
rect 34718 24998 34770 25050
rect 34782 24998 34834 25050
rect 3424 24896 3476 24948
rect 4436 24896 4488 24948
rect 4712 24896 4764 24948
rect 4804 24871 4856 24880
rect 4804 24837 4813 24871
rect 4813 24837 4847 24871
rect 4847 24837 4856 24871
rect 4804 24828 4856 24837
rect 6460 24896 6512 24948
rect 7748 24939 7800 24948
rect 7748 24905 7757 24939
rect 7757 24905 7791 24939
rect 7791 24905 7800 24939
rect 7748 24896 7800 24905
rect 2872 24692 2924 24744
rect 3148 24556 3200 24608
rect 4344 24760 4396 24812
rect 5724 24760 5776 24812
rect 7012 24828 7064 24880
rect 3332 24692 3384 24744
rect 9036 24896 9088 24948
rect 9220 24896 9272 24948
rect 9864 24896 9916 24948
rect 5632 24624 5684 24676
rect 4528 24556 4580 24608
rect 6368 24599 6420 24608
rect 6368 24565 6377 24599
rect 6377 24565 6411 24599
rect 6411 24565 6420 24599
rect 6368 24556 6420 24565
rect 11152 24896 11204 24948
rect 12072 24939 12124 24948
rect 12072 24905 12081 24939
rect 12081 24905 12115 24939
rect 12115 24905 12124 24939
rect 12072 24896 12124 24905
rect 12256 24896 12308 24948
rect 12716 24896 12768 24948
rect 13636 24896 13688 24948
rect 15384 24896 15436 24948
rect 16488 24939 16540 24948
rect 16488 24905 16497 24939
rect 16497 24905 16531 24939
rect 16531 24905 16540 24939
rect 16488 24896 16540 24905
rect 12164 24871 12216 24880
rect 9128 24692 9180 24744
rect 11152 24803 11204 24812
rect 11152 24769 11161 24803
rect 11161 24769 11195 24803
rect 11195 24769 11204 24803
rect 11152 24760 11204 24769
rect 11520 24760 11572 24812
rect 12164 24837 12173 24871
rect 12173 24837 12207 24871
rect 12207 24837 12216 24871
rect 12164 24828 12216 24837
rect 15108 24828 15160 24880
rect 18236 24939 18288 24948
rect 18236 24905 18245 24939
rect 18245 24905 18279 24939
rect 18279 24905 18288 24939
rect 18236 24896 18288 24905
rect 19524 24939 19576 24948
rect 19524 24905 19533 24939
rect 19533 24905 19567 24939
rect 19567 24905 19576 24939
rect 19524 24896 19576 24905
rect 11704 24803 11756 24812
rect 11704 24769 11713 24803
rect 11713 24769 11747 24803
rect 11747 24769 11756 24803
rect 11704 24760 11756 24769
rect 7012 24556 7064 24608
rect 11244 24624 11296 24676
rect 11520 24624 11572 24676
rect 12532 24760 12584 24812
rect 13912 24760 13964 24812
rect 16948 24803 17000 24812
rect 16948 24769 16957 24803
rect 16957 24769 16991 24803
rect 16991 24769 17000 24803
rect 16948 24760 17000 24769
rect 17040 24760 17092 24812
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 19340 24803 19392 24812
rect 19340 24769 19349 24803
rect 19349 24769 19383 24803
rect 19383 24769 19392 24803
rect 19340 24760 19392 24769
rect 15016 24735 15068 24744
rect 15016 24701 15025 24735
rect 15025 24701 15059 24735
rect 15059 24701 15068 24735
rect 15016 24692 15068 24701
rect 20168 24760 20220 24812
rect 21272 24760 21324 24812
rect 20996 24735 21048 24744
rect 20996 24701 21005 24735
rect 21005 24701 21039 24735
rect 21039 24701 21048 24735
rect 20996 24692 21048 24701
rect 9772 24556 9824 24608
rect 11152 24556 11204 24608
rect 11336 24599 11388 24608
rect 11336 24565 11345 24599
rect 11345 24565 11379 24599
rect 11379 24565 11388 24599
rect 11336 24556 11388 24565
rect 12348 24599 12400 24608
rect 12348 24565 12357 24599
rect 12357 24565 12391 24599
rect 12391 24565 12400 24599
rect 12348 24556 12400 24565
rect 21548 24599 21600 24608
rect 21548 24565 21557 24599
rect 21557 24565 21591 24599
rect 21591 24565 21600 24599
rect 21548 24556 21600 24565
rect 23296 24692 23348 24744
rect 23664 24939 23716 24948
rect 23664 24905 23673 24939
rect 23673 24905 23707 24939
rect 23707 24905 23716 24939
rect 23664 24896 23716 24905
rect 24860 24896 24912 24948
rect 30656 24896 30708 24948
rect 31852 24939 31904 24948
rect 31852 24905 31861 24939
rect 31861 24905 31895 24939
rect 31895 24905 31904 24939
rect 31852 24896 31904 24905
rect 25044 24828 25096 24880
rect 26976 24803 27028 24812
rect 26976 24769 26985 24803
rect 26985 24769 27019 24803
rect 27019 24769 27028 24803
rect 26976 24760 27028 24769
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 29000 24828 29052 24880
rect 30196 24828 30248 24880
rect 24400 24735 24452 24744
rect 24400 24701 24409 24735
rect 24409 24701 24443 24735
rect 24443 24701 24452 24735
rect 24400 24692 24452 24701
rect 26516 24692 26568 24744
rect 27068 24735 27120 24744
rect 27068 24701 27077 24735
rect 27077 24701 27111 24735
rect 27111 24701 27120 24735
rect 28264 24760 28316 24812
rect 27068 24692 27120 24701
rect 28632 24692 28684 24744
rect 28816 24735 28868 24744
rect 28816 24701 28825 24735
rect 28825 24701 28859 24735
rect 28859 24701 28868 24735
rect 28816 24692 28868 24701
rect 29460 24803 29512 24812
rect 29460 24769 29469 24803
rect 29469 24769 29503 24803
rect 29503 24769 29512 24803
rect 29460 24760 29512 24769
rect 24860 24624 24912 24676
rect 29184 24667 29236 24676
rect 29184 24633 29193 24667
rect 29193 24633 29227 24667
rect 29227 24633 29236 24667
rect 29184 24624 29236 24633
rect 30012 24624 30064 24676
rect 31300 24803 31352 24812
rect 31300 24769 31309 24803
rect 31309 24769 31343 24803
rect 31343 24769 31352 24803
rect 31300 24760 31352 24769
rect 31392 24803 31444 24812
rect 31392 24769 31401 24803
rect 31401 24769 31435 24803
rect 31435 24769 31444 24803
rect 31392 24760 31444 24769
rect 23112 24556 23164 24608
rect 23388 24556 23440 24608
rect 30656 24556 30708 24608
rect 31576 24556 31628 24608
rect 5147 24454 5199 24506
rect 5211 24454 5263 24506
rect 5275 24454 5327 24506
rect 5339 24454 5391 24506
rect 5403 24454 5455 24506
rect 13541 24454 13593 24506
rect 13605 24454 13657 24506
rect 13669 24454 13721 24506
rect 13733 24454 13785 24506
rect 13797 24454 13849 24506
rect 21935 24454 21987 24506
rect 21999 24454 22051 24506
rect 22063 24454 22115 24506
rect 22127 24454 22179 24506
rect 22191 24454 22243 24506
rect 30329 24454 30381 24506
rect 30393 24454 30445 24506
rect 30457 24454 30509 24506
rect 30521 24454 30573 24506
rect 30585 24454 30637 24506
rect 4344 24352 4396 24404
rect 4712 24395 4764 24404
rect 4712 24361 4721 24395
rect 4721 24361 4755 24395
rect 4755 24361 4764 24395
rect 4712 24352 4764 24361
rect 7196 24352 7248 24404
rect 11336 24352 11388 24404
rect 5724 24216 5776 24268
rect 8484 24216 8536 24268
rect 9220 24216 9272 24268
rect 4896 24191 4948 24200
rect 4896 24157 4905 24191
rect 4905 24157 4939 24191
rect 4939 24157 4948 24191
rect 4896 24148 4948 24157
rect 5080 24191 5132 24200
rect 5080 24157 5089 24191
rect 5089 24157 5123 24191
rect 5123 24157 5132 24191
rect 5080 24148 5132 24157
rect 15016 24352 15068 24404
rect 18420 24352 18472 24404
rect 19340 24352 19392 24404
rect 21272 24395 21324 24404
rect 21272 24361 21281 24395
rect 21281 24361 21315 24395
rect 21315 24361 21324 24395
rect 21272 24352 21324 24361
rect 21548 24352 21600 24404
rect 16580 24284 16632 24336
rect 6552 24123 6604 24132
rect 6552 24089 6561 24123
rect 6561 24089 6595 24123
rect 6595 24089 6604 24123
rect 6552 24080 6604 24089
rect 6644 24080 6696 24132
rect 7012 24080 7064 24132
rect 11888 24080 11940 24132
rect 4344 24055 4396 24064
rect 4344 24021 4353 24055
rect 4353 24021 4387 24055
rect 4387 24021 4396 24055
rect 4344 24012 4396 24021
rect 11244 24055 11296 24064
rect 11244 24021 11253 24055
rect 11253 24021 11287 24055
rect 11287 24021 11296 24055
rect 11244 24012 11296 24021
rect 15844 24148 15896 24200
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 19064 24284 19116 24336
rect 17500 24148 17552 24157
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20168 24148 20220 24200
rect 23112 24216 23164 24268
rect 25412 24216 25464 24268
rect 25872 24148 25924 24200
rect 26148 24148 26200 24200
rect 27068 24216 27120 24268
rect 28540 24284 28592 24336
rect 31576 24395 31628 24404
rect 31576 24361 31585 24395
rect 31585 24361 31619 24395
rect 31619 24361 31628 24395
rect 31576 24352 31628 24361
rect 32588 24395 32640 24404
rect 32588 24361 32597 24395
rect 32597 24361 32631 24395
rect 32631 24361 32640 24395
rect 32588 24352 32640 24361
rect 27160 24191 27212 24200
rect 27160 24157 27169 24191
rect 27169 24157 27203 24191
rect 27203 24157 27212 24191
rect 27160 24148 27212 24157
rect 12072 24012 12124 24064
rect 17316 24012 17368 24064
rect 18788 24080 18840 24132
rect 19708 24080 19760 24132
rect 22468 24080 22520 24132
rect 24860 24123 24912 24132
rect 24860 24089 24869 24123
rect 24869 24089 24903 24123
rect 24903 24089 24912 24123
rect 24860 24080 24912 24089
rect 25320 24080 25372 24132
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 23388 24012 23440 24064
rect 29460 24148 29512 24200
rect 32128 24284 32180 24336
rect 32956 24148 33008 24200
rect 34336 24191 34388 24200
rect 34336 24157 34345 24191
rect 34345 24157 34379 24191
rect 34379 24157 34388 24191
rect 34336 24148 34388 24157
rect 26608 24012 26660 24064
rect 29828 24080 29880 24132
rect 34060 24123 34112 24132
rect 34060 24089 34069 24123
rect 34069 24089 34103 24123
rect 34103 24089 34112 24123
rect 34060 24080 34112 24089
rect 27896 24055 27948 24064
rect 27896 24021 27905 24055
rect 27905 24021 27939 24055
rect 27939 24021 27948 24055
rect 27896 24012 27948 24021
rect 30104 24012 30156 24064
rect 31300 24012 31352 24064
rect 9344 23910 9396 23962
rect 9408 23910 9460 23962
rect 9472 23910 9524 23962
rect 9536 23910 9588 23962
rect 9600 23910 9652 23962
rect 17738 23910 17790 23962
rect 17802 23910 17854 23962
rect 17866 23910 17918 23962
rect 17930 23910 17982 23962
rect 17994 23910 18046 23962
rect 26132 23910 26184 23962
rect 26196 23910 26248 23962
rect 26260 23910 26312 23962
rect 26324 23910 26376 23962
rect 26388 23910 26440 23962
rect 34526 23910 34578 23962
rect 34590 23910 34642 23962
rect 34654 23910 34706 23962
rect 34718 23910 34770 23962
rect 34782 23910 34834 23962
rect 4344 23808 4396 23860
rect 5724 23808 5776 23860
rect 6368 23808 6420 23860
rect 6552 23851 6604 23860
rect 6552 23817 6561 23851
rect 6561 23817 6595 23851
rect 6595 23817 6604 23851
rect 6552 23808 6604 23817
rect 12072 23851 12124 23860
rect 12072 23817 12081 23851
rect 12081 23817 12115 23851
rect 12115 23817 12124 23851
rect 12072 23808 12124 23817
rect 4528 23740 4580 23792
rect 3148 23672 3200 23724
rect 9772 23740 9824 23792
rect 8484 23715 8536 23724
rect 8484 23681 8493 23715
rect 8493 23681 8527 23715
rect 8527 23681 8536 23715
rect 8484 23672 8536 23681
rect 12348 23672 12400 23724
rect 13912 23808 13964 23860
rect 19432 23808 19484 23860
rect 19524 23851 19576 23860
rect 19524 23817 19533 23851
rect 19533 23817 19567 23851
rect 19567 23817 19576 23851
rect 19524 23808 19576 23817
rect 20720 23808 20772 23860
rect 23020 23808 23072 23860
rect 23296 23808 23348 23860
rect 13176 23783 13228 23792
rect 13176 23749 13185 23783
rect 13185 23749 13219 23783
rect 13219 23749 13228 23783
rect 13176 23740 13228 23749
rect 14464 23740 14516 23792
rect 15108 23740 15160 23792
rect 16764 23740 16816 23792
rect 8208 23604 8260 23656
rect 19248 23672 19300 23724
rect 26608 23808 26660 23860
rect 27160 23808 27212 23860
rect 27712 23808 27764 23860
rect 27896 23808 27948 23860
rect 22284 23672 22336 23724
rect 25228 23740 25280 23792
rect 25964 23740 26016 23792
rect 26516 23672 26568 23724
rect 24676 23647 24728 23656
rect 24676 23613 24685 23647
rect 24685 23613 24719 23647
rect 24719 23613 24728 23647
rect 24676 23604 24728 23613
rect 28632 23740 28684 23792
rect 31484 23740 31536 23792
rect 34060 23808 34112 23860
rect 28356 23672 28408 23724
rect 29736 23715 29788 23724
rect 29736 23681 29745 23715
rect 29745 23681 29779 23715
rect 29779 23681 29788 23715
rect 29736 23672 29788 23681
rect 29920 23715 29972 23724
rect 29920 23681 29929 23715
rect 29929 23681 29963 23715
rect 29963 23681 29972 23715
rect 29920 23672 29972 23681
rect 30012 23715 30064 23724
rect 30012 23681 30021 23715
rect 30021 23681 30055 23715
rect 30055 23681 30064 23715
rect 30012 23672 30064 23681
rect 30104 23715 30156 23724
rect 30104 23681 30113 23715
rect 30113 23681 30147 23715
rect 30147 23681 30156 23715
rect 30104 23672 30156 23681
rect 30288 23715 30340 23724
rect 30288 23681 30297 23715
rect 30297 23681 30331 23715
rect 30331 23681 30340 23715
rect 30288 23672 30340 23681
rect 32128 23715 32180 23724
rect 32128 23681 32137 23715
rect 32137 23681 32171 23715
rect 32171 23681 32180 23715
rect 32128 23672 32180 23681
rect 28540 23647 28592 23656
rect 28540 23613 28549 23647
rect 28549 23613 28583 23647
rect 28583 23613 28592 23647
rect 28540 23604 28592 23613
rect 24124 23579 24176 23588
rect 24124 23545 24133 23579
rect 24133 23545 24167 23579
rect 24167 23545 24176 23579
rect 24124 23536 24176 23545
rect 10232 23511 10284 23520
rect 10232 23477 10241 23511
rect 10241 23477 10275 23511
rect 10275 23477 10284 23511
rect 10232 23468 10284 23477
rect 14924 23468 14976 23520
rect 25136 23511 25188 23520
rect 25136 23477 25145 23511
rect 25145 23477 25179 23511
rect 25179 23477 25188 23511
rect 25136 23468 25188 23477
rect 27252 23511 27304 23520
rect 27252 23477 27261 23511
rect 27261 23477 27295 23511
rect 27295 23477 27304 23511
rect 27252 23468 27304 23477
rect 31300 23468 31352 23520
rect 31668 23468 31720 23520
rect 32588 23672 32640 23724
rect 32772 23715 32824 23724
rect 32772 23681 32781 23715
rect 32781 23681 32815 23715
rect 32815 23681 32824 23715
rect 32772 23672 32824 23681
rect 5147 23366 5199 23418
rect 5211 23366 5263 23418
rect 5275 23366 5327 23418
rect 5339 23366 5391 23418
rect 5403 23366 5455 23418
rect 13541 23366 13593 23418
rect 13605 23366 13657 23418
rect 13669 23366 13721 23418
rect 13733 23366 13785 23418
rect 13797 23366 13849 23418
rect 21935 23366 21987 23418
rect 21999 23366 22051 23418
rect 22063 23366 22115 23418
rect 22127 23366 22179 23418
rect 22191 23366 22243 23418
rect 30329 23366 30381 23418
rect 30393 23366 30445 23418
rect 30457 23366 30509 23418
rect 30521 23366 30573 23418
rect 30585 23366 30637 23418
rect 12348 23307 12400 23316
rect 12348 23273 12357 23307
rect 12357 23273 12391 23307
rect 12391 23273 12400 23307
rect 12348 23264 12400 23273
rect 4988 23060 5040 23112
rect 5908 23128 5960 23180
rect 11244 23128 11296 23180
rect 19248 23264 19300 23316
rect 21640 23307 21692 23316
rect 21640 23273 21649 23307
rect 21649 23273 21683 23307
rect 21683 23273 21692 23307
rect 21640 23264 21692 23273
rect 22284 23264 22336 23316
rect 24860 23264 24912 23316
rect 28356 23307 28408 23316
rect 28356 23273 28365 23307
rect 28365 23273 28399 23307
rect 28399 23273 28408 23307
rect 28356 23264 28408 23273
rect 18788 23171 18840 23180
rect 18788 23137 18797 23171
rect 18797 23137 18831 23171
rect 18831 23137 18840 23171
rect 18788 23128 18840 23137
rect 5448 23060 5500 23112
rect 6000 23103 6052 23112
rect 6000 23069 6009 23103
rect 6009 23069 6043 23103
rect 6043 23069 6052 23103
rect 6000 23060 6052 23069
rect 9220 23060 9272 23112
rect 10232 23060 10284 23112
rect 4528 22992 4580 23044
rect 4896 22924 4948 22976
rect 15108 22992 15160 23044
rect 15660 23035 15712 23044
rect 15660 23001 15669 23035
rect 15669 23001 15703 23035
rect 15703 23001 15712 23035
rect 15660 22992 15712 23001
rect 16396 23103 16448 23112
rect 16396 23069 16405 23103
rect 16405 23069 16439 23103
rect 16439 23069 16448 23103
rect 16396 23060 16448 23069
rect 20628 23128 20680 23180
rect 28540 23196 28592 23248
rect 29920 23196 29972 23248
rect 22928 23128 22980 23180
rect 23112 23128 23164 23180
rect 23296 23128 23348 23180
rect 25872 23128 25924 23180
rect 27252 23128 27304 23180
rect 27988 23128 28040 23180
rect 28908 23171 28960 23180
rect 28908 23137 28917 23171
rect 28917 23137 28951 23171
rect 28951 23137 28960 23171
rect 28908 23128 28960 23137
rect 30656 23264 30708 23316
rect 19892 23103 19944 23112
rect 19892 23069 19901 23103
rect 19901 23069 19935 23103
rect 19935 23069 19944 23103
rect 19892 23060 19944 23069
rect 22652 23060 22704 23112
rect 24124 23060 24176 23112
rect 24676 23060 24728 23112
rect 25136 23060 25188 23112
rect 29092 23060 29144 23112
rect 16764 22992 16816 23044
rect 18236 22992 18288 23044
rect 18880 23035 18932 23044
rect 18880 23001 18914 23035
rect 18914 23001 18932 23035
rect 18880 22992 18932 23001
rect 6644 22924 6696 22976
rect 7748 22924 7800 22976
rect 8760 22924 8812 22976
rect 11060 22924 11112 22976
rect 12532 22924 12584 22976
rect 15384 22924 15436 22976
rect 15844 22924 15896 22976
rect 17316 22924 17368 22976
rect 19708 22924 19760 22976
rect 20076 22924 20128 22976
rect 20628 22992 20680 23044
rect 22928 22967 22980 22976
rect 22928 22933 22937 22967
rect 22937 22933 22971 22967
rect 22971 22933 22980 22967
rect 22928 22924 22980 22933
rect 31116 23103 31168 23112
rect 31116 23069 31125 23103
rect 31125 23069 31159 23103
rect 31159 23069 31168 23103
rect 31116 23060 31168 23069
rect 31300 23103 31352 23112
rect 31300 23069 31309 23103
rect 31309 23069 31343 23103
rect 31343 23069 31352 23103
rect 31300 23060 31352 23069
rect 30840 23035 30892 23044
rect 30840 23001 30874 23035
rect 30874 23001 30892 23035
rect 30840 22992 30892 23001
rect 30012 22924 30064 22976
rect 30748 22967 30800 22976
rect 30748 22933 30757 22967
rect 30757 22933 30791 22967
rect 30791 22933 30800 22967
rect 30748 22924 30800 22933
rect 31116 22924 31168 22976
rect 9344 22822 9396 22874
rect 9408 22822 9460 22874
rect 9472 22822 9524 22874
rect 9536 22822 9588 22874
rect 9600 22822 9652 22874
rect 17738 22822 17790 22874
rect 17802 22822 17854 22874
rect 17866 22822 17918 22874
rect 17930 22822 17982 22874
rect 17994 22822 18046 22874
rect 26132 22822 26184 22874
rect 26196 22822 26248 22874
rect 26260 22822 26312 22874
rect 26324 22822 26376 22874
rect 26388 22822 26440 22874
rect 34526 22822 34578 22874
rect 34590 22822 34642 22874
rect 34654 22822 34706 22874
rect 34718 22822 34770 22874
rect 34782 22822 34834 22874
rect 6644 22652 6696 22704
rect 5448 22584 5500 22636
rect 13176 22720 13228 22772
rect 15660 22720 15712 22772
rect 16396 22720 16448 22772
rect 17500 22720 17552 22772
rect 18880 22720 18932 22772
rect 19248 22763 19300 22772
rect 19248 22729 19257 22763
rect 19257 22729 19291 22763
rect 19291 22729 19300 22763
rect 19248 22720 19300 22729
rect 29736 22720 29788 22772
rect 29920 22720 29972 22772
rect 30748 22720 30800 22772
rect 31116 22720 31168 22772
rect 14372 22652 14424 22704
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 7656 22516 7708 22568
rect 12256 22559 12308 22568
rect 12256 22525 12265 22559
rect 12265 22525 12299 22559
rect 12299 22525 12308 22559
rect 12256 22516 12308 22525
rect 12808 22516 12860 22568
rect 8300 22380 8352 22432
rect 9312 22380 9364 22432
rect 16948 22695 17000 22704
rect 16948 22661 16957 22695
rect 16957 22661 16991 22695
rect 16991 22661 17000 22695
rect 16948 22652 17000 22661
rect 17316 22652 17368 22704
rect 16580 22584 16632 22636
rect 18144 22584 18196 22636
rect 21640 22652 21692 22704
rect 18236 22516 18288 22568
rect 20720 22584 20772 22636
rect 20996 22584 21048 22636
rect 24400 22584 24452 22636
rect 28632 22627 28684 22636
rect 28632 22593 28641 22627
rect 28641 22593 28675 22627
rect 28675 22593 28684 22627
rect 28632 22584 28684 22593
rect 32956 22584 33008 22636
rect 24952 22516 25004 22568
rect 29092 22516 29144 22568
rect 30012 22516 30064 22568
rect 32220 22516 32272 22568
rect 18972 22448 19024 22500
rect 21180 22491 21232 22500
rect 21180 22457 21189 22491
rect 21189 22457 21223 22491
rect 21223 22457 21232 22491
rect 21180 22448 21232 22457
rect 32128 22448 32180 22500
rect 23572 22380 23624 22432
rect 23664 22380 23716 22432
rect 29736 22380 29788 22432
rect 32496 22423 32548 22432
rect 32496 22389 32505 22423
rect 32505 22389 32539 22423
rect 32539 22389 32548 22423
rect 32496 22380 32548 22389
rect 34336 22380 34388 22432
rect 5147 22278 5199 22330
rect 5211 22278 5263 22330
rect 5275 22278 5327 22330
rect 5339 22278 5391 22330
rect 5403 22278 5455 22330
rect 13541 22278 13593 22330
rect 13605 22278 13657 22330
rect 13669 22278 13721 22330
rect 13733 22278 13785 22330
rect 13797 22278 13849 22330
rect 21935 22278 21987 22330
rect 21999 22278 22051 22330
rect 22063 22278 22115 22330
rect 22127 22278 22179 22330
rect 22191 22278 22243 22330
rect 30329 22278 30381 22330
rect 30393 22278 30445 22330
rect 30457 22278 30509 22330
rect 30521 22278 30573 22330
rect 30585 22278 30637 22330
rect 6000 22176 6052 22228
rect 12256 22176 12308 22228
rect 24308 22176 24360 22228
rect 24952 22176 25004 22228
rect 12532 22108 12584 22160
rect 14372 22108 14424 22160
rect 1952 21972 2004 22024
rect 5448 21972 5500 22024
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 7748 22015 7800 22024
rect 7748 21981 7757 22015
rect 7757 21981 7791 22015
rect 7791 21981 7800 22015
rect 7748 21972 7800 21981
rect 8208 22083 8260 22092
rect 8208 22049 8217 22083
rect 8217 22049 8251 22083
rect 8251 22049 8260 22083
rect 8208 22040 8260 22049
rect 9312 22083 9364 22092
rect 9312 22049 9321 22083
rect 9321 22049 9355 22083
rect 9355 22049 9364 22083
rect 9312 22040 9364 22049
rect 8392 22015 8444 22024
rect 8392 21981 8402 22015
rect 8402 21981 8436 22015
rect 8436 21981 8444 22015
rect 8392 21972 8444 21981
rect 2688 21904 2740 21956
rect 4344 21904 4396 21956
rect 4528 21904 4580 21956
rect 5356 21904 5408 21956
rect 5816 21947 5868 21956
rect 5816 21913 5825 21947
rect 5825 21913 5859 21947
rect 5859 21913 5868 21947
rect 5816 21904 5868 21913
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 11060 21972 11112 22024
rect 23112 22083 23164 22092
rect 23112 22049 23121 22083
rect 23121 22049 23155 22083
rect 23155 22049 23164 22083
rect 23112 22040 23164 22049
rect 24860 22083 24912 22092
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 14280 21972 14332 22024
rect 9220 21904 9272 21956
rect 11336 21947 11388 21956
rect 11336 21913 11345 21947
rect 11345 21913 11379 21947
rect 11379 21913 11388 21947
rect 11336 21904 11388 21913
rect 9956 21836 10008 21888
rect 12808 21904 12860 21956
rect 12716 21836 12768 21888
rect 14096 21879 14148 21888
rect 14096 21845 14105 21879
rect 14105 21845 14139 21879
rect 14139 21845 14148 21879
rect 14096 21836 14148 21845
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 18236 21972 18288 22024
rect 23020 21972 23072 22024
rect 24860 22049 24869 22083
rect 24869 22049 24903 22083
rect 24903 22049 24912 22083
rect 24860 22040 24912 22049
rect 32220 22219 32272 22228
rect 32220 22185 32229 22219
rect 32229 22185 32263 22219
rect 32263 22185 32272 22219
rect 32220 22176 32272 22185
rect 33416 22108 33468 22160
rect 23664 21972 23716 22024
rect 17500 21904 17552 21956
rect 14740 21836 14792 21888
rect 18604 21836 18656 21888
rect 19708 21836 19760 21888
rect 20628 21836 20680 21888
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 30288 21972 30340 22024
rect 32496 22040 32548 22092
rect 31668 22015 31720 22024
rect 31668 21981 31677 22015
rect 31677 21981 31711 22015
rect 31711 21981 31720 22015
rect 31668 21972 31720 21981
rect 23204 21836 23256 21888
rect 23296 21879 23348 21888
rect 23296 21845 23305 21879
rect 23305 21845 23339 21879
rect 23339 21845 23348 21879
rect 23296 21836 23348 21845
rect 23848 21879 23900 21888
rect 23848 21845 23857 21879
rect 23857 21845 23891 21879
rect 23891 21845 23900 21879
rect 23848 21836 23900 21845
rect 31484 21947 31536 21956
rect 31484 21913 31493 21947
rect 31493 21913 31527 21947
rect 31527 21913 31536 21947
rect 31484 21904 31536 21913
rect 25320 21836 25372 21888
rect 26608 21879 26660 21888
rect 26608 21845 26617 21879
rect 26617 21845 26651 21879
rect 26651 21845 26660 21879
rect 26608 21836 26660 21845
rect 28632 21836 28684 21888
rect 32680 22015 32732 22024
rect 32680 21981 32689 22015
rect 32689 21981 32723 22015
rect 32723 21981 32732 22015
rect 32680 21972 32732 21981
rect 32588 21879 32640 21888
rect 32588 21845 32597 21879
rect 32597 21845 32631 21879
rect 32631 21845 32640 21879
rect 32588 21836 32640 21845
rect 32772 21836 32824 21888
rect 33232 21879 33284 21888
rect 33232 21845 33241 21879
rect 33241 21845 33275 21879
rect 33275 21845 33284 21879
rect 33232 21836 33284 21845
rect 9344 21734 9396 21786
rect 9408 21734 9460 21786
rect 9472 21734 9524 21786
rect 9536 21734 9588 21786
rect 9600 21734 9652 21786
rect 17738 21734 17790 21786
rect 17802 21734 17854 21786
rect 17866 21734 17918 21786
rect 17930 21734 17982 21786
rect 17994 21734 18046 21786
rect 26132 21734 26184 21786
rect 26196 21734 26248 21786
rect 26260 21734 26312 21786
rect 26324 21734 26376 21786
rect 26388 21734 26440 21786
rect 34526 21734 34578 21786
rect 34590 21734 34642 21786
rect 34654 21734 34706 21786
rect 34718 21734 34770 21786
rect 34782 21734 34834 21786
rect 4344 21632 4396 21684
rect 7288 21632 7340 21684
rect 8392 21632 8444 21684
rect 4712 21496 4764 21548
rect 5356 21539 5408 21548
rect 5356 21505 5365 21539
rect 5365 21505 5399 21539
rect 5399 21505 5408 21539
rect 5356 21496 5408 21505
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 7288 21496 7340 21548
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 7564 21428 7616 21480
rect 6000 21360 6052 21412
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 9220 21632 9272 21684
rect 9956 21632 10008 21684
rect 12992 21632 13044 21684
rect 14096 21632 14148 21684
rect 15844 21632 15896 21684
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 17500 21564 17552 21616
rect 17868 21607 17920 21616
rect 17868 21573 17877 21607
rect 17877 21573 17911 21607
rect 17911 21573 17920 21607
rect 17868 21564 17920 21573
rect 18144 21564 18196 21616
rect 18236 21564 18288 21616
rect 10968 21496 11020 21548
rect 4804 21292 4856 21344
rect 5448 21292 5500 21344
rect 12624 21496 12676 21548
rect 12716 21496 12768 21548
rect 12808 21539 12860 21548
rect 12808 21505 12817 21539
rect 12817 21505 12851 21539
rect 12851 21505 12860 21539
rect 12808 21496 12860 21505
rect 16304 21539 16356 21548
rect 16304 21505 16313 21539
rect 16313 21505 16347 21539
rect 16347 21505 16356 21539
rect 16304 21496 16356 21505
rect 13268 21360 13320 21412
rect 17960 21471 18012 21480
rect 17960 21437 17969 21471
rect 17969 21437 18003 21471
rect 18003 21437 18012 21471
rect 17960 21428 18012 21437
rect 18052 21471 18104 21480
rect 18052 21437 18086 21471
rect 18086 21437 18104 21471
rect 18052 21428 18104 21437
rect 19892 21632 19944 21684
rect 18604 21607 18656 21616
rect 18604 21573 18613 21607
rect 18613 21573 18647 21607
rect 18647 21573 18656 21607
rect 18604 21564 18656 21573
rect 19708 21496 19760 21548
rect 19248 21428 19300 21480
rect 22928 21632 22980 21684
rect 24952 21632 25004 21684
rect 26608 21632 26660 21684
rect 30656 21632 30708 21684
rect 31208 21632 31260 21684
rect 33232 21632 33284 21684
rect 21180 21564 21232 21616
rect 21640 21564 21692 21616
rect 25136 21564 25188 21616
rect 27712 21564 27764 21616
rect 31392 21607 31444 21616
rect 31392 21573 31401 21607
rect 31401 21573 31435 21607
rect 31435 21573 31444 21607
rect 31392 21564 31444 21573
rect 20720 21496 20772 21548
rect 22652 21496 22704 21548
rect 25044 21496 25096 21548
rect 25320 21496 25372 21548
rect 26608 21539 26660 21548
rect 26608 21505 26617 21539
rect 26617 21505 26651 21539
rect 26651 21505 26660 21539
rect 26608 21496 26660 21505
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 29920 21539 29972 21548
rect 20812 21360 20864 21412
rect 23020 21428 23072 21480
rect 23848 21428 23900 21480
rect 24584 21428 24636 21480
rect 25228 21428 25280 21480
rect 29920 21505 29929 21539
rect 29929 21505 29963 21539
rect 29963 21505 29972 21539
rect 29920 21496 29972 21505
rect 30932 21496 30984 21548
rect 11152 21292 11204 21344
rect 12440 21292 12492 21344
rect 15936 21292 15988 21344
rect 16948 21292 17000 21344
rect 17868 21292 17920 21344
rect 20628 21292 20680 21344
rect 20720 21335 20772 21344
rect 20720 21301 20729 21335
rect 20729 21301 20763 21335
rect 20763 21301 20772 21335
rect 20720 21292 20772 21301
rect 20904 21335 20956 21344
rect 20904 21301 20913 21335
rect 20913 21301 20947 21335
rect 20947 21301 20956 21335
rect 20904 21292 20956 21301
rect 21640 21335 21692 21344
rect 21640 21301 21649 21335
rect 21649 21301 21683 21335
rect 21683 21301 21692 21335
rect 21640 21292 21692 21301
rect 23204 21292 23256 21344
rect 30748 21471 30800 21480
rect 30748 21437 30757 21471
rect 30757 21437 30791 21471
rect 30791 21437 30800 21471
rect 30748 21428 30800 21437
rect 31116 21428 31168 21480
rect 26516 21292 26568 21344
rect 26884 21292 26936 21344
rect 28816 21335 28868 21344
rect 28816 21301 28825 21335
rect 28825 21301 28859 21335
rect 28859 21301 28868 21335
rect 28816 21292 28868 21301
rect 29828 21292 29880 21344
rect 30104 21292 30156 21344
rect 30288 21292 30340 21344
rect 30564 21335 30616 21344
rect 30564 21301 30573 21335
rect 30573 21301 30607 21335
rect 30607 21301 30616 21335
rect 30564 21292 30616 21301
rect 30840 21292 30892 21344
rect 31300 21292 31352 21344
rect 31484 21292 31536 21344
rect 34796 21496 34848 21548
rect 5147 21190 5199 21242
rect 5211 21190 5263 21242
rect 5275 21190 5327 21242
rect 5339 21190 5391 21242
rect 5403 21190 5455 21242
rect 13541 21190 13593 21242
rect 13605 21190 13657 21242
rect 13669 21190 13721 21242
rect 13733 21190 13785 21242
rect 13797 21190 13849 21242
rect 21935 21190 21987 21242
rect 21999 21190 22051 21242
rect 22063 21190 22115 21242
rect 22127 21190 22179 21242
rect 22191 21190 22243 21242
rect 30329 21190 30381 21242
rect 30393 21190 30445 21242
rect 30457 21190 30509 21242
rect 30521 21190 30573 21242
rect 30585 21190 30637 21242
rect 9680 21088 9732 21140
rect 12348 21088 12400 21140
rect 13268 21088 13320 21140
rect 15936 21088 15988 21140
rect 16304 21088 16356 21140
rect 18052 21088 18104 21140
rect 20628 21088 20680 21140
rect 20812 21088 20864 21140
rect 20904 21088 20956 21140
rect 21732 21088 21784 21140
rect 22468 21088 22520 21140
rect 26608 21088 26660 21140
rect 28816 21088 28868 21140
rect 29920 21088 29972 21140
rect 30748 21088 30800 21140
rect 30840 21131 30892 21140
rect 30840 21097 30849 21131
rect 30849 21097 30883 21131
rect 30883 21097 30892 21131
rect 30840 21088 30892 21097
rect 30932 21088 30984 21140
rect 31116 21088 31168 21140
rect 12440 20952 12492 21004
rect 13176 20952 13228 21004
rect 15844 20952 15896 21004
rect 5540 20884 5592 20936
rect 6736 20884 6788 20936
rect 7104 20884 7156 20936
rect 11336 20927 11388 20936
rect 11336 20893 11345 20927
rect 11345 20893 11379 20927
rect 11379 20893 11388 20927
rect 11336 20884 11388 20893
rect 11520 20927 11572 20936
rect 11520 20893 11529 20927
rect 11529 20893 11563 20927
rect 11563 20893 11572 20927
rect 11520 20884 11572 20893
rect 12532 20884 12584 20936
rect 14740 20884 14792 20936
rect 17500 20884 17552 20936
rect 18236 20884 18288 20936
rect 20168 20927 20220 20936
rect 20168 20893 20177 20927
rect 20177 20893 20211 20927
rect 20211 20893 20220 20927
rect 20168 20884 20220 20893
rect 23112 21020 23164 21072
rect 4988 20859 5040 20868
rect 4988 20825 4997 20859
rect 4997 20825 5031 20859
rect 5031 20825 5040 20859
rect 4988 20816 5040 20825
rect 6276 20816 6328 20868
rect 7472 20816 7524 20868
rect 17868 20859 17920 20868
rect 17868 20825 17877 20859
rect 17877 20825 17911 20859
rect 17911 20825 17920 20859
rect 17868 20816 17920 20825
rect 18788 20859 18840 20868
rect 18788 20825 18797 20859
rect 18797 20825 18831 20859
rect 18831 20825 18840 20859
rect 18788 20816 18840 20825
rect 19248 20816 19300 20868
rect 21548 20884 21600 20936
rect 21824 20884 21876 20936
rect 22744 20884 22796 20936
rect 22928 20927 22980 20936
rect 22928 20893 22937 20927
rect 22937 20893 22971 20927
rect 22971 20893 22980 20927
rect 22928 20884 22980 20893
rect 22376 20816 22428 20868
rect 4804 20748 4856 20800
rect 5540 20748 5592 20800
rect 17316 20791 17368 20800
rect 17316 20757 17325 20791
rect 17325 20757 17359 20791
rect 17359 20757 17368 20791
rect 17316 20748 17368 20757
rect 17592 20748 17644 20800
rect 17960 20748 18012 20800
rect 18512 20748 18564 20800
rect 20352 20748 20404 20800
rect 22652 20748 22704 20800
rect 22928 20748 22980 20800
rect 24400 20791 24452 20800
rect 24400 20757 24409 20791
rect 24409 20757 24443 20791
rect 24443 20757 24452 20791
rect 24400 20748 24452 20757
rect 25412 20791 25464 20800
rect 25412 20757 25421 20791
rect 25421 20757 25455 20791
rect 25455 20757 25464 20791
rect 25412 20748 25464 20757
rect 25596 20927 25648 20936
rect 25596 20893 25605 20927
rect 25605 20893 25639 20927
rect 25639 20893 25648 20927
rect 25596 20884 25648 20893
rect 26884 20952 26936 21004
rect 30104 21020 30156 21072
rect 28724 20927 28776 20936
rect 28724 20893 28733 20927
rect 28733 20893 28767 20927
rect 28767 20893 28776 20927
rect 28724 20884 28776 20893
rect 30656 20952 30708 21004
rect 34336 20995 34388 21004
rect 34336 20961 34345 20995
rect 34345 20961 34379 20995
rect 34379 20961 34388 20995
rect 34336 20952 34388 20961
rect 32036 20884 32088 20936
rect 32588 20884 32640 20936
rect 32956 20884 33008 20936
rect 28172 20791 28224 20800
rect 28172 20757 28181 20791
rect 28181 20757 28215 20791
rect 28215 20757 28224 20791
rect 28172 20748 28224 20757
rect 30932 20816 30984 20868
rect 9344 20646 9396 20698
rect 9408 20646 9460 20698
rect 9472 20646 9524 20698
rect 9536 20646 9588 20698
rect 9600 20646 9652 20698
rect 17738 20646 17790 20698
rect 17802 20646 17854 20698
rect 17866 20646 17918 20698
rect 17930 20646 17982 20698
rect 17994 20646 18046 20698
rect 26132 20646 26184 20698
rect 26196 20646 26248 20698
rect 26260 20646 26312 20698
rect 26324 20646 26376 20698
rect 26388 20646 26440 20698
rect 34526 20646 34578 20698
rect 34590 20646 34642 20698
rect 34654 20646 34706 20698
rect 34718 20646 34770 20698
rect 34782 20646 34834 20698
rect 4988 20587 5040 20596
rect 4988 20553 4997 20587
rect 4997 20553 5031 20587
rect 5031 20553 5040 20587
rect 4988 20544 5040 20553
rect 6368 20544 6420 20596
rect 6920 20544 6972 20596
rect 8668 20544 8720 20596
rect 10600 20544 10652 20596
rect 11520 20544 11572 20596
rect 15844 20544 15896 20596
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 18144 20587 18196 20596
rect 18144 20553 18153 20587
rect 18153 20553 18187 20587
rect 18187 20553 18196 20587
rect 18144 20544 18196 20553
rect 21548 20544 21600 20596
rect 2688 20476 2740 20528
rect 4896 20476 4948 20528
rect 4528 20451 4580 20460
rect 4528 20417 4537 20451
rect 4537 20417 4571 20451
rect 4571 20417 4580 20451
rect 4528 20408 4580 20417
rect 5908 20476 5960 20528
rect 1400 20340 1452 20392
rect 1952 20383 2004 20392
rect 1952 20349 1961 20383
rect 1961 20349 1995 20383
rect 1995 20349 2004 20383
rect 1952 20340 2004 20349
rect 2320 20383 2372 20392
rect 2320 20349 2329 20383
rect 2329 20349 2363 20383
rect 2363 20349 2372 20383
rect 2320 20340 2372 20349
rect 4620 20383 4672 20392
rect 4620 20349 4629 20383
rect 4629 20349 4663 20383
rect 4663 20349 4672 20383
rect 4620 20340 4672 20349
rect 4804 20383 4856 20392
rect 4804 20349 4813 20383
rect 4813 20349 4847 20383
rect 4847 20349 4856 20383
rect 4804 20340 4856 20349
rect 5632 20451 5684 20460
rect 5632 20417 5641 20451
rect 5641 20417 5675 20451
rect 5675 20417 5684 20451
rect 5632 20408 5684 20417
rect 5724 20408 5776 20460
rect 5816 20408 5868 20460
rect 6276 20408 6328 20460
rect 6552 20451 6604 20460
rect 6552 20417 6561 20451
rect 6561 20417 6595 20451
rect 6595 20417 6604 20451
rect 6552 20408 6604 20417
rect 6920 20451 6972 20460
rect 6920 20417 6929 20451
rect 6929 20417 6963 20451
rect 6963 20417 6972 20451
rect 6920 20408 6972 20417
rect 7104 20408 7156 20460
rect 7288 20451 7340 20460
rect 7288 20417 7297 20451
rect 7297 20417 7331 20451
rect 7331 20417 7340 20451
rect 7288 20408 7340 20417
rect 7748 20476 7800 20528
rect 7472 20451 7524 20460
rect 7472 20417 7481 20451
rect 7481 20417 7515 20451
rect 7515 20417 7524 20451
rect 7472 20408 7524 20417
rect 8392 20408 8444 20460
rect 8944 20451 8996 20460
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 9680 20476 9732 20528
rect 10232 20476 10284 20528
rect 9864 20340 9916 20392
rect 10416 20451 10468 20460
rect 10416 20417 10425 20451
rect 10425 20417 10459 20451
rect 10459 20417 10468 20451
rect 10416 20408 10468 20417
rect 10600 20408 10652 20460
rect 10508 20340 10560 20392
rect 4988 20272 5040 20324
rect 4160 20247 4212 20256
rect 4160 20213 4169 20247
rect 4169 20213 4203 20247
rect 4203 20213 4212 20247
rect 4160 20204 4212 20213
rect 6000 20204 6052 20256
rect 8668 20272 8720 20324
rect 12256 20451 12308 20460
rect 12256 20417 12265 20451
rect 12265 20417 12299 20451
rect 12299 20417 12308 20451
rect 12256 20408 12308 20417
rect 12440 20451 12492 20460
rect 12440 20417 12461 20451
rect 12461 20417 12492 20451
rect 12440 20408 12492 20417
rect 12900 20408 12952 20460
rect 14740 20408 14792 20460
rect 17224 20476 17276 20528
rect 18788 20476 18840 20528
rect 21640 20476 21692 20528
rect 17040 20408 17092 20460
rect 17316 20451 17368 20460
rect 17316 20417 17325 20451
rect 17325 20417 17359 20451
rect 17359 20417 17368 20451
rect 17316 20408 17368 20417
rect 17868 20408 17920 20460
rect 26976 20544 27028 20596
rect 21732 20408 21784 20460
rect 22468 20451 22520 20460
rect 22468 20417 22477 20451
rect 22477 20417 22511 20451
rect 22511 20417 22520 20451
rect 22468 20408 22520 20417
rect 23112 20476 23164 20528
rect 25412 20476 25464 20528
rect 27712 20476 27764 20528
rect 24860 20408 24912 20460
rect 29736 20544 29788 20596
rect 30932 20544 30984 20596
rect 31392 20544 31444 20596
rect 32680 20544 32732 20596
rect 28080 20476 28132 20528
rect 30748 20476 30800 20528
rect 31116 20476 31168 20528
rect 33048 20408 33100 20460
rect 21548 20272 21600 20324
rect 7288 20204 7340 20256
rect 7564 20247 7616 20256
rect 7564 20213 7573 20247
rect 7573 20213 7607 20247
rect 7607 20213 7616 20247
rect 7564 20204 7616 20213
rect 7748 20247 7800 20256
rect 7748 20213 7757 20247
rect 7757 20213 7791 20247
rect 7791 20213 7800 20247
rect 7748 20204 7800 20213
rect 10324 20204 10376 20256
rect 10968 20204 11020 20256
rect 12624 20204 12676 20256
rect 14372 20247 14424 20256
rect 14372 20213 14381 20247
rect 14381 20213 14415 20247
rect 14415 20213 14424 20247
rect 14372 20204 14424 20213
rect 17868 20204 17920 20256
rect 21180 20204 21232 20256
rect 22376 20204 22428 20256
rect 22928 20204 22980 20256
rect 25688 20204 25740 20256
rect 30012 20272 30064 20324
rect 33416 20383 33468 20392
rect 33416 20349 33425 20383
rect 33425 20349 33459 20383
rect 33459 20349 33468 20383
rect 33416 20340 33468 20349
rect 27712 20204 27764 20256
rect 27988 20204 28040 20256
rect 28172 20247 28224 20256
rect 28172 20213 28202 20247
rect 28202 20213 28224 20247
rect 28172 20204 28224 20213
rect 29920 20204 29972 20256
rect 5147 20102 5199 20154
rect 5211 20102 5263 20154
rect 5275 20102 5327 20154
rect 5339 20102 5391 20154
rect 5403 20102 5455 20154
rect 13541 20102 13593 20154
rect 13605 20102 13657 20154
rect 13669 20102 13721 20154
rect 13733 20102 13785 20154
rect 13797 20102 13849 20154
rect 21935 20102 21987 20154
rect 21999 20102 22051 20154
rect 22063 20102 22115 20154
rect 22127 20102 22179 20154
rect 22191 20102 22243 20154
rect 30329 20102 30381 20154
rect 30393 20102 30445 20154
rect 30457 20102 30509 20154
rect 30521 20102 30573 20154
rect 30585 20102 30637 20154
rect 2320 20000 2372 20052
rect 4160 20000 4212 20052
rect 4620 20000 4672 20052
rect 4712 20000 4764 20052
rect 5540 20000 5592 20052
rect 7104 20043 7156 20052
rect 7104 20009 7113 20043
rect 7113 20009 7147 20043
rect 7147 20009 7156 20043
rect 7104 20000 7156 20009
rect 7748 20000 7800 20052
rect 9864 20000 9916 20052
rect 10416 20000 10468 20052
rect 12256 20000 12308 20052
rect 12532 20000 12584 20052
rect 940 19796 992 19848
rect 4620 19796 4672 19848
rect 4804 19796 4856 19848
rect 6644 19864 6696 19916
rect 7288 19864 7340 19916
rect 4160 19728 4212 19780
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 3608 19660 3660 19712
rect 5724 19839 5776 19848
rect 5724 19805 5733 19839
rect 5733 19805 5767 19839
rect 5767 19805 5776 19839
rect 5724 19796 5776 19805
rect 5908 19839 5960 19848
rect 5908 19805 5917 19839
rect 5917 19805 5951 19839
rect 5951 19805 5960 19839
rect 5908 19796 5960 19805
rect 7196 19839 7248 19848
rect 7196 19805 7205 19839
rect 7205 19805 7239 19839
rect 7239 19805 7248 19839
rect 7196 19796 7248 19805
rect 6000 19771 6052 19780
rect 6000 19737 6009 19771
rect 6009 19737 6043 19771
rect 6043 19737 6052 19771
rect 6000 19728 6052 19737
rect 6828 19728 6880 19780
rect 8392 19796 8444 19848
rect 9036 19796 9088 19848
rect 9680 19796 9732 19848
rect 10232 19932 10284 19984
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 11060 19864 11112 19916
rect 11336 19796 11388 19848
rect 17224 20000 17276 20052
rect 18236 20000 18288 20052
rect 22468 20000 22520 20052
rect 25596 20000 25648 20052
rect 28724 20000 28776 20052
rect 29920 20000 29972 20052
rect 30012 20043 30064 20052
rect 30012 20009 30021 20043
rect 30021 20009 30055 20043
rect 30055 20009 30064 20043
rect 30012 20000 30064 20009
rect 21180 19932 21232 19984
rect 19616 19864 19668 19916
rect 23020 19864 23072 19916
rect 5448 19703 5500 19712
rect 5448 19669 5457 19703
rect 5457 19669 5491 19703
rect 5491 19669 5500 19703
rect 5448 19660 5500 19669
rect 5540 19660 5592 19712
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 13452 19728 13504 19780
rect 17040 19728 17092 19780
rect 18512 19796 18564 19848
rect 19708 19796 19760 19848
rect 22560 19839 22612 19848
rect 22560 19805 22569 19839
rect 22569 19805 22603 19839
rect 22603 19805 22612 19839
rect 22560 19796 22612 19805
rect 22744 19839 22796 19848
rect 22744 19805 22753 19839
rect 22753 19805 22787 19839
rect 22787 19805 22796 19839
rect 23756 19932 23808 19984
rect 23204 19864 23256 19916
rect 22744 19796 22796 19805
rect 23296 19796 23348 19848
rect 23756 19796 23808 19848
rect 17592 19728 17644 19780
rect 26884 19864 26936 19916
rect 10508 19703 10560 19712
rect 10508 19669 10517 19703
rect 10517 19669 10551 19703
rect 10551 19669 10560 19703
rect 10508 19660 10560 19669
rect 11060 19660 11112 19712
rect 17132 19703 17184 19712
rect 17132 19669 17157 19703
rect 17157 19669 17184 19703
rect 17132 19660 17184 19669
rect 17316 19660 17368 19712
rect 17500 19660 17552 19712
rect 18144 19660 18196 19712
rect 19340 19703 19392 19712
rect 19340 19669 19349 19703
rect 19349 19669 19383 19703
rect 19383 19669 19392 19703
rect 19340 19660 19392 19669
rect 22284 19660 22336 19712
rect 23664 19660 23716 19712
rect 25688 19839 25740 19848
rect 25688 19805 25697 19839
rect 25697 19805 25731 19839
rect 25731 19805 25740 19839
rect 25688 19796 25740 19805
rect 26792 19839 26844 19848
rect 26792 19805 26801 19839
rect 26801 19805 26835 19839
rect 26835 19805 26844 19839
rect 26792 19796 26844 19805
rect 27804 19864 27856 19916
rect 28448 19907 28500 19916
rect 28448 19873 28457 19907
rect 28457 19873 28491 19907
rect 28491 19873 28500 19907
rect 28448 19864 28500 19873
rect 28172 19728 28224 19780
rect 29368 19796 29420 19848
rect 24400 19703 24452 19712
rect 24400 19669 24409 19703
rect 24409 19669 24443 19703
rect 24443 19669 24452 19703
rect 24400 19660 24452 19669
rect 30380 19703 30432 19712
rect 30380 19669 30389 19703
rect 30389 19669 30423 19703
rect 30423 19669 30432 19703
rect 30380 19660 30432 19669
rect 9344 19558 9396 19610
rect 9408 19558 9460 19610
rect 9472 19558 9524 19610
rect 9536 19558 9588 19610
rect 9600 19558 9652 19610
rect 17738 19558 17790 19610
rect 17802 19558 17854 19610
rect 17866 19558 17918 19610
rect 17930 19558 17982 19610
rect 17994 19558 18046 19610
rect 26132 19558 26184 19610
rect 26196 19558 26248 19610
rect 26260 19558 26312 19610
rect 26324 19558 26376 19610
rect 26388 19558 26440 19610
rect 34526 19558 34578 19610
rect 34590 19558 34642 19610
rect 34654 19558 34706 19610
rect 34718 19558 34770 19610
rect 34782 19558 34834 19610
rect 3148 19499 3200 19508
rect 3148 19465 3157 19499
rect 3157 19465 3191 19499
rect 3191 19465 3200 19499
rect 3148 19456 3200 19465
rect 4160 19456 4212 19508
rect 4712 19456 4764 19508
rect 4804 19456 4856 19508
rect 4988 19456 5040 19508
rect 5632 19456 5684 19508
rect 6828 19456 6880 19508
rect 12808 19456 12860 19508
rect 13452 19456 13504 19508
rect 15292 19456 15344 19508
rect 17224 19456 17276 19508
rect 17592 19456 17644 19508
rect 19340 19456 19392 19508
rect 1584 19388 1636 19440
rect 2688 19388 2740 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 3884 19320 3936 19372
rect 7104 19388 7156 19440
rect 8392 19388 8444 19440
rect 14740 19388 14792 19440
rect 4896 19320 4948 19372
rect 5908 19320 5960 19372
rect 6920 19320 6972 19372
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 11704 19320 11756 19372
rect 11796 19363 11848 19372
rect 11796 19329 11805 19363
rect 11805 19329 11839 19363
rect 11839 19329 11848 19363
rect 11796 19320 11848 19329
rect 11980 19320 12032 19372
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 4712 19252 4764 19304
rect 5172 19252 5224 19304
rect 5724 19252 5776 19304
rect 8484 19295 8536 19304
rect 8484 19261 8493 19295
rect 8493 19261 8527 19295
rect 8527 19261 8536 19295
rect 8484 19252 8536 19261
rect 9772 19252 9824 19304
rect 13176 19320 13228 19372
rect 17316 19320 17368 19372
rect 31392 19499 31444 19508
rect 31392 19465 31401 19499
rect 31401 19465 31435 19499
rect 31435 19465 31444 19499
rect 31392 19456 31444 19465
rect 22560 19388 22612 19440
rect 23756 19388 23808 19440
rect 25044 19388 25096 19440
rect 12348 19184 12400 19236
rect 17132 19252 17184 19304
rect 20260 19320 20312 19372
rect 17592 19184 17644 19236
rect 20352 19295 20404 19304
rect 20352 19261 20361 19295
rect 20361 19261 20395 19295
rect 20395 19261 20404 19295
rect 20352 19252 20404 19261
rect 20628 19320 20680 19372
rect 20904 19252 20956 19304
rect 23480 19295 23532 19304
rect 23480 19261 23489 19295
rect 23489 19261 23523 19295
rect 23523 19261 23532 19295
rect 23480 19252 23532 19261
rect 24400 19252 24452 19304
rect 26792 19388 26844 19440
rect 26516 19363 26568 19372
rect 26516 19329 26525 19363
rect 26525 19329 26559 19363
rect 26559 19329 26568 19363
rect 26516 19320 26568 19329
rect 27344 19388 27396 19440
rect 30380 19388 30432 19440
rect 31024 19388 31076 19440
rect 5632 19116 5684 19168
rect 7564 19159 7616 19168
rect 7564 19125 7573 19159
rect 7573 19125 7607 19159
rect 7607 19125 7616 19159
rect 7564 19116 7616 19125
rect 13268 19116 13320 19168
rect 13912 19116 13964 19168
rect 23388 19184 23440 19236
rect 24952 19184 25004 19236
rect 26976 19363 27028 19372
rect 26976 19329 26985 19363
rect 26985 19329 27019 19363
rect 27019 19329 27028 19363
rect 26976 19320 27028 19329
rect 33048 19456 33100 19508
rect 28724 19295 28776 19304
rect 28724 19261 28733 19295
rect 28733 19261 28767 19295
rect 28767 19261 28776 19295
rect 28724 19252 28776 19261
rect 25136 19116 25188 19168
rect 30656 19184 30708 19236
rect 32496 19320 32548 19372
rect 31392 19252 31444 19304
rect 32680 19295 32732 19304
rect 32680 19261 32689 19295
rect 32689 19261 32723 19295
rect 32723 19261 32732 19295
rect 32680 19252 32732 19261
rect 32128 19184 32180 19236
rect 26792 19116 26844 19168
rect 30196 19159 30248 19168
rect 30196 19125 30205 19159
rect 30205 19125 30239 19159
rect 30239 19125 30248 19159
rect 30196 19116 30248 19125
rect 31576 19116 31628 19168
rect 5147 19014 5199 19066
rect 5211 19014 5263 19066
rect 5275 19014 5327 19066
rect 5339 19014 5391 19066
rect 5403 19014 5455 19066
rect 13541 19014 13593 19066
rect 13605 19014 13657 19066
rect 13669 19014 13721 19066
rect 13733 19014 13785 19066
rect 13797 19014 13849 19066
rect 21935 19014 21987 19066
rect 21999 19014 22051 19066
rect 22063 19014 22115 19066
rect 22127 19014 22179 19066
rect 22191 19014 22243 19066
rect 30329 19014 30381 19066
rect 30393 19014 30445 19066
rect 30457 19014 30509 19066
rect 30521 19014 30573 19066
rect 30585 19014 30637 19066
rect 1860 18912 1912 18964
rect 9772 18912 9824 18964
rect 12992 18912 13044 18964
rect 19616 18912 19668 18964
rect 6368 18844 6420 18896
rect 7288 18844 7340 18896
rect 1400 18776 1452 18828
rect 8300 18776 8352 18828
rect 2964 18708 3016 18760
rect 5264 18708 5316 18760
rect 5724 18708 5776 18760
rect 6920 18708 6972 18760
rect 7380 18751 7432 18760
rect 7380 18717 7389 18751
rect 7389 18717 7423 18751
rect 7423 18717 7432 18751
rect 7380 18708 7432 18717
rect 7564 18708 7616 18760
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 3700 18640 3752 18692
rect 8300 18640 8352 18692
rect 9588 18844 9640 18896
rect 9864 18844 9916 18896
rect 10324 18844 10376 18896
rect 8760 18776 8812 18828
rect 8576 18708 8628 18760
rect 9680 18708 9732 18760
rect 9772 18751 9824 18760
rect 20260 18844 20312 18896
rect 9772 18717 9799 18751
rect 9799 18717 9824 18751
rect 9772 18708 9824 18717
rect 11060 18751 11112 18760
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 11336 18708 11388 18760
rect 12808 18751 12860 18760
rect 10048 18640 10100 18692
rect 7104 18572 7156 18624
rect 7840 18572 7892 18624
rect 8576 18572 8628 18624
rect 9772 18572 9824 18624
rect 10140 18615 10192 18624
rect 10140 18581 10149 18615
rect 10149 18581 10183 18615
rect 10183 18581 10192 18615
rect 10140 18572 10192 18581
rect 12072 18640 12124 18692
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13452 18708 13504 18760
rect 13268 18640 13320 18692
rect 14096 18708 14148 18760
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 18144 18776 18196 18828
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 21824 18887 21876 18896
rect 21824 18853 21833 18887
rect 21833 18853 21867 18887
rect 21867 18853 21876 18887
rect 21824 18844 21876 18853
rect 22468 18844 22520 18896
rect 23204 18955 23256 18964
rect 23204 18921 23213 18955
rect 23213 18921 23247 18955
rect 23247 18921 23256 18955
rect 23204 18912 23256 18921
rect 26516 18912 26568 18964
rect 29368 18912 29420 18964
rect 30840 18912 30892 18964
rect 24952 18844 25004 18896
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 22560 18751 22612 18760
rect 22560 18717 22569 18751
rect 22569 18717 22603 18751
rect 22603 18717 22612 18751
rect 22560 18708 22612 18717
rect 22744 18708 22796 18760
rect 26884 18819 26936 18828
rect 26884 18785 26893 18819
rect 26893 18785 26927 18819
rect 26927 18785 26936 18819
rect 26884 18776 26936 18785
rect 28724 18776 28776 18828
rect 18880 18615 18932 18624
rect 18880 18581 18889 18615
rect 18889 18581 18923 18615
rect 18923 18581 18932 18615
rect 18880 18572 18932 18581
rect 19616 18640 19668 18692
rect 20444 18572 20496 18624
rect 22284 18640 22336 18692
rect 24400 18751 24452 18760
rect 24400 18717 24409 18751
rect 24409 18717 24443 18751
rect 24443 18717 24452 18751
rect 24400 18708 24452 18717
rect 28632 18751 28684 18760
rect 28632 18717 28641 18751
rect 28641 18717 28675 18751
rect 28675 18717 28684 18751
rect 28632 18708 28684 18717
rect 29000 18708 29052 18760
rect 28264 18640 28316 18692
rect 30196 18683 30248 18692
rect 30196 18649 30205 18683
rect 30205 18649 30239 18683
rect 30239 18649 30248 18683
rect 30196 18640 30248 18649
rect 22928 18572 22980 18624
rect 23020 18572 23072 18624
rect 23112 18572 23164 18624
rect 23296 18572 23348 18624
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 29368 18572 29420 18624
rect 30564 18751 30616 18760
rect 30564 18717 30573 18751
rect 30573 18717 30607 18751
rect 30607 18717 30616 18751
rect 30564 18708 30616 18717
rect 30656 18751 30708 18760
rect 30656 18717 30665 18751
rect 30665 18717 30699 18751
rect 30699 18717 30708 18751
rect 30656 18708 30708 18717
rect 32312 18844 32364 18896
rect 32680 18912 32732 18964
rect 31576 18751 31628 18760
rect 31576 18717 31585 18751
rect 31585 18717 31619 18751
rect 31619 18717 31628 18751
rect 31576 18708 31628 18717
rect 31668 18751 31720 18760
rect 31668 18717 31677 18751
rect 31677 18717 31711 18751
rect 31711 18717 31720 18751
rect 31668 18708 31720 18717
rect 32220 18708 32272 18760
rect 32956 18751 33008 18760
rect 32956 18717 32965 18751
rect 32965 18717 32999 18751
rect 32999 18717 33008 18751
rect 32956 18708 33008 18717
rect 32680 18640 32732 18692
rect 31392 18572 31444 18624
rect 31576 18572 31628 18624
rect 31852 18615 31904 18624
rect 31852 18581 31861 18615
rect 31861 18581 31895 18615
rect 31895 18581 31904 18615
rect 31852 18572 31904 18581
rect 32864 18572 32916 18624
rect 9344 18470 9396 18522
rect 9408 18470 9460 18522
rect 9472 18470 9524 18522
rect 9536 18470 9588 18522
rect 9600 18470 9652 18522
rect 17738 18470 17790 18522
rect 17802 18470 17854 18522
rect 17866 18470 17918 18522
rect 17930 18470 17982 18522
rect 17994 18470 18046 18522
rect 26132 18470 26184 18522
rect 26196 18470 26248 18522
rect 26260 18470 26312 18522
rect 26324 18470 26376 18522
rect 26388 18470 26440 18522
rect 34526 18470 34578 18522
rect 34590 18470 34642 18522
rect 34654 18470 34706 18522
rect 34718 18470 34770 18522
rect 34782 18470 34834 18522
rect 1860 18368 1912 18420
rect 3700 18368 3752 18420
rect 3608 18275 3660 18284
rect 3608 18241 3617 18275
rect 3617 18241 3651 18275
rect 3651 18241 3660 18275
rect 3608 18232 3660 18241
rect 3884 18300 3936 18352
rect 3976 18275 4028 18284
rect 3976 18241 3985 18275
rect 3985 18241 4019 18275
rect 4019 18241 4028 18275
rect 3976 18232 4028 18241
rect 4528 18232 4580 18284
rect 4988 18368 5040 18420
rect 5724 18368 5776 18420
rect 6920 18368 6972 18420
rect 4804 18300 4856 18352
rect 5540 18232 5592 18284
rect 5816 18232 5868 18284
rect 6368 18232 6420 18284
rect 9864 18368 9916 18420
rect 12348 18368 12400 18420
rect 8116 18343 8168 18352
rect 8116 18309 8125 18343
rect 8125 18309 8159 18343
rect 8159 18309 8168 18343
rect 8116 18300 8168 18309
rect 8300 18300 8352 18352
rect 6000 18164 6052 18216
rect 8668 18232 8720 18284
rect 8852 18300 8904 18352
rect 9128 18275 9180 18284
rect 9128 18241 9137 18275
rect 9137 18241 9171 18275
rect 9171 18241 9180 18275
rect 9128 18232 9180 18241
rect 9312 18232 9364 18284
rect 9772 18275 9824 18284
rect 9772 18241 9781 18275
rect 9781 18241 9815 18275
rect 9815 18241 9824 18275
rect 9772 18232 9824 18241
rect 10140 18232 10192 18284
rect 15752 18368 15804 18420
rect 17500 18368 17552 18420
rect 18696 18368 18748 18420
rect 11152 18232 11204 18284
rect 8484 18164 8536 18216
rect 9680 18164 9732 18216
rect 5816 18096 5868 18148
rect 8668 18096 8720 18148
rect 11980 18164 12032 18216
rect 12716 18275 12768 18284
rect 12716 18241 12725 18275
rect 12725 18241 12759 18275
rect 12759 18241 12768 18275
rect 12716 18232 12768 18241
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 4988 18028 5040 18080
rect 5264 18028 5316 18080
rect 5448 18028 5500 18080
rect 8944 18028 8996 18080
rect 12992 18164 13044 18216
rect 13728 18232 13780 18284
rect 18512 18300 18564 18352
rect 18880 18368 18932 18420
rect 23296 18368 23348 18420
rect 19524 18300 19576 18352
rect 21732 18300 21784 18352
rect 14556 18232 14608 18284
rect 15108 18275 15160 18284
rect 15108 18241 15117 18275
rect 15117 18241 15151 18275
rect 15151 18241 15160 18275
rect 15108 18232 15160 18241
rect 14740 18164 14792 18216
rect 14832 18164 14884 18216
rect 17684 18232 17736 18284
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 22928 18275 22980 18284
rect 22928 18241 22937 18275
rect 22937 18241 22971 18275
rect 22971 18241 22980 18275
rect 22928 18232 22980 18241
rect 24584 18368 24636 18420
rect 26792 18368 26844 18420
rect 23480 18232 23532 18284
rect 18052 18207 18104 18216
rect 18052 18173 18086 18207
rect 18086 18173 18104 18207
rect 18052 18164 18104 18173
rect 18236 18164 18288 18216
rect 23020 18164 23072 18216
rect 15476 18096 15528 18148
rect 15844 18096 15896 18148
rect 20260 18139 20312 18148
rect 20260 18105 20269 18139
rect 20269 18105 20303 18139
rect 20303 18105 20312 18139
rect 20260 18096 20312 18105
rect 9956 18028 10008 18080
rect 11980 18028 12032 18080
rect 12716 18028 12768 18080
rect 14740 18028 14792 18080
rect 15108 18028 15160 18080
rect 15200 18028 15252 18080
rect 15568 18028 15620 18080
rect 16304 18071 16356 18080
rect 16304 18037 16313 18071
rect 16313 18037 16347 18071
rect 16347 18037 16356 18071
rect 16304 18028 16356 18037
rect 18512 18028 18564 18080
rect 22284 18096 22336 18148
rect 23112 18096 23164 18148
rect 23664 18275 23716 18284
rect 23664 18241 23673 18275
rect 23673 18241 23707 18275
rect 23707 18241 23716 18275
rect 23664 18232 23716 18241
rect 23480 18028 23532 18080
rect 24124 18164 24176 18216
rect 24952 18300 25004 18352
rect 28356 18232 28408 18284
rect 29736 18275 29788 18284
rect 29736 18241 29745 18275
rect 29745 18241 29779 18275
rect 29779 18241 29788 18275
rect 29736 18232 29788 18241
rect 32864 18368 32916 18420
rect 31576 18300 31628 18352
rect 31852 18232 31904 18284
rect 32588 18232 32640 18284
rect 32956 18300 33008 18352
rect 23848 18071 23900 18080
rect 23848 18037 23857 18071
rect 23857 18037 23891 18071
rect 23891 18037 23900 18071
rect 23848 18028 23900 18037
rect 27804 18071 27856 18080
rect 27804 18037 27813 18071
rect 27813 18037 27847 18071
rect 27847 18037 27856 18071
rect 27804 18028 27856 18037
rect 28264 18028 28316 18080
rect 29368 18028 29420 18080
rect 32220 18028 32272 18080
rect 32864 18028 32916 18080
rect 5147 17926 5199 17978
rect 5211 17926 5263 17978
rect 5275 17926 5327 17978
rect 5339 17926 5391 17978
rect 5403 17926 5455 17978
rect 13541 17926 13593 17978
rect 13605 17926 13657 17978
rect 13669 17926 13721 17978
rect 13733 17926 13785 17978
rect 13797 17926 13849 17978
rect 21935 17926 21987 17978
rect 21999 17926 22051 17978
rect 22063 17926 22115 17978
rect 22127 17926 22179 17978
rect 22191 17926 22243 17978
rect 30329 17926 30381 17978
rect 30393 17926 30445 17978
rect 30457 17926 30509 17978
rect 30521 17926 30573 17978
rect 30585 17926 30637 17978
rect 3884 17824 3936 17876
rect 3976 17824 4028 17876
rect 3424 17756 3476 17808
rect 3608 17663 3660 17672
rect 3608 17629 3617 17663
rect 3617 17629 3651 17663
rect 3651 17629 3660 17663
rect 3608 17620 3660 17629
rect 3700 17620 3752 17672
rect 7380 17799 7432 17808
rect 7380 17765 7389 17799
rect 7389 17765 7423 17799
rect 7423 17765 7432 17799
rect 7380 17756 7432 17765
rect 4712 17688 4764 17740
rect 4804 17688 4856 17740
rect 3516 17552 3568 17604
rect 3792 17527 3844 17536
rect 3792 17493 3801 17527
rect 3801 17493 3835 17527
rect 3835 17493 3844 17527
rect 3792 17484 3844 17493
rect 4252 17552 4304 17604
rect 4528 17620 4580 17672
rect 5540 17688 5592 17740
rect 6920 17688 6972 17740
rect 5816 17620 5868 17672
rect 5908 17620 5960 17672
rect 6276 17620 6328 17672
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 7656 17552 7708 17604
rect 8116 17484 8168 17536
rect 9772 17824 9824 17876
rect 8944 17756 8996 17808
rect 8300 17688 8352 17740
rect 9128 17688 9180 17740
rect 14832 17867 14884 17876
rect 14832 17833 14841 17867
rect 14841 17833 14875 17867
rect 14875 17833 14884 17867
rect 14832 17824 14884 17833
rect 10324 17688 10376 17740
rect 12348 17688 12400 17740
rect 12716 17688 12768 17740
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 8852 17620 8904 17672
rect 8944 17663 8996 17672
rect 8944 17629 8953 17663
rect 8953 17629 8987 17663
rect 8987 17629 8996 17663
rect 8944 17620 8996 17629
rect 9036 17620 9088 17672
rect 9680 17663 9732 17672
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 10692 17620 10744 17629
rect 11336 17620 11388 17672
rect 11428 17663 11480 17672
rect 11428 17629 11437 17663
rect 11437 17629 11471 17663
rect 11471 17629 11480 17663
rect 11428 17620 11480 17629
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 11612 17663 11664 17672
rect 11612 17629 11621 17663
rect 11621 17629 11655 17663
rect 11655 17629 11664 17663
rect 11612 17620 11664 17629
rect 13360 17620 13412 17672
rect 13912 17663 13964 17672
rect 13912 17629 13921 17663
rect 13921 17629 13955 17663
rect 13955 17629 13964 17663
rect 13912 17620 13964 17629
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 14556 17620 14608 17629
rect 15476 17620 15528 17672
rect 16396 17756 16448 17808
rect 16948 17756 17000 17808
rect 17684 17756 17736 17808
rect 19340 17824 19392 17876
rect 20628 17824 20680 17876
rect 22284 17824 22336 17876
rect 22560 17867 22612 17876
rect 22560 17833 22569 17867
rect 22569 17833 22603 17867
rect 22603 17833 22612 17867
rect 22560 17824 22612 17833
rect 23204 17824 23256 17876
rect 19892 17756 19944 17808
rect 12072 17552 12124 17604
rect 16304 17620 16356 17672
rect 8760 17484 8812 17536
rect 9220 17484 9272 17536
rect 11152 17484 11204 17536
rect 13084 17484 13136 17536
rect 14648 17527 14700 17536
rect 14648 17493 14657 17527
rect 14657 17493 14691 17527
rect 14691 17493 14700 17527
rect 14648 17484 14700 17493
rect 16028 17484 16080 17536
rect 16948 17620 17000 17672
rect 18052 17663 18104 17672
rect 18052 17629 18061 17663
rect 18061 17629 18095 17663
rect 18095 17629 18104 17663
rect 18052 17620 18104 17629
rect 20168 17663 20220 17672
rect 20168 17629 20177 17663
rect 20177 17629 20211 17663
rect 20211 17629 20220 17663
rect 20168 17620 20220 17629
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 17592 17552 17644 17604
rect 20260 17552 20312 17604
rect 23572 17824 23624 17876
rect 23940 17824 23992 17876
rect 18144 17484 18196 17536
rect 18696 17484 18748 17536
rect 20996 17484 21048 17536
rect 21640 17663 21692 17672
rect 21640 17629 21649 17663
rect 21649 17629 21683 17663
rect 21683 17629 21692 17663
rect 21640 17620 21692 17629
rect 23480 17756 23532 17808
rect 24400 17867 24452 17876
rect 24400 17833 24409 17867
rect 24409 17833 24443 17867
rect 24443 17833 24452 17867
rect 24400 17824 24452 17833
rect 28540 17824 28592 17876
rect 28632 17824 28684 17876
rect 31484 17824 31536 17876
rect 32588 17867 32640 17876
rect 32588 17833 32597 17867
rect 32597 17833 32631 17867
rect 32631 17833 32640 17867
rect 32588 17824 32640 17833
rect 24768 17756 24820 17808
rect 26884 17756 26936 17808
rect 30012 17756 30064 17808
rect 30656 17756 30708 17808
rect 23480 17620 23532 17672
rect 23572 17663 23624 17672
rect 23572 17629 23581 17663
rect 23581 17629 23615 17663
rect 23615 17629 23624 17663
rect 23572 17620 23624 17629
rect 23848 17663 23900 17672
rect 23848 17629 23857 17663
rect 23857 17629 23891 17663
rect 23891 17629 23900 17663
rect 23848 17620 23900 17629
rect 27804 17688 27856 17740
rect 26608 17620 26660 17672
rect 27988 17663 28040 17672
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 28172 17663 28224 17672
rect 28172 17629 28181 17663
rect 28181 17629 28215 17663
rect 28215 17629 28224 17663
rect 28172 17620 28224 17629
rect 28264 17663 28316 17672
rect 28264 17629 28273 17663
rect 28273 17629 28307 17663
rect 28307 17629 28316 17663
rect 28264 17620 28316 17629
rect 22560 17484 22612 17536
rect 22928 17595 22980 17604
rect 22928 17561 22937 17595
rect 22937 17561 22971 17595
rect 22971 17561 22980 17595
rect 22928 17552 22980 17561
rect 23480 17527 23532 17536
rect 23480 17493 23489 17527
rect 23489 17493 23523 17527
rect 23523 17493 23532 17527
rect 23480 17484 23532 17493
rect 23664 17552 23716 17604
rect 27620 17552 27672 17604
rect 27896 17552 27948 17604
rect 28448 17620 28500 17672
rect 31116 17688 31168 17740
rect 31576 17688 31628 17740
rect 31852 17620 31904 17672
rect 32128 17663 32180 17672
rect 32128 17629 32137 17663
rect 32137 17629 32171 17663
rect 32171 17629 32180 17663
rect 32128 17620 32180 17629
rect 24860 17484 24912 17536
rect 26608 17527 26660 17536
rect 26608 17493 26617 17527
rect 26617 17493 26651 17527
rect 26651 17493 26660 17527
rect 26608 17484 26660 17493
rect 26700 17527 26752 17536
rect 26700 17493 26709 17527
rect 26709 17493 26743 17527
rect 26743 17493 26752 17527
rect 26700 17484 26752 17493
rect 29552 17484 29604 17536
rect 30932 17484 30984 17536
rect 32220 17484 32272 17536
rect 32496 17620 32548 17672
rect 32772 17552 32824 17604
rect 33508 17527 33560 17536
rect 33508 17493 33517 17527
rect 33517 17493 33551 17527
rect 33551 17493 33560 17527
rect 33508 17484 33560 17493
rect 9344 17382 9396 17434
rect 9408 17382 9460 17434
rect 9472 17382 9524 17434
rect 9536 17382 9588 17434
rect 9600 17382 9652 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 17930 17382 17982 17434
rect 17994 17382 18046 17434
rect 26132 17382 26184 17434
rect 26196 17382 26248 17434
rect 26260 17382 26312 17434
rect 26324 17382 26376 17434
rect 26388 17382 26440 17434
rect 34526 17382 34578 17434
rect 34590 17382 34642 17434
rect 34654 17382 34706 17434
rect 34718 17382 34770 17434
rect 34782 17382 34834 17434
rect 3424 17280 3476 17332
rect 3608 17280 3660 17332
rect 4252 17280 4304 17332
rect 2964 17144 3016 17196
rect 3516 17187 3568 17196
rect 3516 17153 3525 17187
rect 3525 17153 3559 17187
rect 3559 17153 3568 17187
rect 3516 17144 3568 17153
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 3700 17144 3752 17196
rect 5080 17212 5132 17264
rect 5724 17144 5776 17196
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 4804 17076 4856 17128
rect 3148 16983 3200 16992
rect 3148 16949 3157 16983
rect 3157 16949 3191 16983
rect 3191 16949 3200 16983
rect 3148 16940 3200 16949
rect 4988 16940 5040 16992
rect 9036 17280 9088 17332
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 7656 17187 7708 17196
rect 7656 17153 7665 17187
rect 7665 17153 7699 17187
rect 7699 17153 7708 17187
rect 7656 17144 7708 17153
rect 7748 17144 7800 17196
rect 8300 17144 8352 17196
rect 9680 17212 9732 17264
rect 9772 17212 9824 17264
rect 7656 17008 7708 17060
rect 7748 16940 7800 16992
rect 8484 17008 8536 17060
rect 11520 17280 11572 17332
rect 11244 17212 11296 17264
rect 12440 17280 12492 17332
rect 9772 17076 9824 17128
rect 11612 17144 11664 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 8300 16940 8352 16992
rect 9128 16940 9180 16992
rect 9220 16940 9272 16992
rect 9680 16940 9732 16992
rect 10416 16940 10468 16992
rect 10876 16983 10928 16992
rect 10876 16949 10885 16983
rect 10885 16949 10919 16983
rect 10919 16949 10928 16983
rect 10876 16940 10928 16949
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 12348 17144 12400 17196
rect 14648 17280 14700 17332
rect 17500 17280 17552 17332
rect 18144 17280 18196 17332
rect 27988 17280 28040 17332
rect 11612 16940 11664 16992
rect 11980 16940 12032 16992
rect 12992 17144 13044 17196
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 13452 17144 13504 17196
rect 13544 17144 13596 17196
rect 17592 17255 17644 17264
rect 17592 17221 17601 17255
rect 17601 17221 17635 17255
rect 17635 17221 17644 17255
rect 17592 17212 17644 17221
rect 12532 17051 12584 17060
rect 12532 17017 12541 17051
rect 12541 17017 12575 17051
rect 12575 17017 12584 17051
rect 12532 17008 12584 17017
rect 12716 17008 12768 17060
rect 14924 17187 14976 17196
rect 14924 17153 14933 17187
rect 14933 17153 14967 17187
rect 14967 17153 14976 17187
rect 14924 17144 14976 17153
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 13912 17008 13964 17060
rect 18788 17212 18840 17264
rect 18512 17144 18564 17196
rect 18328 17076 18380 17128
rect 18696 17144 18748 17196
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 21640 17144 21692 17196
rect 29000 17280 29052 17332
rect 29552 17212 29604 17264
rect 19340 17076 19392 17128
rect 19984 17076 20036 17128
rect 22284 17076 22336 17128
rect 28816 17187 28868 17196
rect 28816 17153 28825 17187
rect 28825 17153 28859 17187
rect 28859 17153 28868 17187
rect 28816 17144 28868 17153
rect 28908 17144 28960 17196
rect 29276 17144 29328 17196
rect 31668 17280 31720 17332
rect 32680 17280 32732 17332
rect 33416 17280 33468 17332
rect 30932 17212 30984 17264
rect 31024 17187 31076 17196
rect 31024 17153 31033 17187
rect 31033 17153 31067 17187
rect 31067 17153 31076 17187
rect 31024 17144 31076 17153
rect 31116 17187 31168 17196
rect 31116 17153 31125 17187
rect 31125 17153 31159 17187
rect 31159 17153 31168 17187
rect 31116 17144 31168 17153
rect 31208 17144 31260 17196
rect 31576 17144 31628 17196
rect 32772 17144 32824 17196
rect 32956 17187 33008 17196
rect 32956 17153 32965 17187
rect 32965 17153 32999 17187
rect 32999 17153 33008 17187
rect 32956 17144 33008 17153
rect 33140 17187 33192 17196
rect 33140 17153 33149 17187
rect 33149 17153 33183 17187
rect 33183 17153 33192 17187
rect 33140 17144 33192 17153
rect 33692 17187 33744 17196
rect 33692 17153 33701 17187
rect 33701 17153 33735 17187
rect 33735 17153 33744 17187
rect 33692 17144 33744 17153
rect 27620 17008 27672 17060
rect 30932 17008 30984 17060
rect 14188 16940 14240 16992
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 15660 16983 15712 16992
rect 15660 16949 15669 16983
rect 15669 16949 15703 16983
rect 15703 16949 15712 16983
rect 15660 16940 15712 16949
rect 18144 16940 18196 16992
rect 18420 16940 18472 16992
rect 21180 16983 21232 16992
rect 21180 16949 21189 16983
rect 21189 16949 21223 16983
rect 21223 16949 21232 16983
rect 21180 16940 21232 16949
rect 30656 16940 30708 16992
rect 5147 16838 5199 16890
rect 5211 16838 5263 16890
rect 5275 16838 5327 16890
rect 5339 16838 5391 16890
rect 5403 16838 5455 16890
rect 13541 16838 13593 16890
rect 13605 16838 13657 16890
rect 13669 16838 13721 16890
rect 13733 16838 13785 16890
rect 13797 16838 13849 16890
rect 21935 16838 21987 16890
rect 21999 16838 22051 16890
rect 22063 16838 22115 16890
rect 22127 16838 22179 16890
rect 22191 16838 22243 16890
rect 30329 16838 30381 16890
rect 30393 16838 30445 16890
rect 30457 16838 30509 16890
rect 30521 16838 30573 16890
rect 30585 16838 30637 16890
rect 3976 16736 4028 16788
rect 5632 16779 5684 16788
rect 5632 16745 5656 16779
rect 5656 16745 5684 16779
rect 5632 16736 5684 16745
rect 5816 16736 5868 16788
rect 3148 16532 3200 16584
rect 4068 16600 4120 16652
rect 7840 16736 7892 16788
rect 9772 16736 9824 16788
rect 13912 16779 13964 16788
rect 13912 16745 13921 16779
rect 13921 16745 13955 16779
rect 13955 16745 13964 16779
rect 13912 16736 13964 16745
rect 15108 16736 15160 16788
rect 15384 16736 15436 16788
rect 15752 16736 15804 16788
rect 16028 16736 16080 16788
rect 21180 16736 21232 16788
rect 22744 16736 22796 16788
rect 23664 16736 23716 16788
rect 24768 16736 24820 16788
rect 26700 16736 26752 16788
rect 27620 16779 27672 16788
rect 27620 16745 27629 16779
rect 27629 16745 27663 16779
rect 27663 16745 27672 16779
rect 27620 16736 27672 16745
rect 29276 16779 29328 16788
rect 29276 16745 29285 16779
rect 29285 16745 29319 16779
rect 29319 16745 29328 16779
rect 29276 16736 29328 16745
rect 31024 16736 31076 16788
rect 31208 16736 31260 16788
rect 31300 16779 31352 16788
rect 31300 16745 31309 16779
rect 31309 16745 31343 16779
rect 31343 16745 31352 16779
rect 31300 16736 31352 16745
rect 33140 16736 33192 16788
rect 33508 16736 33560 16788
rect 33692 16736 33744 16788
rect 10876 16668 10928 16720
rect 11888 16668 11940 16720
rect 5540 16532 5592 16584
rect 6000 16532 6052 16584
rect 6276 16575 6328 16584
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 3056 16507 3108 16516
rect 3056 16473 3065 16507
rect 3065 16473 3099 16507
rect 3099 16473 3108 16507
rect 3056 16464 3108 16473
rect 3884 16464 3936 16516
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 6828 16575 6880 16584
rect 6828 16541 6837 16575
rect 6837 16541 6871 16575
rect 6871 16541 6880 16575
rect 6828 16532 6880 16541
rect 8668 16600 8720 16652
rect 12440 16600 12492 16652
rect 13544 16600 13596 16652
rect 15292 16600 15344 16652
rect 20168 16668 20220 16720
rect 7380 16532 7432 16584
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 7748 16575 7800 16584
rect 7748 16541 7757 16575
rect 7757 16541 7791 16575
rect 7791 16541 7800 16575
rect 7748 16532 7800 16541
rect 7840 16575 7892 16584
rect 7840 16541 7849 16575
rect 7849 16541 7883 16575
rect 7883 16541 7892 16575
rect 7840 16532 7892 16541
rect 7564 16464 7616 16516
rect 9404 16532 9456 16584
rect 9680 16532 9732 16584
rect 9312 16464 9364 16516
rect 11244 16532 11296 16584
rect 12256 16532 12308 16584
rect 13360 16507 13412 16516
rect 13360 16473 13369 16507
rect 13369 16473 13403 16507
rect 13403 16473 13412 16507
rect 13360 16464 13412 16473
rect 9772 16396 9824 16448
rect 10692 16396 10744 16448
rect 13544 16464 13596 16516
rect 14372 16532 14424 16584
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 15200 16532 15252 16584
rect 15476 16532 15528 16584
rect 15844 16532 15896 16584
rect 19892 16600 19944 16652
rect 16120 16575 16172 16584
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 16120 16532 16172 16541
rect 18144 16532 18196 16584
rect 18236 16532 18288 16584
rect 24860 16643 24912 16652
rect 24860 16609 24869 16643
rect 24869 16609 24903 16643
rect 24903 16609 24912 16643
rect 24860 16600 24912 16609
rect 26884 16600 26936 16652
rect 30656 16600 30708 16652
rect 20260 16575 20312 16584
rect 20260 16541 20269 16575
rect 20269 16541 20303 16575
rect 20303 16541 20312 16575
rect 20260 16532 20312 16541
rect 20444 16575 20496 16584
rect 20444 16541 20453 16575
rect 20453 16541 20487 16575
rect 20487 16541 20496 16575
rect 20444 16532 20496 16541
rect 21640 16575 21692 16584
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 22928 16532 22980 16584
rect 28264 16575 28316 16584
rect 28264 16541 28273 16575
rect 28273 16541 28307 16575
rect 28307 16541 28316 16575
rect 28264 16532 28316 16541
rect 14280 16396 14332 16448
rect 15568 16464 15620 16516
rect 24124 16464 24176 16516
rect 26792 16464 26844 16516
rect 30932 16575 30984 16584
rect 30932 16541 30941 16575
rect 30941 16541 30975 16575
rect 30975 16541 30984 16575
rect 30932 16532 30984 16541
rect 31024 16575 31076 16584
rect 31024 16541 31033 16575
rect 31033 16541 31067 16575
rect 31067 16541 31076 16575
rect 31024 16532 31076 16541
rect 33140 16532 33192 16584
rect 32772 16464 32824 16516
rect 15384 16396 15436 16448
rect 15660 16396 15712 16448
rect 18420 16396 18472 16448
rect 24400 16439 24452 16448
rect 24400 16405 24409 16439
rect 24409 16405 24443 16439
rect 24443 16405 24452 16439
rect 24400 16396 24452 16405
rect 24768 16439 24820 16448
rect 24768 16405 24777 16439
rect 24777 16405 24811 16439
rect 24811 16405 24820 16439
rect 24768 16396 24820 16405
rect 27712 16439 27764 16448
rect 27712 16405 27721 16439
rect 27721 16405 27755 16439
rect 27755 16405 27764 16439
rect 27712 16396 27764 16405
rect 28908 16396 28960 16448
rect 31392 16396 31444 16448
rect 31852 16396 31904 16448
rect 32588 16396 32640 16448
rect 32956 16396 33008 16448
rect 9344 16294 9396 16346
rect 9408 16294 9460 16346
rect 9472 16294 9524 16346
rect 9536 16294 9588 16346
rect 9600 16294 9652 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 17930 16294 17982 16346
rect 17994 16294 18046 16346
rect 26132 16294 26184 16346
rect 26196 16294 26248 16346
rect 26260 16294 26312 16346
rect 26324 16294 26376 16346
rect 26388 16294 26440 16346
rect 34526 16294 34578 16346
rect 34590 16294 34642 16346
rect 34654 16294 34706 16346
rect 34718 16294 34770 16346
rect 34782 16294 34834 16346
rect 3608 16192 3660 16244
rect 4804 16235 4856 16244
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 5172 16192 5224 16244
rect 7932 16192 7984 16244
rect 8208 16192 8260 16244
rect 8300 16192 8352 16244
rect 4620 16124 4672 16176
rect 8576 16235 8628 16244
rect 8576 16201 8585 16235
rect 8585 16201 8619 16235
rect 8619 16201 8628 16235
rect 8576 16192 8628 16201
rect 9128 16192 9180 16244
rect 11152 16192 11204 16244
rect 12532 16192 12584 16244
rect 18420 16192 18472 16244
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 22284 16192 22336 16244
rect 23204 16192 23256 16244
rect 1492 16056 1544 16108
rect 4068 16056 4120 16108
rect 4712 16099 4764 16108
rect 3056 15988 3108 16040
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 4712 16056 4764 16065
rect 4804 15988 4856 16040
rect 5448 16056 5500 16108
rect 8300 16056 8352 16108
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 9864 16099 9916 16108
rect 9864 16065 9873 16099
rect 9873 16065 9907 16099
rect 9907 16065 9916 16099
rect 9864 16056 9916 16065
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 11336 16056 11388 16108
rect 12808 16056 12860 16108
rect 8852 15988 8904 16040
rect 10416 15988 10468 16040
rect 11888 15988 11940 16040
rect 15016 16056 15068 16108
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 15384 16099 15436 16108
rect 15384 16065 15393 16099
rect 15393 16065 15427 16099
rect 15427 16065 15436 16099
rect 15384 16056 15436 16065
rect 22744 16124 22796 16176
rect 23756 16192 23808 16244
rect 24400 16192 24452 16244
rect 24768 16192 24820 16244
rect 26792 16235 26844 16244
rect 26792 16201 26801 16235
rect 26801 16201 26835 16235
rect 26835 16201 26844 16235
rect 26792 16192 26844 16201
rect 15568 16056 15620 16108
rect 16212 16056 16264 16108
rect 19616 16056 19668 16108
rect 22928 16056 22980 16108
rect 15752 15988 15804 16040
rect 18236 16031 18288 16040
rect 18236 15997 18245 16031
rect 18245 15997 18279 16031
rect 18279 15997 18288 16031
rect 18236 15988 18288 15997
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 22744 15988 22796 16040
rect 1952 15920 2004 15972
rect 6920 15920 6972 15972
rect 8024 15920 8076 15972
rect 8116 15920 8168 15972
rect 10784 15920 10836 15972
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6092 15852 6144 15904
rect 6368 15852 6420 15904
rect 11704 15920 11756 15972
rect 13268 15920 13320 15972
rect 13544 15920 13596 15972
rect 22652 15920 22704 15972
rect 23112 16099 23164 16108
rect 23112 16065 23121 16099
rect 23121 16065 23155 16099
rect 23155 16065 23164 16099
rect 23112 16056 23164 16065
rect 23296 16056 23348 16108
rect 26700 16124 26752 16176
rect 27712 16192 27764 16244
rect 30012 16192 30064 16244
rect 28172 16124 28224 16176
rect 24124 16099 24176 16108
rect 24124 16065 24133 16099
rect 24133 16065 24167 16099
rect 24167 16065 24176 16099
rect 24124 16056 24176 16065
rect 32588 16192 32640 16244
rect 23480 15920 23532 15972
rect 25596 15988 25648 16040
rect 26884 16056 26936 16108
rect 29000 16056 29052 16108
rect 29368 16056 29420 16108
rect 32864 16167 32916 16176
rect 32864 16133 32873 16167
rect 32873 16133 32907 16167
rect 32907 16133 32916 16167
rect 32864 16124 32916 16133
rect 27436 15988 27488 16040
rect 28172 15988 28224 16040
rect 13084 15852 13136 15904
rect 15384 15852 15436 15904
rect 20260 15852 20312 15904
rect 23296 15852 23348 15904
rect 28172 15852 28224 15904
rect 28908 15895 28960 15904
rect 28908 15861 28917 15895
rect 28917 15861 28951 15895
rect 28951 15861 28960 15895
rect 28908 15852 28960 15861
rect 29460 15895 29512 15904
rect 29460 15861 29469 15895
rect 29469 15861 29503 15895
rect 29503 15861 29512 15895
rect 29460 15852 29512 15861
rect 31024 16056 31076 16108
rect 31392 16056 31444 16108
rect 32220 16056 32272 16108
rect 31024 15920 31076 15972
rect 32772 15920 32824 15972
rect 32956 15852 33008 15904
rect 5147 15750 5199 15802
rect 5211 15750 5263 15802
rect 5275 15750 5327 15802
rect 5339 15750 5391 15802
rect 5403 15750 5455 15802
rect 13541 15750 13593 15802
rect 13605 15750 13657 15802
rect 13669 15750 13721 15802
rect 13733 15750 13785 15802
rect 13797 15750 13849 15802
rect 21935 15750 21987 15802
rect 21999 15750 22051 15802
rect 22063 15750 22115 15802
rect 22127 15750 22179 15802
rect 22191 15750 22243 15802
rect 30329 15750 30381 15802
rect 30393 15750 30445 15802
rect 30457 15750 30509 15802
rect 30521 15750 30573 15802
rect 30585 15750 30637 15802
rect 3792 15648 3844 15700
rect 6368 15648 6420 15700
rect 1400 15512 1452 15564
rect 6828 15580 6880 15632
rect 7564 15648 7616 15700
rect 8024 15648 8076 15700
rect 8576 15691 8628 15700
rect 8576 15657 8585 15691
rect 8585 15657 8619 15691
rect 8619 15657 8628 15691
rect 8576 15648 8628 15657
rect 6276 15512 6328 15564
rect 7380 15512 7432 15564
rect 1492 15487 1544 15496
rect 1492 15453 1501 15487
rect 1501 15453 1535 15487
rect 1535 15453 1544 15487
rect 1492 15444 1544 15453
rect 5632 15444 5684 15496
rect 2964 15376 3016 15428
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6092 15308 6144 15360
rect 8392 15580 8444 15632
rect 8944 15580 8996 15632
rect 7564 15376 7616 15428
rect 8024 15487 8076 15496
rect 8024 15453 8034 15487
rect 8034 15453 8068 15487
rect 8068 15453 8076 15487
rect 8024 15444 8076 15453
rect 8116 15444 8168 15496
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 10048 15648 10100 15700
rect 10508 15648 10560 15700
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 13268 15691 13320 15700
rect 13268 15657 13277 15691
rect 13277 15657 13311 15691
rect 13311 15657 13320 15691
rect 13268 15648 13320 15657
rect 15200 15648 15252 15700
rect 15844 15648 15896 15700
rect 10692 15555 10744 15564
rect 10692 15521 10701 15555
rect 10701 15521 10735 15555
rect 10735 15521 10744 15555
rect 10692 15512 10744 15521
rect 11520 15580 11572 15632
rect 12072 15580 12124 15632
rect 9588 15487 9640 15496
rect 9588 15453 9597 15487
rect 9597 15453 9631 15487
rect 9631 15453 9640 15487
rect 9588 15444 9640 15453
rect 9864 15444 9916 15496
rect 10784 15444 10836 15496
rect 10876 15487 10928 15496
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 11152 15444 11204 15496
rect 11796 15512 11848 15564
rect 15108 15580 15160 15632
rect 16304 15580 16356 15632
rect 8208 15419 8260 15428
rect 8208 15385 8217 15419
rect 8217 15385 8251 15419
rect 8251 15385 8260 15419
rect 8208 15376 8260 15385
rect 7748 15308 7800 15360
rect 7932 15308 7984 15360
rect 9680 15376 9732 15428
rect 10692 15376 10744 15428
rect 12164 15419 12216 15428
rect 12164 15385 12173 15419
rect 12173 15385 12207 15419
rect 12207 15385 12216 15419
rect 12164 15376 12216 15385
rect 8944 15308 8996 15360
rect 9588 15308 9640 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 10048 15308 10100 15360
rect 10876 15308 10928 15360
rect 11888 15308 11940 15360
rect 12992 15419 13044 15428
rect 12992 15385 13001 15419
rect 13001 15385 13035 15419
rect 13035 15385 13044 15419
rect 12992 15376 13044 15385
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 16028 15444 16080 15496
rect 16672 15487 16724 15496
rect 16672 15453 16681 15487
rect 16681 15453 16715 15487
rect 16715 15453 16724 15487
rect 16672 15444 16724 15453
rect 19432 15512 19484 15564
rect 20904 15648 20956 15700
rect 21640 15648 21692 15700
rect 22928 15691 22980 15700
rect 22928 15657 22937 15691
rect 22937 15657 22971 15691
rect 22971 15657 22980 15691
rect 22928 15648 22980 15657
rect 26792 15648 26844 15700
rect 22744 15580 22796 15632
rect 23480 15580 23532 15632
rect 22284 15512 22336 15564
rect 23296 15512 23348 15564
rect 13176 15308 13228 15360
rect 19248 15376 19300 15428
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 20168 15444 20220 15496
rect 20628 15444 20680 15496
rect 20444 15376 20496 15428
rect 20996 15376 21048 15428
rect 21640 15487 21692 15496
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 21732 15487 21784 15496
rect 21732 15453 21741 15487
rect 21741 15453 21775 15487
rect 21775 15453 21784 15487
rect 21732 15444 21784 15453
rect 24124 15512 24176 15564
rect 22008 15419 22060 15428
rect 22008 15385 22017 15419
rect 22017 15385 22051 15419
rect 22051 15385 22060 15419
rect 22008 15376 22060 15385
rect 16488 15308 16540 15360
rect 18144 15308 18196 15360
rect 19524 15308 19576 15360
rect 19984 15308 20036 15360
rect 20352 15308 20404 15360
rect 22284 15376 22336 15428
rect 22836 15376 22888 15428
rect 22928 15308 22980 15360
rect 23204 15419 23256 15428
rect 23204 15385 23213 15419
rect 23213 15385 23247 15419
rect 23247 15385 23256 15419
rect 23204 15376 23256 15385
rect 23296 15376 23348 15428
rect 25504 15487 25556 15496
rect 25504 15453 25513 15487
rect 25513 15453 25547 15487
rect 25547 15453 25556 15487
rect 25504 15444 25556 15453
rect 28264 15648 28316 15700
rect 29460 15648 29512 15700
rect 27896 15580 27948 15632
rect 28080 15580 28132 15632
rect 28172 15555 28224 15564
rect 28172 15521 28181 15555
rect 28181 15521 28215 15555
rect 28215 15521 28224 15555
rect 28172 15512 28224 15521
rect 29552 15487 29604 15496
rect 29552 15453 29561 15487
rect 29561 15453 29595 15487
rect 29595 15453 29604 15487
rect 29552 15444 29604 15453
rect 29736 15648 29788 15700
rect 31392 15648 31444 15700
rect 31024 15580 31076 15632
rect 24952 15308 25004 15360
rect 27436 15376 27488 15428
rect 27528 15351 27580 15360
rect 27528 15317 27537 15351
rect 27537 15317 27571 15351
rect 27571 15317 27580 15351
rect 27528 15308 27580 15317
rect 29000 15308 29052 15360
rect 31944 15308 31996 15360
rect 33416 15308 33468 15360
rect 9344 15206 9396 15258
rect 9408 15206 9460 15258
rect 9472 15206 9524 15258
rect 9536 15206 9588 15258
rect 9600 15206 9652 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 17930 15206 17982 15258
rect 17994 15206 18046 15258
rect 26132 15206 26184 15258
rect 26196 15206 26248 15258
rect 26260 15206 26312 15258
rect 26324 15206 26376 15258
rect 26388 15206 26440 15258
rect 34526 15206 34578 15258
rect 34590 15206 34642 15258
rect 34654 15206 34706 15258
rect 34718 15206 34770 15258
rect 34782 15206 34834 15258
rect 4804 15104 4856 15156
rect 5816 15104 5868 15156
rect 6920 15147 6972 15156
rect 6920 15113 6929 15147
rect 6929 15113 6963 15147
rect 6963 15113 6972 15147
rect 6920 15104 6972 15113
rect 7104 15104 7156 15156
rect 7840 15104 7892 15156
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 10784 15104 10836 15156
rect 12624 15104 12676 15156
rect 13084 15104 13136 15156
rect 3056 14968 3108 15020
rect 3332 15011 3384 15020
rect 3332 14977 3341 15011
rect 3341 14977 3375 15011
rect 3375 14977 3384 15011
rect 3332 14968 3384 14977
rect 3976 14968 4028 15020
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 4528 15036 4580 15088
rect 6828 15036 6880 15088
rect 5540 14968 5592 15020
rect 4344 14832 4396 14884
rect 4712 14832 4764 14884
rect 5540 14832 5592 14884
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 7472 14968 7524 15020
rect 8668 14968 8720 15020
rect 8944 14968 8996 15020
rect 9680 14968 9732 15020
rect 10416 14968 10468 15020
rect 11888 14968 11940 15020
rect 11980 14968 12032 15020
rect 12348 14968 12400 15020
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 7288 14900 7340 14952
rect 8024 14900 8076 14952
rect 9036 14900 9088 14952
rect 9772 14900 9824 14952
rect 9864 14900 9916 14952
rect 13912 14968 13964 15020
rect 14096 14968 14148 15020
rect 16488 15079 16540 15088
rect 16488 15045 16497 15079
rect 16497 15045 16531 15079
rect 16531 15045 16540 15079
rect 16488 15036 16540 15045
rect 19248 15104 19300 15156
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 16028 14968 16080 15020
rect 16304 15011 16356 15020
rect 16304 14977 16313 15011
rect 16313 14977 16347 15011
rect 16347 14977 16356 15011
rect 16856 15011 16908 15020
rect 16304 14968 16356 14977
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 3884 14764 3936 14816
rect 11796 14832 11848 14884
rect 13084 14832 13136 14884
rect 16580 14900 16632 14952
rect 18144 14968 18196 15020
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 20168 15104 20220 15156
rect 20352 15104 20404 15156
rect 19524 15036 19576 15088
rect 14096 14875 14148 14884
rect 14096 14841 14105 14875
rect 14105 14841 14139 14875
rect 14139 14841 14148 14875
rect 14096 14832 14148 14841
rect 14740 14832 14792 14884
rect 5724 14764 5776 14816
rect 7104 14764 7156 14816
rect 8944 14764 8996 14816
rect 10324 14764 10376 14816
rect 11428 14764 11480 14816
rect 13452 14764 13504 14816
rect 15108 14764 15160 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 16304 14832 16356 14884
rect 17132 14900 17184 14952
rect 19708 15011 19760 15020
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 21732 15104 21784 15156
rect 24952 15104 25004 15156
rect 25504 15104 25556 15156
rect 27528 15104 27580 15156
rect 22744 15036 22796 15088
rect 20536 14968 20588 15020
rect 20812 14968 20864 15020
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 22836 14968 22888 15020
rect 23020 15011 23072 15020
rect 23020 14977 23029 15011
rect 23029 14977 23063 15011
rect 23063 14977 23072 15011
rect 23020 14968 23072 14977
rect 23296 14968 23348 15020
rect 28080 15036 28132 15088
rect 30104 15036 30156 15088
rect 30932 15036 30984 15088
rect 31576 15036 31628 15088
rect 33416 15036 33468 15088
rect 29368 14968 29420 15020
rect 31208 15011 31260 15020
rect 31208 14977 31217 15011
rect 31217 14977 31251 15011
rect 31251 14977 31260 15011
rect 31208 14968 31260 14977
rect 31668 15011 31720 15020
rect 31668 14977 31677 15011
rect 31677 14977 31711 15011
rect 31711 14977 31720 15011
rect 31668 14968 31720 14977
rect 32864 14968 32916 15020
rect 17592 14832 17644 14884
rect 19340 14900 19392 14952
rect 21548 14900 21600 14952
rect 18420 14875 18472 14884
rect 18420 14841 18429 14875
rect 18429 14841 18463 14875
rect 18463 14841 18472 14875
rect 18420 14832 18472 14841
rect 19156 14832 19208 14884
rect 20076 14875 20128 14884
rect 20076 14841 20085 14875
rect 20085 14841 20119 14875
rect 20119 14841 20128 14875
rect 20076 14832 20128 14841
rect 20720 14832 20772 14884
rect 22928 14900 22980 14952
rect 25964 14900 26016 14952
rect 27344 14900 27396 14952
rect 30748 14900 30800 14952
rect 31852 14943 31904 14952
rect 31852 14909 31861 14943
rect 31861 14909 31895 14943
rect 31895 14909 31904 14943
rect 31852 14900 31904 14909
rect 28632 14807 28684 14816
rect 28632 14773 28641 14807
rect 28641 14773 28675 14807
rect 28675 14773 28684 14807
rect 28632 14764 28684 14773
rect 31300 14764 31352 14816
rect 31484 14807 31536 14816
rect 31484 14773 31493 14807
rect 31493 14773 31527 14807
rect 31527 14773 31536 14807
rect 31484 14764 31536 14773
rect 31852 14807 31904 14816
rect 31852 14773 31861 14807
rect 31861 14773 31895 14807
rect 31895 14773 31904 14807
rect 31852 14764 31904 14773
rect 34152 14807 34204 14816
rect 34152 14773 34161 14807
rect 34161 14773 34195 14807
rect 34195 14773 34204 14807
rect 34152 14764 34204 14773
rect 5147 14662 5199 14714
rect 5211 14662 5263 14714
rect 5275 14662 5327 14714
rect 5339 14662 5391 14714
rect 5403 14662 5455 14714
rect 13541 14662 13593 14714
rect 13605 14662 13657 14714
rect 13669 14662 13721 14714
rect 13733 14662 13785 14714
rect 13797 14662 13849 14714
rect 21935 14662 21987 14714
rect 21999 14662 22051 14714
rect 22063 14662 22115 14714
rect 22127 14662 22179 14714
rect 22191 14662 22243 14714
rect 30329 14662 30381 14714
rect 30393 14662 30445 14714
rect 30457 14662 30509 14714
rect 30521 14662 30573 14714
rect 30585 14662 30637 14714
rect 7012 14603 7064 14612
rect 7012 14569 7021 14603
rect 7021 14569 7055 14603
rect 7055 14569 7064 14603
rect 7012 14560 7064 14569
rect 8852 14560 8904 14612
rect 10324 14560 10376 14612
rect 10968 14560 11020 14612
rect 12532 14560 12584 14612
rect 14096 14560 14148 14612
rect 15108 14560 15160 14612
rect 15200 14603 15252 14612
rect 15200 14569 15209 14603
rect 15209 14569 15243 14603
rect 15243 14569 15252 14603
rect 15200 14560 15252 14569
rect 16856 14560 16908 14612
rect 17132 14560 17184 14612
rect 18328 14560 18380 14612
rect 19340 14560 19392 14612
rect 19984 14603 20036 14612
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 21088 14560 21140 14612
rect 3792 14492 3844 14544
rect 4252 14492 4304 14544
rect 6184 14492 6236 14544
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 4804 14356 4856 14408
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 7564 14492 7616 14544
rect 9864 14492 9916 14544
rect 7748 14424 7800 14476
rect 13084 14492 13136 14544
rect 11152 14424 11204 14476
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 7564 14356 7616 14408
rect 9128 14356 9180 14408
rect 9956 14356 10008 14408
rect 11060 14356 11112 14408
rect 4528 14263 4580 14272
rect 4528 14229 4537 14263
rect 4537 14229 4571 14263
rect 4571 14229 4580 14263
rect 4528 14220 4580 14229
rect 4896 14220 4948 14272
rect 5448 14220 5500 14272
rect 5540 14220 5592 14272
rect 5816 14220 5868 14272
rect 8116 14288 8168 14340
rect 8392 14288 8444 14340
rect 7012 14220 7064 14272
rect 7196 14220 7248 14272
rect 9128 14220 9180 14272
rect 10232 14220 10284 14272
rect 11244 14356 11296 14408
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 12440 14356 12492 14408
rect 12532 14356 12584 14408
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 16028 14424 16080 14476
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 11336 14220 11388 14272
rect 12072 14220 12124 14272
rect 13452 14356 13504 14408
rect 13636 14288 13688 14340
rect 14280 14356 14332 14408
rect 15384 14399 15436 14408
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 15568 14356 15620 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 16856 14424 16908 14476
rect 13360 14220 13412 14272
rect 14096 14220 14148 14272
rect 15936 14220 15988 14272
rect 16304 14356 16356 14408
rect 18144 14399 18196 14408
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 17592 14288 17644 14340
rect 19156 14288 19208 14340
rect 20628 14467 20680 14476
rect 20628 14433 20637 14467
rect 20637 14433 20671 14467
rect 20671 14433 20680 14467
rect 20628 14424 20680 14433
rect 19432 14356 19484 14408
rect 19708 14356 19760 14408
rect 20352 14399 20404 14408
rect 20352 14365 20361 14399
rect 20361 14365 20395 14399
rect 20395 14365 20404 14399
rect 20352 14356 20404 14365
rect 20260 14288 20312 14340
rect 21180 14492 21232 14544
rect 21824 14424 21876 14476
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 23020 14424 23072 14476
rect 21640 14288 21692 14340
rect 22744 14399 22796 14408
rect 22744 14365 22753 14399
rect 22753 14365 22787 14399
rect 22787 14365 22796 14399
rect 22744 14356 22796 14365
rect 22928 14399 22980 14408
rect 22928 14365 22937 14399
rect 22937 14365 22971 14399
rect 22971 14365 22980 14399
rect 22928 14356 22980 14365
rect 23296 14399 23348 14408
rect 23296 14365 23305 14399
rect 23305 14365 23339 14399
rect 23339 14365 23348 14399
rect 23296 14356 23348 14365
rect 29368 14603 29420 14612
rect 29368 14569 29377 14603
rect 29377 14569 29411 14603
rect 29411 14569 29420 14603
rect 29368 14560 29420 14569
rect 32220 14560 32272 14612
rect 25964 14467 26016 14476
rect 25964 14433 25973 14467
rect 25973 14433 26007 14467
rect 26007 14433 26016 14467
rect 25964 14424 26016 14433
rect 26884 14492 26936 14544
rect 31944 14492 31996 14544
rect 27620 14467 27672 14476
rect 27620 14433 27629 14467
rect 27629 14433 27663 14467
rect 27663 14433 27672 14467
rect 27620 14424 27672 14433
rect 25688 14356 25740 14408
rect 31392 14356 31444 14408
rect 34704 14492 34756 14544
rect 27528 14331 27580 14340
rect 18420 14220 18472 14272
rect 19892 14220 19944 14272
rect 20536 14220 20588 14272
rect 20812 14220 20864 14272
rect 22560 14220 22612 14272
rect 27528 14297 27537 14331
rect 27537 14297 27571 14331
rect 27571 14297 27580 14331
rect 27528 14288 27580 14297
rect 27896 14331 27948 14340
rect 27896 14297 27905 14331
rect 27905 14297 27939 14331
rect 27939 14297 27948 14331
rect 27896 14288 27948 14297
rect 29368 14288 29420 14340
rect 31116 14288 31168 14340
rect 26056 14220 26108 14272
rect 26516 14220 26568 14272
rect 26608 14263 26660 14272
rect 26608 14229 26617 14263
rect 26617 14229 26651 14263
rect 26651 14229 26660 14263
rect 26608 14220 26660 14229
rect 31576 14263 31628 14272
rect 31576 14229 31585 14263
rect 31585 14229 31619 14263
rect 31619 14229 31628 14263
rect 31576 14220 31628 14229
rect 31852 14331 31904 14340
rect 31852 14297 31861 14331
rect 31861 14297 31895 14331
rect 31895 14297 31904 14331
rect 31852 14288 31904 14297
rect 31944 14331 31996 14340
rect 31944 14297 31953 14331
rect 31953 14297 31987 14331
rect 31987 14297 31996 14331
rect 31944 14288 31996 14297
rect 32864 14356 32916 14408
rect 34152 14356 34204 14408
rect 32220 14220 32272 14272
rect 32312 14263 32364 14272
rect 32312 14229 32321 14263
rect 32321 14229 32355 14263
rect 32355 14229 32364 14263
rect 32312 14220 32364 14229
rect 9344 14118 9396 14170
rect 9408 14118 9460 14170
rect 9472 14118 9524 14170
rect 9536 14118 9588 14170
rect 9600 14118 9652 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 17930 14118 17982 14170
rect 17994 14118 18046 14170
rect 26132 14118 26184 14170
rect 26196 14118 26248 14170
rect 26260 14118 26312 14170
rect 26324 14118 26376 14170
rect 26388 14118 26440 14170
rect 34526 14118 34578 14170
rect 34590 14118 34642 14170
rect 34654 14118 34706 14170
rect 34718 14118 34770 14170
rect 34782 14118 34834 14170
rect 3976 14016 4028 14068
rect 4620 14016 4672 14068
rect 5448 14059 5500 14068
rect 5448 14025 5457 14059
rect 5457 14025 5491 14059
rect 5491 14025 5500 14059
rect 5448 14016 5500 14025
rect 3884 13948 3936 14000
rect 3332 13880 3384 13932
rect 3608 13880 3660 13932
rect 3792 13812 3844 13864
rect 4620 13923 4672 13932
rect 4620 13889 4629 13923
rect 4629 13889 4663 13923
rect 4663 13889 4672 13923
rect 4620 13880 4672 13889
rect 4712 13880 4764 13932
rect 5816 13948 5868 14000
rect 5724 13880 5776 13932
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 7288 14016 7340 14068
rect 7380 14016 7432 14068
rect 9864 14016 9916 14068
rect 10416 14016 10468 14068
rect 6552 13948 6604 14000
rect 7012 13948 7064 14000
rect 4344 13676 4396 13728
rect 5080 13676 5132 13728
rect 6092 13812 6144 13864
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 5356 13676 5408 13728
rect 6000 13676 6052 13728
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 8668 13855 8720 13864
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 9496 13880 9548 13932
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 9680 13880 9732 13889
rect 9772 13923 9824 13932
rect 9772 13889 9781 13923
rect 9781 13889 9815 13923
rect 9815 13889 9824 13923
rect 9772 13880 9824 13889
rect 9864 13880 9916 13932
rect 10232 13948 10284 14000
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 9220 13855 9272 13864
rect 9220 13821 9229 13855
rect 9229 13821 9263 13855
rect 9263 13821 9272 13855
rect 9220 13812 9272 13821
rect 9404 13744 9456 13796
rect 9864 13787 9916 13796
rect 9864 13753 9873 13787
rect 9873 13753 9907 13787
rect 9907 13753 9916 13787
rect 9864 13744 9916 13753
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 11612 14016 11664 14068
rect 13084 14016 13136 14068
rect 13176 14016 13228 14068
rect 16672 14016 16724 14068
rect 12992 13880 13044 13932
rect 13360 13948 13412 14000
rect 13636 13948 13688 14000
rect 15384 13948 15436 14000
rect 12164 13744 12216 13796
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 12716 13744 12768 13796
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 13912 13880 13964 13932
rect 14188 13880 14240 13932
rect 15292 13880 15344 13932
rect 15752 13880 15804 13932
rect 16028 13923 16080 13932
rect 16028 13889 16037 13923
rect 16037 13889 16071 13923
rect 16071 13889 16080 13923
rect 16028 13880 16080 13889
rect 18144 13948 18196 14000
rect 20720 14016 20772 14068
rect 24124 14016 24176 14068
rect 25688 14059 25740 14068
rect 25688 14025 25697 14059
rect 25697 14025 25731 14059
rect 25731 14025 25740 14059
rect 25688 14016 25740 14025
rect 26608 14016 26660 14068
rect 18328 13880 18380 13932
rect 18420 13923 18472 13932
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 16304 13812 16356 13864
rect 16028 13744 16080 13796
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 20812 13880 20864 13932
rect 23664 13923 23716 13932
rect 23664 13889 23673 13923
rect 23673 13889 23707 13923
rect 23707 13889 23716 13923
rect 23664 13880 23716 13889
rect 25596 13948 25648 14000
rect 26516 13948 26568 14000
rect 26884 13948 26936 14000
rect 25504 13880 25556 13932
rect 27528 14016 27580 14068
rect 27896 14059 27948 14068
rect 27896 14025 27905 14059
rect 27905 14025 27939 14059
rect 27939 14025 27948 14059
rect 27896 14016 27948 14025
rect 31116 14016 31168 14068
rect 31944 14016 31996 14068
rect 19432 13812 19484 13864
rect 21732 13812 21784 13864
rect 21456 13744 21508 13796
rect 22928 13744 22980 13796
rect 26700 13812 26752 13864
rect 28356 13923 28408 13932
rect 28356 13889 28365 13923
rect 28365 13889 28399 13923
rect 28399 13889 28408 13923
rect 28356 13880 28408 13889
rect 28632 13923 28684 13932
rect 28632 13889 28641 13923
rect 28641 13889 28675 13923
rect 28675 13889 28684 13923
rect 28632 13880 28684 13889
rect 32312 13991 32364 14000
rect 32312 13957 32321 13991
rect 32321 13957 32355 13991
rect 32355 13957 32364 13991
rect 32312 13948 32364 13957
rect 30656 13880 30708 13932
rect 31116 13880 31168 13932
rect 31484 13923 31536 13932
rect 31484 13889 31493 13923
rect 31493 13889 31527 13923
rect 31527 13889 31536 13923
rect 31484 13880 31536 13889
rect 31576 13880 31628 13932
rect 31944 13880 31996 13932
rect 32220 13880 32272 13932
rect 27988 13744 28040 13796
rect 28816 13744 28868 13796
rect 8852 13676 8904 13728
rect 10784 13676 10836 13728
rect 10876 13676 10928 13728
rect 12900 13676 12952 13728
rect 27252 13676 27304 13728
rect 30196 13676 30248 13728
rect 31852 13676 31904 13728
rect 5147 13574 5199 13626
rect 5211 13574 5263 13626
rect 5275 13574 5327 13626
rect 5339 13574 5391 13626
rect 5403 13574 5455 13626
rect 13541 13574 13593 13626
rect 13605 13574 13657 13626
rect 13669 13574 13721 13626
rect 13733 13574 13785 13626
rect 13797 13574 13849 13626
rect 21935 13574 21987 13626
rect 21999 13574 22051 13626
rect 22063 13574 22115 13626
rect 22127 13574 22179 13626
rect 22191 13574 22243 13626
rect 30329 13574 30381 13626
rect 30393 13574 30445 13626
rect 30457 13574 30509 13626
rect 30521 13574 30573 13626
rect 30585 13574 30637 13626
rect 4712 13472 4764 13524
rect 6828 13472 6880 13524
rect 7196 13472 7248 13524
rect 7840 13472 7892 13524
rect 7932 13472 7984 13524
rect 8208 13472 8260 13524
rect 4344 13404 4396 13456
rect 8116 13404 8168 13456
rect 940 13268 992 13320
rect 3332 13268 3384 13320
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 6184 13336 6236 13388
rect 3792 13268 3844 13277
rect 4252 13311 4304 13320
rect 4252 13277 4261 13311
rect 4261 13277 4295 13311
rect 4295 13277 4304 13311
rect 4252 13268 4304 13277
rect 1676 13132 1728 13184
rect 3976 13132 4028 13184
rect 5724 13268 5776 13320
rect 5816 13268 5868 13320
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 8024 13336 8076 13388
rect 7656 13311 7708 13320
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 7656 13268 7708 13277
rect 5632 13200 5684 13252
rect 6828 13200 6880 13252
rect 8208 13268 8260 13320
rect 9496 13472 9548 13524
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 12256 13472 12308 13524
rect 12716 13515 12768 13524
rect 12716 13481 12725 13515
rect 12725 13481 12759 13515
rect 12759 13481 12768 13515
rect 12716 13472 12768 13481
rect 13360 13472 13412 13524
rect 15660 13472 15712 13524
rect 9220 13404 9272 13456
rect 11428 13404 11480 13456
rect 13084 13404 13136 13456
rect 9404 13268 9456 13320
rect 10416 13268 10468 13320
rect 10876 13268 10928 13320
rect 11152 13268 11204 13320
rect 11244 13268 11296 13320
rect 11520 13311 11572 13320
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 12072 13311 12124 13320
rect 6000 13132 6052 13184
rect 6276 13132 6328 13184
rect 6552 13132 6604 13184
rect 8852 13132 8904 13184
rect 8944 13132 8996 13184
rect 9128 13132 9180 13184
rect 11152 13132 11204 13184
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12164 13311 12216 13320
rect 12164 13277 12174 13311
rect 12174 13277 12208 13311
rect 12208 13277 12216 13311
rect 12164 13268 12216 13277
rect 12716 13268 12768 13320
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 12900 13268 12952 13320
rect 20536 13472 20588 13524
rect 20352 13404 20404 13456
rect 21640 13404 21692 13456
rect 22744 13515 22796 13524
rect 22744 13481 22753 13515
rect 22753 13481 22787 13515
rect 22787 13481 22796 13515
rect 22744 13472 22796 13481
rect 23112 13472 23164 13524
rect 23664 13472 23716 13524
rect 26700 13472 26752 13524
rect 13360 13200 13412 13252
rect 15476 13268 15528 13320
rect 15660 13311 15712 13320
rect 15660 13277 15669 13311
rect 15669 13277 15703 13311
rect 15703 13277 15712 13311
rect 15660 13268 15712 13277
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 21548 13336 21600 13388
rect 20536 13243 20588 13252
rect 20536 13209 20545 13243
rect 20545 13209 20579 13243
rect 20579 13209 20588 13243
rect 20536 13200 20588 13209
rect 21456 13268 21508 13320
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22652 13404 22704 13456
rect 22836 13404 22888 13456
rect 30656 13472 30708 13524
rect 31300 13515 31352 13524
rect 31300 13481 31309 13515
rect 31309 13481 31343 13515
rect 31343 13481 31352 13515
rect 31300 13472 31352 13481
rect 24124 13379 24176 13388
rect 24124 13345 24133 13379
rect 24133 13345 24167 13379
rect 24167 13345 24176 13379
rect 24124 13336 24176 13345
rect 24676 13336 24728 13388
rect 24952 13379 25004 13388
rect 24952 13345 24961 13379
rect 24961 13345 24995 13379
rect 24995 13345 25004 13379
rect 24952 13336 25004 13345
rect 27252 13336 27304 13388
rect 27620 13379 27672 13388
rect 27620 13345 27629 13379
rect 27629 13345 27663 13379
rect 27663 13345 27672 13379
rect 27620 13336 27672 13345
rect 31484 13472 31536 13524
rect 31668 13515 31720 13524
rect 31668 13481 31677 13515
rect 31677 13481 31711 13515
rect 31711 13481 31720 13515
rect 31668 13472 31720 13481
rect 22928 13311 22980 13320
rect 22928 13277 22937 13311
rect 22937 13277 22971 13311
rect 22971 13277 22980 13311
rect 22928 13268 22980 13277
rect 12532 13132 12584 13184
rect 12900 13132 12952 13184
rect 15752 13132 15804 13184
rect 20352 13175 20404 13184
rect 20352 13141 20361 13175
rect 20361 13141 20395 13175
rect 20395 13141 20404 13175
rect 20352 13132 20404 13141
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 21916 13200 21968 13252
rect 23388 13268 23440 13320
rect 26056 13268 26108 13320
rect 28172 13268 28224 13320
rect 31116 13336 31168 13388
rect 23664 13200 23716 13252
rect 27436 13200 27488 13252
rect 29552 13200 29604 13252
rect 30196 13243 30248 13252
rect 30196 13209 30205 13243
rect 30205 13209 30239 13243
rect 30239 13209 30248 13243
rect 30196 13200 30248 13209
rect 30656 13200 30708 13252
rect 22284 13132 22336 13184
rect 23296 13132 23348 13184
rect 23572 13132 23624 13184
rect 27896 13175 27948 13184
rect 27896 13141 27905 13175
rect 27905 13141 27939 13175
rect 27939 13141 27948 13175
rect 27896 13132 27948 13141
rect 32680 13132 32732 13184
rect 9344 13030 9396 13082
rect 9408 13030 9460 13082
rect 9472 13030 9524 13082
rect 9536 13030 9588 13082
rect 9600 13030 9652 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 17930 13030 17982 13082
rect 17994 13030 18046 13082
rect 26132 13030 26184 13082
rect 26196 13030 26248 13082
rect 26260 13030 26312 13082
rect 26324 13030 26376 13082
rect 26388 13030 26440 13082
rect 34526 13030 34578 13082
rect 34590 13030 34642 13082
rect 34654 13030 34706 13082
rect 34718 13030 34770 13082
rect 34782 13030 34834 13082
rect 6276 12928 6328 12980
rect 7472 12928 7524 12980
rect 9220 12928 9272 12980
rect 11980 12928 12032 12980
rect 12164 12928 12216 12980
rect 12440 12928 12492 12980
rect 12808 12928 12860 12980
rect 16120 12928 16172 12980
rect 20352 12928 20404 12980
rect 21916 12928 21968 12980
rect 23296 12928 23348 12980
rect 31300 12928 31352 12980
rect 31944 12971 31996 12980
rect 31944 12937 31953 12971
rect 31953 12937 31987 12971
rect 31987 12937 31996 12971
rect 31944 12928 31996 12937
rect 8300 12860 8352 12912
rect 9588 12860 9640 12912
rect 11888 12860 11940 12912
rect 16212 12860 16264 12912
rect 22284 12860 22336 12912
rect 6552 12792 6604 12844
rect 8760 12792 8812 12844
rect 9128 12792 9180 12844
rect 11336 12724 11388 12776
rect 6828 12656 6880 12708
rect 8208 12656 8260 12708
rect 14096 12656 14148 12708
rect 15016 12656 15068 12708
rect 15752 12724 15804 12776
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 18328 12792 18380 12844
rect 23388 12860 23440 12912
rect 25504 12860 25556 12912
rect 22928 12835 22980 12844
rect 22928 12801 22937 12835
rect 22937 12801 22971 12835
rect 22971 12801 22980 12835
rect 22928 12792 22980 12801
rect 24860 12835 24912 12844
rect 24860 12801 24869 12835
rect 24869 12801 24903 12835
rect 24903 12801 24912 12835
rect 24860 12792 24912 12801
rect 25044 12792 25096 12844
rect 27344 12835 27396 12844
rect 27344 12801 27353 12835
rect 27353 12801 27387 12835
rect 27387 12801 27396 12835
rect 27344 12792 27396 12801
rect 27896 12792 27948 12844
rect 31484 12835 31536 12844
rect 31484 12801 31493 12835
rect 31493 12801 31527 12835
rect 31527 12801 31536 12835
rect 31484 12792 31536 12801
rect 23480 12724 23532 12776
rect 23572 12724 23624 12776
rect 24216 12724 24268 12776
rect 27528 12724 27580 12776
rect 27988 12767 28040 12776
rect 27988 12733 27997 12767
rect 27997 12733 28031 12767
rect 28031 12733 28040 12767
rect 27988 12724 28040 12733
rect 31760 12835 31812 12844
rect 31760 12801 31769 12835
rect 31769 12801 31803 12835
rect 31803 12801 31812 12835
rect 31760 12792 31812 12801
rect 32680 12835 32732 12844
rect 32680 12801 32689 12835
rect 32689 12801 32723 12835
rect 32723 12801 32732 12835
rect 32680 12792 32732 12801
rect 33416 12724 33468 12776
rect 33692 12767 33744 12776
rect 33692 12733 33701 12767
rect 33701 12733 33735 12767
rect 33735 12733 33744 12767
rect 33692 12724 33744 12733
rect 33876 12792 33928 12844
rect 33968 12835 34020 12844
rect 33968 12801 33977 12835
rect 33977 12801 34011 12835
rect 34011 12801 34020 12835
rect 33968 12792 34020 12801
rect 34152 12835 34204 12844
rect 34152 12801 34161 12835
rect 34161 12801 34195 12835
rect 34195 12801 34204 12835
rect 34152 12792 34204 12801
rect 7288 12588 7340 12640
rect 7656 12588 7708 12640
rect 8760 12588 8812 12640
rect 8944 12588 8996 12640
rect 10968 12588 11020 12640
rect 15476 12588 15528 12640
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 22284 12588 22336 12640
rect 24676 12631 24728 12640
rect 24676 12597 24685 12631
rect 24685 12597 24719 12631
rect 24719 12597 24728 12631
rect 24676 12588 24728 12597
rect 26976 12631 27028 12640
rect 26976 12597 26985 12631
rect 26985 12597 27019 12631
rect 27019 12597 27028 12631
rect 26976 12588 27028 12597
rect 32036 12588 32088 12640
rect 5147 12486 5199 12538
rect 5211 12486 5263 12538
rect 5275 12486 5327 12538
rect 5339 12486 5391 12538
rect 5403 12486 5455 12538
rect 13541 12486 13593 12538
rect 13605 12486 13657 12538
rect 13669 12486 13721 12538
rect 13733 12486 13785 12538
rect 13797 12486 13849 12538
rect 21935 12486 21987 12538
rect 21999 12486 22051 12538
rect 22063 12486 22115 12538
rect 22127 12486 22179 12538
rect 22191 12486 22243 12538
rect 30329 12486 30381 12538
rect 30393 12486 30445 12538
rect 30457 12486 30509 12538
rect 30521 12486 30573 12538
rect 30585 12486 30637 12538
rect 3792 12384 3844 12436
rect 7104 12384 7156 12436
rect 3424 12316 3476 12368
rect 3332 12248 3384 12300
rect 3608 12223 3660 12232
rect 3608 12189 3617 12223
rect 3617 12189 3651 12223
rect 3651 12189 3660 12223
rect 3608 12180 3660 12189
rect 3884 12180 3936 12232
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 6276 12248 6328 12300
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 4068 12112 4120 12164
rect 5540 12180 5592 12232
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 5448 12155 5500 12164
rect 5448 12121 5457 12155
rect 5457 12121 5491 12155
rect 5491 12121 5500 12155
rect 5448 12112 5500 12121
rect 4252 12044 4304 12096
rect 5080 12087 5132 12096
rect 5080 12053 5089 12087
rect 5089 12053 5123 12087
rect 5123 12053 5132 12087
rect 5080 12044 5132 12053
rect 5816 12044 5868 12096
rect 6184 12044 6236 12096
rect 6460 12223 6512 12232
rect 6460 12189 6466 12223
rect 6466 12189 6500 12223
rect 6500 12189 6512 12223
rect 9036 12384 9088 12436
rect 11060 12427 11112 12436
rect 11060 12393 11069 12427
rect 11069 12393 11103 12427
rect 11103 12393 11112 12427
rect 11060 12384 11112 12393
rect 11980 12384 12032 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 7472 12248 7524 12300
rect 7656 12248 7708 12300
rect 8392 12316 8444 12368
rect 9312 12316 9364 12368
rect 9956 12316 10008 12368
rect 6460 12180 6512 12189
rect 7748 12180 7800 12232
rect 8208 12180 8260 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9588 12248 9640 12300
rect 8300 12112 8352 12164
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 11152 12180 11204 12232
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 12532 12180 12584 12232
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 9864 12112 9916 12164
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 7012 12044 7064 12096
rect 7840 12087 7892 12096
rect 7840 12053 7849 12087
rect 7849 12053 7883 12087
rect 7883 12053 7892 12087
rect 7840 12044 7892 12053
rect 8484 12044 8536 12096
rect 9404 12044 9456 12096
rect 10324 12112 10376 12164
rect 11428 12155 11480 12164
rect 11428 12121 11437 12155
rect 11437 12121 11471 12155
rect 11471 12121 11480 12155
rect 11428 12112 11480 12121
rect 13452 12359 13504 12368
rect 13452 12325 13461 12359
rect 13461 12325 13495 12359
rect 13495 12325 13504 12359
rect 13452 12316 13504 12325
rect 17592 12384 17644 12436
rect 18420 12384 18472 12436
rect 18696 12384 18748 12436
rect 20444 12384 20496 12436
rect 21548 12384 21600 12436
rect 22376 12384 22428 12436
rect 23480 12384 23532 12436
rect 19708 12316 19760 12368
rect 17500 12248 17552 12300
rect 18144 12248 18196 12300
rect 13360 12180 13412 12232
rect 16856 12180 16908 12232
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 17040 12112 17092 12164
rect 10692 12044 10744 12096
rect 11888 12044 11940 12096
rect 12992 12044 13044 12096
rect 16488 12087 16540 12096
rect 16488 12053 16497 12087
rect 16497 12053 16531 12087
rect 16531 12053 16540 12087
rect 16488 12044 16540 12053
rect 17408 12044 17460 12096
rect 17592 12087 17644 12096
rect 17592 12053 17601 12087
rect 17601 12053 17635 12087
rect 17635 12053 17644 12087
rect 17592 12044 17644 12053
rect 18788 12180 18840 12232
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20260 12180 20312 12189
rect 18328 12155 18380 12164
rect 18328 12121 18337 12155
rect 18337 12121 18371 12155
rect 18371 12121 18380 12155
rect 18328 12112 18380 12121
rect 19708 12112 19760 12164
rect 21548 12223 21600 12232
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 22560 12248 22612 12300
rect 22284 12180 22336 12232
rect 23296 12316 23348 12368
rect 22836 12248 22888 12300
rect 25044 12384 25096 12436
rect 23572 12291 23624 12300
rect 23572 12257 23581 12291
rect 23581 12257 23615 12291
rect 23615 12257 23624 12291
rect 23572 12248 23624 12257
rect 26516 12291 26568 12300
rect 26516 12257 26525 12291
rect 26525 12257 26559 12291
rect 26559 12257 26568 12291
rect 26516 12248 26568 12257
rect 26792 12291 26844 12300
rect 26792 12257 26801 12291
rect 26801 12257 26835 12291
rect 26835 12257 26844 12291
rect 26792 12248 26844 12257
rect 27436 12248 27488 12300
rect 29736 12384 29788 12436
rect 30932 12384 30984 12436
rect 22376 12112 22428 12164
rect 23756 12180 23808 12232
rect 23664 12112 23716 12164
rect 25688 12180 25740 12232
rect 29000 12248 29052 12300
rect 29552 12223 29604 12232
rect 29552 12189 29561 12223
rect 29561 12189 29595 12223
rect 29595 12189 29604 12223
rect 29552 12180 29604 12189
rect 24676 12155 24728 12164
rect 24676 12121 24685 12155
rect 24685 12121 24719 12155
rect 24719 12121 24728 12155
rect 24676 12112 24728 12121
rect 18144 12087 18196 12096
rect 18144 12053 18171 12087
rect 18171 12053 18196 12087
rect 18144 12044 18196 12053
rect 18604 12044 18656 12096
rect 20168 12087 20220 12096
rect 20168 12053 20177 12087
rect 20177 12053 20211 12087
rect 20211 12053 20220 12087
rect 20168 12044 20220 12053
rect 20996 12044 21048 12096
rect 21088 12044 21140 12096
rect 24032 12044 24084 12096
rect 24952 12044 25004 12096
rect 30012 12180 30064 12232
rect 31024 12316 31076 12368
rect 31392 12384 31444 12436
rect 31576 12384 31628 12436
rect 31760 12384 31812 12436
rect 33876 12384 33928 12436
rect 34152 12384 34204 12436
rect 29736 12155 29788 12164
rect 29736 12121 29745 12155
rect 29745 12121 29779 12155
rect 29779 12121 29788 12155
rect 29736 12112 29788 12121
rect 28172 12044 28224 12096
rect 30196 12087 30248 12096
rect 30196 12053 30205 12087
rect 30205 12053 30239 12087
rect 30239 12053 30248 12087
rect 30196 12044 30248 12053
rect 30564 12087 30616 12096
rect 30564 12053 30573 12087
rect 30573 12053 30607 12087
rect 30607 12053 30616 12087
rect 30564 12044 30616 12053
rect 31208 12180 31260 12232
rect 31300 12223 31352 12232
rect 31300 12189 31309 12223
rect 31309 12189 31343 12223
rect 31343 12189 31352 12223
rect 31300 12180 31352 12189
rect 31484 12155 31536 12164
rect 31484 12121 31493 12155
rect 31493 12121 31527 12155
rect 31527 12121 31536 12155
rect 31484 12112 31536 12121
rect 31668 12223 31720 12232
rect 31668 12189 31677 12223
rect 31677 12189 31711 12223
rect 31711 12189 31720 12223
rect 31668 12180 31720 12189
rect 31760 12223 31812 12232
rect 31760 12189 31769 12223
rect 31769 12189 31803 12223
rect 31803 12189 31812 12223
rect 31760 12180 31812 12189
rect 32036 12112 32088 12164
rect 33968 12087 34020 12096
rect 33968 12053 33977 12087
rect 33977 12053 34011 12087
rect 34011 12053 34020 12087
rect 33968 12044 34020 12053
rect 9344 11942 9396 11994
rect 9408 11942 9460 11994
rect 9472 11942 9524 11994
rect 9536 11942 9588 11994
rect 9600 11942 9652 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 17930 11942 17982 11994
rect 17994 11942 18046 11994
rect 26132 11942 26184 11994
rect 26196 11942 26248 11994
rect 26260 11942 26312 11994
rect 26324 11942 26376 11994
rect 26388 11942 26440 11994
rect 34526 11942 34578 11994
rect 34590 11942 34642 11994
rect 34654 11942 34706 11994
rect 34718 11942 34770 11994
rect 34782 11942 34834 11994
rect 3240 11840 3292 11892
rect 4068 11840 4120 11892
rect 5080 11840 5132 11892
rect 6460 11840 6512 11892
rect 6552 11840 6604 11892
rect 6736 11840 6788 11892
rect 7564 11840 7616 11892
rect 8484 11840 8536 11892
rect 9036 11840 9088 11892
rect 9220 11840 9272 11892
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 3700 11704 3752 11756
rect 3884 11704 3936 11756
rect 4252 11747 4304 11756
rect 4252 11713 4261 11747
rect 4261 11713 4295 11747
rect 4295 11713 4304 11747
rect 4252 11704 4304 11713
rect 4436 11636 4488 11688
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 6184 11704 6236 11756
rect 7472 11772 7524 11824
rect 8116 11772 8168 11824
rect 9772 11772 9824 11824
rect 6368 11679 6420 11688
rect 6368 11645 6377 11679
rect 6377 11645 6411 11679
rect 6411 11645 6420 11679
rect 6368 11636 6420 11645
rect 6920 11704 6972 11756
rect 7012 11636 7064 11688
rect 7748 11704 7800 11756
rect 8208 11636 8260 11688
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 3976 11500 4028 11552
rect 8116 11568 8168 11620
rect 9036 11747 9088 11756
rect 9036 11713 9046 11747
rect 9046 11713 9080 11747
rect 9080 11713 9088 11747
rect 9036 11704 9088 11713
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 10416 11772 10468 11824
rect 8760 11636 8812 11688
rect 10232 11704 10284 11756
rect 10324 11704 10376 11756
rect 10784 11840 10836 11892
rect 10692 11772 10744 11824
rect 11428 11772 11480 11824
rect 9496 11679 9548 11680
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11628 9548 11645
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11244 11704 11296 11756
rect 11888 11840 11940 11892
rect 12072 11840 12124 11892
rect 12900 11840 12952 11892
rect 13268 11840 13320 11892
rect 13452 11840 13504 11892
rect 16488 11840 16540 11892
rect 17040 11840 17092 11892
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 13636 11772 13688 11824
rect 13544 11747 13596 11756
rect 13544 11713 13553 11747
rect 13553 11713 13587 11747
rect 13587 11713 13596 11747
rect 13544 11704 13596 11713
rect 13728 11747 13780 11756
rect 13728 11713 13737 11747
rect 13737 11713 13771 11747
rect 13771 11713 13780 11747
rect 13728 11704 13780 11713
rect 17408 11772 17460 11824
rect 18144 11840 18196 11892
rect 18420 11840 18472 11892
rect 16764 11747 16816 11756
rect 16764 11713 16773 11747
rect 16773 11713 16807 11747
rect 16807 11713 16816 11747
rect 16764 11704 16816 11713
rect 17224 11704 17276 11756
rect 18236 11772 18288 11824
rect 19708 11883 19760 11892
rect 19708 11849 19717 11883
rect 19717 11849 19751 11883
rect 19751 11849 19760 11883
rect 19708 11840 19760 11849
rect 21088 11840 21140 11892
rect 21548 11840 21600 11892
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 8392 11500 8444 11552
rect 10324 11568 10376 11620
rect 16856 11636 16908 11688
rect 17040 11679 17092 11688
rect 17040 11645 17049 11679
rect 17049 11645 17083 11679
rect 17083 11645 17092 11679
rect 17040 11636 17092 11645
rect 19616 11704 19668 11756
rect 19984 11704 20036 11756
rect 20076 11747 20128 11756
rect 20076 11713 20085 11747
rect 20085 11713 20119 11747
rect 20119 11713 20128 11747
rect 20076 11704 20128 11713
rect 20168 11704 20220 11756
rect 20444 11747 20496 11756
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 20444 11704 20496 11713
rect 21548 11704 21600 11756
rect 22376 11840 22428 11892
rect 22468 11883 22520 11892
rect 22468 11849 22477 11883
rect 22477 11849 22511 11883
rect 22511 11849 22520 11883
rect 22468 11840 22520 11849
rect 21732 11772 21784 11824
rect 22652 11772 22704 11824
rect 24032 11840 24084 11892
rect 24860 11840 24912 11892
rect 24952 11883 25004 11892
rect 24952 11849 24961 11883
rect 24961 11849 24995 11883
rect 24995 11849 25004 11883
rect 24952 11840 25004 11849
rect 27988 11772 28040 11824
rect 30196 11772 30248 11824
rect 18604 11636 18656 11688
rect 9956 11500 10008 11552
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 10508 11500 10560 11552
rect 11152 11500 11204 11552
rect 11336 11543 11388 11552
rect 11336 11509 11345 11543
rect 11345 11509 11379 11543
rect 11379 11509 11388 11543
rect 11336 11500 11388 11509
rect 15200 11500 15252 11552
rect 20168 11568 20220 11620
rect 20904 11636 20956 11688
rect 21640 11636 21692 11688
rect 22560 11704 22612 11756
rect 22744 11735 22754 11756
rect 22754 11735 22788 11756
rect 22788 11735 22796 11756
rect 22744 11704 22796 11735
rect 17960 11500 18012 11552
rect 18420 11500 18472 11552
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 29000 11704 29052 11756
rect 30564 11840 30616 11892
rect 31300 11772 31352 11824
rect 22836 11568 22888 11620
rect 22928 11568 22980 11620
rect 24308 11636 24360 11688
rect 25044 11636 25096 11688
rect 29552 11636 29604 11688
rect 31392 11568 31444 11620
rect 31944 11568 31996 11620
rect 27528 11500 27580 11552
rect 30012 11500 30064 11552
rect 31208 11500 31260 11552
rect 31668 11543 31720 11552
rect 31668 11509 31677 11543
rect 31677 11509 31711 11543
rect 31711 11509 31720 11543
rect 31668 11500 31720 11509
rect 32496 11500 32548 11552
rect 5147 11398 5199 11450
rect 5211 11398 5263 11450
rect 5275 11398 5327 11450
rect 5339 11398 5391 11450
rect 5403 11398 5455 11450
rect 13541 11398 13593 11450
rect 13605 11398 13657 11450
rect 13669 11398 13721 11450
rect 13733 11398 13785 11450
rect 13797 11398 13849 11450
rect 21935 11398 21987 11450
rect 21999 11398 22051 11450
rect 22063 11398 22115 11450
rect 22127 11398 22179 11450
rect 22191 11398 22243 11450
rect 30329 11398 30381 11450
rect 30393 11398 30445 11450
rect 30457 11398 30509 11450
rect 30521 11398 30573 11450
rect 30585 11398 30637 11450
rect 3424 11296 3476 11348
rect 4436 11296 4488 11348
rect 5540 11296 5592 11348
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 8116 11296 8168 11348
rect 9036 11296 9088 11348
rect 9956 11339 10008 11348
rect 9956 11305 9965 11339
rect 9965 11305 9999 11339
rect 9999 11305 10008 11339
rect 9956 11296 10008 11305
rect 10324 11296 10376 11348
rect 11244 11296 11296 11348
rect 11336 11296 11388 11348
rect 12348 11296 12400 11348
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 1676 11203 1728 11212
rect 1676 11169 1685 11203
rect 1685 11169 1719 11203
rect 1719 11169 1728 11203
rect 1676 11160 1728 11169
rect 2964 11092 3016 11144
rect 3240 11092 3292 11144
rect 6184 11160 6236 11212
rect 6460 11203 6512 11212
rect 6460 11169 6469 11203
rect 6469 11169 6503 11203
rect 6503 11169 6512 11203
rect 6460 11160 6512 11169
rect 6828 11271 6880 11280
rect 6828 11237 6837 11271
rect 6837 11237 6871 11271
rect 6871 11237 6880 11271
rect 6828 11228 6880 11237
rect 7472 11160 7524 11212
rect 8944 11228 8996 11280
rect 3976 11024 4028 11076
rect 6736 11092 6788 11144
rect 7288 11092 7340 11144
rect 3148 10999 3200 11008
rect 3148 10965 3157 10999
rect 3157 10965 3191 10999
rect 3191 10965 3200 10999
rect 3148 10956 3200 10965
rect 4712 11024 4764 11076
rect 7932 11092 7984 11144
rect 8208 11092 8260 11144
rect 8852 11092 8904 11144
rect 12900 11228 12952 11280
rect 9772 11160 9824 11212
rect 13084 11296 13136 11348
rect 13912 11296 13964 11348
rect 17960 11296 18012 11348
rect 20904 11296 20956 11348
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 21456 11296 21508 11348
rect 21548 11296 21600 11348
rect 30656 11296 30708 11348
rect 31300 11296 31352 11348
rect 31576 11296 31628 11348
rect 8576 11024 8628 11076
rect 8760 11024 8812 11076
rect 6828 10956 6880 11008
rect 8024 10956 8076 11008
rect 9956 10956 10008 11008
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 12532 11092 12584 11144
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 17040 11228 17092 11280
rect 17592 11228 17644 11280
rect 18512 11228 18564 11280
rect 14004 11160 14056 11212
rect 14556 11160 14608 11212
rect 15200 11160 15252 11212
rect 12532 10956 12584 11008
rect 13268 11024 13320 11076
rect 13360 10956 13412 11008
rect 15936 10956 15988 11008
rect 26516 11228 26568 11280
rect 30012 11228 30064 11280
rect 31760 11228 31812 11280
rect 20076 11024 20128 11076
rect 22928 11160 22980 11212
rect 22652 11092 22704 11144
rect 22744 11092 22796 11144
rect 27620 11160 27672 11212
rect 22560 11067 22612 11076
rect 22560 11033 22569 11067
rect 22569 11033 22603 11067
rect 22603 11033 22612 11067
rect 22560 11024 22612 11033
rect 26700 11135 26752 11144
rect 26700 11101 26709 11135
rect 26709 11101 26743 11135
rect 26743 11101 26752 11135
rect 26700 11092 26752 11101
rect 29000 11160 29052 11212
rect 30932 11160 30984 11212
rect 32036 11203 32088 11212
rect 28540 11092 28592 11144
rect 30288 11135 30340 11144
rect 25688 11024 25740 11076
rect 30288 11101 30297 11135
rect 30297 11101 30331 11135
rect 30331 11101 30340 11135
rect 30288 11092 30340 11101
rect 32036 11169 32045 11203
rect 32045 11169 32079 11203
rect 32079 11169 32088 11203
rect 32036 11160 32088 11169
rect 31300 11135 31352 11144
rect 31300 11101 31309 11135
rect 31309 11101 31343 11135
rect 31343 11101 31352 11135
rect 31300 11092 31352 11101
rect 31668 11092 31720 11144
rect 28724 10999 28776 11008
rect 28724 10965 28733 10999
rect 28733 10965 28767 10999
rect 28767 10965 28776 10999
rect 28724 10956 28776 10965
rect 31208 10956 31260 11008
rect 33048 10956 33100 11008
rect 9344 10854 9396 10906
rect 9408 10854 9460 10906
rect 9472 10854 9524 10906
rect 9536 10854 9588 10906
rect 9600 10854 9652 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 17930 10854 17982 10906
rect 17994 10854 18046 10906
rect 26132 10854 26184 10906
rect 26196 10854 26248 10906
rect 26260 10854 26312 10906
rect 26324 10854 26376 10906
rect 26388 10854 26440 10906
rect 34526 10854 34578 10906
rect 34590 10854 34642 10906
rect 34654 10854 34706 10906
rect 34718 10854 34770 10906
rect 34782 10854 34834 10906
rect 9680 10752 9732 10804
rect 17500 10752 17552 10804
rect 3148 10616 3200 10668
rect 4620 10616 4672 10668
rect 6276 10684 6328 10736
rect 6368 10684 6420 10736
rect 4988 10659 5040 10668
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 7748 10684 7800 10736
rect 12808 10684 12860 10736
rect 4712 10591 4764 10600
rect 4712 10557 4721 10591
rect 4721 10557 4755 10591
rect 4755 10557 4764 10591
rect 4712 10548 4764 10557
rect 3332 10480 3384 10532
rect 5816 10548 5868 10600
rect 6920 10548 6972 10600
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3056 10412 3108 10421
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 6828 10480 6880 10532
rect 7564 10616 7616 10668
rect 11060 10616 11112 10668
rect 12716 10616 12768 10668
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 17592 10616 17644 10668
rect 20168 10795 20220 10804
rect 20168 10761 20177 10795
rect 20177 10761 20211 10795
rect 20211 10761 20220 10795
rect 20168 10752 20220 10761
rect 25688 10752 25740 10804
rect 25136 10684 25188 10736
rect 26700 10752 26752 10804
rect 30288 10727 30340 10736
rect 30288 10693 30297 10727
rect 30297 10693 30331 10727
rect 30331 10693 30340 10727
rect 30288 10684 30340 10693
rect 30932 10684 30984 10736
rect 19984 10616 20036 10668
rect 23112 10659 23164 10668
rect 23112 10625 23121 10659
rect 23121 10625 23155 10659
rect 23155 10625 23164 10659
rect 23112 10616 23164 10625
rect 24124 10616 24176 10668
rect 24492 10659 24544 10668
rect 24492 10625 24501 10659
rect 24501 10625 24535 10659
rect 24535 10625 24544 10659
rect 24492 10616 24544 10625
rect 28724 10659 28776 10668
rect 28724 10625 28733 10659
rect 28733 10625 28767 10659
rect 28767 10625 28776 10659
rect 28724 10616 28776 10625
rect 11244 10548 11296 10600
rect 13084 10548 13136 10600
rect 13176 10548 13228 10600
rect 13360 10548 13412 10600
rect 17868 10591 17920 10600
rect 17868 10557 17902 10591
rect 17902 10557 17920 10591
rect 17868 10548 17920 10557
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 27528 10591 27580 10600
rect 27528 10557 27537 10591
rect 27537 10557 27571 10591
rect 27571 10557 27580 10591
rect 27528 10548 27580 10557
rect 31576 10659 31628 10668
rect 31576 10625 31585 10659
rect 31585 10625 31619 10659
rect 31619 10625 31628 10659
rect 31576 10616 31628 10625
rect 31760 10659 31812 10668
rect 31760 10625 31769 10659
rect 31769 10625 31803 10659
rect 31803 10625 31812 10659
rect 31760 10616 31812 10625
rect 32496 10659 32548 10668
rect 32496 10625 32505 10659
rect 32505 10625 32539 10659
rect 32539 10625 32548 10659
rect 32496 10616 32548 10625
rect 33048 10795 33100 10804
rect 33048 10761 33057 10795
rect 33057 10761 33091 10795
rect 33091 10761 33100 10795
rect 33048 10752 33100 10761
rect 33048 10616 33100 10668
rect 8576 10480 8628 10532
rect 7104 10412 7156 10464
rect 28172 10480 28224 10532
rect 30656 10523 30708 10532
rect 30656 10489 30665 10523
rect 30665 10489 30699 10523
rect 30699 10489 30708 10523
rect 30656 10480 30708 10489
rect 31300 10480 31352 10532
rect 32220 10548 32272 10600
rect 33784 10548 33836 10600
rect 33876 10480 33928 10532
rect 12348 10412 12400 10464
rect 12624 10412 12676 10464
rect 22928 10455 22980 10464
rect 22928 10421 22937 10455
rect 22937 10421 22971 10455
rect 22971 10421 22980 10455
rect 22928 10412 22980 10421
rect 26608 10412 26660 10464
rect 28540 10412 28592 10464
rect 31208 10412 31260 10464
rect 31760 10412 31812 10464
rect 31944 10412 31996 10464
rect 32128 10455 32180 10464
rect 32128 10421 32137 10455
rect 32137 10421 32171 10455
rect 32171 10421 32180 10455
rect 32128 10412 32180 10421
rect 5147 10310 5199 10362
rect 5211 10310 5263 10362
rect 5275 10310 5327 10362
rect 5339 10310 5391 10362
rect 5403 10310 5455 10362
rect 13541 10310 13593 10362
rect 13605 10310 13657 10362
rect 13669 10310 13721 10362
rect 13733 10310 13785 10362
rect 13797 10310 13849 10362
rect 21935 10310 21987 10362
rect 21999 10310 22051 10362
rect 22063 10310 22115 10362
rect 22127 10310 22179 10362
rect 22191 10310 22243 10362
rect 30329 10310 30381 10362
rect 30393 10310 30445 10362
rect 30457 10310 30509 10362
rect 30521 10310 30573 10362
rect 30585 10310 30637 10362
rect 6368 10208 6420 10260
rect 6644 10208 6696 10260
rect 5816 10072 5868 10124
rect 7748 10208 7800 10260
rect 8576 10208 8628 10260
rect 8668 10208 8720 10260
rect 8208 10140 8260 10192
rect 8484 10140 8536 10192
rect 5540 10004 5592 10056
rect 11060 10208 11112 10260
rect 13452 10208 13504 10260
rect 17408 10208 17460 10260
rect 17868 10251 17920 10260
rect 17868 10217 17877 10251
rect 17877 10217 17911 10251
rect 17911 10217 17920 10251
rect 17868 10208 17920 10217
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 19064 10208 19116 10260
rect 22928 10208 22980 10260
rect 24492 10208 24544 10260
rect 27620 10208 27672 10260
rect 11152 10140 11204 10192
rect 13176 10140 13228 10192
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 4528 9936 4580 9988
rect 7196 10004 7248 10056
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 7932 10004 7984 10056
rect 8392 10004 8444 10056
rect 11244 10072 11296 10124
rect 11428 10072 11480 10124
rect 11704 10072 11756 10124
rect 9220 10004 9272 10056
rect 7012 9936 7064 9988
rect 7104 9979 7156 9988
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 7104 9936 7156 9945
rect 7472 9936 7524 9988
rect 9680 10004 9732 10056
rect 10876 10004 10928 10056
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 11796 10004 11848 10056
rect 12072 10004 12124 10056
rect 12256 10004 12308 10056
rect 12532 10072 12584 10124
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 12900 10004 12952 10056
rect 7656 9868 7708 9920
rect 24400 10140 24452 10192
rect 23480 10072 23532 10124
rect 24124 10072 24176 10124
rect 24308 10072 24360 10124
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 17408 9936 17460 9988
rect 10324 9868 10376 9920
rect 10416 9868 10468 9920
rect 11060 9868 11112 9920
rect 12992 9868 13044 9920
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 14096 9868 14148 9920
rect 17316 9868 17368 9920
rect 20168 9936 20220 9988
rect 19984 9868 20036 9920
rect 25136 10004 25188 10056
rect 26608 10115 26660 10124
rect 26608 10081 26617 10115
rect 26617 10081 26651 10115
rect 26651 10081 26660 10115
rect 26608 10072 26660 10081
rect 25044 9936 25096 9988
rect 28264 10004 28316 10056
rect 28172 9979 28224 9988
rect 28172 9945 28181 9979
rect 28181 9945 28215 9979
rect 28215 9945 28224 9979
rect 28172 9936 28224 9945
rect 28816 10047 28868 10056
rect 28816 10013 28825 10047
rect 28825 10013 28859 10047
rect 28859 10013 28868 10047
rect 28816 10004 28868 10013
rect 28356 9868 28408 9920
rect 31300 10251 31352 10260
rect 31300 10217 31309 10251
rect 31309 10217 31343 10251
rect 31343 10217 31352 10251
rect 31300 10208 31352 10217
rect 31024 10140 31076 10192
rect 31576 10140 31628 10192
rect 32128 10208 32180 10260
rect 33876 10208 33928 10260
rect 32220 10140 32272 10192
rect 32220 9936 32272 9988
rect 34336 10004 34388 10056
rect 32956 9868 33008 9920
rect 9344 9766 9396 9818
rect 9408 9766 9460 9818
rect 9472 9766 9524 9818
rect 9536 9766 9588 9818
rect 9600 9766 9652 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 17930 9766 17982 9818
rect 17994 9766 18046 9818
rect 26132 9766 26184 9818
rect 26196 9766 26248 9818
rect 26260 9766 26312 9818
rect 26324 9766 26376 9818
rect 26388 9766 26440 9818
rect 34526 9766 34578 9818
rect 34590 9766 34642 9818
rect 34654 9766 34706 9818
rect 34718 9766 34770 9818
rect 34782 9766 34834 9818
rect 6184 9664 6236 9716
rect 8760 9664 8812 9716
rect 9220 9664 9272 9716
rect 9496 9664 9548 9716
rect 9588 9664 9640 9716
rect 9680 9664 9732 9716
rect 3056 9596 3108 9648
rect 3240 9596 3292 9648
rect 1400 9528 1452 9580
rect 2688 9571 2740 9580
rect 2688 9537 2697 9571
rect 2697 9537 2731 9571
rect 2731 9537 2740 9571
rect 2688 9528 2740 9537
rect 8024 9528 8076 9580
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 9312 9596 9364 9648
rect 8944 9392 8996 9444
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 7012 9324 7064 9376
rect 9864 9571 9916 9580
rect 9864 9537 9873 9571
rect 9873 9537 9907 9571
rect 9907 9537 9916 9571
rect 9864 9528 9916 9537
rect 10048 9707 10100 9716
rect 10048 9673 10057 9707
rect 10057 9673 10091 9707
rect 10091 9673 10100 9707
rect 10048 9664 10100 9673
rect 10324 9664 10376 9716
rect 10508 9596 10560 9648
rect 10600 9596 10652 9648
rect 11060 9596 11112 9648
rect 11428 9664 11480 9716
rect 11612 9664 11664 9716
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11704 9596 11756 9648
rect 11244 9528 11296 9580
rect 11428 9528 11480 9580
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 12624 9596 12676 9648
rect 13084 9664 13136 9716
rect 17224 9664 17276 9716
rect 17592 9664 17644 9716
rect 13176 9596 13228 9648
rect 13268 9596 13320 9648
rect 14648 9596 14700 9648
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 12440 9528 12492 9580
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 13360 9528 13412 9580
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 13728 9571 13780 9580
rect 13728 9537 13737 9571
rect 13737 9537 13771 9571
rect 13771 9537 13780 9571
rect 13728 9528 13780 9537
rect 9404 9392 9456 9444
rect 11704 9392 11756 9444
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 15476 9596 15528 9648
rect 15844 9596 15896 9648
rect 17316 9596 17368 9648
rect 18144 9596 18196 9648
rect 21640 9639 21692 9648
rect 21640 9605 21649 9639
rect 21649 9605 21683 9639
rect 21683 9605 21692 9639
rect 21640 9596 21692 9605
rect 21732 9596 21784 9648
rect 21824 9634 21876 9686
rect 23112 9664 23164 9716
rect 27896 9664 27948 9716
rect 28816 9664 28868 9716
rect 14740 9460 14792 9469
rect 15016 9435 15068 9444
rect 15016 9401 15025 9435
rect 15025 9401 15059 9435
rect 15059 9401 15068 9435
rect 15016 9392 15068 9401
rect 15108 9392 15160 9444
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 15844 9460 15896 9512
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 19984 9528 20036 9580
rect 17408 9460 17460 9512
rect 11244 9324 11296 9376
rect 12440 9324 12492 9376
rect 12992 9324 13044 9376
rect 14464 9324 14516 9376
rect 15200 9367 15252 9376
rect 15200 9333 15209 9367
rect 15209 9333 15243 9367
rect 15243 9333 15252 9367
rect 15200 9324 15252 9333
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 16120 9324 16172 9376
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16212 9324 16264 9333
rect 17500 9324 17552 9376
rect 18696 9503 18748 9512
rect 18696 9469 18705 9503
rect 18705 9469 18739 9503
rect 18739 9469 18748 9503
rect 18696 9460 18748 9469
rect 19064 9460 19116 9512
rect 20168 9503 20220 9512
rect 20168 9469 20177 9503
rect 20177 9469 20211 9503
rect 20211 9469 20220 9503
rect 20168 9460 20220 9469
rect 20536 9460 20588 9512
rect 21180 9571 21232 9580
rect 21180 9537 21189 9571
rect 21189 9537 21223 9571
rect 21223 9537 21232 9571
rect 21180 9528 21232 9537
rect 21364 9571 21416 9580
rect 21364 9537 21373 9571
rect 21373 9537 21407 9571
rect 21407 9537 21416 9571
rect 21364 9528 21416 9537
rect 22560 9596 22612 9648
rect 26516 9596 26568 9648
rect 19892 9392 19944 9444
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 22008 9503 22060 9512
rect 22008 9469 22017 9503
rect 22017 9469 22051 9503
rect 22051 9469 22060 9503
rect 22008 9460 22060 9469
rect 24400 9571 24452 9580
rect 24400 9537 24409 9571
rect 24409 9537 24443 9571
rect 24443 9537 24452 9571
rect 24400 9528 24452 9537
rect 22284 9460 22336 9512
rect 25044 9460 25096 9512
rect 22560 9392 22612 9444
rect 27804 9528 27856 9580
rect 29552 9528 29604 9580
rect 30840 9528 30892 9580
rect 31668 9528 31720 9580
rect 27160 9460 27212 9512
rect 27528 9503 27580 9512
rect 27528 9469 27537 9503
rect 27537 9469 27571 9503
rect 27571 9469 27580 9503
rect 27528 9460 27580 9469
rect 29920 9503 29972 9512
rect 29920 9469 29929 9503
rect 29929 9469 29963 9503
rect 29963 9469 29972 9503
rect 29920 9460 29972 9469
rect 31300 9460 31352 9512
rect 20628 9324 20680 9376
rect 20904 9324 20956 9376
rect 20996 9324 21048 9376
rect 31116 9392 31168 9444
rect 31484 9392 31536 9444
rect 26332 9324 26384 9376
rect 26516 9324 26568 9376
rect 29828 9367 29880 9376
rect 29828 9333 29837 9367
rect 29837 9333 29871 9367
rect 29871 9333 29880 9367
rect 29828 9324 29880 9333
rect 31208 9367 31260 9376
rect 31208 9333 31217 9367
rect 31217 9333 31251 9367
rect 31251 9333 31260 9367
rect 31208 9324 31260 9333
rect 5147 9222 5199 9274
rect 5211 9222 5263 9274
rect 5275 9222 5327 9274
rect 5339 9222 5391 9274
rect 5403 9222 5455 9274
rect 13541 9222 13593 9274
rect 13605 9222 13657 9274
rect 13669 9222 13721 9274
rect 13733 9222 13785 9274
rect 13797 9222 13849 9274
rect 21935 9222 21987 9274
rect 21999 9222 22051 9274
rect 22063 9222 22115 9274
rect 22127 9222 22179 9274
rect 22191 9222 22243 9274
rect 30329 9222 30381 9274
rect 30393 9222 30445 9274
rect 30457 9222 30509 9274
rect 30521 9222 30573 9274
rect 30585 9222 30637 9274
rect 4436 9120 4488 9172
rect 8024 9120 8076 9172
rect 8852 9120 8904 9172
rect 9588 9120 9640 9172
rect 10968 9120 11020 9172
rect 11520 9120 11572 9172
rect 12348 9120 12400 9172
rect 9496 8984 9548 9036
rect 9956 8984 10008 9036
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 12256 8916 12308 8968
rect 14464 9120 14516 9172
rect 15752 9120 15804 9172
rect 16212 9120 16264 9172
rect 16304 9120 16356 9172
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 17408 9163 17460 9172
rect 17408 9129 17417 9163
rect 17417 9129 17451 9163
rect 17451 9129 17460 9163
rect 17408 9120 17460 9129
rect 14740 8916 14792 8968
rect 14648 8848 14700 8900
rect 13912 8780 13964 8832
rect 15108 8916 15160 8968
rect 15568 8916 15620 8968
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 16120 8984 16172 9036
rect 16488 8959 16540 8968
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 15844 8848 15896 8900
rect 15660 8780 15712 8832
rect 16672 8848 16724 8900
rect 17592 8823 17644 8832
rect 17592 8789 17619 8823
rect 17619 8789 17644 8823
rect 17592 8780 17644 8789
rect 18144 9120 18196 9172
rect 18696 9120 18748 9172
rect 20904 9163 20956 9172
rect 20904 9129 20913 9163
rect 20913 9129 20947 9163
rect 20947 9129 20956 9163
rect 20904 9120 20956 9129
rect 21180 9120 21232 9172
rect 20628 8916 20680 8968
rect 21640 8984 21692 9036
rect 21916 9027 21968 9036
rect 21916 8993 21925 9027
rect 21925 8993 21959 9027
rect 21959 8993 21968 9027
rect 21916 8984 21968 8993
rect 22376 8984 22428 9036
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 18052 8848 18104 8900
rect 20536 8848 20588 8900
rect 18144 8780 18196 8832
rect 21732 8848 21784 8900
rect 22468 8916 22520 8968
rect 23756 9120 23808 9172
rect 26332 9027 26384 9036
rect 26332 8993 26341 9027
rect 26341 8993 26375 9027
rect 26375 8993 26384 9027
rect 26332 8984 26384 8993
rect 26056 8959 26108 8968
rect 26056 8925 26065 8959
rect 26065 8925 26099 8959
rect 26099 8925 26108 8959
rect 26056 8916 26108 8925
rect 27804 9163 27856 9172
rect 27804 9129 27813 9163
rect 27813 9129 27847 9163
rect 27847 9129 27856 9163
rect 27804 9120 27856 9129
rect 30840 9163 30892 9172
rect 30840 9129 30849 9163
rect 30849 9129 30883 9163
rect 30883 9129 30892 9163
rect 30840 9120 30892 9129
rect 31760 9163 31812 9172
rect 28264 9027 28316 9036
rect 28264 8993 28273 9027
rect 28273 8993 28307 9027
rect 28307 8993 28316 9027
rect 28264 8984 28316 8993
rect 27896 8959 27948 8968
rect 27896 8925 27905 8959
rect 27905 8925 27939 8959
rect 27939 8925 27948 8959
rect 27896 8916 27948 8925
rect 26608 8848 26660 8900
rect 29828 8848 29880 8900
rect 31760 9129 31769 9163
rect 31769 9129 31803 9163
rect 31803 9129 31812 9163
rect 31760 9120 31812 9129
rect 32036 9163 32088 9172
rect 32036 9129 32045 9163
rect 32045 9129 32079 9163
rect 32079 9129 32088 9163
rect 32036 9120 32088 9129
rect 32220 9120 32272 9172
rect 31576 9052 31628 9104
rect 31668 8984 31720 9036
rect 32404 8984 32456 9036
rect 33048 8984 33100 9036
rect 31484 8848 31536 8900
rect 23756 8823 23808 8832
rect 23756 8789 23765 8823
rect 23765 8789 23799 8823
rect 23799 8789 23808 8823
rect 23756 8780 23808 8789
rect 25596 8780 25648 8832
rect 27344 8780 27396 8832
rect 28356 8780 28408 8832
rect 28724 8823 28776 8832
rect 28724 8789 28733 8823
rect 28733 8789 28767 8823
rect 28767 8789 28776 8823
rect 28724 8780 28776 8789
rect 31392 8823 31444 8832
rect 31392 8789 31401 8823
rect 31401 8789 31435 8823
rect 31435 8789 31444 8823
rect 31392 8780 31444 8789
rect 31760 8780 31812 8832
rect 33048 8823 33100 8832
rect 33048 8789 33057 8823
rect 33057 8789 33091 8823
rect 33091 8789 33100 8823
rect 33048 8780 33100 8789
rect 9344 8678 9396 8730
rect 9408 8678 9460 8730
rect 9472 8678 9524 8730
rect 9536 8678 9588 8730
rect 9600 8678 9652 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 17930 8678 17982 8730
rect 17994 8678 18046 8730
rect 26132 8678 26184 8730
rect 26196 8678 26248 8730
rect 26260 8678 26312 8730
rect 26324 8678 26376 8730
rect 26388 8678 26440 8730
rect 34526 8678 34578 8730
rect 34590 8678 34642 8730
rect 34654 8678 34706 8730
rect 34718 8678 34770 8730
rect 34782 8678 34834 8730
rect 15752 8576 15804 8628
rect 16488 8576 16540 8628
rect 17316 8576 17368 8628
rect 17592 8576 17644 8628
rect 18972 8508 19024 8560
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 21916 8576 21968 8628
rect 18236 8440 18288 8492
rect 21824 8508 21876 8560
rect 18052 8372 18104 8424
rect 20996 8440 21048 8492
rect 21456 8440 21508 8492
rect 22560 8440 22612 8492
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 25596 8576 25648 8628
rect 26608 8508 26660 8560
rect 29000 8576 29052 8628
rect 29828 8619 29880 8628
rect 29828 8585 29837 8619
rect 29837 8585 29871 8619
rect 29871 8585 29880 8619
rect 29828 8576 29880 8585
rect 33048 8576 33100 8628
rect 31484 8508 31536 8560
rect 23480 8483 23532 8492
rect 23480 8449 23489 8483
rect 23489 8449 23523 8483
rect 23523 8449 23532 8483
rect 23480 8440 23532 8449
rect 24860 8440 24912 8492
rect 26056 8440 26108 8492
rect 26516 8440 26568 8492
rect 30840 8440 30892 8492
rect 31392 8483 31444 8492
rect 31392 8449 31401 8483
rect 31401 8449 31435 8483
rect 31435 8449 31444 8483
rect 31392 8440 31444 8449
rect 32956 8508 33008 8560
rect 23756 8415 23808 8424
rect 23756 8381 23765 8415
rect 23765 8381 23799 8415
rect 23799 8381 23808 8415
rect 23756 8372 23808 8381
rect 24952 8372 25004 8424
rect 27620 8372 27672 8424
rect 28356 8415 28408 8424
rect 28356 8381 28365 8415
rect 28365 8381 28399 8415
rect 28399 8381 28408 8415
rect 28356 8372 28408 8381
rect 31024 8372 31076 8424
rect 31576 8372 31628 8424
rect 19248 8236 19300 8288
rect 21732 8304 21784 8356
rect 22376 8304 22428 8356
rect 23480 8304 23532 8356
rect 27712 8304 27764 8356
rect 34796 8304 34848 8356
rect 20444 8236 20496 8288
rect 22928 8279 22980 8288
rect 22928 8245 22937 8279
rect 22937 8245 22971 8279
rect 22971 8245 22980 8279
rect 22928 8236 22980 8245
rect 27068 8279 27120 8288
rect 27068 8245 27077 8279
rect 27077 8245 27111 8279
rect 27111 8245 27120 8279
rect 27068 8236 27120 8245
rect 31484 8236 31536 8288
rect 34060 8236 34112 8288
rect 5147 8134 5199 8186
rect 5211 8134 5263 8186
rect 5275 8134 5327 8186
rect 5339 8134 5391 8186
rect 5403 8134 5455 8186
rect 13541 8134 13593 8186
rect 13605 8134 13657 8186
rect 13669 8134 13721 8186
rect 13733 8134 13785 8186
rect 13797 8134 13849 8186
rect 21935 8134 21987 8186
rect 21999 8134 22051 8186
rect 22063 8134 22115 8186
rect 22127 8134 22179 8186
rect 22191 8134 22243 8186
rect 30329 8134 30381 8186
rect 30393 8134 30445 8186
rect 30457 8134 30509 8186
rect 30521 8134 30573 8186
rect 30585 8134 30637 8186
rect 13912 8075 13964 8084
rect 13912 8041 13921 8075
rect 13921 8041 13955 8075
rect 13955 8041 13964 8075
rect 13912 8032 13964 8041
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 17224 8032 17276 8084
rect 17592 8032 17644 8084
rect 19892 8032 19944 8084
rect 23112 8032 23164 8084
rect 17408 7964 17460 8016
rect 18236 7964 18288 8016
rect 19708 7964 19760 8016
rect 12164 7939 12216 7948
rect 12164 7905 12173 7939
rect 12173 7905 12207 7939
rect 12207 7905 12216 7939
rect 12164 7896 12216 7905
rect 17316 7896 17368 7948
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 16212 7828 16264 7880
rect 17500 7828 17552 7880
rect 19616 7896 19668 7948
rect 22284 7939 22336 7948
rect 22284 7905 22293 7939
rect 22293 7905 22327 7939
rect 22327 7905 22336 7939
rect 22284 7896 22336 7905
rect 22652 7896 22704 7948
rect 23480 7896 23532 7948
rect 24952 7896 25004 7948
rect 28356 8032 28408 8084
rect 31392 8032 31444 8084
rect 12440 7803 12492 7812
rect 12440 7769 12449 7803
rect 12449 7769 12483 7803
rect 12483 7769 12492 7803
rect 12440 7760 12492 7769
rect 13912 7760 13964 7812
rect 16396 7760 16448 7812
rect 17500 7735 17552 7744
rect 17500 7701 17509 7735
rect 17509 7701 17543 7735
rect 17543 7701 17552 7735
rect 17500 7692 17552 7701
rect 18972 7828 19024 7880
rect 18052 7803 18104 7812
rect 18052 7769 18061 7803
rect 18061 7769 18095 7803
rect 18095 7769 18104 7803
rect 18052 7760 18104 7769
rect 18788 7760 18840 7812
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 23756 7871 23808 7880
rect 23756 7837 23765 7871
rect 23765 7837 23799 7871
rect 23799 7837 23808 7871
rect 27068 7896 27120 7948
rect 27160 7896 27212 7948
rect 27896 7896 27948 7948
rect 28448 7939 28500 7948
rect 28448 7905 28457 7939
rect 28457 7905 28491 7939
rect 28491 7905 28500 7939
rect 28448 7896 28500 7905
rect 34060 7939 34112 7948
rect 34060 7905 34069 7939
rect 34069 7905 34103 7939
rect 34103 7905 34112 7939
rect 34060 7896 34112 7905
rect 23756 7828 23808 7837
rect 27252 7871 27304 7880
rect 27252 7837 27253 7871
rect 27253 7837 27287 7871
rect 27287 7837 27304 7871
rect 27252 7828 27304 7837
rect 27712 7828 27764 7880
rect 28540 7871 28592 7880
rect 28540 7837 28549 7871
rect 28549 7837 28583 7871
rect 28583 7837 28592 7871
rect 28540 7828 28592 7837
rect 28724 7871 28776 7880
rect 28724 7837 28733 7871
rect 28733 7837 28767 7871
rect 28767 7837 28776 7871
rect 28724 7828 28776 7837
rect 32956 7828 33008 7880
rect 34336 7871 34388 7880
rect 34336 7837 34345 7871
rect 34345 7837 34379 7871
rect 34379 7837 34388 7871
rect 34336 7828 34388 7837
rect 27804 7760 27856 7812
rect 29736 7760 29788 7812
rect 31300 7760 31352 7812
rect 19800 7735 19852 7744
rect 19800 7701 19809 7735
rect 19809 7701 19843 7735
rect 19843 7701 19852 7735
rect 19800 7692 19852 7701
rect 19892 7735 19944 7744
rect 19892 7701 19901 7735
rect 19901 7701 19935 7735
rect 19935 7701 19944 7735
rect 19892 7692 19944 7701
rect 21456 7692 21508 7744
rect 21640 7692 21692 7744
rect 24400 7735 24452 7744
rect 24400 7701 24409 7735
rect 24409 7701 24443 7735
rect 24443 7701 24452 7735
rect 24400 7692 24452 7701
rect 24768 7735 24820 7744
rect 24768 7701 24777 7735
rect 24777 7701 24811 7735
rect 24811 7701 24820 7735
rect 24768 7692 24820 7701
rect 26976 7735 27028 7744
rect 26976 7701 26985 7735
rect 26985 7701 27019 7735
rect 27019 7701 27028 7735
rect 26976 7692 27028 7701
rect 27068 7735 27120 7744
rect 27068 7701 27077 7735
rect 27077 7701 27111 7735
rect 27111 7701 27120 7735
rect 27068 7692 27120 7701
rect 30840 7735 30892 7744
rect 30840 7701 30865 7735
rect 30865 7701 30892 7735
rect 30840 7692 30892 7701
rect 9344 7590 9396 7642
rect 9408 7590 9460 7642
rect 9472 7590 9524 7642
rect 9536 7590 9588 7642
rect 9600 7590 9652 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 17930 7590 17982 7642
rect 17994 7590 18046 7642
rect 26132 7590 26184 7642
rect 26196 7590 26248 7642
rect 26260 7590 26312 7642
rect 26324 7590 26376 7642
rect 26388 7590 26440 7642
rect 34526 7590 34578 7642
rect 34590 7590 34642 7642
rect 34654 7590 34706 7642
rect 34718 7590 34770 7642
rect 34782 7590 34834 7642
rect 12440 7488 12492 7540
rect 13912 7420 13964 7472
rect 14832 7420 14884 7472
rect 15844 7488 15896 7540
rect 16396 7488 16448 7540
rect 16672 7488 16724 7540
rect 17408 7488 17460 7540
rect 18972 7488 19024 7540
rect 19708 7488 19760 7540
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 12164 7284 12216 7336
rect 13268 7284 13320 7336
rect 13360 7284 13412 7336
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 16212 7352 16264 7404
rect 16120 7284 16172 7336
rect 18236 7352 18288 7404
rect 18420 7352 18472 7404
rect 19248 7420 19300 7472
rect 18972 7395 19024 7404
rect 18972 7361 18981 7395
rect 18981 7361 19015 7395
rect 19015 7361 19024 7395
rect 18972 7352 19024 7361
rect 20444 7488 20496 7540
rect 21640 7531 21692 7540
rect 21640 7497 21649 7531
rect 21649 7497 21683 7531
rect 21683 7497 21692 7531
rect 21640 7488 21692 7497
rect 22100 7420 22152 7472
rect 22928 7488 22980 7540
rect 23756 7488 23808 7540
rect 24400 7488 24452 7540
rect 24768 7488 24820 7540
rect 19248 7284 19300 7336
rect 19616 7216 19668 7268
rect 16028 7148 16080 7200
rect 17408 7191 17460 7200
rect 17408 7157 17417 7191
rect 17417 7157 17451 7191
rect 17451 7157 17460 7191
rect 17408 7148 17460 7157
rect 19524 7148 19576 7200
rect 22192 7284 22244 7336
rect 23756 7352 23808 7404
rect 24216 7352 24268 7404
rect 26976 7488 27028 7540
rect 27252 7488 27304 7540
rect 31852 7531 31904 7540
rect 31852 7497 31861 7531
rect 31861 7497 31895 7531
rect 31895 7497 31904 7531
rect 31852 7488 31904 7497
rect 30840 7420 30892 7472
rect 22284 7148 22336 7200
rect 24860 7148 24912 7200
rect 31484 7395 31536 7404
rect 31484 7361 31493 7395
rect 31493 7361 31527 7395
rect 31527 7361 31536 7395
rect 31484 7352 31536 7361
rect 31576 7327 31628 7336
rect 31576 7293 31585 7327
rect 31585 7293 31619 7327
rect 31619 7293 31628 7327
rect 31576 7284 31628 7293
rect 29828 7148 29880 7200
rect 32588 7216 32640 7268
rect 30932 7148 30984 7200
rect 31484 7191 31536 7200
rect 31484 7157 31493 7191
rect 31493 7157 31527 7191
rect 31527 7157 31536 7191
rect 31484 7148 31536 7157
rect 5147 7046 5199 7098
rect 5211 7046 5263 7098
rect 5275 7046 5327 7098
rect 5339 7046 5391 7098
rect 5403 7046 5455 7098
rect 13541 7046 13593 7098
rect 13605 7046 13657 7098
rect 13669 7046 13721 7098
rect 13733 7046 13785 7098
rect 13797 7046 13849 7098
rect 21935 7046 21987 7098
rect 21999 7046 22051 7098
rect 22063 7046 22115 7098
rect 22127 7046 22179 7098
rect 22191 7046 22243 7098
rect 30329 7046 30381 7098
rect 30393 7046 30445 7098
rect 30457 7046 30509 7098
rect 30521 7046 30573 7098
rect 30585 7046 30637 7098
rect 7932 6944 7984 6996
rect 16396 6944 16448 6996
rect 17408 6944 17460 6996
rect 18420 6944 18472 6996
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 27068 6944 27120 6996
rect 27804 6987 27856 6996
rect 27804 6953 27813 6987
rect 27813 6953 27847 6987
rect 27847 6953 27856 6987
rect 27804 6944 27856 6953
rect 31024 6987 31076 6996
rect 31024 6953 31033 6987
rect 31033 6953 31067 6987
rect 31067 6953 31076 6987
rect 31024 6944 31076 6953
rect 16120 6851 16172 6860
rect 16120 6817 16129 6851
rect 16129 6817 16163 6851
rect 16163 6817 16172 6851
rect 16120 6808 16172 6817
rect 19800 6919 19852 6928
rect 19800 6885 19809 6919
rect 19809 6885 19843 6919
rect 19843 6885 19852 6919
rect 19800 6876 19852 6885
rect 2688 6740 2740 6792
rect 3240 6740 3292 6792
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 19892 6740 19944 6792
rect 26056 6851 26108 6860
rect 26056 6817 26065 6851
rect 26065 6817 26099 6851
rect 26099 6817 26108 6851
rect 26056 6808 26108 6817
rect 26976 6808 27028 6860
rect 27528 6808 27580 6860
rect 23572 6783 23624 6792
rect 23572 6749 23581 6783
rect 23581 6749 23615 6783
rect 23615 6749 23624 6783
rect 23572 6740 23624 6749
rect 29920 6808 29972 6860
rect 32404 6851 32456 6860
rect 32404 6817 32413 6851
rect 32413 6817 32447 6851
rect 32447 6817 32456 6851
rect 32404 6808 32456 6817
rect 32588 6851 32640 6860
rect 32588 6817 32597 6851
rect 32597 6817 32631 6851
rect 32631 6817 32640 6851
rect 32588 6808 32640 6817
rect 30748 6783 30800 6792
rect 30748 6749 30757 6783
rect 30757 6749 30791 6783
rect 30791 6749 30800 6783
rect 30748 6740 30800 6749
rect 30840 6783 30892 6792
rect 30840 6749 30849 6783
rect 30849 6749 30883 6783
rect 30883 6749 30892 6783
rect 30840 6740 30892 6749
rect 31576 6740 31628 6792
rect 1676 6715 1728 6724
rect 1676 6681 1685 6715
rect 1685 6681 1719 6715
rect 1719 6681 1728 6715
rect 1676 6672 1728 6681
rect 15200 6672 15252 6724
rect 16212 6715 16264 6724
rect 16212 6681 16221 6715
rect 16221 6681 16255 6715
rect 16255 6681 16264 6715
rect 16212 6672 16264 6681
rect 19156 6672 19208 6724
rect 19984 6672 20036 6724
rect 26608 6672 26660 6724
rect 28816 6672 28868 6724
rect 15568 6604 15620 6656
rect 19340 6604 19392 6656
rect 23388 6647 23440 6656
rect 23388 6613 23397 6647
rect 23397 6613 23431 6647
rect 23431 6613 23440 6647
rect 23388 6604 23440 6613
rect 29644 6647 29696 6656
rect 29644 6613 29653 6647
rect 29653 6613 29687 6647
rect 29687 6613 29696 6647
rect 29644 6604 29696 6613
rect 30196 6672 30248 6724
rect 30932 6672 30984 6724
rect 33048 6647 33100 6656
rect 33048 6613 33057 6647
rect 33057 6613 33091 6647
rect 33091 6613 33100 6647
rect 33048 6604 33100 6613
rect 9344 6502 9396 6554
rect 9408 6502 9460 6554
rect 9472 6502 9524 6554
rect 9536 6502 9588 6554
rect 9600 6502 9652 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 17930 6502 17982 6554
rect 17994 6502 18046 6554
rect 26132 6502 26184 6554
rect 26196 6502 26248 6554
rect 26260 6502 26312 6554
rect 26324 6502 26376 6554
rect 26388 6502 26440 6554
rect 34526 6502 34578 6554
rect 34590 6502 34642 6554
rect 34654 6502 34706 6554
rect 34718 6502 34770 6554
rect 34782 6502 34834 6554
rect 1676 6400 1728 6452
rect 3240 6332 3292 6384
rect 10692 6400 10744 6452
rect 11796 6375 11848 6384
rect 11796 6341 11805 6375
rect 11805 6341 11839 6375
rect 11839 6341 11848 6375
rect 11796 6332 11848 6341
rect 13268 6400 13320 6452
rect 13360 6332 13412 6384
rect 940 6264 992 6316
rect 2688 6264 2740 6316
rect 14556 6400 14608 6452
rect 15200 6443 15252 6452
rect 15200 6409 15209 6443
rect 15209 6409 15243 6443
rect 15243 6409 15252 6443
rect 15200 6400 15252 6409
rect 19156 6400 19208 6452
rect 19340 6400 19392 6452
rect 22468 6400 22520 6452
rect 23572 6400 23624 6452
rect 27344 6400 27396 6452
rect 29552 6443 29604 6452
rect 18972 6332 19024 6384
rect 19064 6375 19116 6384
rect 19064 6341 19073 6375
rect 19073 6341 19107 6375
rect 19107 6341 19116 6375
rect 19064 6332 19116 6341
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 12808 6196 12860 6248
rect 14832 6264 14884 6316
rect 29552 6409 29561 6443
rect 29561 6409 29595 6443
rect 29595 6409 29604 6443
rect 29552 6400 29604 6409
rect 29736 6443 29788 6452
rect 29736 6409 29745 6443
rect 29745 6409 29779 6443
rect 29779 6409 29788 6443
rect 29736 6400 29788 6409
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 22468 6264 22520 6316
rect 14096 6196 14148 6248
rect 22652 6239 22704 6248
rect 22652 6205 22661 6239
rect 22661 6205 22695 6239
rect 22695 6205 22704 6239
rect 22652 6196 22704 6205
rect 24952 6196 25004 6248
rect 25872 6239 25924 6248
rect 25872 6205 25881 6239
rect 25881 6205 25915 6239
rect 25915 6205 25924 6239
rect 25872 6196 25924 6205
rect 27344 6196 27396 6248
rect 27804 6332 27856 6384
rect 30748 6400 30800 6452
rect 31760 6400 31812 6452
rect 27528 6307 27580 6316
rect 27528 6273 27537 6307
rect 27537 6273 27571 6307
rect 27571 6273 27580 6307
rect 27528 6264 27580 6273
rect 29920 6307 29972 6316
rect 29920 6273 29929 6307
rect 29929 6273 29963 6307
rect 29963 6273 29972 6307
rect 29920 6264 29972 6273
rect 13268 6103 13320 6112
rect 13268 6069 13277 6103
rect 13277 6069 13311 6103
rect 13311 6069 13320 6103
rect 13268 6060 13320 6069
rect 19524 6103 19576 6112
rect 19524 6069 19533 6103
rect 19533 6069 19567 6103
rect 19567 6069 19576 6103
rect 19524 6060 19576 6069
rect 20260 6060 20312 6112
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 24124 6060 24176 6112
rect 26792 6128 26844 6180
rect 27896 6128 27948 6180
rect 29828 6196 29880 6248
rect 30196 6307 30248 6316
rect 30196 6273 30205 6307
rect 30205 6273 30239 6307
rect 30239 6273 30248 6307
rect 30196 6264 30248 6273
rect 30104 6196 30156 6248
rect 30380 6307 30432 6316
rect 30380 6273 30389 6307
rect 30389 6273 30423 6307
rect 30423 6273 30432 6307
rect 30380 6264 30432 6273
rect 24860 6103 24912 6112
rect 24860 6069 24869 6103
rect 24869 6069 24903 6103
rect 24903 6069 24912 6103
rect 24860 6060 24912 6069
rect 25320 6103 25372 6112
rect 25320 6069 25329 6103
rect 25329 6069 25363 6103
rect 25363 6069 25372 6103
rect 25320 6060 25372 6069
rect 27804 6103 27856 6112
rect 27804 6069 27813 6103
rect 27813 6069 27847 6103
rect 27847 6069 27856 6103
rect 27804 6060 27856 6069
rect 29368 6171 29420 6180
rect 29368 6137 29377 6171
rect 29377 6137 29411 6171
rect 29411 6137 29420 6171
rect 29368 6128 29420 6137
rect 32496 6332 32548 6384
rect 32128 6264 32180 6316
rect 32956 6264 33008 6316
rect 34336 6307 34388 6316
rect 34336 6273 34345 6307
rect 34345 6273 34379 6307
rect 34379 6273 34388 6307
rect 34336 6264 34388 6273
rect 34060 6239 34112 6248
rect 34060 6205 34069 6239
rect 34069 6205 34103 6239
rect 34103 6205 34112 6239
rect 34060 6196 34112 6205
rect 5147 5958 5199 6010
rect 5211 5958 5263 6010
rect 5275 5958 5327 6010
rect 5339 5958 5391 6010
rect 5403 5958 5455 6010
rect 13541 5958 13593 6010
rect 13605 5958 13657 6010
rect 13669 5958 13721 6010
rect 13733 5958 13785 6010
rect 13797 5958 13849 6010
rect 21935 5958 21987 6010
rect 21999 5958 22051 6010
rect 22063 5958 22115 6010
rect 22127 5958 22179 6010
rect 22191 5958 22243 6010
rect 30329 5958 30381 6010
rect 30393 5958 30445 6010
rect 30457 5958 30509 6010
rect 30521 5958 30573 6010
rect 30585 5958 30637 6010
rect 13268 5856 13320 5908
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 20536 5856 20588 5908
rect 21824 5856 21876 5908
rect 22560 5856 22612 5908
rect 23388 5856 23440 5908
rect 26700 5899 26752 5908
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 19524 5763 19576 5772
rect 19524 5729 19533 5763
rect 19533 5729 19567 5763
rect 19567 5729 19576 5763
rect 19524 5720 19576 5729
rect 26700 5865 26709 5899
rect 26709 5865 26743 5899
rect 26743 5865 26752 5899
rect 26700 5856 26752 5865
rect 29368 5856 29420 5908
rect 29644 5856 29696 5908
rect 29828 5856 29880 5908
rect 30196 5856 30248 5908
rect 31760 5856 31812 5908
rect 34060 5856 34112 5908
rect 24768 5788 24820 5840
rect 22284 5720 22336 5772
rect 24216 5720 24268 5772
rect 25320 5720 25372 5772
rect 26608 5720 26660 5772
rect 27620 5720 27672 5772
rect 28816 5720 28868 5772
rect 17132 5584 17184 5636
rect 19984 5584 20036 5636
rect 21456 5584 21508 5636
rect 21824 5559 21876 5568
rect 21824 5525 21833 5559
rect 21833 5525 21867 5559
rect 21867 5525 21876 5559
rect 21824 5516 21876 5525
rect 23756 5584 23808 5636
rect 23480 5516 23532 5568
rect 24124 5516 24176 5568
rect 26700 5584 26752 5636
rect 27896 5627 27948 5636
rect 27896 5593 27905 5627
rect 27905 5593 27939 5627
rect 27939 5593 27948 5627
rect 27896 5584 27948 5593
rect 31852 5695 31904 5704
rect 31852 5661 31861 5695
rect 31861 5661 31895 5695
rect 31895 5661 31904 5695
rect 31852 5652 31904 5661
rect 26884 5516 26936 5568
rect 27804 5559 27856 5568
rect 27804 5525 27813 5559
rect 27813 5525 27847 5559
rect 27847 5525 27856 5559
rect 27804 5516 27856 5525
rect 30380 5516 30432 5568
rect 31116 5516 31168 5568
rect 32496 5652 32548 5704
rect 33048 5652 33100 5704
rect 9344 5414 9396 5466
rect 9408 5414 9460 5466
rect 9472 5414 9524 5466
rect 9536 5414 9588 5466
rect 9600 5414 9652 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 17930 5414 17982 5466
rect 17994 5414 18046 5466
rect 26132 5414 26184 5466
rect 26196 5414 26248 5466
rect 26260 5414 26312 5466
rect 26324 5414 26376 5466
rect 26388 5414 26440 5466
rect 34526 5414 34578 5466
rect 34590 5414 34642 5466
rect 34654 5414 34706 5466
rect 34718 5414 34770 5466
rect 34782 5414 34834 5466
rect 19984 5312 20036 5364
rect 15752 5244 15804 5296
rect 17132 5244 17184 5296
rect 20260 5244 20312 5296
rect 12808 5176 12860 5228
rect 14832 5176 14884 5228
rect 16488 5219 16540 5228
rect 16488 5185 16497 5219
rect 16497 5185 16531 5219
rect 16531 5185 16540 5219
rect 16488 5176 16540 5185
rect 13176 5151 13228 5160
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 15752 5108 15804 5160
rect 16212 5151 16264 5160
rect 16212 5117 16221 5151
rect 16221 5117 16255 5151
rect 16255 5117 16264 5151
rect 16212 5108 16264 5117
rect 19892 5151 19944 5160
rect 19892 5117 19901 5151
rect 19901 5117 19935 5151
rect 19935 5117 19944 5151
rect 19892 5108 19944 5117
rect 21180 5108 21232 5160
rect 22468 5312 22520 5364
rect 23480 5312 23532 5364
rect 24860 5312 24912 5364
rect 24952 5312 25004 5364
rect 21456 5244 21508 5296
rect 25872 5312 25924 5364
rect 26792 5312 26844 5364
rect 26884 5312 26936 5364
rect 23664 5219 23716 5228
rect 23664 5185 23673 5219
rect 23673 5185 23707 5219
rect 23707 5185 23716 5219
rect 23664 5176 23716 5185
rect 22560 5108 22612 5160
rect 23756 5040 23808 5092
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 24860 5219 24912 5228
rect 24860 5185 24870 5219
rect 24870 5185 24904 5219
rect 24904 5185 24912 5219
rect 24860 5176 24912 5185
rect 25044 5219 25096 5228
rect 25044 5185 25053 5219
rect 25053 5185 25087 5219
rect 25087 5185 25096 5219
rect 25044 5176 25096 5185
rect 25228 5219 25280 5228
rect 25228 5185 25242 5219
rect 25242 5185 25276 5219
rect 25276 5185 25280 5219
rect 25228 5176 25280 5185
rect 28540 5312 28592 5364
rect 30380 5312 30432 5364
rect 31484 5312 31536 5364
rect 27160 5219 27212 5228
rect 27160 5185 27169 5219
rect 27169 5185 27203 5219
rect 27203 5185 27212 5219
rect 27160 5176 27212 5185
rect 28908 5219 28960 5228
rect 28908 5185 28917 5219
rect 28917 5185 28951 5219
rect 28951 5185 28960 5219
rect 28908 5176 28960 5185
rect 30656 5219 30708 5228
rect 30656 5185 30665 5219
rect 30665 5185 30699 5219
rect 30699 5185 30708 5219
rect 30656 5176 30708 5185
rect 28816 5108 28868 5160
rect 29368 5108 29420 5160
rect 30196 5108 30248 5160
rect 26792 5083 26844 5092
rect 26792 5049 26801 5083
rect 26801 5049 26835 5083
rect 26835 5049 26844 5083
rect 26792 5040 26844 5049
rect 27344 5040 27396 5092
rect 29920 5040 29972 5092
rect 30196 4972 30248 5024
rect 5147 4870 5199 4922
rect 5211 4870 5263 4922
rect 5275 4870 5327 4922
rect 5339 4870 5391 4922
rect 5403 4870 5455 4922
rect 13541 4870 13593 4922
rect 13605 4870 13657 4922
rect 13669 4870 13721 4922
rect 13733 4870 13785 4922
rect 13797 4870 13849 4922
rect 21935 4870 21987 4922
rect 21999 4870 22051 4922
rect 22063 4870 22115 4922
rect 22127 4870 22179 4922
rect 22191 4870 22243 4922
rect 30329 4870 30381 4922
rect 30393 4870 30445 4922
rect 30457 4870 30509 4922
rect 30521 4870 30573 4922
rect 30585 4870 30637 4922
rect 13176 4768 13228 4820
rect 16212 4768 16264 4820
rect 23664 4811 23716 4820
rect 23664 4777 23673 4811
rect 23673 4777 23707 4811
rect 23707 4777 23716 4811
rect 23664 4768 23716 4777
rect 25044 4768 25096 4820
rect 27344 4768 27396 4820
rect 28908 4768 28960 4820
rect 21180 4632 21232 4684
rect 22284 4632 22336 4684
rect 25228 4700 25280 4752
rect 27160 4700 27212 4752
rect 29368 4743 29420 4752
rect 29368 4709 29377 4743
rect 29377 4709 29411 4743
rect 29411 4709 29420 4743
rect 29368 4700 29420 4709
rect 30104 4768 30156 4820
rect 30656 4768 30708 4820
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 14648 4607 14700 4616
rect 14648 4573 14657 4607
rect 14657 4573 14691 4607
rect 14691 4573 14700 4607
rect 14648 4564 14700 4573
rect 18144 4607 18196 4616
rect 18144 4573 18153 4607
rect 18153 4573 18187 4607
rect 18187 4573 18196 4607
rect 18144 4564 18196 4573
rect 21824 4564 21876 4616
rect 23756 4564 23808 4616
rect 24492 4564 24544 4616
rect 14372 4428 14424 4480
rect 16764 4428 16816 4480
rect 19432 4428 19484 4480
rect 23480 4496 23532 4548
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 25964 4428 26016 4480
rect 9344 4326 9396 4378
rect 9408 4326 9460 4378
rect 9472 4326 9524 4378
rect 9536 4326 9588 4378
rect 9600 4326 9652 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 17930 4326 17982 4378
rect 17994 4326 18046 4378
rect 26132 4326 26184 4378
rect 26196 4326 26248 4378
rect 26260 4326 26312 4378
rect 26324 4326 26376 4378
rect 26388 4326 26440 4378
rect 34526 4326 34578 4378
rect 34590 4326 34642 4378
rect 34654 4326 34706 4378
rect 34718 4326 34770 4378
rect 34782 4326 34834 4378
rect 12808 4224 12860 4276
rect 14648 4224 14700 4276
rect 23480 4224 23532 4276
rect 24400 4224 24452 4276
rect 25964 4267 26016 4276
rect 25964 4233 25973 4267
rect 25973 4233 26007 4267
rect 26007 4233 26016 4267
rect 25964 4224 26016 4233
rect 14372 4156 14424 4208
rect 17132 4156 17184 4208
rect 19984 4156 20036 4208
rect 19892 4088 19944 4140
rect 24492 4156 24544 4208
rect 26608 4156 26660 4208
rect 26792 4156 26844 4208
rect 28908 4224 28960 4276
rect 30196 4267 30248 4276
rect 30196 4233 30205 4267
rect 30205 4233 30239 4267
rect 30239 4233 30248 4267
rect 30196 4224 30248 4233
rect 32128 4156 32180 4208
rect 12164 4063 12216 4072
rect 12164 4029 12173 4063
rect 12173 4029 12207 4063
rect 12207 4029 12216 4063
rect 12164 4020 12216 4029
rect 12808 4020 12860 4072
rect 13820 4020 13872 4072
rect 15660 4063 15712 4072
rect 15660 4029 15669 4063
rect 15669 4029 15703 4063
rect 15703 4029 15712 4063
rect 15660 4020 15712 4029
rect 16488 4020 16540 4072
rect 18236 4020 18288 4072
rect 19432 4063 19484 4072
rect 19432 4029 19441 4063
rect 19441 4029 19475 4063
rect 19475 4029 19484 4063
rect 19432 4020 19484 4029
rect 24216 4131 24268 4140
rect 24216 4097 24225 4131
rect 24225 4097 24259 4131
rect 24259 4097 24268 4131
rect 24216 4088 24268 4097
rect 26976 4131 27028 4140
rect 26976 4097 26985 4131
rect 26985 4097 27019 4131
rect 27019 4097 27028 4131
rect 26976 4088 27028 4097
rect 34336 4088 34388 4140
rect 22376 4020 22428 4072
rect 31668 4063 31720 4072
rect 31668 4029 31677 4063
rect 31677 4029 31711 4063
rect 31711 4029 31720 4063
rect 31668 4020 31720 4029
rect 5147 3782 5199 3834
rect 5211 3782 5263 3834
rect 5275 3782 5327 3834
rect 5339 3782 5391 3834
rect 5403 3782 5455 3834
rect 13541 3782 13593 3834
rect 13605 3782 13657 3834
rect 13669 3782 13721 3834
rect 13733 3782 13785 3834
rect 13797 3782 13849 3834
rect 21935 3782 21987 3834
rect 21999 3782 22051 3834
rect 22063 3782 22115 3834
rect 22127 3782 22179 3834
rect 22191 3782 22243 3834
rect 30329 3782 30381 3834
rect 30393 3782 30445 3834
rect 30457 3782 30509 3834
rect 30521 3782 30573 3834
rect 30585 3782 30637 3834
rect 18144 3680 18196 3732
rect 19340 3544 19392 3596
rect 17132 3476 17184 3528
rect 24584 3408 24636 3460
rect 9344 3238 9396 3290
rect 9408 3238 9460 3290
rect 9472 3238 9524 3290
rect 9536 3238 9588 3290
rect 9600 3238 9652 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 17930 3238 17982 3290
rect 17994 3238 18046 3290
rect 26132 3238 26184 3290
rect 26196 3238 26248 3290
rect 26260 3238 26312 3290
rect 26324 3238 26376 3290
rect 26388 3238 26440 3290
rect 34526 3238 34578 3290
rect 34590 3238 34642 3290
rect 34654 3238 34706 3290
rect 34718 3238 34770 3290
rect 34782 3238 34834 3290
rect 5147 2694 5199 2746
rect 5211 2694 5263 2746
rect 5275 2694 5327 2746
rect 5339 2694 5391 2746
rect 5403 2694 5455 2746
rect 13541 2694 13593 2746
rect 13605 2694 13657 2746
rect 13669 2694 13721 2746
rect 13733 2694 13785 2746
rect 13797 2694 13849 2746
rect 21935 2694 21987 2746
rect 21999 2694 22051 2746
rect 22063 2694 22115 2746
rect 22127 2694 22179 2746
rect 22191 2694 22243 2746
rect 30329 2694 30381 2746
rect 30393 2694 30445 2746
rect 30457 2694 30509 2746
rect 30521 2694 30573 2746
rect 30585 2694 30637 2746
rect 7472 2592 7524 2644
rect 12164 2592 12216 2644
rect 24584 2635 24636 2644
rect 24584 2601 24593 2635
rect 24593 2601 24627 2635
rect 24627 2601 24636 2635
rect 24584 2592 24636 2601
rect 31668 2592 31720 2644
rect 15660 2456 15712 2508
rect 20 2388 72 2440
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 12256 2388 12308 2440
rect 16948 2388 17000 2440
rect 24492 2388 24544 2440
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 11796 2252 11848 2304
rect 19064 2252 19116 2304
rect 34428 2252 34480 2304
rect 9344 2150 9396 2202
rect 9408 2150 9460 2202
rect 9472 2150 9524 2202
rect 9536 2150 9588 2202
rect 9600 2150 9652 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
rect 17930 2150 17982 2202
rect 17994 2150 18046 2202
rect 26132 2150 26184 2202
rect 26196 2150 26248 2202
rect 26260 2150 26312 2202
rect 26324 2150 26376 2202
rect 26388 2150 26440 2202
rect 34526 2150 34578 2202
rect 34590 2150 34642 2202
rect 34654 2150 34706 2202
rect 34718 2150 34770 2202
rect 34782 2150 34834 2202
<< metal2 >>
rect 1306 37217 1362 38017
rect 7746 37217 7802 38017
rect 13542 37346 13598 38017
rect 13542 37318 13768 37346
rect 13542 37217 13598 37318
rect 1320 35290 1348 37217
rect 5147 35388 5455 35397
rect 5147 35386 5153 35388
rect 5209 35386 5233 35388
rect 5289 35386 5313 35388
rect 5369 35386 5393 35388
rect 5449 35386 5455 35388
rect 5209 35334 5211 35386
rect 5391 35334 5393 35386
rect 5147 35332 5153 35334
rect 5209 35332 5233 35334
rect 5289 35332 5313 35334
rect 5369 35332 5393 35334
rect 5449 35332 5455 35334
rect 5147 35323 5455 35332
rect 1308 35284 1360 35290
rect 1308 35226 1360 35232
rect 7760 35086 7788 37217
rect 13740 35850 13768 37318
rect 19982 37217 20038 38017
rect 26422 37217 26478 38017
rect 32862 37217 32918 38017
rect 13740 35822 13952 35850
rect 13541 35388 13849 35397
rect 13541 35386 13547 35388
rect 13603 35386 13627 35388
rect 13683 35386 13707 35388
rect 13763 35386 13787 35388
rect 13843 35386 13849 35388
rect 13603 35334 13605 35386
rect 13785 35334 13787 35386
rect 13541 35332 13547 35334
rect 13603 35332 13627 35334
rect 13683 35332 13707 35334
rect 13763 35332 13787 35334
rect 13843 35332 13849 35334
rect 13541 35323 13849 35332
rect 9220 35216 9272 35222
rect 9220 35158 9272 35164
rect 7748 35080 7800 35086
rect 7748 35022 7800 35028
rect 8116 35080 8168 35086
rect 8116 35022 8168 35028
rect 1768 35012 1820 35018
rect 1768 34954 1820 34960
rect 940 32904 992 32910
rect 940 32846 992 32852
rect 952 32745 980 32846
rect 938 32736 994 32745
rect 938 32671 994 32680
rect 1400 26308 1452 26314
rect 1400 26250 1452 26256
rect 1412 26217 1440 26250
rect 1398 26208 1454 26217
rect 1398 26143 1454 26152
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 940 19848 992 19854
rect 938 19816 940 19825
rect 992 19816 994 19825
rect 938 19751 994 19760
rect 1412 19378 1440 20334
rect 1780 20074 1808 34954
rect 7932 34944 7984 34950
rect 7932 34886 7984 34892
rect 7944 34678 7972 34886
rect 7932 34672 7984 34678
rect 7932 34614 7984 34620
rect 5724 34604 5776 34610
rect 5724 34546 5776 34552
rect 3608 34536 3660 34542
rect 3608 34478 3660 34484
rect 3516 32768 3568 32774
rect 3516 32710 3568 32716
rect 2136 32360 2188 32366
rect 2136 32302 2188 32308
rect 2148 32026 2176 32302
rect 2780 32224 2832 32230
rect 2780 32166 2832 32172
rect 3528 32178 3556 32710
rect 3620 32366 3648 34478
rect 4620 34400 4672 34406
rect 4620 34342 4672 34348
rect 5632 34400 5684 34406
rect 5632 34342 5684 34348
rect 4632 34202 4660 34342
rect 5147 34300 5455 34309
rect 5147 34298 5153 34300
rect 5209 34298 5233 34300
rect 5289 34298 5313 34300
rect 5369 34298 5393 34300
rect 5449 34298 5455 34300
rect 5209 34246 5211 34298
rect 5391 34246 5393 34298
rect 5147 34244 5153 34246
rect 5209 34244 5233 34246
rect 5289 34244 5313 34246
rect 5369 34244 5393 34246
rect 5449 34244 5455 34246
rect 5147 34235 5455 34244
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 4160 34128 4212 34134
rect 4160 34070 4212 34076
rect 3976 33992 4028 33998
rect 3976 33934 4028 33940
rect 3988 33318 4016 33934
rect 3976 33312 4028 33318
rect 3976 33254 4028 33260
rect 3988 32910 4016 33254
rect 3976 32904 4028 32910
rect 3976 32846 4028 32852
rect 3884 32768 3936 32774
rect 3884 32710 3936 32716
rect 3896 32570 3924 32710
rect 3884 32564 3936 32570
rect 3884 32506 3936 32512
rect 3608 32360 3660 32366
rect 3608 32302 3660 32308
rect 3608 32224 3660 32230
rect 3528 32172 3608 32178
rect 3528 32166 3660 32172
rect 3700 32224 3752 32230
rect 3700 32166 3752 32172
rect 2136 32020 2188 32026
rect 2136 31962 2188 31968
rect 2792 31346 2820 32166
rect 3528 32150 3648 32166
rect 3620 31890 3648 32150
rect 3712 32026 3740 32166
rect 3700 32020 3752 32026
rect 3700 31962 3752 31968
rect 3608 31884 3660 31890
rect 3608 31826 3660 31832
rect 3988 31822 4016 32846
rect 4172 32230 4200 34070
rect 4344 33856 4396 33862
rect 4344 33798 4396 33804
rect 4356 33658 4384 33798
rect 4344 33652 4396 33658
rect 4344 33594 4396 33600
rect 5644 33318 5672 34342
rect 5736 33998 5764 34546
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5724 33992 5776 33998
rect 5724 33934 5776 33940
rect 5632 33312 5684 33318
rect 5632 33254 5684 33260
rect 5147 33212 5455 33221
rect 5147 33210 5153 33212
rect 5209 33210 5233 33212
rect 5289 33210 5313 33212
rect 5369 33210 5393 33212
rect 5449 33210 5455 33212
rect 5209 33158 5211 33210
rect 5391 33158 5393 33210
rect 5147 33156 5153 33158
rect 5209 33156 5233 33158
rect 5289 33156 5313 33158
rect 5369 33156 5393 33158
rect 5449 33156 5455 33158
rect 5147 33147 5455 33156
rect 4896 32768 4948 32774
rect 4896 32710 4948 32716
rect 4344 32496 4396 32502
rect 4344 32438 4396 32444
rect 4160 32224 4212 32230
rect 4160 32166 4212 32172
rect 4252 32224 4304 32230
rect 4252 32166 4304 32172
rect 4264 32026 4292 32166
rect 4252 32020 4304 32026
rect 4252 31962 4304 31968
rect 3976 31816 4028 31822
rect 3976 31758 4028 31764
rect 4356 31414 4384 32438
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4632 32042 4660 32370
rect 4448 32014 4660 32042
rect 4908 32026 4936 32710
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 4896 32020 4948 32026
rect 4448 31754 4476 32014
rect 4896 31962 4948 31968
rect 5000 31754 5028 32166
rect 5147 32124 5455 32133
rect 5147 32122 5153 32124
rect 5209 32122 5233 32124
rect 5289 32122 5313 32124
rect 5369 32122 5393 32124
rect 5449 32122 5455 32124
rect 5209 32070 5211 32122
rect 5391 32070 5393 32122
rect 5147 32068 5153 32070
rect 5209 32068 5233 32070
rect 5289 32068 5313 32070
rect 5369 32068 5393 32070
rect 5449 32068 5455 32070
rect 5147 32059 5455 32068
rect 5540 31816 5592 31822
rect 5540 31758 5592 31764
rect 4436 31748 4488 31754
rect 4436 31690 4488 31696
rect 4988 31748 5040 31754
rect 4988 31690 5040 31696
rect 4448 31482 4476 31690
rect 4804 31680 4856 31686
rect 4804 31622 4856 31628
rect 4436 31476 4488 31482
rect 4436 31418 4488 31424
rect 4344 31408 4396 31414
rect 4344 31350 4396 31356
rect 2780 31340 2832 31346
rect 2780 31282 2832 31288
rect 2792 30734 2820 31282
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 3068 30938 3096 31214
rect 3056 30932 3108 30938
rect 3056 30874 3108 30880
rect 4816 30734 4844 31622
rect 5552 31498 5580 31758
rect 5644 31754 5672 33254
rect 5632 31748 5684 31754
rect 5632 31690 5684 31696
rect 5736 31686 5764 33934
rect 5920 33862 5948 34478
rect 7012 34400 7064 34406
rect 7012 34342 7064 34348
rect 7656 34400 7708 34406
rect 7656 34342 7708 34348
rect 6828 33924 6880 33930
rect 6828 33866 6880 33872
rect 5908 33856 5960 33862
rect 5908 33798 5960 33804
rect 5920 33658 5948 33798
rect 6840 33658 6868 33866
rect 5908 33652 5960 33658
rect 5908 33594 5960 33600
rect 6828 33652 6880 33658
rect 6828 33594 6880 33600
rect 5816 33584 5868 33590
rect 5816 33526 5868 33532
rect 5828 33454 5856 33526
rect 5920 33454 5948 33594
rect 7024 33522 7052 34342
rect 7668 34066 7696 34342
rect 8128 34202 8156 35022
rect 9232 34678 9260 35158
rect 13924 35154 13952 35822
rect 15752 35216 15804 35222
rect 15752 35158 15804 35164
rect 13912 35148 13964 35154
rect 13912 35090 13964 35096
rect 12532 35012 12584 35018
rect 12532 34954 12584 34960
rect 9772 34944 9824 34950
rect 9772 34886 9824 34892
rect 9344 34844 9652 34853
rect 9344 34842 9350 34844
rect 9406 34842 9430 34844
rect 9486 34842 9510 34844
rect 9566 34842 9590 34844
rect 9646 34842 9652 34844
rect 9406 34790 9408 34842
rect 9588 34790 9590 34842
rect 9344 34788 9350 34790
rect 9406 34788 9430 34790
rect 9486 34788 9510 34790
rect 9566 34788 9590 34790
rect 9646 34788 9652 34790
rect 9344 34779 9652 34788
rect 9784 34678 9812 34886
rect 12544 34746 12572 34954
rect 13636 34944 13688 34950
rect 13636 34886 13688 34892
rect 13912 34944 13964 34950
rect 13912 34886 13964 34892
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 13648 34746 13676 34886
rect 12532 34740 12584 34746
rect 12532 34682 12584 34688
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 13924 34678 13952 34886
rect 9220 34672 9272 34678
rect 9220 34614 9272 34620
rect 9588 34672 9640 34678
rect 9588 34614 9640 34620
rect 9772 34672 9824 34678
rect 9772 34614 9824 34620
rect 13912 34672 13964 34678
rect 13912 34614 13964 34620
rect 8944 34400 8996 34406
rect 8944 34342 8996 34348
rect 9404 34400 9456 34406
rect 9404 34342 9456 34348
rect 7932 34196 7984 34202
rect 7932 34138 7984 34144
rect 8116 34196 8168 34202
rect 8116 34138 8168 34144
rect 7656 34060 7708 34066
rect 7656 34002 7708 34008
rect 7104 33856 7156 33862
rect 7104 33798 7156 33804
rect 6552 33516 6604 33522
rect 6552 33458 6604 33464
rect 7012 33516 7064 33522
rect 7012 33458 7064 33464
rect 5816 33448 5868 33454
rect 5816 33390 5868 33396
rect 5908 33448 5960 33454
rect 5908 33390 5960 33396
rect 6000 33448 6052 33454
rect 6052 33396 6224 33402
rect 6000 33390 6224 33396
rect 5828 32910 5856 33390
rect 5920 33318 5948 33390
rect 6012 33386 6224 33390
rect 6012 33380 6236 33386
rect 6012 33374 6184 33380
rect 6184 33322 6236 33328
rect 5908 33312 5960 33318
rect 5908 33254 5960 33260
rect 6196 33266 6224 33322
rect 6368 33312 6420 33318
rect 6196 33238 6316 33266
rect 6368 33254 6420 33260
rect 6184 33040 6236 33046
rect 6184 32982 6236 32988
rect 6196 32910 6224 32982
rect 6288 32910 6316 33238
rect 6380 32910 6408 33254
rect 6564 33114 6592 33458
rect 7116 33454 7144 33798
rect 7104 33448 7156 33454
rect 7104 33390 7156 33396
rect 7944 33114 7972 34138
rect 8024 33924 8076 33930
rect 8024 33866 8076 33872
rect 8300 33924 8352 33930
rect 8300 33866 8352 33872
rect 6552 33108 6604 33114
rect 6552 33050 6604 33056
rect 7932 33108 7984 33114
rect 7932 33050 7984 33056
rect 8036 32910 8064 33866
rect 8312 33522 8340 33866
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 8852 33516 8904 33522
rect 8852 33458 8904 33464
rect 8864 33114 8892 33458
rect 8300 33108 8352 33114
rect 8300 33050 8352 33056
rect 8852 33108 8904 33114
rect 8852 33050 8904 33056
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 6184 32904 6236 32910
rect 6184 32846 6236 32852
rect 6276 32904 6328 32910
rect 6276 32846 6328 32852
rect 6368 32904 6420 32910
rect 6368 32846 6420 32852
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5724 31680 5776 31686
rect 5724 31622 5776 31628
rect 5552 31470 5764 31498
rect 5736 31346 5764 31470
rect 5724 31340 5776 31346
rect 5724 31282 5776 31288
rect 5147 31036 5455 31045
rect 5147 31034 5153 31036
rect 5209 31034 5233 31036
rect 5289 31034 5313 31036
rect 5369 31034 5393 31036
rect 5449 31034 5455 31036
rect 5209 30982 5211 31034
rect 5391 30982 5393 31034
rect 5147 30980 5153 30982
rect 5209 30980 5233 30982
rect 5289 30980 5313 30982
rect 5369 30980 5393 30982
rect 5449 30980 5455 30982
rect 5147 30971 5455 30980
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 2792 29714 2820 30670
rect 5147 29948 5455 29957
rect 5147 29946 5153 29948
rect 5209 29946 5233 29948
rect 5289 29946 5313 29948
rect 5369 29946 5393 29948
rect 5449 29946 5455 29948
rect 5209 29894 5211 29946
rect 5391 29894 5393 29946
rect 5147 29892 5153 29894
rect 5209 29892 5233 29894
rect 5289 29892 5313 29894
rect 5369 29892 5393 29894
rect 5449 29892 5455 29894
rect 5147 29883 5455 29892
rect 2780 29708 2832 29714
rect 2780 29650 2832 29656
rect 4068 29572 4120 29578
rect 4068 29514 4120 29520
rect 4080 29306 4108 29514
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 5540 29504 5592 29510
rect 5540 29446 5592 29452
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3884 29164 3936 29170
rect 3884 29106 3936 29112
rect 4436 29164 4488 29170
rect 4436 29106 4488 29112
rect 3252 28558 3280 29106
rect 3896 28762 3924 29106
rect 4160 28960 4212 28966
rect 4160 28902 4212 28908
rect 3884 28756 3936 28762
rect 3884 28698 3936 28704
rect 3608 28620 3660 28626
rect 3608 28562 3660 28568
rect 3240 28552 3292 28558
rect 3240 28494 3292 28500
rect 3252 28422 3280 28494
rect 2504 28416 2556 28422
rect 2504 28358 2556 28364
rect 3240 28416 3292 28422
rect 3240 28358 3292 28364
rect 2516 28218 2544 28358
rect 3620 28218 3648 28562
rect 3976 28552 4028 28558
rect 4172 28506 4200 28902
rect 4028 28500 4200 28506
rect 3976 28494 4200 28500
rect 4344 28552 4396 28558
rect 4344 28494 4396 28500
rect 3700 28484 3752 28490
rect 3988 28478 4200 28494
rect 3700 28426 3752 28432
rect 3712 28218 3740 28426
rect 2504 28212 2556 28218
rect 2504 28154 2556 28160
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 3700 28212 3752 28218
rect 3700 28154 3752 28160
rect 4172 28082 4200 28478
rect 4160 28076 4212 28082
rect 4160 28018 4212 28024
rect 3976 28008 4028 28014
rect 3976 27950 4028 27956
rect 3240 27872 3292 27878
rect 3240 27814 3292 27820
rect 3252 27470 3280 27814
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 3252 26450 3280 27406
rect 3240 26444 3292 26450
rect 3240 26386 3292 26392
rect 1860 26308 1912 26314
rect 1860 26250 1912 26256
rect 1872 20210 1900 26250
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2884 24750 2912 25094
rect 3252 24936 3280 26386
rect 3424 26376 3476 26382
rect 3424 26318 3476 26324
rect 3436 26042 3464 26318
rect 3988 26042 4016 27950
rect 3424 26036 3476 26042
rect 3424 25978 3476 25984
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 4172 25906 4200 28018
rect 4356 27946 4384 28494
rect 4448 28490 4476 29106
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4908 28694 4936 28970
rect 4896 28688 4948 28694
rect 4896 28630 4948 28636
rect 4908 28558 4936 28630
rect 4896 28552 4948 28558
rect 4896 28494 4948 28500
rect 4436 28484 4488 28490
rect 4436 28426 4488 28432
rect 4344 27940 4396 27946
rect 4344 27882 4396 27888
rect 4160 25900 4212 25906
rect 4160 25842 4212 25848
rect 4172 25498 4200 25842
rect 4160 25492 4212 25498
rect 4160 25434 4212 25440
rect 3332 25288 3384 25294
rect 3332 25230 3384 25236
rect 3424 25288 3476 25294
rect 3424 25230 3476 25236
rect 3160 24908 3280 24936
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 3160 24614 3188 24908
rect 3344 24750 3372 25230
rect 3436 24954 3464 25230
rect 3424 24948 3476 24954
rect 3424 24890 3476 24896
rect 4356 24818 4384 27882
rect 5000 27878 5028 29446
rect 5552 29170 5580 29446
rect 5540 29164 5592 29170
rect 5540 29106 5592 29112
rect 5147 28860 5455 28869
rect 5147 28858 5153 28860
rect 5209 28858 5233 28860
rect 5289 28858 5313 28860
rect 5369 28858 5393 28860
rect 5449 28858 5455 28860
rect 5209 28806 5211 28858
rect 5391 28806 5393 28858
rect 5147 28804 5153 28806
rect 5209 28804 5233 28806
rect 5289 28804 5313 28806
rect 5369 28804 5393 28806
rect 5449 28804 5455 28806
rect 5147 28795 5455 28804
rect 5552 28626 5580 29106
rect 5632 29096 5684 29102
rect 5632 29038 5684 29044
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5644 28558 5672 29038
rect 5724 28960 5776 28966
rect 5724 28902 5776 28908
rect 5736 28558 5764 28902
rect 5828 28762 5856 31826
rect 5908 31680 5960 31686
rect 5908 31622 5960 31628
rect 6092 31680 6144 31686
rect 6092 31622 6144 31628
rect 5920 31414 5948 31622
rect 6104 31414 6132 31622
rect 5908 31408 5960 31414
rect 5908 31350 5960 31356
rect 6092 31408 6144 31414
rect 6092 31350 6144 31356
rect 5920 30666 5948 31350
rect 6000 31136 6052 31142
rect 6000 31078 6052 31084
rect 6012 30938 6040 31078
rect 6000 30932 6052 30938
rect 6000 30874 6052 30880
rect 5908 30660 5960 30666
rect 5908 30602 5960 30608
rect 6000 29096 6052 29102
rect 6000 29038 6052 29044
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5632 28552 5684 28558
rect 5632 28494 5684 28500
rect 5724 28552 5776 28558
rect 5724 28494 5776 28500
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5460 28218 5488 28358
rect 5448 28212 5500 28218
rect 5448 28154 5500 28160
rect 5828 28082 5856 28698
rect 6012 28558 6040 29038
rect 6000 28552 6052 28558
rect 6000 28494 6052 28500
rect 5816 28076 5868 28082
rect 5816 28018 5868 28024
rect 5908 28076 5960 28082
rect 5908 28018 5960 28024
rect 4988 27872 5040 27878
rect 4988 27814 5040 27820
rect 5540 27872 5592 27878
rect 5540 27814 5592 27820
rect 5000 27402 5028 27814
rect 5147 27772 5455 27781
rect 5147 27770 5153 27772
rect 5209 27770 5233 27772
rect 5289 27770 5313 27772
rect 5369 27770 5393 27772
rect 5449 27770 5455 27772
rect 5209 27718 5211 27770
rect 5391 27718 5393 27770
rect 5147 27716 5153 27718
rect 5209 27716 5233 27718
rect 5289 27716 5313 27718
rect 5369 27716 5393 27718
rect 5449 27716 5455 27718
rect 5147 27707 5455 27716
rect 5552 27674 5580 27814
rect 5540 27668 5592 27674
rect 5540 27610 5592 27616
rect 5920 27402 5948 28018
rect 6196 28014 6224 32846
rect 6288 32502 6316 32846
rect 6276 32496 6328 32502
rect 6276 32438 6328 32444
rect 6380 32298 6408 32846
rect 8036 32570 8064 32846
rect 8024 32564 8076 32570
rect 8024 32506 8076 32512
rect 8208 32496 8260 32502
rect 8208 32438 8260 32444
rect 6920 32360 6972 32366
rect 6920 32302 6972 32308
rect 6368 32292 6420 32298
rect 6368 32234 6420 32240
rect 6552 32224 6604 32230
rect 6552 32166 6604 32172
rect 6276 31952 6328 31958
rect 6276 31894 6328 31900
rect 6288 30190 6316 31894
rect 6368 31816 6420 31822
rect 6368 31758 6420 31764
rect 6380 31482 6408 31758
rect 6368 31476 6420 31482
rect 6368 31418 6420 31424
rect 6564 30326 6592 32166
rect 6932 31346 6960 32302
rect 8220 32026 8248 32438
rect 8208 32020 8260 32026
rect 8208 31962 8260 31968
rect 8312 31822 8340 33050
rect 8956 32910 8984 34342
rect 9416 33998 9444 34342
rect 9600 34134 9628 34614
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 10600 34536 10652 34542
rect 10600 34478 10652 34484
rect 11336 34536 11388 34542
rect 11336 34478 11388 34484
rect 9588 34128 9640 34134
rect 9588 34070 9640 34076
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 9600 33946 9628 34070
rect 9600 33918 9720 33946
rect 9344 33756 9652 33765
rect 9344 33754 9350 33756
rect 9406 33754 9430 33756
rect 9486 33754 9510 33756
rect 9566 33754 9590 33756
rect 9646 33754 9652 33756
rect 9406 33702 9408 33754
rect 9588 33702 9590 33754
rect 9344 33700 9350 33702
rect 9406 33700 9430 33702
rect 9486 33700 9510 33702
rect 9566 33700 9590 33702
rect 9646 33700 9652 33702
rect 9344 33691 9652 33700
rect 9128 33312 9180 33318
rect 9128 33254 9180 33260
rect 8944 32904 8996 32910
rect 8944 32846 8996 32852
rect 8484 32768 8536 32774
rect 8484 32710 8536 32716
rect 8496 32570 8524 32710
rect 8484 32564 8536 32570
rect 8484 32506 8536 32512
rect 8576 31884 8628 31890
rect 8576 31826 8628 31832
rect 8300 31816 8352 31822
rect 8300 31758 8352 31764
rect 8116 31680 8168 31686
rect 8116 31622 8168 31628
rect 8128 31346 8156 31622
rect 8588 31482 8616 31826
rect 8576 31476 8628 31482
rect 8576 31418 8628 31424
rect 6920 31340 6972 31346
rect 6920 31282 6972 31288
rect 8116 31340 8168 31346
rect 8116 31282 8168 31288
rect 6932 30938 6960 31282
rect 8760 31272 8812 31278
rect 8760 31214 8812 31220
rect 7380 31136 7432 31142
rect 7380 31078 7432 31084
rect 7392 30938 7420 31078
rect 6920 30932 6972 30938
rect 6920 30874 6972 30880
rect 7380 30932 7432 30938
rect 7380 30874 7432 30880
rect 8772 30598 8800 31214
rect 8956 30802 8984 32846
rect 9140 32842 9168 33254
rect 9692 32842 9720 33918
rect 9128 32836 9180 32842
rect 9128 32778 9180 32784
rect 9680 32836 9732 32842
rect 9680 32778 9732 32784
rect 9344 32668 9652 32677
rect 9344 32666 9350 32668
rect 9406 32666 9430 32668
rect 9486 32666 9510 32668
rect 9566 32666 9590 32668
rect 9646 32666 9652 32668
rect 9406 32614 9408 32666
rect 9588 32614 9590 32666
rect 9344 32612 9350 32614
rect 9406 32612 9430 32614
rect 9486 32612 9510 32614
rect 9566 32612 9590 32614
rect 9646 32612 9652 32614
rect 9344 32603 9652 32612
rect 9692 32570 9720 32778
rect 9864 32768 9916 32774
rect 9864 32710 9916 32716
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9036 32496 9088 32502
rect 9036 32438 9088 32444
rect 9048 32178 9076 32438
rect 9128 32360 9180 32366
rect 9680 32360 9732 32366
rect 9180 32320 9260 32348
rect 9128 32302 9180 32308
rect 9128 32224 9180 32230
rect 9048 32172 9128 32178
rect 9048 32166 9180 32172
rect 9048 32150 9168 32166
rect 9140 31686 9168 32150
rect 9232 31958 9260 32320
rect 9680 32302 9732 32308
rect 9220 31952 9272 31958
rect 9220 31894 9272 31900
rect 9128 31680 9180 31686
rect 9128 31622 9180 31628
rect 9140 31278 9168 31622
rect 9232 31414 9260 31894
rect 9692 31822 9720 32302
rect 9876 32026 9904 32710
rect 10324 32564 10376 32570
rect 10324 32506 10376 32512
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 9680 31816 9732 31822
rect 9680 31758 9732 31764
rect 9344 31580 9652 31589
rect 9344 31578 9350 31580
rect 9406 31578 9430 31580
rect 9486 31578 9510 31580
rect 9566 31578 9590 31580
rect 9646 31578 9652 31580
rect 9406 31526 9408 31578
rect 9588 31526 9590 31578
rect 9344 31524 9350 31526
rect 9406 31524 9430 31526
rect 9486 31524 9510 31526
rect 9566 31524 9590 31526
rect 9646 31524 9652 31526
rect 9344 31515 9652 31524
rect 9220 31408 9272 31414
rect 9220 31350 9272 31356
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 8944 30796 8996 30802
rect 8944 30738 8996 30744
rect 8760 30592 8812 30598
rect 8760 30534 8812 30540
rect 8772 30326 8800 30534
rect 6552 30320 6604 30326
rect 6552 30262 6604 30268
rect 8760 30320 8812 30326
rect 8760 30262 8812 30268
rect 6276 30184 6328 30190
rect 6276 30126 6328 30132
rect 6736 30184 6788 30190
rect 6736 30126 6788 30132
rect 6748 29306 6776 30126
rect 6920 30048 6972 30054
rect 6920 29990 6972 29996
rect 6736 29300 6788 29306
rect 6736 29242 6788 29248
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 6184 28008 6236 28014
rect 6184 27950 6236 27956
rect 6472 27606 6500 28494
rect 6460 27600 6512 27606
rect 6460 27542 6512 27548
rect 4988 27396 5040 27402
rect 4988 27338 5040 27344
rect 5908 27396 5960 27402
rect 5908 27338 5960 27344
rect 5000 26364 5028 27338
rect 5147 26684 5455 26693
rect 5147 26682 5153 26684
rect 5209 26682 5233 26684
rect 5289 26682 5313 26684
rect 5369 26682 5393 26684
rect 5449 26682 5455 26684
rect 5209 26630 5211 26682
rect 5391 26630 5393 26682
rect 5147 26628 5153 26630
rect 5209 26628 5233 26630
rect 5289 26628 5313 26630
rect 5369 26628 5393 26630
rect 5449 26628 5455 26630
rect 5147 26619 5455 26628
rect 5080 26376 5132 26382
rect 5000 26336 5080 26364
rect 5080 26318 5132 26324
rect 5632 26376 5684 26382
rect 5632 26318 5684 26324
rect 5540 26240 5592 26246
rect 5540 26182 5592 26188
rect 5552 25974 5580 26182
rect 5540 25968 5592 25974
rect 5540 25910 5592 25916
rect 4712 25832 4764 25838
rect 4712 25774 4764 25780
rect 4436 25356 4488 25362
rect 4436 25298 4488 25304
rect 4448 24954 4476 25298
rect 4724 24954 4752 25774
rect 4988 25764 5040 25770
rect 4988 25706 5040 25712
rect 5000 25226 5028 25706
rect 5147 25596 5455 25605
rect 5147 25594 5153 25596
rect 5209 25594 5233 25596
rect 5289 25594 5313 25596
rect 5369 25594 5393 25596
rect 5449 25594 5455 25596
rect 5209 25542 5211 25594
rect 5391 25542 5393 25594
rect 5147 25540 5153 25542
rect 5209 25540 5233 25542
rect 5289 25540 5313 25542
rect 5369 25540 5393 25542
rect 5449 25540 5455 25542
rect 5147 25531 5455 25540
rect 5552 25498 5580 25910
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 4988 25220 5040 25226
rect 4988 25162 5040 25168
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4436 24948 4488 24954
rect 4436 24890 4488 24896
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 4344 24812 4396 24818
rect 4344 24754 4396 24760
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 3148 24608 3200 24614
rect 3148 24550 3200 24556
rect 3160 23730 3188 24550
rect 4356 24410 4384 24754
rect 4528 24608 4580 24614
rect 4528 24550 4580 24556
rect 4344 24404 4396 24410
rect 4344 24346 4396 24352
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4356 23866 4384 24006
rect 4344 23860 4396 23866
rect 4344 23802 4396 23808
rect 4540 23798 4568 24550
rect 4724 24410 4752 24890
rect 4816 24886 4844 25094
rect 4804 24880 4856 24886
rect 4856 24828 4936 24834
rect 4804 24822 4936 24828
rect 4816 24806 4936 24822
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4908 24206 4936 24806
rect 5644 24682 5672 26318
rect 5908 26240 5960 26246
rect 5908 26182 5960 26188
rect 5724 25900 5776 25906
rect 5724 25842 5776 25848
rect 5736 24818 5764 25842
rect 5920 25702 5948 26182
rect 6932 25974 6960 29990
rect 8576 29708 8628 29714
rect 8576 29650 8628 29656
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7668 29238 7696 29446
rect 7656 29232 7708 29238
rect 7656 29174 7708 29180
rect 8484 29232 8536 29238
rect 8588 29220 8616 29650
rect 8956 29238 8984 30738
rect 9232 30258 9260 31350
rect 9692 31346 9720 31758
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 9344 30492 9652 30501
rect 9344 30490 9350 30492
rect 9406 30490 9430 30492
rect 9486 30490 9510 30492
rect 9566 30490 9590 30492
rect 9646 30490 9652 30492
rect 9406 30438 9408 30490
rect 9588 30438 9590 30490
rect 9344 30436 9350 30438
rect 9406 30436 9430 30438
rect 9486 30436 9510 30438
rect 9566 30436 9590 30438
rect 9646 30436 9652 30438
rect 9344 30427 9652 30436
rect 9220 30252 9272 30258
rect 9220 30194 9272 30200
rect 9036 30116 9088 30122
rect 9036 30058 9088 30064
rect 9048 29850 9076 30058
rect 9128 30048 9180 30054
rect 9128 29990 9180 29996
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 9140 29617 9168 29990
rect 9232 29866 9260 30194
rect 9692 30190 9720 31282
rect 9772 30592 9824 30598
rect 9772 30534 9824 30540
rect 9680 30184 9732 30190
rect 9680 30126 9732 30132
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9232 29838 9352 29866
rect 9692 29850 9720 29990
rect 9324 29782 9352 29838
rect 9680 29844 9732 29850
rect 9680 29786 9732 29792
rect 9312 29776 9364 29782
rect 9312 29718 9364 29724
rect 9588 29708 9640 29714
rect 9640 29668 9720 29696
rect 9588 29650 9640 29656
rect 9126 29608 9182 29617
rect 9126 29543 9128 29552
rect 9180 29543 9182 29552
rect 9220 29572 9272 29578
rect 9128 29514 9180 29520
rect 9220 29514 9272 29520
rect 8536 29192 8616 29220
rect 8944 29232 8996 29238
rect 8484 29174 8536 29180
rect 8944 29174 8996 29180
rect 7012 29164 7064 29170
rect 7012 29106 7064 29112
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 7024 28218 7052 29106
rect 7196 28960 7248 28966
rect 7196 28902 7248 28908
rect 7380 28960 7432 28966
rect 7380 28902 7432 28908
rect 7208 28694 7236 28902
rect 7288 28756 7340 28762
rect 7288 28698 7340 28704
rect 7196 28688 7248 28694
rect 7196 28630 7248 28636
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 7012 26920 7064 26926
rect 7012 26862 7064 26868
rect 6920 25968 6972 25974
rect 6920 25910 6972 25916
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5908 25696 5960 25702
rect 5908 25638 5960 25644
rect 5828 25362 5856 25638
rect 5816 25356 5868 25362
rect 5816 25298 5868 25304
rect 5724 24812 5776 24818
rect 5724 24754 5776 24760
rect 5632 24676 5684 24682
rect 5632 24618 5684 24624
rect 5147 24508 5455 24517
rect 5147 24506 5153 24508
rect 5209 24506 5233 24508
rect 5289 24506 5313 24508
rect 5369 24506 5393 24508
rect 5449 24506 5455 24508
rect 5209 24454 5211 24506
rect 5391 24454 5393 24506
rect 5147 24452 5153 24454
rect 5209 24452 5233 24454
rect 5289 24452 5313 24454
rect 5369 24452 5393 24454
rect 5449 24452 5455 24454
rect 5147 24443 5455 24452
rect 5736 24274 5764 24754
rect 5724 24268 5776 24274
rect 5724 24210 5776 24216
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 5080 24200 5132 24206
rect 5080 24142 5132 24148
rect 4528 23792 4580 23798
rect 4528 23734 4580 23740
rect 3148 23724 3200 23730
rect 3148 23666 3200 23672
rect 4540 23050 4568 23734
rect 5092 23474 5120 24142
rect 5736 23866 5764 24210
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 5000 23446 5120 23474
rect 5000 23118 5028 23446
rect 5147 23420 5455 23429
rect 5147 23418 5153 23420
rect 5209 23418 5233 23420
rect 5289 23418 5313 23420
rect 5369 23418 5393 23420
rect 5449 23418 5455 23420
rect 5209 23366 5211 23418
rect 5391 23366 5393 23418
rect 5147 23364 5153 23366
rect 5209 23364 5233 23366
rect 5289 23364 5313 23366
rect 5369 23364 5393 23366
rect 5449 23364 5455 23366
rect 5147 23355 5455 23364
rect 5920 23186 5948 25638
rect 6932 25158 6960 25774
rect 7024 25702 7052 26862
rect 7300 26858 7328 28698
rect 7392 28490 7420 28902
rect 8864 28490 8892 29106
rect 8956 28626 8984 29174
rect 9232 29170 9260 29514
rect 9344 29404 9652 29413
rect 9344 29402 9350 29404
rect 9406 29402 9430 29404
rect 9486 29402 9510 29404
rect 9566 29402 9590 29404
rect 9646 29402 9652 29404
rect 9406 29350 9408 29402
rect 9588 29350 9590 29402
rect 9344 29348 9350 29350
rect 9406 29348 9430 29350
rect 9486 29348 9510 29350
rect 9566 29348 9590 29350
rect 9646 29348 9652 29350
rect 9344 29339 9652 29348
rect 9692 29238 9720 29668
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9220 29164 9272 29170
rect 9220 29106 9272 29112
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 8944 28620 8996 28626
rect 8944 28562 8996 28568
rect 9140 28490 9168 28902
rect 9784 28490 9812 30534
rect 9876 30054 9904 31962
rect 9956 31680 10008 31686
rect 9956 31622 10008 31628
rect 9968 31482 9996 31622
rect 9956 31476 10008 31482
rect 9956 31418 10008 31424
rect 10336 30734 10364 32506
rect 10612 31822 10640 34478
rect 10692 32768 10744 32774
rect 10692 32710 10744 32716
rect 10704 32570 10732 32710
rect 10692 32564 10744 32570
rect 10692 32506 10744 32512
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10416 31680 10468 31686
rect 10416 31622 10468 31628
rect 10428 31346 10456 31622
rect 10416 31340 10468 31346
rect 10416 31282 10468 31288
rect 10324 30728 10376 30734
rect 10324 30670 10376 30676
rect 10612 30598 10640 31758
rect 10600 30592 10652 30598
rect 10600 30534 10652 30540
rect 9864 30048 9916 30054
rect 10048 30048 10100 30054
rect 9916 29996 9996 30002
rect 9864 29990 9996 29996
rect 10048 29990 10100 29996
rect 9876 29974 9996 29990
rect 7380 28484 7432 28490
rect 7380 28426 7432 28432
rect 7656 28484 7708 28490
rect 7656 28426 7708 28432
rect 8852 28484 8904 28490
rect 8852 28426 8904 28432
rect 9128 28484 9180 28490
rect 9128 28426 9180 28432
rect 9772 28484 9824 28490
rect 9772 28426 9824 28432
rect 7668 28218 7696 28426
rect 8576 28416 8628 28422
rect 8576 28358 8628 28364
rect 7656 28212 7708 28218
rect 7656 28154 7708 28160
rect 7668 26926 7696 28154
rect 8588 28150 8616 28358
rect 8576 28144 8628 28150
rect 8576 28086 8628 28092
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7288 26852 7340 26858
rect 7288 26794 7340 26800
rect 7300 26586 7328 26794
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7196 26308 7248 26314
rect 7196 26250 7248 26256
rect 7208 26042 7236 26250
rect 7484 26042 7512 26726
rect 7668 26450 7696 26862
rect 7656 26444 7708 26450
rect 7656 26386 7708 26392
rect 8668 26240 8720 26246
rect 8668 26182 8720 26188
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7472 26036 7524 26042
rect 7472 25978 7524 25984
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7840 25696 7892 25702
rect 7840 25638 7892 25644
rect 7208 25498 7236 25638
rect 7852 25498 7880 25638
rect 8680 25498 8708 26182
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 8668 25492 8720 25498
rect 8668 25434 8720 25440
rect 7196 25356 7248 25362
rect 7196 25298 7248 25304
rect 7208 25158 7236 25298
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 7012 25152 7064 25158
rect 7012 25094 7064 25100
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 6472 24954 6500 25094
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 7024 24886 7052 25094
rect 7012 24880 7064 24886
rect 7012 24822 7064 24828
rect 6368 24608 6420 24614
rect 6368 24550 6420 24556
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 6380 23866 6408 24550
rect 7024 24138 7052 24550
rect 7208 24410 7236 25094
rect 7760 24954 7788 25230
rect 7748 24948 7800 24954
rect 7748 24890 7800 24896
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 8484 24268 8536 24274
rect 8484 24210 8536 24216
rect 6552 24132 6604 24138
rect 6552 24074 6604 24080
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 6564 23866 6592 24074
rect 6368 23860 6420 23866
rect 6368 23802 6420 23808
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 5908 23180 5960 23186
rect 5908 23122 5960 23128
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 4528 23044 4580 23050
rect 4528 22986 4580 22992
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1964 20398 1992 21966
rect 4540 21962 4568 22986
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 2688 21956 2740 21962
rect 2688 21898 2740 21904
rect 4344 21956 4396 21962
rect 4344 21898 4396 21904
rect 4528 21956 4580 21962
rect 4528 21898 4580 21904
rect 2700 20534 2728 21898
rect 4356 21690 4384 21898
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 2688 20528 2740 20534
rect 2688 20470 2740 20476
rect 1952 20392 2004 20398
rect 1952 20334 2004 20340
rect 2320 20392 2372 20398
rect 2320 20334 2372 20340
rect 1872 20182 1992 20210
rect 1780 20046 1900 20074
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1596 19446 1624 19654
rect 1584 19440 1636 19446
rect 1584 19382 1636 19388
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 18834 1440 19314
rect 1872 18970 1900 20046
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1872 18426 1900 18634
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1412 15570 1440 17070
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 952 13025 980 13262
rect 938 13016 994 13025
rect 938 12951 994 12960
rect 1412 11218 1440 15506
rect 1504 15502 1532 16050
rect 1964 15978 1992 20182
rect 2332 20058 2360 20334
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2700 19446 2728 20470
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4172 20058 4200 20198
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 2688 19440 2740 19446
rect 3160 19417 3188 19450
rect 2688 19382 2740 19388
rect 3146 19408 3202 19417
rect 3146 19343 3202 19352
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2976 17202 3004 18702
rect 3620 18290 3648 19654
rect 4172 19514 4200 19722
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3700 18692 3752 18698
rect 3700 18634 3752 18640
rect 3712 18426 3740 18634
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3896 18358 3924 19314
rect 3884 18352 3936 18358
rect 3884 18294 3936 18300
rect 3608 18284 3660 18290
rect 3660 18244 3740 18272
rect 3608 18226 3660 18232
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 3436 17338 3464 17750
rect 3712 17678 3740 18244
rect 3896 17882 3924 18294
rect 4540 18290 4568 20402
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4632 20058 4660 20334
rect 4724 20058 4752 21490
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4816 20806 4844 21286
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4816 20398 4844 20742
rect 4908 20534 4936 22918
rect 5460 22642 5488 23054
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 5147 22332 5455 22341
rect 5147 22330 5153 22332
rect 5209 22330 5233 22332
rect 5289 22330 5313 22332
rect 5369 22330 5393 22332
rect 5449 22330 5455 22332
rect 5209 22278 5211 22330
rect 5391 22278 5393 22330
rect 5147 22276 5153 22278
rect 5209 22276 5233 22278
rect 5289 22276 5313 22278
rect 5369 22276 5393 22278
rect 5449 22276 5455 22278
rect 5147 22267 5455 22276
rect 6012 22234 6040 23054
rect 6656 22982 6684 24074
rect 8496 23730 8524 24210
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 6656 22710 6684 22918
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 6000 22228 6052 22234
rect 6000 22170 6052 22176
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 5368 21554 5396 21898
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5460 21350 5488 21966
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5147 21244 5455 21253
rect 5147 21242 5153 21244
rect 5209 21242 5233 21244
rect 5289 21242 5313 21244
rect 5369 21242 5393 21244
rect 5449 21242 5455 21244
rect 5209 21190 5211 21242
rect 5391 21190 5393 21242
rect 5147 21188 5153 21190
rect 5209 21188 5233 21190
rect 5289 21188 5313 21190
rect 5369 21188 5393 21190
rect 5449 21188 5455 21190
rect 5147 21179 5455 21188
rect 5552 20942 5580 21490
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 5000 20602 5028 20810
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 4896 20528 4948 20534
rect 4896 20470 4948 20476
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4908 19938 4936 20470
rect 4988 20324 5040 20330
rect 4988 20266 5040 20272
rect 4816 19910 4936 19938
rect 4816 19854 4844 19910
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4632 18873 4660 19790
rect 4816 19514 4844 19790
rect 5000 19514 5028 20266
rect 5147 20156 5455 20165
rect 5147 20154 5153 20156
rect 5209 20154 5233 20156
rect 5289 20154 5313 20156
rect 5369 20154 5393 20156
rect 5449 20154 5455 20156
rect 5209 20102 5211 20154
rect 5391 20102 5393 20154
rect 5147 20100 5153 20102
rect 5209 20100 5233 20102
rect 5289 20100 5313 20102
rect 5369 20100 5393 20102
rect 5449 20100 5455 20102
rect 5147 20091 5455 20100
rect 5552 20058 5580 20742
rect 5828 20466 5856 21898
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 5908 20528 5960 20534
rect 5908 20470 5960 20476
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5184 19774 5580 19802
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4724 19310 4752 19450
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4618 18864 4674 18873
rect 4618 18799 4674 18808
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 3988 17882 4016 18226
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 4724 17746 4752 19246
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 4816 17746 4844 18294
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3700 17672 3752 17678
rect 4528 17672 4580 17678
rect 3700 17614 3752 17620
rect 4448 17632 4528 17660
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3528 17202 3556 17546
rect 3620 17338 3648 17614
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3606 17232 3662 17241
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 3516 17196 3568 17202
rect 3712 17202 3740 17614
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3606 17167 3608 17176
rect 3516 17138 3568 17144
rect 3660 17167 3662 17176
rect 3700 17196 3752 17202
rect 3608 17138 3660 17144
rect 3700 17138 3752 17144
rect 1952 15972 2004 15978
rect 1952 15914 2004 15920
rect 1492 15496 1544 15502
rect 1492 15438 1544 15444
rect 2976 15434 3004 17138
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 3160 16590 3188 16934
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 3068 16046 3096 16458
rect 3620 16250 3648 17138
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 11218 1716 13126
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1412 9586 1440 11154
rect 2976 11150 3004 15370
rect 3068 15026 3096 15982
rect 3804 15706 3832 17478
rect 4264 17338 4292 17546
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3896 16522 3924 17070
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3988 15026 4016 16730
rect 4448 16697 4476 17632
rect 4528 17614 4580 17620
rect 4816 17134 4844 17682
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4434 16688 4490 16697
rect 4068 16652 4120 16658
rect 4434 16623 4490 16632
rect 4068 16594 4120 16600
rect 4080 16114 4108 16594
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 15026 4108 16050
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 3344 13938 3372 14962
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3344 13326 3372 13874
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12306 3372 13262
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3252 11898 3280 12038
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3436 11762 3464 12310
rect 3620 12238 3648 13874
rect 3804 13870 3832 14486
rect 3896 14006 3924 14758
rect 3988 14074 4016 14962
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3884 14000 3936 14006
rect 4264 13977 4292 14486
rect 3884 13942 3936 13948
rect 4250 13968 4306 13977
rect 4250 13903 4306 13912
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 4264 13326 4292 13903
rect 4356 13734 4384 14826
rect 4448 14260 4476 16623
rect 4816 16250 4844 17070
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15094 4568 15846
rect 4528 15088 4580 15094
rect 4528 15030 4580 15036
rect 4528 14272 4580 14278
rect 4448 14232 4528 14260
rect 4528 14214 4580 14220
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4356 13462 4384 13670
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 3804 12442 3832 13262
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3792 12436 3844 12442
rect 3844 12396 3924 12424
rect 3792 12378 3844 12384
rect 3896 12238 3924 12396
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3424 11756 3476 11762
rect 3620 11744 3648 12174
rect 3896 11762 3924 12174
rect 3700 11756 3752 11762
rect 3620 11716 3700 11744
rect 3424 11698 3476 11704
rect 3700 11698 3752 11704
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10674 3188 10950
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3068 9654 3096 10406
rect 3252 9654 3280 11086
rect 3344 10538 3372 11494
rect 3436 11354 3464 11698
rect 3988 11558 4016 13126
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4080 11898 4108 12106
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4264 11762 4292 12038
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4448 11694 4476 12174
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3988 11082 4016 11494
rect 4448 11354 4476 11630
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 4540 9994 4568 14214
rect 4632 14074 4660 16118
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4724 14890 4752 16050
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4816 15162 4844 15982
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4724 14414 4752 14826
rect 4816 14414 4844 15098
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4908 14278 4936 19314
rect 5000 18426 5028 19450
rect 5184 19310 5212 19774
rect 5552 19718 5580 19774
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5460 19258 5488 19654
rect 5644 19514 5672 20402
rect 5736 20369 5764 20402
rect 5722 20360 5778 20369
rect 5722 20295 5778 20304
rect 5736 19854 5764 20295
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5460 19230 5580 19258
rect 5147 19068 5455 19077
rect 5147 19066 5153 19068
rect 5209 19066 5233 19068
rect 5289 19066 5313 19068
rect 5369 19066 5393 19068
rect 5449 19066 5455 19068
rect 5209 19014 5211 19066
rect 5391 19014 5393 19066
rect 5147 19012 5153 19014
rect 5209 19012 5233 19014
rect 5289 19012 5313 19014
rect 5369 19012 5393 19014
rect 5449 19012 5455 19014
rect 5147 19003 5455 19012
rect 5552 18850 5580 19230
rect 5644 19174 5672 19450
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5460 18822 5580 18850
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 5276 18086 5304 18702
rect 5460 18086 5488 18822
rect 5736 18766 5764 19246
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5540 18284 5592 18290
rect 5592 18244 5672 18272
rect 5540 18226 5592 18232
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5000 17252 5028 18022
rect 5147 17980 5455 17989
rect 5147 17978 5153 17980
rect 5209 17978 5233 17980
rect 5289 17978 5313 17980
rect 5369 17978 5393 17980
rect 5449 17978 5455 17980
rect 5209 17926 5211 17978
rect 5391 17926 5393 17978
rect 5147 17924 5153 17926
rect 5209 17924 5233 17926
rect 5289 17924 5313 17926
rect 5369 17924 5393 17926
rect 5449 17924 5455 17926
rect 5147 17915 5455 17924
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5080 17264 5132 17270
rect 5000 17224 5080 17252
rect 5080 17206 5132 17212
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4618 13968 4674 13977
rect 4618 13903 4620 13912
rect 4672 13903 4674 13912
rect 4712 13932 4764 13938
rect 4620 13874 4672 13880
rect 4712 13874 4764 13880
rect 4724 13530 4752 13874
rect 4712 13524 4764 13530
rect 4632 13484 4712 13512
rect 4632 10674 4660 13484
rect 4712 13466 4764 13472
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4724 10606 4752 11018
rect 5000 10674 5028 16934
rect 5147 16892 5455 16901
rect 5147 16890 5153 16892
rect 5209 16890 5233 16892
rect 5289 16890 5313 16892
rect 5369 16890 5393 16892
rect 5449 16890 5455 16892
rect 5209 16838 5211 16890
rect 5391 16838 5393 16890
rect 5147 16836 5153 16838
rect 5209 16836 5233 16838
rect 5289 16836 5313 16838
rect 5369 16836 5393 16838
rect 5449 16836 5455 16838
rect 5147 16827 5455 16836
rect 5552 16674 5580 17682
rect 5644 16794 5672 18244
rect 5736 17202 5764 18362
rect 5828 18290 5856 20402
rect 5920 19854 5948 20470
rect 6012 20262 6040 21354
rect 6276 20868 6328 20874
rect 6276 20810 6328 20816
rect 6288 20466 6316 20810
rect 6380 20602 6408 21966
rect 7300 21690 7328 22510
rect 7668 22094 7696 22510
rect 7576 22066 7696 22094
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6564 20466 6684 20482
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6552 20460 6684 20466
rect 6604 20454 6684 20460
rect 6552 20402 6604 20408
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6656 19922 6684 20454
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5998 19816 6054 19825
rect 5920 19378 5948 19790
rect 5998 19751 6000 19760
rect 6052 19751 6054 19760
rect 6000 19722 6052 19728
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 6748 19334 6776 20878
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6932 20466 6960 20538
rect 7116 20466 7144 20878
rect 7300 20466 7328 21490
rect 7576 21486 7604 22066
rect 7760 22030 7788 22918
rect 8220 22098 8248 23598
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7472 20868 7524 20874
rect 7472 20810 7524 20816
rect 7484 20466 7512 20810
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7116 20058 7144 20402
rect 7576 20262 7604 21422
rect 7760 20534 7788 21966
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7300 19922 7328 20198
rect 7760 20058 7788 20198
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6840 19514 6868 19722
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 7104 19440 7156 19446
rect 7208 19394 7236 19790
rect 7156 19388 7236 19394
rect 7104 19382 7236 19388
rect 6920 19372 6972 19378
rect 6748 19306 6868 19334
rect 7116 19366 7236 19382
rect 6920 19314 6972 19320
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6380 18290 6408 18838
rect 5816 18284 5868 18290
rect 6368 18284 6420 18290
rect 5868 18244 5948 18272
rect 5816 18226 5868 18232
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5828 17678 5856 18090
rect 5920 17678 5948 18244
rect 6368 18226 6420 18232
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5828 16794 5856 17614
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5460 16646 5580 16674
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5184 15910 5212 16186
rect 5460 16114 5488 16646
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5147 15804 5455 15813
rect 5147 15802 5153 15804
rect 5209 15802 5233 15804
rect 5289 15802 5313 15804
rect 5369 15802 5393 15804
rect 5449 15802 5455 15804
rect 5209 15750 5211 15802
rect 5391 15750 5393 15802
rect 5147 15748 5153 15750
rect 5209 15748 5233 15750
rect 5289 15748 5313 15750
rect 5369 15748 5393 15750
rect 5449 15748 5455 15750
rect 5147 15739 5455 15748
rect 5552 15026 5580 16526
rect 5644 15502 5672 16730
rect 6012 16590 6040 18158
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6288 16590 6316 17614
rect 6840 16590 6868 19306
rect 6932 18766 6960 19314
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6932 18426 6960 18702
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 7116 17785 7144 18566
rect 7102 17776 7158 17785
rect 6920 17740 6972 17746
rect 7102 17711 7158 17720
rect 6920 17682 6972 17688
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6276 16584 6328 16590
rect 6828 16584 6880 16590
rect 6276 16526 6328 16532
rect 6826 16552 6828 16561
rect 6880 16552 6882 16561
rect 6826 16487 6882 16496
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 15910 6408 16390
rect 6932 16096 6960 17682
rect 6840 16068 6960 16096
rect 6092 15904 6144 15910
rect 6368 15904 6420 15910
rect 6092 15846 6144 15852
rect 6288 15852 6368 15858
rect 6288 15846 6420 15852
rect 6104 15502 6132 15846
rect 6288 15830 6408 15846
rect 6288 15570 6316 15830
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 5814 15192 5870 15201
rect 5814 15127 5816 15136
rect 5868 15127 5870 15136
rect 5816 15098 5868 15104
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5552 14890 5580 14962
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5147 14716 5455 14725
rect 5147 14714 5153 14716
rect 5209 14714 5233 14716
rect 5289 14714 5313 14716
rect 5369 14714 5393 14716
rect 5449 14714 5455 14716
rect 5209 14662 5211 14714
rect 5391 14662 5393 14714
rect 5147 14660 5153 14662
rect 5209 14660 5233 14662
rect 5289 14660 5313 14662
rect 5369 14660 5393 14662
rect 5449 14660 5455 14662
rect 5147 14651 5455 14660
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5460 14074 5488 14214
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5080 13728 5132 13734
rect 5356 13728 5408 13734
rect 5132 13688 5356 13716
rect 5080 13670 5132 13676
rect 5356 13670 5408 13676
rect 5147 13628 5455 13637
rect 5147 13626 5153 13628
rect 5209 13626 5233 13628
rect 5289 13626 5313 13628
rect 5369 13626 5393 13628
rect 5449 13626 5455 13628
rect 5209 13574 5211 13626
rect 5391 13574 5393 13626
rect 5147 13572 5153 13574
rect 5209 13572 5233 13574
rect 5289 13572 5313 13574
rect 5369 13572 5393 13574
rect 5449 13572 5455 13574
rect 5147 13563 5455 13572
rect 5147 12540 5455 12549
rect 5147 12538 5153 12540
rect 5209 12538 5233 12540
rect 5289 12538 5313 12540
rect 5369 12538 5393 12540
rect 5449 12538 5455 12540
rect 5209 12486 5211 12538
rect 5391 12486 5393 12538
rect 5147 12484 5153 12486
rect 5209 12484 5233 12486
rect 5289 12484 5313 12486
rect 5369 12484 5393 12486
rect 5449 12484 5455 12486
rect 5147 12475 5455 12484
rect 5552 12238 5580 14214
rect 5736 13938 5764 14758
rect 5828 14278 5856 15098
rect 6104 14414 6132 15302
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5644 13258 5672 13806
rect 5736 13326 5764 13874
rect 5828 13326 5856 13942
rect 6104 13870 6132 14350
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6000 13728 6052 13734
rect 6196 13716 6224 14486
rect 6000 13670 6052 13676
rect 6104 13688 6224 13716
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 6012 13190 6040 13670
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6104 12238 6132 13688
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 5540 12232 5592 12238
rect 5446 12200 5502 12209
rect 5540 12174 5592 12180
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 5446 12135 5448 12144
rect 5500 12135 5502 12144
rect 5448 12106 5500 12112
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5092 11898 5120 12038
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5078 11792 5134 11801
rect 5078 11727 5080 11736
rect 5132 11727 5134 11736
rect 5080 11698 5132 11704
rect 5147 11452 5455 11461
rect 5147 11450 5153 11452
rect 5209 11450 5233 11452
rect 5289 11450 5313 11452
rect 5369 11450 5393 11452
rect 5449 11450 5455 11452
rect 5209 11398 5211 11450
rect 5391 11398 5393 11450
rect 5147 11396 5153 11398
rect 5209 11396 5233 11398
rect 5289 11396 5313 11398
rect 5369 11396 5393 11398
rect 5449 11396 5455 11398
rect 5147 11387 5455 11396
rect 5552 11354 5580 12174
rect 6196 12102 6224 13330
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12986 6316 13126
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6288 12306 6316 12922
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5828 10606 5856 12038
rect 6196 11762 6224 12038
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6196 11218 6224 11698
rect 6380 11694 6408 15642
rect 6840 15638 6868 16068
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6932 15473 6960 15914
rect 6918 15464 6974 15473
rect 6918 15399 6974 15408
rect 6932 15162 6960 15399
rect 7116 15162 7144 17711
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12238 6500 13262
rect 6564 13190 6592 13942
rect 6840 13530 6868 15030
rect 7010 14920 7066 14929
rect 7010 14855 7066 14864
rect 7024 14618 7052 14855
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 14006 7052 14214
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7116 13938 7144 14758
rect 7208 14278 7236 19366
rect 7300 18902 7328 19858
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7300 17678 7328 18838
rect 7392 18766 7420 19314
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 18766 7604 19110
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7392 17814 7420 18702
rect 7380 17808 7432 17814
rect 7380 17750 7432 17756
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7300 14958 7328 17614
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7378 17232 7434 17241
rect 7668 17202 7696 17546
rect 7760 17202 7788 19994
rect 7852 18630 7880 21490
rect 8312 18850 8340 22374
rect 8772 22030 8800 22918
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8404 21690 8432 21966
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8404 19854 8432 20402
rect 8680 20330 8708 20538
rect 8668 20324 8720 20330
rect 8668 20266 8720 20272
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8404 19446 8432 19790
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8482 19408 8538 19417
rect 8128 18834 8340 18850
rect 8128 18828 8352 18834
rect 8128 18822 8300 18828
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 8128 18358 8156 18822
rect 8300 18770 8352 18776
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8312 18358 8340 18634
rect 8116 18352 8168 18358
rect 8300 18352 8352 18358
rect 8116 18294 8168 18300
rect 8220 18312 8300 18340
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 7378 17167 7380 17176
rect 7432 17167 7434 17176
rect 7656 17196 7708 17202
rect 7380 17138 7432 17144
rect 7656 17138 7708 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7668 17066 7696 17138
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7760 16776 7788 16934
rect 7930 16824 7986 16833
rect 7668 16748 7788 16776
rect 7840 16788 7892 16794
rect 7668 16590 7696 16748
rect 7930 16759 7986 16768
rect 7840 16730 7892 16736
rect 7746 16688 7802 16697
rect 7746 16623 7802 16632
rect 7760 16590 7788 16623
rect 7852 16590 7880 16730
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7392 15570 7420 16526
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7576 15706 7604 16458
rect 7852 15994 7880 16526
rect 7944 16250 7972 16759
rect 8128 16289 8156 17478
rect 8114 16280 8170 16289
rect 7932 16244 7984 16250
rect 8220 16250 8248 18312
rect 8300 18294 8352 18300
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8312 17202 8340 17682
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8312 16998 8340 17138
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8298 16416 8354 16425
rect 8298 16351 8354 16360
rect 8312 16250 8340 16351
rect 8114 16215 8170 16224
rect 8208 16244 8260 16250
rect 7932 16186 7984 16192
rect 8208 16186 8260 16192
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 7668 15966 7880 15994
rect 8024 15972 8076 15978
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7564 15428 7616 15434
rect 7564 15370 7616 15376
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7300 14074 7328 14350
rect 7392 14074 7420 14962
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6472 11898 6500 12174
rect 6564 11898 6592 12786
rect 6840 12714 6868 13194
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6840 12356 6868 12650
rect 7024 12434 7052 13806
rect 7116 12442 7144 13874
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 6748 12328 6868 12356
rect 6932 12406 7052 12434
rect 7104 12436 7156 12442
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6380 11354 6408 11630
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6274 10976 6330 10985
rect 6274 10911 6330 10920
rect 6288 10742 6316 10911
rect 6380 10742 6408 11290
rect 6472 11218 6500 11834
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5147 10364 5455 10373
rect 5147 10362 5153 10364
rect 5209 10362 5233 10364
rect 5289 10362 5313 10364
rect 5369 10362 5393 10364
rect 5449 10362 5455 10364
rect 5209 10310 5211 10362
rect 5391 10310 5393 10362
rect 5147 10308 5153 10310
rect 5209 10308 5233 10310
rect 5289 10308 5313 10310
rect 5369 10308 5393 10310
rect 5449 10308 5455 10310
rect 5147 10299 5455 10308
rect 5552 10062 5580 10406
rect 5828 10130 5856 10542
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 10266 6408 10406
rect 6656 10266 6684 12038
rect 6748 11898 6776 12328
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6748 11150 6776 11834
rect 6932 11762 6960 12406
rect 7104 12378 7156 12384
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6736 11144 6788 11150
rect 6840 11121 6868 11222
rect 6736 11086 6788 11092
rect 6826 11112 6882 11121
rect 6826 11047 6882 11056
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10538 6868 10950
rect 6932 10606 6960 11698
rect 7024 11694 7052 12038
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6828 10532 6880 10538
rect 6828 10474 6880 10480
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 6196 9722 6224 9998
rect 7116 9994 7144 10406
rect 7208 10062 7236 13466
rect 7484 12986 7512 14962
rect 7576 14550 7604 15370
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 11150 7328 12582
rect 7470 12472 7526 12481
rect 7470 12407 7526 12416
rect 7484 12306 7512 12407
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7484 11830 7512 12242
rect 7576 11898 7604 14350
rect 7668 13410 7696 15966
rect 8024 15914 8076 15920
rect 8116 15972 8168 15978
rect 8116 15914 8168 15920
rect 8036 15706 8064 15914
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8128 15502 8156 15914
rect 8024 15496 8076 15502
rect 7852 15456 8024 15484
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7760 14482 7788 15302
rect 7852 15162 7880 15456
rect 8024 15438 8076 15444
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 7932 15360 7984 15366
rect 8220 15314 8248 15370
rect 7932 15302 7984 15308
rect 7944 15201 7972 15302
rect 8036 15286 8248 15314
rect 7930 15192 7986 15201
rect 7840 15156 7892 15162
rect 7930 15127 7986 15136
rect 7840 15098 7892 15104
rect 8036 15076 8064 15286
rect 8312 15178 8340 16050
rect 8404 15638 8432 19382
rect 8482 19343 8538 19352
rect 8496 19310 8524 19343
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8576 18760 8628 18766
rect 8496 18720 8576 18748
rect 8496 18222 8524 18720
rect 8576 18702 8628 18708
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 7944 15048 8064 15076
rect 8220 15150 8340 15178
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7944 14362 7972 15048
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7852 14334 7972 14362
rect 7852 13530 7880 14334
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7668 13382 7880 13410
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7668 12646 7696 13262
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7668 12306 7696 12582
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7564 11892 7616 11898
rect 7616 11852 7696 11880
rect 7564 11834 7616 11840
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7484 9994 7512 11154
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10062 7604 10610
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2700 6798 2728 9522
rect 3252 6798 3280 9590
rect 7024 9382 7052 9930
rect 7668 9926 7696 11852
rect 7760 11762 7788 12174
rect 7852 12102 7880 13382
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7944 11150 7972 13466
rect 8036 13394 8064 14894
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8128 13462 8156 14282
rect 8220 13530 8248 15150
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 8404 13938 8432 14282
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8298 13424 8354 13433
rect 8024 13388 8076 13394
rect 8354 13382 8432 13410
rect 8298 13359 8354 13368
rect 8024 13330 8076 13336
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7760 10266 7788 10678
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7944 10062 7972 11086
rect 8036 11014 8064 13330
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12714 8248 13262
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8128 11626 8156 11766
rect 8220 11694 8248 12174
rect 8312 12170 8340 12854
rect 8404 12374 8432 13382
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8496 12220 8524 17002
rect 8588 16250 8616 18566
rect 8680 18290 8708 20266
rect 8758 18864 8814 18873
rect 8758 18799 8760 18808
rect 8812 18799 8814 18808
rect 8760 18770 8812 18776
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8680 16658 8708 18090
rect 8772 17542 8800 18770
rect 8864 18358 8892 28426
rect 9344 28316 9652 28325
rect 9344 28314 9350 28316
rect 9406 28314 9430 28316
rect 9486 28314 9510 28316
rect 9566 28314 9590 28316
rect 9646 28314 9652 28316
rect 9406 28262 9408 28314
rect 9588 28262 9590 28314
rect 9344 28260 9350 28262
rect 9406 28260 9430 28262
rect 9486 28260 9510 28262
rect 9566 28260 9590 28262
rect 9646 28260 9652 28262
rect 9344 28251 9652 28260
rect 9784 28150 9812 28426
rect 9772 28144 9824 28150
rect 9772 28086 9824 28092
rect 9344 27228 9652 27237
rect 9344 27226 9350 27228
rect 9406 27226 9430 27228
rect 9486 27226 9510 27228
rect 9566 27226 9590 27228
rect 9646 27226 9652 27228
rect 9406 27174 9408 27226
rect 9588 27174 9590 27226
rect 9344 27172 9350 27174
rect 9406 27172 9430 27174
rect 9486 27172 9510 27174
rect 9566 27172 9590 27174
rect 9646 27172 9652 27174
rect 9344 27163 9652 27172
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 9036 25152 9088 25158
rect 9036 25094 9088 25100
rect 9048 24954 9076 25094
rect 9036 24948 9088 24954
rect 9036 24890 9088 24896
rect 9140 24750 9168 25638
rect 9232 25498 9260 26862
rect 9784 26382 9812 28086
rect 9968 26586 9996 29974
rect 10060 29238 10088 29990
rect 10612 29646 10640 30534
rect 10692 29776 10744 29782
rect 10692 29718 10744 29724
rect 10600 29640 10652 29646
rect 10230 29608 10286 29617
rect 10600 29582 10652 29588
rect 10230 29543 10286 29552
rect 10244 29510 10272 29543
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 10048 29232 10100 29238
rect 10048 29174 10100 29180
rect 10704 29102 10732 29718
rect 11244 29708 11296 29714
rect 11244 29650 11296 29656
rect 11256 29170 11284 29650
rect 11244 29164 11296 29170
rect 11244 29106 11296 29112
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10704 28762 10732 29038
rect 10692 28756 10744 28762
rect 10692 28698 10744 28704
rect 11256 28014 11284 29106
rect 11348 28626 11376 34478
rect 14096 34400 14148 34406
rect 14096 34342 14148 34348
rect 13541 34300 13849 34309
rect 13541 34298 13547 34300
rect 13603 34298 13627 34300
rect 13683 34298 13707 34300
rect 13763 34298 13787 34300
rect 13843 34298 13849 34300
rect 13603 34246 13605 34298
rect 13785 34246 13787 34298
rect 13541 34244 13547 34246
rect 13603 34244 13627 34246
rect 13683 34244 13707 34246
rect 13763 34244 13787 34246
rect 13843 34244 13849 34246
rect 13541 34235 13849 34244
rect 14108 34066 14136 34342
rect 14200 34066 14228 34546
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 14476 34202 14504 34478
rect 14464 34196 14516 34202
rect 14464 34138 14516 34144
rect 14096 34060 14148 34066
rect 14096 34002 14148 34008
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 15108 34060 15160 34066
rect 15108 34002 15160 34008
rect 13452 33380 13504 33386
rect 13452 33322 13504 33328
rect 13464 32978 13492 33322
rect 13541 33212 13849 33221
rect 13541 33210 13547 33212
rect 13603 33210 13627 33212
rect 13683 33210 13707 33212
rect 13763 33210 13787 33212
rect 13843 33210 13849 33212
rect 13603 33158 13605 33210
rect 13785 33158 13787 33210
rect 13541 33156 13547 33158
rect 13603 33156 13627 33158
rect 13683 33156 13707 33158
rect 13763 33156 13787 33158
rect 13843 33156 13849 33158
rect 13541 33147 13849 33156
rect 15120 32978 15148 34002
rect 15672 33930 15700 34886
rect 15764 34610 15792 35158
rect 19996 35086 20024 37217
rect 21935 35388 22243 35397
rect 21935 35386 21941 35388
rect 21997 35386 22021 35388
rect 22077 35386 22101 35388
rect 22157 35386 22181 35388
rect 22237 35386 22243 35388
rect 21997 35334 21999 35386
rect 22179 35334 22181 35386
rect 21935 35332 21941 35334
rect 21997 35332 22021 35334
rect 22077 35332 22101 35334
rect 22157 35332 22181 35334
rect 22237 35332 22243 35334
rect 21935 35323 22243 35332
rect 26436 35290 26464 37217
rect 30329 35388 30637 35397
rect 30329 35386 30335 35388
rect 30391 35386 30415 35388
rect 30471 35386 30495 35388
rect 30551 35386 30575 35388
rect 30631 35386 30637 35388
rect 30391 35334 30393 35386
rect 30573 35334 30575 35386
rect 30329 35332 30335 35334
rect 30391 35332 30415 35334
rect 30471 35332 30495 35334
rect 30551 35332 30575 35334
rect 30631 35332 30637 35334
rect 30329 35323 30637 35332
rect 26424 35284 26476 35290
rect 26424 35226 26476 35232
rect 32876 35086 32904 37217
rect 16580 35080 16632 35086
rect 16580 35022 16632 35028
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 19984 35080 20036 35086
rect 19984 35022 20036 35028
rect 32864 35080 32916 35086
rect 32864 35022 32916 35028
rect 16592 34610 16620 35022
rect 15752 34604 15804 34610
rect 15752 34546 15804 34552
rect 16580 34604 16632 34610
rect 16580 34546 16632 34552
rect 15660 33924 15712 33930
rect 15660 33866 15712 33872
rect 13452 32972 13504 32978
rect 13452 32914 13504 32920
rect 15108 32972 15160 32978
rect 15108 32914 15160 32920
rect 12808 32904 12860 32910
rect 12808 32846 12860 32852
rect 12348 32428 12400 32434
rect 12348 32370 12400 32376
rect 12360 31890 12388 32370
rect 12716 32360 12768 32366
rect 12716 32302 12768 32308
rect 12728 32026 12756 32302
rect 12716 32020 12768 32026
rect 12716 31962 12768 31968
rect 12348 31884 12400 31890
rect 12348 31826 12400 31832
rect 11704 31748 11756 31754
rect 11704 31690 11756 31696
rect 11716 31482 11744 31690
rect 11704 31476 11756 31482
rect 11704 31418 11756 31424
rect 12360 30802 12388 31826
rect 12820 31686 12848 32846
rect 12808 31680 12860 31686
rect 12808 31622 12860 31628
rect 12348 30796 12400 30802
rect 12348 30738 12400 30744
rect 12360 29714 12388 30738
rect 11704 29708 11756 29714
rect 11704 29650 11756 29656
rect 12348 29708 12400 29714
rect 12348 29650 12400 29656
rect 11428 29572 11480 29578
rect 11428 29514 11480 29520
rect 11440 29238 11468 29514
rect 11520 29504 11572 29510
rect 11520 29446 11572 29452
rect 11428 29232 11480 29238
rect 11428 29174 11480 29180
rect 11532 29034 11560 29446
rect 11716 29238 11744 29650
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11520 29028 11572 29034
rect 11520 28970 11572 28976
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11980 28076 12032 28082
rect 11980 28018 12032 28024
rect 11244 28008 11296 28014
rect 11244 27950 11296 27956
rect 11992 27470 12020 28018
rect 12164 28008 12216 28014
rect 12164 27950 12216 27956
rect 10324 27464 10376 27470
rect 10324 27406 10376 27412
rect 11244 27464 11296 27470
rect 11244 27406 11296 27412
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 10152 27130 10180 27270
rect 10140 27124 10192 27130
rect 10140 27066 10192 27072
rect 10336 26586 10364 27406
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 10876 26920 10928 26926
rect 10876 26862 10928 26868
rect 9956 26580 10008 26586
rect 9956 26522 10008 26528
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 9772 26376 9824 26382
rect 9772 26318 9824 26324
rect 9344 26140 9652 26149
rect 9344 26138 9350 26140
rect 9406 26138 9430 26140
rect 9486 26138 9510 26140
rect 9566 26138 9590 26140
rect 9646 26138 9652 26140
rect 9406 26086 9408 26138
rect 9588 26086 9590 26138
rect 9344 26084 9350 26086
rect 9406 26084 9430 26086
rect 9486 26084 9510 26086
rect 9566 26084 9590 26086
rect 9646 26084 9652 26086
rect 9344 26075 9652 26084
rect 9220 25492 9272 25498
rect 9220 25434 9272 25440
rect 9232 24954 9260 25434
rect 9344 25052 9652 25061
rect 9344 25050 9350 25052
rect 9406 25050 9430 25052
rect 9486 25050 9510 25052
rect 9566 25050 9590 25052
rect 9646 25050 9652 25052
rect 9406 24998 9408 25050
rect 9588 24998 9590 25050
rect 9344 24996 9350 24998
rect 9406 24996 9430 24998
rect 9486 24996 9510 24998
rect 9566 24996 9590 24998
rect 9646 24996 9652 24998
rect 9344 24987 9652 24996
rect 9220 24948 9272 24954
rect 9220 24890 9272 24896
rect 9128 24744 9180 24750
rect 9128 24686 9180 24692
rect 9232 24274 9260 24890
rect 9784 24614 9812 26318
rect 9968 25702 9996 26522
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 9864 25220 9916 25226
rect 9864 25162 9916 25168
rect 9876 24954 9904 25162
rect 9968 25158 9996 25638
rect 10888 25294 10916 26862
rect 11072 26450 11100 27270
rect 11256 27130 11284 27406
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 11900 27062 11928 27270
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 11992 26790 12020 27406
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11532 26518 11560 26726
rect 11520 26512 11572 26518
rect 11520 26454 11572 26460
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9864 24948 9916 24954
rect 10888 24936 10916 25230
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 11244 25152 11296 25158
rect 11244 25094 11296 25100
rect 11164 24954 11192 25094
rect 11152 24948 11204 24954
rect 10888 24908 11008 24936
rect 9864 24890 9916 24896
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 9344 23964 9652 23973
rect 9344 23962 9350 23964
rect 9406 23962 9430 23964
rect 9486 23962 9510 23964
rect 9566 23962 9590 23964
rect 9646 23962 9652 23964
rect 9406 23910 9408 23962
rect 9588 23910 9590 23962
rect 9344 23908 9350 23910
rect 9406 23908 9430 23910
rect 9486 23908 9510 23910
rect 9566 23908 9590 23910
rect 9646 23908 9652 23910
rect 9344 23899 9652 23908
rect 9784 23798 9812 24550
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10980 23474 11008 24908
rect 11152 24890 11204 24896
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 11164 24614 11192 24754
rect 11256 24682 11284 25094
rect 11244 24676 11296 24682
rect 11244 24618 11296 24624
rect 11348 24614 11376 25230
rect 11532 24818 11560 26454
rect 12072 25968 12124 25974
rect 12072 25910 12124 25916
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 11716 24818 11744 25230
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11532 24682 11560 24754
rect 11520 24676 11572 24682
rect 11520 24618 11572 24624
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11336 24608 11388 24614
rect 11336 24550 11388 24556
rect 11348 24410 11376 24550
rect 11336 24404 11388 24410
rect 11336 24346 11388 24352
rect 11992 24154 12020 25230
rect 12084 24954 12112 25910
rect 12176 25294 12204 27950
rect 12268 26586 12296 29446
rect 12348 29096 12400 29102
rect 12348 29038 12400 29044
rect 12360 28218 12388 29038
rect 12348 28212 12400 28218
rect 12348 28154 12400 28160
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12360 27130 12388 28018
rect 12532 27872 12584 27878
rect 12532 27814 12584 27820
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12360 26450 12388 27066
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 12544 26382 12572 27814
rect 12820 26772 12848 31622
rect 13464 30258 13492 32914
rect 14740 32904 14792 32910
rect 14740 32846 14792 32852
rect 14752 32502 14780 32846
rect 15120 32570 15148 32914
rect 15384 32836 15436 32842
rect 15384 32778 15436 32784
rect 15396 32570 15424 32778
rect 15108 32564 15160 32570
rect 15108 32506 15160 32512
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 14096 32496 14148 32502
rect 14096 32438 14148 32444
rect 14740 32496 14792 32502
rect 14740 32438 14792 32444
rect 13820 32428 13872 32434
rect 13872 32388 13952 32416
rect 13820 32370 13872 32376
rect 13541 32124 13849 32133
rect 13541 32122 13547 32124
rect 13603 32122 13627 32124
rect 13683 32122 13707 32124
rect 13763 32122 13787 32124
rect 13843 32122 13849 32124
rect 13603 32070 13605 32122
rect 13785 32070 13787 32122
rect 13541 32068 13547 32070
rect 13603 32068 13627 32070
rect 13683 32068 13707 32070
rect 13763 32068 13787 32070
rect 13843 32068 13849 32070
rect 13541 32059 13849 32068
rect 13541 31036 13849 31045
rect 13541 31034 13547 31036
rect 13603 31034 13627 31036
rect 13683 31034 13707 31036
rect 13763 31034 13787 31036
rect 13843 31034 13849 31036
rect 13603 30982 13605 31034
rect 13785 30982 13787 31034
rect 13541 30980 13547 30982
rect 13603 30980 13627 30982
rect 13683 30980 13707 30982
rect 13763 30980 13787 30982
rect 13843 30980 13849 30982
rect 13541 30971 13849 30980
rect 13924 30734 13952 32388
rect 14004 32292 14056 32298
rect 14004 32234 14056 32240
rect 14016 31958 14044 32234
rect 14108 32026 14136 32438
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 14188 32224 14240 32230
rect 14188 32166 14240 32172
rect 14280 32224 14332 32230
rect 14280 32166 14332 32172
rect 14096 32020 14148 32026
rect 14096 31962 14148 31968
rect 14004 31952 14056 31958
rect 14004 31894 14056 31900
rect 14016 31142 14044 31894
rect 14200 31822 14228 32166
rect 14292 32026 14320 32166
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 15028 31822 15056 32370
rect 14188 31816 14240 31822
rect 14188 31758 14240 31764
rect 15016 31816 15068 31822
rect 15016 31758 15068 31764
rect 15028 31346 15056 31758
rect 15120 31754 15148 32506
rect 15764 31754 15792 34546
rect 16488 34536 16540 34542
rect 16488 34478 16540 34484
rect 16764 34536 16816 34542
rect 16764 34478 16816 34484
rect 16500 33862 16528 34478
rect 16776 34202 16804 34478
rect 16764 34196 16816 34202
rect 16764 34138 16816 34144
rect 16488 33856 16540 33862
rect 16488 33798 16540 33804
rect 16500 33130 16528 33798
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16500 33102 16620 33130
rect 16592 32978 16620 33102
rect 16684 33046 16712 33458
rect 17040 33312 17092 33318
rect 17040 33254 17092 33260
rect 16672 33040 16724 33046
rect 16672 32982 16724 32988
rect 16580 32972 16632 32978
rect 16580 32914 16632 32920
rect 16592 31754 16620 32914
rect 16684 32570 16712 32982
rect 17052 32570 17080 33254
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 17040 32564 17092 32570
rect 17040 32506 17092 32512
rect 17144 31906 17172 35022
rect 22284 35012 22336 35018
rect 22284 34954 22336 34960
rect 24216 35012 24268 35018
rect 24216 34954 24268 34960
rect 27068 35012 27120 35018
rect 27068 34954 27120 34960
rect 17738 34844 18046 34853
rect 17738 34842 17744 34844
rect 17800 34842 17824 34844
rect 17880 34842 17904 34844
rect 17960 34842 17984 34844
rect 18040 34842 18046 34844
rect 17800 34790 17802 34842
rect 17982 34790 17984 34842
rect 17738 34788 17744 34790
rect 17800 34788 17824 34790
rect 17880 34788 17904 34790
rect 17960 34788 17984 34790
rect 18040 34788 18046 34790
rect 17738 34779 18046 34788
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 17328 34066 17356 34546
rect 19352 34542 19380 34682
rect 22296 34610 22324 34954
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 19616 34604 19668 34610
rect 19616 34546 19668 34552
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 17592 34536 17644 34542
rect 17592 34478 17644 34484
rect 19340 34536 19392 34542
rect 19340 34478 19392 34484
rect 17604 34202 17632 34478
rect 18788 34400 18840 34406
rect 18788 34342 18840 34348
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 17592 34196 17644 34202
rect 17592 34138 17644 34144
rect 18800 34066 18828 34342
rect 17316 34060 17368 34066
rect 17316 34002 17368 34008
rect 18788 34060 18840 34066
rect 18788 34002 18840 34008
rect 19352 33998 19380 34342
rect 19628 34202 19656 34546
rect 22376 34536 22428 34542
rect 22572 34524 22600 34682
rect 23112 34672 23164 34678
rect 23112 34614 23164 34620
rect 23124 34542 23152 34614
rect 22428 34496 22600 34524
rect 22652 34536 22704 34542
rect 22376 34478 22428 34484
rect 22652 34478 22704 34484
rect 23112 34536 23164 34542
rect 23112 34478 23164 34484
rect 21824 34468 21876 34474
rect 21824 34410 21876 34416
rect 19984 34400 20036 34406
rect 19984 34342 20036 34348
rect 21640 34400 21692 34406
rect 21640 34342 21692 34348
rect 19616 34196 19668 34202
rect 19616 34138 19668 34144
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 19352 33862 19380 33934
rect 19340 33856 19392 33862
rect 19340 33798 19392 33804
rect 17738 33756 18046 33765
rect 17738 33754 17744 33756
rect 17800 33754 17824 33756
rect 17880 33754 17904 33756
rect 17960 33754 17984 33756
rect 18040 33754 18046 33756
rect 17800 33702 17802 33754
rect 17982 33702 17984 33754
rect 17738 33700 17744 33702
rect 17800 33700 17824 33702
rect 17880 33700 17904 33702
rect 17960 33700 17984 33702
rect 18040 33700 18046 33702
rect 17738 33691 18046 33700
rect 17500 33652 17552 33658
rect 17500 33594 17552 33600
rect 17224 33448 17276 33454
rect 17224 33390 17276 33396
rect 17236 32978 17264 33390
rect 17224 32972 17276 32978
rect 17224 32914 17276 32920
rect 17512 32416 17540 33594
rect 19248 33516 19300 33522
rect 19248 33458 19300 33464
rect 19260 32910 19288 33458
rect 19352 33386 19380 33798
rect 19996 33658 20024 34342
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20180 33658 20208 33798
rect 19984 33652 20036 33658
rect 19984 33594 20036 33600
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 19708 33584 19760 33590
rect 19708 33526 19760 33532
rect 19340 33380 19392 33386
rect 19340 33322 19392 33328
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19352 32842 19380 33322
rect 19524 33312 19576 33318
rect 19524 33254 19576 33260
rect 19340 32836 19392 32842
rect 19340 32778 19392 32784
rect 17592 32768 17644 32774
rect 17592 32710 17644 32716
rect 17604 32570 17632 32710
rect 17738 32668 18046 32677
rect 17738 32666 17744 32668
rect 17800 32666 17824 32668
rect 17880 32666 17904 32668
rect 17960 32666 17984 32668
rect 18040 32666 18046 32668
rect 17800 32614 17802 32666
rect 17982 32614 17984 32666
rect 17738 32612 17744 32614
rect 17800 32612 17824 32614
rect 17880 32612 17904 32614
rect 17960 32612 17984 32614
rect 18040 32612 18046 32614
rect 17738 32603 18046 32612
rect 17592 32564 17644 32570
rect 17592 32506 17644 32512
rect 17592 32428 17644 32434
rect 17512 32388 17592 32416
rect 17592 32370 17644 32376
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17408 32360 17460 32366
rect 17408 32302 17460 32308
rect 17420 32026 17448 32302
rect 17592 32292 17644 32298
rect 17592 32234 17644 32240
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17144 31878 17264 31906
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 15120 31726 15332 31754
rect 15764 31726 15884 31754
rect 16592 31726 16712 31754
rect 15200 31408 15252 31414
rect 15200 31350 15252 31356
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 15016 31340 15068 31346
rect 15016 31282 15068 31288
rect 14004 31136 14056 31142
rect 14004 31078 14056 31084
rect 14372 31136 14424 31142
rect 14372 31078 14424 31084
rect 13912 30728 13964 30734
rect 13912 30670 13964 30676
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 13820 30592 13872 30598
rect 13820 30534 13872 30540
rect 13832 30258 13860 30534
rect 14292 30394 14320 30670
rect 14280 30388 14332 30394
rect 14280 30330 14332 30336
rect 13452 30252 13504 30258
rect 13452 30194 13504 30200
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 13912 30252 13964 30258
rect 13912 30194 13964 30200
rect 12992 29504 13044 29510
rect 12992 29446 13044 29452
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 12912 27402 12940 29106
rect 13004 29102 13032 29446
rect 12992 29096 13044 29102
rect 12992 29038 13044 29044
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 12912 26926 12940 27338
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 13084 26920 13136 26926
rect 13084 26862 13136 26868
rect 12820 26744 12940 26772
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12532 25764 12584 25770
rect 12532 25706 12584 25712
rect 12716 25764 12768 25770
rect 12716 25706 12768 25712
rect 12164 25288 12216 25294
rect 12164 25230 12216 25236
rect 12256 25220 12308 25226
rect 12256 25162 12308 25168
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 12072 24948 12124 24954
rect 12072 24890 12124 24896
rect 12176 24886 12204 25094
rect 12268 24954 12296 25162
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 12544 24818 12572 25706
rect 12728 24954 12756 25706
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 11900 24138 12020 24154
rect 11888 24132 12020 24138
rect 11940 24126 12020 24132
rect 11888 24074 11940 24080
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 10244 23118 10272 23462
rect 10980 23446 11100 23474
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 9232 22658 9260 23054
rect 9344 22876 9652 22885
rect 9344 22874 9350 22876
rect 9406 22874 9430 22876
rect 9486 22874 9510 22876
rect 9566 22874 9590 22876
rect 9646 22874 9652 22876
rect 9406 22822 9408 22874
rect 9588 22822 9590 22874
rect 9344 22820 9350 22822
rect 9406 22820 9430 22822
rect 9486 22820 9510 22822
rect 9566 22820 9590 22822
rect 9646 22820 9652 22822
rect 9344 22811 9652 22820
rect 9232 22630 9352 22658
rect 9324 22438 9352 22630
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9324 22098 9352 22374
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9232 21690 9260 21898
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9344 21788 9652 21797
rect 9344 21786 9350 21788
rect 9406 21786 9430 21788
rect 9486 21786 9510 21788
rect 9566 21786 9590 21788
rect 9646 21786 9652 21788
rect 9406 21734 9408 21786
rect 9588 21734 9590 21786
rect 9344 21732 9350 21734
rect 9406 21732 9430 21734
rect 9486 21732 9510 21734
rect 9566 21732 9590 21734
rect 9646 21732 9652 21734
rect 9344 21723 9652 21732
rect 9968 21690 9996 21830
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8956 18986 8984 20402
rect 9048 19854 9076 21490
rect 9692 21146 9720 21490
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9344 20700 9652 20709
rect 9344 20698 9350 20700
rect 9406 20698 9430 20700
rect 9486 20698 9510 20700
rect 9566 20698 9590 20700
rect 9646 20698 9652 20700
rect 9406 20646 9408 20698
rect 9588 20646 9590 20698
rect 9344 20644 9350 20646
rect 9406 20644 9430 20646
rect 9486 20644 9510 20646
rect 9566 20644 9590 20646
rect 9646 20644 9652 20646
rect 9344 20635 9652 20644
rect 10244 20534 10272 23054
rect 11072 22982 11100 23446
rect 11256 23186 11284 24006
rect 12084 23866 12112 24006
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12360 23730 12388 24550
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12360 23322 12388 23666
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 11072 22030 11100 22918
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12268 22234 12296 22510
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12544 22166 12572 22918
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 9692 19854 9720 20470
rect 10612 20466 10640 20538
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9876 20058 9904 20334
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 8956 18958 9076 18986
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 8864 17678 8892 18294
rect 8944 18080 8996 18086
rect 9048 18068 9076 18958
rect 9140 18290 9168 19654
rect 9344 19612 9652 19621
rect 9344 19610 9350 19612
rect 9406 19610 9430 19612
rect 9486 19610 9510 19612
rect 9566 19610 9590 19612
rect 9646 19610 9652 19612
rect 9406 19558 9408 19610
rect 9588 19558 9590 19610
rect 9344 19556 9350 19558
rect 9406 19556 9430 19558
rect 9486 19556 9510 19558
rect 9566 19556 9590 19558
rect 9646 19556 9652 19558
rect 9344 19547 9652 19556
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9784 18970 9812 19246
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9588 18896 9640 18902
rect 9864 18896 9916 18902
rect 9640 18844 9864 18850
rect 9588 18838 9916 18844
rect 9600 18822 9904 18838
rect 9680 18760 9732 18766
rect 9678 18728 9680 18737
rect 9772 18760 9824 18766
rect 9732 18728 9734 18737
rect 9824 18720 9904 18748
rect 9772 18702 9824 18708
rect 9678 18663 9734 18672
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9344 18524 9652 18533
rect 9344 18522 9350 18524
rect 9406 18522 9430 18524
rect 9486 18522 9510 18524
rect 9566 18522 9590 18524
rect 9646 18522 9652 18524
rect 9406 18470 9408 18522
rect 9588 18470 9590 18522
rect 9344 18468 9350 18470
rect 9406 18468 9430 18470
rect 9486 18468 9510 18470
rect 9566 18468 9590 18470
rect 9646 18468 9652 18470
rect 9344 18459 9652 18468
rect 9784 18408 9812 18566
rect 9876 18426 9904 18720
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 9692 18380 9812 18408
rect 9864 18420 9916 18426
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 8996 18040 9076 18068
rect 8944 18022 8996 18028
rect 8944 17808 8996 17814
rect 8942 17776 8944 17785
rect 8996 17776 8998 17785
rect 8942 17711 8998 17720
rect 9048 17678 9076 18040
rect 9140 17746 9168 18226
rect 9324 17785 9352 18226
rect 9692 18222 9720 18380
rect 9864 18362 9916 18368
rect 9772 18284 9824 18290
rect 10060 18272 10088 18634
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10152 18290 10180 18566
rect 9824 18244 10088 18272
rect 10140 18284 10192 18290
rect 9772 18226 9824 18232
rect 10140 18226 10192 18232
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9310 17776 9366 17785
rect 9128 17740 9180 17746
rect 9310 17711 9366 17720
rect 9128 17682 9180 17688
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8772 16425 8800 17478
rect 8850 16688 8906 16697
rect 8956 16674 8984 17614
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8906 16646 8984 16674
rect 8850 16623 8906 16632
rect 8758 16416 8814 16425
rect 8758 16351 8814 16360
rect 8758 16280 8814 16289
rect 8576 16244 8628 16250
rect 8628 16204 8708 16232
rect 8758 16215 8814 16224
rect 8576 16186 8628 16192
rect 8574 16144 8630 16153
rect 8574 16079 8630 16088
rect 8588 15706 8616 16079
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8680 15026 8708 16204
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8574 14784 8630 14793
rect 8574 14719 8630 14728
rect 8404 12192 8524 12220
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8208 11688 8260 11694
rect 8404 11665 8432 12192
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11898 8524 12038
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8208 11630 8260 11636
rect 8390 11656 8446 11665
rect 8116 11620 8168 11626
rect 8446 11614 8524 11642
rect 8390 11591 8446 11600
rect 8116 11562 8168 11568
rect 8128 11354 8156 11562
rect 8208 11552 8260 11558
rect 8392 11552 8444 11558
rect 8208 11494 8260 11500
rect 8390 11520 8392 11529
rect 8444 11520 8446 11529
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8220 11150 8248 11494
rect 8390 11455 8446 11464
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8220 10282 8248 11086
rect 8220 10254 8432 10282
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7668 9674 7696 9862
rect 7668 9646 8064 9674
rect 8036 9586 8064 9646
rect 8220 9586 8248 10134
rect 8404 10062 8432 10254
rect 8496 10198 8524 11614
rect 8588 11082 8616 14719
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8588 10985 8616 11018
rect 8574 10976 8630 10985
rect 8574 10911 8630 10920
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8588 10266 8616 10474
rect 8680 10266 8708 13806
rect 8772 12850 8800 16215
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8864 14618 8892 15982
rect 8956 15638 8984 16646
rect 8944 15632 8996 15638
rect 8944 15574 8996 15580
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 15026 8984 15302
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8956 14822 8984 14962
rect 9048 14958 9076 17274
rect 9232 16998 9260 17478
rect 9344 17436 9652 17445
rect 9344 17434 9350 17436
rect 9406 17434 9430 17436
rect 9486 17434 9510 17436
rect 9566 17434 9590 17436
rect 9646 17434 9652 17436
rect 9406 17382 9408 17434
rect 9588 17382 9590 17434
rect 9344 17380 9350 17382
rect 9406 17380 9430 17382
rect 9486 17380 9510 17382
rect 9566 17380 9590 17382
rect 9646 17380 9652 17382
rect 9344 17371 9652 17380
rect 9692 17270 9720 17614
rect 9784 17270 9812 17818
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9140 16250 9168 16934
rect 9310 16824 9366 16833
rect 9310 16759 9366 16768
rect 9324 16522 9352 16759
rect 9692 16590 9720 16934
rect 9784 16794 9812 17070
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9404 16584 9456 16590
rect 9402 16552 9404 16561
rect 9680 16584 9732 16590
rect 9456 16552 9458 16561
rect 9312 16516 9364 16522
rect 9680 16526 9732 16532
rect 9402 16487 9458 16496
rect 9312 16458 9364 16464
rect 9416 16436 9444 16487
rect 9772 16448 9824 16454
rect 9416 16408 9720 16436
rect 9344 16348 9652 16357
rect 9344 16346 9350 16348
rect 9406 16346 9430 16348
rect 9486 16346 9510 16348
rect 9566 16346 9590 16348
rect 9646 16346 9652 16348
rect 9406 16294 9408 16346
rect 9588 16294 9590 16346
rect 9344 16292 9350 16294
rect 9406 16292 9430 16294
rect 9486 16292 9510 16294
rect 9566 16292 9590 16294
rect 9646 16292 9652 16294
rect 9344 16283 9652 16292
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8864 13818 8892 14554
rect 9140 14414 9168 16186
rect 9692 16114 9720 16408
rect 9772 16390 9824 16396
rect 9680 16108 9732 16114
rect 9416 16068 9680 16096
rect 9218 16008 9274 16017
rect 9218 15943 9274 15952
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 13870 9168 14214
rect 9232 13870 9260 15943
rect 9416 15502 9444 16068
rect 9680 16050 9732 16056
rect 9678 15600 9734 15609
rect 9678 15535 9734 15544
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9600 15366 9628 15438
rect 9692 15434 9720 15535
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9588 15360 9640 15366
rect 9784 15337 9812 16390
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9876 15502 9904 16050
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9864 15360 9916 15366
rect 9588 15302 9640 15308
rect 9770 15328 9826 15337
rect 9864 15302 9916 15308
rect 9344 15260 9652 15269
rect 9770 15263 9826 15272
rect 9344 15258 9350 15260
rect 9406 15258 9430 15260
rect 9486 15258 9510 15260
rect 9566 15258 9590 15260
rect 9646 15258 9652 15260
rect 9406 15206 9408 15258
rect 9588 15206 9590 15258
rect 9344 15204 9350 15206
rect 9406 15204 9430 15206
rect 9486 15204 9510 15206
rect 9566 15204 9590 15206
rect 9646 15204 9652 15206
rect 9344 15195 9652 15204
rect 9784 15162 9812 15263
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9344 14172 9652 14181
rect 9344 14170 9350 14172
rect 9406 14170 9430 14172
rect 9486 14170 9510 14172
rect 9566 14170 9590 14172
rect 9646 14170 9652 14172
rect 9406 14118 9408 14170
rect 9588 14118 9590 14170
rect 9344 14116 9350 14118
rect 9406 14116 9430 14118
rect 9486 14116 9510 14118
rect 9566 14116 9590 14118
rect 9646 14116 9652 14118
rect 9344 14107 9652 14116
rect 9692 13938 9720 14962
rect 9876 14958 9904 15302
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9784 13938 9812 14894
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9876 14074 9904 14486
rect 9968 14414 9996 18022
rect 10244 17728 10272 19926
rect 10336 19854 10364 20198
rect 10428 20058 10456 20402
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10336 18902 10364 19790
rect 10520 19718 10548 20334
rect 10980 20262 11008 21490
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10324 17740 10376 17746
rect 10244 17700 10324 17728
rect 10324 17682 10376 17688
rect 10336 16114 10364 17682
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10324 16108 10376 16114
rect 10244 16068 10324 16096
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10060 15366 10088 15642
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 10244 14278 10272 16068
rect 10324 16050 10376 16056
rect 10428 16046 10456 16934
rect 10704 16538 10732 17614
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16726 10916 16934
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10612 16510 10732 16538
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10520 15706 10548 16050
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10336 14618 10364 14758
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 13938 9904 14010
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9036 13864 9088 13870
rect 8864 13790 8984 13818
rect 9036 13806 9088 13812
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8864 13190 8892 13670
rect 8956 13190 8984 13790
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 11694 8800 12582
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8772 11082 8800 11630
rect 8864 11150 8892 13126
rect 8956 12646 8984 13126
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 9048 12442 9076 13806
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9140 12850 9168 13126
rect 9232 12986 9260 13398
rect 9416 13326 9444 13738
rect 9508 13530 9536 13874
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9344 13084 9652 13093
rect 9344 13082 9350 13084
rect 9406 13082 9430 13084
rect 9486 13082 9510 13084
rect 9566 13082 9590 13084
rect 9646 13082 9652 13084
rect 9406 13030 9408 13082
rect 9588 13030 9590 13082
rect 9344 13028 9350 13030
rect 9406 13028 9430 13030
rect 9486 13028 9510 13030
rect 9566 13028 9590 13030
rect 9646 13028 9652 13030
rect 9344 13019 9652 13028
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9140 12322 9168 12786
rect 8956 12294 9168 12322
rect 8956 11286 8984 12294
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9036 11892 9088 11898
rect 9140 11880 9168 12174
rect 9232 11898 9260 12922
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9310 12472 9366 12481
rect 9310 12407 9366 12416
rect 9324 12374 9352 12407
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9600 12306 9628 12854
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9416 12102 9444 12174
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9344 11996 9652 12005
rect 9344 11994 9350 11996
rect 9406 11994 9430 11996
rect 9486 11994 9510 11996
rect 9566 11994 9590 11996
rect 9646 11994 9652 11996
rect 9406 11942 9408 11994
rect 9588 11942 9590 11994
rect 9344 11940 9350 11942
rect 9406 11940 9430 11942
rect 9486 11940 9510 11942
rect 9566 11940 9590 11942
rect 9646 11940 9652 11942
rect 9344 11931 9652 11940
rect 9088 11852 9168 11880
rect 9220 11892 9272 11898
rect 9036 11834 9088 11840
rect 9220 11834 9272 11840
rect 9784 11830 9812 13874
rect 9864 13796 9916 13802
rect 9916 13756 9996 13784
rect 9864 13738 9916 13744
rect 9968 12374 9996 13756
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9048 11354 9076 11698
rect 9140 11393 9168 11698
rect 9496 11680 9548 11686
rect 9402 11656 9458 11665
rect 9458 11628 9496 11642
rect 9458 11622 9548 11628
rect 9458 11614 9536 11622
rect 9402 11591 9458 11600
rect 9784 11529 9812 11766
rect 9770 11520 9826 11529
rect 9770 11455 9826 11464
rect 9126 11384 9182 11393
rect 9036 11348 9088 11354
rect 9126 11319 9182 11328
rect 9036 11290 9088 11296
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8772 9722 8800 11018
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 4448 9178 4476 9318
rect 5147 9276 5455 9285
rect 5147 9274 5153 9276
rect 5209 9274 5233 9276
rect 5289 9274 5313 9276
rect 5369 9274 5393 9276
rect 5449 9274 5455 9276
rect 5209 9222 5211 9274
rect 5391 9222 5393 9274
rect 5147 9220 5153 9222
rect 5209 9220 5233 9222
rect 5289 9220 5313 9222
rect 5369 9220 5393 9222
rect 5449 9220 5455 9222
rect 5147 9211 5455 9220
rect 8036 9178 8064 9522
rect 8864 9178 8892 11086
rect 8956 9450 8984 11222
rect 9784 11218 9812 11455
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9344 10908 9652 10917
rect 9344 10906 9350 10908
rect 9406 10906 9430 10908
rect 9486 10906 9510 10908
rect 9566 10906 9590 10908
rect 9646 10906 9652 10908
rect 9406 10854 9408 10906
rect 9588 10854 9590 10906
rect 9344 10852 9350 10854
rect 9406 10852 9430 10854
rect 9486 10852 9510 10854
rect 9566 10852 9590 10854
rect 9646 10852 9652 10854
rect 9344 10843 9652 10852
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9692 10062 9720 10746
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9232 9722 9260 9998
rect 9344 9820 9652 9829
rect 9344 9818 9350 9820
rect 9406 9818 9430 9820
rect 9486 9818 9510 9820
rect 9566 9818 9590 9820
rect 9646 9818 9652 9820
rect 9406 9766 9408 9818
rect 9588 9766 9590 9818
rect 9344 9764 9350 9766
rect 9406 9764 9430 9766
rect 9486 9764 9510 9766
rect 9566 9764 9590 9766
rect 9646 9764 9652 9766
rect 9344 9755 9652 9764
rect 9692 9722 9720 9998
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9312 9648 9364 9654
rect 9364 9608 9444 9636
rect 9312 9590 9364 9596
rect 9416 9450 9444 9608
rect 8944 9444 8996 9450
rect 8944 9386 8996 9392
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8956 8974 8984 9386
rect 9508 9042 9536 9658
rect 9600 9178 9628 9658
rect 9876 9586 9904 12106
rect 9968 11558 9996 12310
rect 10244 11762 10272 13942
rect 10336 13870 10364 14554
rect 10428 14074 10456 14962
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10336 11937 10364 12106
rect 10322 11928 10378 11937
rect 10322 11863 10378 11872
rect 10336 11762 10364 11863
rect 10428 11830 10456 13262
rect 10416 11824 10468 11830
rect 10414 11792 10416 11801
rect 10468 11792 10470 11801
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10324 11756 10376 11762
rect 10414 11727 10470 11736
rect 10324 11698 10376 11704
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9968 11354 9996 11494
rect 10060 11393 10088 11494
rect 10046 11384 10102 11393
rect 9956 11348 10008 11354
rect 10046 11319 10102 11328
rect 9956 11290 10008 11296
rect 10244 11150 10272 11698
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10336 11354 10364 11562
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9968 9042 9996 10950
rect 10428 10010 10456 11727
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10060 9982 10456 10010
rect 10060 9722 10088 9982
rect 10428 9926 10456 9982
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10336 9722 10364 9862
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10520 9654 10548 11494
rect 10612 9654 10640 16510
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 16114 10732 16390
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10796 15706 10824 15914
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10704 15434 10732 15506
rect 10888 15502 10916 16662
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10704 13716 10732 15370
rect 10796 15162 10824 15438
rect 10888 15366 10916 15438
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10888 13734 10916 15302
rect 10980 14618 11008 20198
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11072 19718 11100 19858
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 18766 11100 19654
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 15502 11100 18702
rect 11164 18290 11192 21286
rect 11348 20942 11376 21898
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11348 19854 11376 20878
rect 11532 20602 11560 20878
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12268 20369 12296 20402
rect 12254 20360 12310 20369
rect 12254 20295 12310 20304
rect 12268 20058 12296 20295
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11978 19816 12034 19825
rect 11978 19751 12034 19760
rect 11702 19408 11758 19417
rect 11992 19378 12020 19751
rect 11702 19343 11704 19352
rect 11756 19343 11758 19352
rect 11796 19372 11848 19378
rect 11704 19314 11756 19320
rect 11796 19314 11848 19320
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12360 19334 12388 21082
rect 12452 21010 12480 21286
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12452 20466 12480 20946
rect 12544 20942 12572 22102
rect 12820 21962 12848 22510
rect 12808 21956 12860 21962
rect 12808 21898 12860 21904
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12728 21554 12756 21830
rect 12820 21554 12848 21898
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12636 20262 12664 21490
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11164 17542 11192 18226
rect 11348 17678 11376 18702
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11244 17264 11296 17270
rect 11244 17206 11296 17212
rect 11256 16590 11284 17206
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11164 15502 11192 16186
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11164 14482 11192 15438
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10784 13728 10836 13734
rect 10704 13688 10784 13716
rect 10784 13670 10836 13676
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11830 10732 12038
rect 10796 11898 10824 13670
rect 10888 13326 10916 13670
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 12322 11008 12582
rect 11072 12442 11100 14350
rect 11164 13326 11192 14418
rect 11256 14414 11284 16526
rect 11348 16114 11376 17614
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11348 14278 11376 16050
rect 11440 14822 11468 17614
rect 11532 17338 11560 17614
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11624 17202 11652 17614
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11520 15632 11572 15638
rect 11518 15600 11520 15609
rect 11572 15600 11574 15609
rect 11518 15535 11574 15544
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11256 13977 11284 14214
rect 11242 13968 11298 13977
rect 11242 13903 11298 13912
rect 11256 13433 11284 13903
rect 11440 13462 11468 14350
rect 11428 13456 11480 13462
rect 11242 13424 11298 13433
rect 11428 13398 11480 13404
rect 11242 13359 11298 13368
rect 11256 13326 11284 13359
rect 11532 13326 11560 15535
rect 11624 14074 11652 16934
rect 11716 15978 11744 17138
rect 11808 16153 11836 19314
rect 11992 18222 12020 19314
rect 12360 19306 12480 19334
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12070 18728 12126 18737
rect 12070 18663 12072 18672
rect 12124 18663 12126 18672
rect 12072 18634 12124 18640
rect 12360 18426 12388 19178
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11900 16726 11928 17138
rect 11992 16998 12020 18022
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 11794 16144 11850 16153
rect 11794 16079 11850 16088
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11624 13530 11652 14010
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10980 12294 11100 12322
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 11072 11762 11100 12294
rect 11164 12238 11192 13126
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11348 12434 11376 12718
rect 11256 12406 11376 12434
rect 11256 12238 11284 12406
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11440 11830 11468 12106
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11072 10826 11100 11698
rect 11164 11558 11192 11698
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11256 11354 11284 11698
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11354 11376 11494
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11072 10798 11376 10826
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11072 10266 11100 10610
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9761 10916 9998
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10874 9752 10930 9761
rect 10874 9687 10930 9696
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10888 9586 10916 9687
rect 11072 9654 11100 9862
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 10244 8974 10272 9454
rect 10980 9178 11008 9522
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11164 9042 11192 10134
rect 11256 10130 11284 10542
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11256 9586 11284 10066
rect 11244 9580 11296 9586
rect 11348 9568 11376 10798
rect 11716 10130 11744 15914
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11808 14890 11836 15506
rect 11900 15366 11928 15982
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11900 15065 11928 15302
rect 11886 15056 11942 15065
rect 11992 15026 12020 16934
rect 12084 15638 12112 17546
rect 12360 17202 12388 17682
rect 12452 17338 12480 19306
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12268 16590 12296 17138
rect 12452 16658 12480 17274
rect 12544 17184 12572 19994
rect 12636 19378 12664 20198
rect 12820 19514 12848 21490
rect 12912 20584 12940 26744
rect 13096 26586 13124 26862
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 13188 23798 13216 28358
rect 13464 28150 13492 30194
rect 13541 29948 13849 29957
rect 13541 29946 13547 29948
rect 13603 29946 13627 29948
rect 13683 29946 13707 29948
rect 13763 29946 13787 29948
rect 13843 29946 13849 29948
rect 13603 29894 13605 29946
rect 13785 29894 13787 29946
rect 13541 29892 13547 29894
rect 13603 29892 13627 29894
rect 13683 29892 13707 29894
rect 13763 29892 13787 29894
rect 13843 29892 13849 29894
rect 13541 29883 13849 29892
rect 13924 29578 13952 30194
rect 14004 30184 14056 30190
rect 14004 30126 14056 30132
rect 14016 29646 14044 30126
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 14004 29640 14056 29646
rect 14004 29582 14056 29588
rect 13912 29572 13964 29578
rect 13912 29514 13964 29520
rect 13924 29322 13952 29514
rect 13832 29294 13952 29322
rect 13832 29238 13860 29294
rect 13820 29232 13872 29238
rect 13820 29174 13872 29180
rect 14016 29170 14044 29582
rect 14004 29164 14056 29170
rect 14004 29106 14056 29112
rect 13541 28860 13849 28869
rect 13541 28858 13547 28860
rect 13603 28858 13627 28860
rect 13683 28858 13707 28860
rect 13763 28858 13787 28860
rect 13843 28858 13849 28860
rect 13603 28806 13605 28858
rect 13785 28806 13787 28858
rect 13541 28804 13547 28806
rect 13603 28804 13627 28806
rect 13683 28804 13707 28806
rect 13763 28804 13787 28806
rect 13843 28804 13849 28806
rect 13541 28795 13849 28804
rect 14108 28626 14136 29650
rect 14384 29034 14412 31078
rect 14844 30938 14872 31282
rect 14832 30932 14884 30938
rect 14832 30874 14884 30880
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 14568 29850 14596 30670
rect 15212 30394 15240 31350
rect 15304 30802 15332 31726
rect 15568 31136 15620 31142
rect 15568 31078 15620 31084
rect 15580 30802 15608 31078
rect 15292 30796 15344 30802
rect 15292 30738 15344 30744
rect 15568 30796 15620 30802
rect 15568 30738 15620 30744
rect 15660 30660 15712 30666
rect 15660 30602 15712 30608
rect 15568 30592 15620 30598
rect 15568 30534 15620 30540
rect 15580 30394 15608 30534
rect 15672 30394 15700 30602
rect 15200 30388 15252 30394
rect 15200 30330 15252 30336
rect 15568 30388 15620 30394
rect 15568 30330 15620 30336
rect 15660 30388 15712 30394
rect 15660 30330 15712 30336
rect 15752 30184 15804 30190
rect 15752 30126 15804 30132
rect 14556 29844 14608 29850
rect 14556 29786 14608 29792
rect 14568 29102 14596 29786
rect 15476 29640 15528 29646
rect 15476 29582 15528 29588
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 15028 29306 15056 29446
rect 15488 29306 15516 29582
rect 15016 29300 15068 29306
rect 15016 29242 15068 29248
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 14556 29096 14608 29102
rect 14556 29038 14608 29044
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14372 29028 14424 29034
rect 14372 28970 14424 28976
rect 14280 28960 14332 28966
rect 14280 28902 14332 28908
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 14292 28490 14320 28902
rect 14280 28484 14332 28490
rect 14280 28426 14332 28432
rect 13452 28144 13504 28150
rect 13452 28086 13504 28092
rect 13541 27772 13849 27781
rect 13541 27770 13547 27772
rect 13603 27770 13627 27772
rect 13683 27770 13707 27772
rect 13763 27770 13787 27772
rect 13843 27770 13849 27772
rect 13603 27718 13605 27770
rect 13785 27718 13787 27770
rect 13541 27716 13547 27718
rect 13603 27716 13627 27718
rect 13683 27716 13707 27718
rect 13763 27716 13787 27718
rect 13843 27716 13849 27718
rect 13541 27707 13849 27716
rect 13912 27464 13964 27470
rect 13912 27406 13964 27412
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 13372 27130 13400 27338
rect 13360 27124 13412 27130
rect 13360 27066 13412 27072
rect 13924 26790 13952 27406
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 13541 26684 13849 26693
rect 13541 26682 13547 26684
rect 13603 26682 13627 26684
rect 13683 26682 13707 26684
rect 13763 26682 13787 26684
rect 13843 26682 13849 26684
rect 13603 26630 13605 26682
rect 13785 26630 13787 26682
rect 13541 26628 13547 26630
rect 13603 26628 13627 26630
rect 13683 26628 13707 26630
rect 13763 26628 13787 26630
rect 13843 26628 13849 26630
rect 13541 26619 13849 26628
rect 13924 26382 13952 26726
rect 14108 26586 14136 27406
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14292 27130 14320 27270
rect 14280 27124 14332 27130
rect 14280 27066 14332 27072
rect 14384 26874 14412 28970
rect 14660 27538 14688 29038
rect 15764 28762 15792 30126
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 14648 27532 14700 27538
rect 14648 27474 14700 27480
rect 15856 27470 15884 31726
rect 16684 30734 16712 31726
rect 17144 31482 17172 31758
rect 17132 31476 17184 31482
rect 17132 31418 17184 31424
rect 17040 30864 17092 30870
rect 17040 30806 17092 30812
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16592 29034 16620 30126
rect 16684 29510 16712 30670
rect 17052 30394 17080 30806
rect 17040 30388 17092 30394
rect 17040 30330 17092 30336
rect 16672 29504 16724 29510
rect 17132 29504 17184 29510
rect 16672 29446 16724 29452
rect 17052 29464 17132 29492
rect 16580 29028 16632 29034
rect 16580 28970 16632 28976
rect 16592 28762 16620 28970
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16580 28484 16632 28490
rect 16684 28472 16712 29446
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 16960 28694 16988 29106
rect 17052 29034 17080 29464
rect 17132 29446 17184 29452
rect 17040 29028 17092 29034
rect 17040 28970 17092 28976
rect 16948 28688 17000 28694
rect 16948 28630 17000 28636
rect 16632 28444 16712 28472
rect 16580 28426 16632 28432
rect 16028 27600 16080 27606
rect 16028 27542 16080 27548
rect 15384 27464 15436 27470
rect 15384 27406 15436 27412
rect 15844 27464 15896 27470
rect 15844 27406 15896 27412
rect 15396 27062 15424 27406
rect 16040 27130 16068 27542
rect 16028 27124 16080 27130
rect 16028 27066 16080 27072
rect 15384 27056 15436 27062
rect 15384 26998 15436 27004
rect 14464 26920 14516 26926
rect 14384 26868 14464 26874
rect 14384 26862 14516 26868
rect 14384 26846 14504 26862
rect 14384 26586 14412 26846
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 14372 26580 14424 26586
rect 14372 26522 14424 26528
rect 14844 26382 14872 26726
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14832 26376 14884 26382
rect 14832 26318 14884 26324
rect 13541 25596 13849 25605
rect 13541 25594 13547 25596
rect 13603 25594 13627 25596
rect 13683 25594 13707 25596
rect 13763 25594 13787 25596
rect 13843 25594 13849 25596
rect 13603 25542 13605 25594
rect 13785 25542 13787 25594
rect 13541 25540 13547 25542
rect 13603 25540 13627 25542
rect 13683 25540 13707 25542
rect 13763 25540 13787 25542
rect 13843 25540 13849 25542
rect 13541 25531 13849 25540
rect 13924 25294 13952 26318
rect 14568 25702 14596 26318
rect 14740 26308 14792 26314
rect 14740 26250 14792 26256
rect 14752 25906 14780 26250
rect 14844 25906 14872 26318
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14556 25696 14608 25702
rect 14556 25638 14608 25644
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13636 25220 13688 25226
rect 13636 25162 13688 25168
rect 13648 24954 13676 25162
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13924 24818 13952 25230
rect 14568 25226 14596 25638
rect 14556 25220 14608 25226
rect 14556 25162 14608 25168
rect 15396 24954 15424 26998
rect 16212 26920 16264 26926
rect 16212 26862 16264 26868
rect 16224 25226 16252 26862
rect 16488 26784 16540 26790
rect 16488 26726 16540 26732
rect 16500 26586 16528 26726
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16592 26314 16620 28426
rect 16856 27464 16908 27470
rect 16856 27406 16908 27412
rect 16672 27396 16724 27402
rect 16672 27338 16724 27344
rect 16684 27130 16712 27338
rect 16868 27130 16896 27406
rect 16960 27130 16988 28630
rect 17052 28490 17080 28970
rect 17040 28484 17092 28490
rect 17040 28426 17092 28432
rect 17040 28144 17092 28150
rect 17040 28086 17092 28092
rect 17052 27334 17080 28086
rect 17040 27328 17092 27334
rect 17040 27270 17092 27276
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16776 26450 16804 26862
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16776 25362 16804 26386
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16212 25220 16264 25226
rect 16212 25162 16264 25168
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15108 24880 15160 24886
rect 15108 24822 15160 24828
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13541 24508 13849 24517
rect 13541 24506 13547 24508
rect 13603 24506 13627 24508
rect 13683 24506 13707 24508
rect 13763 24506 13787 24508
rect 13843 24506 13849 24508
rect 13603 24454 13605 24506
rect 13785 24454 13787 24506
rect 13541 24452 13547 24454
rect 13603 24452 13627 24454
rect 13683 24452 13707 24454
rect 13763 24452 13787 24454
rect 13843 24452 13849 24454
rect 13541 24443 13849 24452
rect 13924 23866 13952 24754
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 15028 24410 15056 24686
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 15120 23798 15148 24822
rect 15856 24206 15884 25094
rect 16500 24954 16528 25230
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16948 25220 17000 25226
rect 16948 25162 17000 25168
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 16592 24342 16620 25162
rect 16960 24818 16988 25162
rect 17052 24818 17080 27270
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 16580 24336 16632 24342
rect 16580 24278 16632 24284
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 13176 23792 13228 23798
rect 14464 23792 14516 23798
rect 13176 23734 13228 23740
rect 14384 23752 14464 23780
rect 13541 23420 13849 23429
rect 13541 23418 13547 23420
rect 13603 23418 13627 23420
rect 13683 23418 13707 23420
rect 13763 23418 13787 23420
rect 13843 23418 13849 23420
rect 13603 23366 13605 23418
rect 13785 23366 13787 23418
rect 13541 23364 13547 23366
rect 13603 23364 13627 23366
rect 13683 23364 13707 23366
rect 13763 23364 13787 23366
rect 13843 23364 13849 23366
rect 13541 23355 13849 23364
rect 13176 22772 13228 22778
rect 13176 22714 13228 22720
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13004 21690 13032 21966
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 13188 21010 13216 22714
rect 14384 22710 14412 23752
rect 14464 23734 14516 23740
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 14924 23520 14976 23526
rect 14924 23462 14976 23468
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 13541 22332 13849 22341
rect 13541 22330 13547 22332
rect 13603 22330 13627 22332
rect 13683 22330 13707 22332
rect 13763 22330 13787 22332
rect 13843 22330 13849 22332
rect 13603 22278 13605 22330
rect 13785 22278 13787 22330
rect 13541 22276 13547 22278
rect 13603 22276 13627 22278
rect 13683 22276 13707 22278
rect 13763 22276 13787 22278
rect 13843 22276 13849 22278
rect 13541 22267 13849 22276
rect 14384 22166 14412 22646
rect 14372 22160 14424 22166
rect 14292 22108 14372 22114
rect 14292 22102 14424 22108
rect 14292 22086 14412 22102
rect 14292 22030 14320 22086
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14108 21690 14136 21830
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 13280 21146 13308 21354
rect 13541 21244 13849 21253
rect 13541 21242 13547 21244
rect 13603 21242 13627 21244
rect 13683 21242 13707 21244
rect 13763 21242 13787 21244
rect 13843 21242 13849 21244
rect 13603 21190 13605 21242
rect 13785 21190 13787 21242
rect 13541 21188 13547 21190
rect 13603 21188 13627 21190
rect 13683 21188 13707 21190
rect 13763 21188 13787 21190
rect 13843 21188 13849 21190
rect 13541 21179 13849 21188
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 12912 20556 13032 20584
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12912 19417 12940 20402
rect 12898 19408 12954 19417
rect 12624 19372 12676 19378
rect 12898 19343 12954 19352
rect 12624 19314 12676 19320
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12820 18290 12848 18702
rect 12912 18290 12940 19343
rect 13004 18970 13032 20556
rect 13188 19378 13216 20946
rect 14752 20942 14780 21830
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14752 20466 14780 20878
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 13541 20156 13849 20165
rect 13541 20154 13547 20156
rect 13603 20154 13627 20156
rect 13683 20154 13707 20156
rect 13763 20154 13787 20156
rect 13843 20154 13849 20156
rect 13603 20102 13605 20154
rect 13785 20102 13787 20154
rect 13541 20100 13547 20102
rect 13603 20100 13627 20102
rect 13683 20100 13707 20102
rect 13763 20100 13787 20102
rect 13843 20100 13849 20102
rect 13541 20091 13849 20100
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13464 19514 13492 19722
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12728 18170 12756 18226
rect 12992 18216 13044 18222
rect 12728 18142 12848 18170
rect 12992 18158 13044 18164
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17746 12756 18022
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12544 17156 12664 17184
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 12164 15428 12216 15434
rect 12164 15370 12216 15376
rect 12176 15337 12204 15370
rect 12162 15328 12218 15337
rect 12218 15286 12388 15314
rect 12162 15263 12218 15272
rect 12360 15026 12388 15286
rect 11886 14991 11888 15000
rect 11940 14991 11942 15000
rect 11980 15020 12032 15026
rect 11888 14962 11940 14968
rect 11980 14962 12032 14968
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 11900 12918 11928 14962
rect 11992 12986 12020 14962
rect 12452 14414 12480 16594
rect 12544 16250 12572 17002
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12636 15162 12664 17156
rect 12728 17066 12756 17682
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12820 16946 12848 18142
rect 13004 17202 13032 18158
rect 13188 17746 13216 19314
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13280 18698 13308 19110
rect 13464 18850 13492 19450
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13541 19068 13849 19077
rect 13541 19066 13547 19068
rect 13603 19066 13627 19068
rect 13683 19066 13707 19068
rect 13763 19066 13787 19068
rect 13843 19066 13849 19068
rect 13603 19014 13605 19066
rect 13785 19014 13787 19066
rect 13541 19012 13547 19014
rect 13603 19012 13627 19014
rect 13683 19012 13707 19014
rect 13763 19012 13787 19014
rect 13843 19012 13849 19014
rect 13541 19003 13849 19012
rect 13464 18822 13584 18850
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13280 18290 13308 18634
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17202 13124 17478
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13084 17196 13136 17202
rect 13268 17196 13320 17202
rect 13084 17138 13136 17144
rect 13188 17156 13268 17184
rect 13188 16946 13216 17156
rect 13268 17138 13320 17144
rect 12820 16918 13216 16946
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12820 14929 12848 16050
rect 12806 14920 12862 14929
rect 12806 14855 12862 14864
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12544 14414 12572 14554
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12532 14408 12584 14414
rect 12584 14368 12664 14396
rect 12532 14350 12584 14356
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12084 13326 12112 14214
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12176 13326 12204 13738
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11900 11937 11928 12038
rect 11886 11928 11942 11937
rect 11886 11863 11888 11872
rect 11940 11863 11942 11872
rect 11888 11834 11940 11840
rect 11886 11792 11942 11801
rect 11886 11727 11888 11736
rect 11940 11727 11942 11736
rect 11888 11698 11940 11704
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11440 9722 11468 10066
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11428 9580 11480 9586
rect 11348 9540 11428 9568
rect 11244 9522 11296 9528
rect 11428 9522 11480 9528
rect 11256 9382 11284 9522
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11532 9178 11560 9998
rect 11624 9722 11652 9998
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11716 9450 11744 9590
rect 11808 9586 11836 9998
rect 11992 9602 12020 12378
rect 12084 11898 12112 13262
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12176 11234 12204 12922
rect 12084 11206 12204 11234
rect 12084 10062 12112 11206
rect 12268 10062 12296 13466
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12360 11354 12388 11698
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12162 9616 12218 9625
rect 11992 9586 12162 9602
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11980 9580 12162 9586
rect 12032 9574 12162 9580
rect 12162 9551 12218 9560
rect 11980 9522 12032 9528
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 12268 9058 12296 9998
rect 12360 9178 12388 10406
rect 12452 9761 12480 12922
rect 12544 12442 12572 13126
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12544 11150 12572 12174
rect 12636 11744 12664 14368
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12728 13530 12756 13738
rect 12912 13734 12940 16918
rect 13372 16522 13400 17614
rect 13464 17202 13492 18702
rect 13556 18272 13584 18822
rect 13728 18284 13780 18290
rect 13556 18244 13728 18272
rect 13728 18226 13780 18232
rect 13541 17980 13849 17989
rect 13541 17978 13547 17980
rect 13603 17978 13627 17980
rect 13683 17978 13707 17980
rect 13763 17978 13787 17980
rect 13843 17978 13849 17980
rect 13603 17926 13605 17978
rect 13785 17926 13787 17978
rect 13541 17924 13547 17926
rect 13603 17924 13627 17926
rect 13683 17924 13707 17926
rect 13763 17924 13787 17926
rect 13843 17924 13849 17926
rect 13541 17915 13849 17924
rect 13924 17678 13952 19110
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13556 16980 13584 17138
rect 13912 17060 13964 17066
rect 13912 17002 13964 17008
rect 13464 16952 13584 16980
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 13004 13938 13032 15370
rect 13096 15162 13124 15846
rect 13280 15706 13308 15914
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 13096 14550 13124 14826
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13096 14074 13124 14350
rect 13188 14074 13216 15302
rect 13464 15144 13492 16952
rect 13541 16892 13849 16901
rect 13541 16890 13547 16892
rect 13603 16890 13627 16892
rect 13683 16890 13707 16892
rect 13763 16890 13787 16892
rect 13843 16890 13849 16892
rect 13603 16838 13605 16890
rect 13785 16838 13787 16890
rect 13541 16836 13547 16838
rect 13603 16836 13627 16838
rect 13683 16836 13707 16838
rect 13763 16836 13787 16838
rect 13843 16836 13849 16838
rect 13541 16827 13849 16836
rect 13924 16794 13952 17002
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13544 16652 13596 16658
rect 13596 16612 14044 16640
rect 13544 16594 13596 16600
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13556 15978 13584 16458
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13541 15804 13849 15813
rect 13541 15802 13547 15804
rect 13603 15802 13627 15804
rect 13683 15802 13707 15804
rect 13763 15802 13787 15804
rect 13843 15802 13849 15804
rect 13603 15750 13605 15802
rect 13785 15750 13787 15802
rect 13541 15748 13547 15750
rect 13603 15748 13627 15750
rect 13683 15748 13707 15750
rect 13763 15748 13787 15750
rect 13843 15748 13849 15750
rect 13541 15739 13849 15748
rect 13280 15116 13492 15144
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12728 12434 12756 13262
rect 12820 12986 12848 13262
rect 12912 13190 12940 13262
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12728 12406 12848 12434
rect 12716 12232 12768 12238
rect 12714 12200 12716 12209
rect 12768 12200 12770 12209
rect 12714 12135 12770 12144
rect 12716 11756 12768 11762
rect 12636 11716 12716 11744
rect 12716 11698 12768 11704
rect 12532 11144 12584 11150
rect 12530 11112 12532 11121
rect 12624 11144 12676 11150
rect 12584 11112 12586 11121
rect 12624 11086 12676 11092
rect 12530 11047 12586 11056
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10130 12572 10950
rect 12636 10470 12664 11086
rect 12728 10674 12756 11698
rect 12820 10742 12848 12406
rect 12912 11898 12940 13126
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12900 11280 12952 11286
rect 13004 11268 13032 12038
rect 13096 11354 13124 13398
rect 13174 11928 13230 11937
rect 13280 11898 13308 15116
rect 13450 15056 13506 15065
rect 13360 15020 13412 15026
rect 13450 14991 13452 15000
rect 13360 14962 13412 14968
rect 13504 14991 13506 15000
rect 13912 15020 13964 15026
rect 13452 14962 13504 14968
rect 13912 14962 13964 14968
rect 13372 14278 13400 14962
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14414 13492 14758
rect 13541 14716 13849 14725
rect 13541 14714 13547 14716
rect 13603 14714 13627 14716
rect 13683 14714 13707 14716
rect 13763 14714 13787 14716
rect 13843 14714 13849 14716
rect 13603 14662 13605 14714
rect 13785 14662 13787 14714
rect 13541 14660 13547 14662
rect 13603 14660 13627 14662
rect 13683 14660 13707 14662
rect 13763 14660 13787 14662
rect 13843 14660 13849 14662
rect 13541 14651 13849 14660
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13360 14000 13412 14006
rect 13358 13968 13360 13977
rect 13412 13968 13414 13977
rect 13358 13903 13414 13912
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13372 13530 13400 13806
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13372 12238 13400 13194
rect 13464 12434 13492 14350
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13648 14006 13676 14282
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13924 13938 13952 14962
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13832 13784 13860 13874
rect 13832 13756 13952 13784
rect 13541 13628 13849 13637
rect 13541 13626 13547 13628
rect 13603 13626 13627 13628
rect 13683 13626 13707 13628
rect 13763 13626 13787 13628
rect 13843 13626 13849 13628
rect 13603 13574 13605 13626
rect 13785 13574 13787 13626
rect 13541 13572 13547 13574
rect 13603 13572 13627 13574
rect 13683 13572 13707 13574
rect 13763 13572 13787 13574
rect 13843 13572 13849 13574
rect 13541 13563 13849 13572
rect 13541 12540 13849 12549
rect 13541 12538 13547 12540
rect 13603 12538 13627 12540
rect 13683 12538 13707 12540
rect 13763 12538 13787 12540
rect 13843 12538 13849 12540
rect 13603 12486 13605 12538
rect 13785 12486 13787 12538
rect 13541 12484 13547 12486
rect 13603 12484 13627 12486
rect 13683 12484 13707 12486
rect 13763 12484 13787 12486
rect 13843 12484 13849 12486
rect 13541 12475 13849 12484
rect 13464 12406 13676 12434
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13174 11863 13230 11872
rect 13268 11892 13320 11898
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12952 11240 13032 11268
rect 12900 11222 12952 11228
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12912 10062 12940 11222
rect 13096 10606 13124 11290
rect 13188 10606 13216 11863
rect 13268 11834 13320 11840
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12438 9752 12494 9761
rect 12438 9687 12494 9696
rect 12452 9586 12480 9687
rect 12636 9654 12664 9998
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12452 9058 12480 9318
rect 11152 9036 11204 9042
rect 12268 9030 12480 9058
rect 11152 8978 11204 8984
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 12256 8968 12308 8974
rect 12544 8956 12572 9522
rect 13004 9382 13032 9862
rect 13096 9722 13124 9862
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13188 9654 13216 10134
rect 13280 9654 13308 11018
rect 13372 11014 13400 12174
rect 13464 11898 13492 12310
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13648 11830 13676 12406
rect 13726 11928 13782 11937
rect 13726 11863 13782 11872
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13740 11762 13768 11863
rect 13544 11756 13596 11762
rect 13464 11716 13544 11744
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13372 9586 13400 10542
rect 13464 10266 13492 11716
rect 13544 11698 13596 11704
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13541 11452 13849 11461
rect 13541 11450 13547 11452
rect 13603 11450 13627 11452
rect 13683 11450 13707 11452
rect 13763 11450 13787 11452
rect 13843 11450 13849 11452
rect 13603 11398 13605 11450
rect 13785 11398 13787 11450
rect 13541 11396 13547 11398
rect 13603 11396 13627 11398
rect 13683 11396 13707 11398
rect 13763 11396 13787 11398
rect 13843 11396 13849 11398
rect 13541 11387 13849 11396
rect 13924 11354 13952 13756
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14016 11218 14044 16612
rect 14108 15026 14136 18702
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 14618 14136 14826
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 12714 14136 14214
rect 14200 13938 14228 16934
rect 14384 16590 14412 20198
rect 14752 19446 14780 20402
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14568 17678 14596 18226
rect 14740 18216 14792 18222
rect 14660 18164 14740 18170
rect 14660 18158 14792 18164
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14660 18142 14780 18158
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14660 17542 14688 18142
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14660 17338 14688 17478
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 14414 14320 16390
rect 14752 14890 14780 18022
rect 14844 17882 14872 18158
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14936 17202 14964 23462
rect 15120 23050 15148 23734
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 15108 23044 15160 23050
rect 15108 22986 15160 22992
rect 15660 23044 15712 23050
rect 15660 22986 15712 22992
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15108 18284 15160 18290
rect 15160 18244 15240 18272
rect 15108 18226 15160 18232
rect 15212 18086 15240 18244
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 15120 16794 15148 18022
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15028 16114 15056 16526
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15120 15638 15148 16730
rect 15212 16590 15240 17070
rect 15304 16998 15332 19450
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15396 16794 15424 22918
rect 15672 22778 15700 22986
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15856 22030 15884 22918
rect 16408 22778 16436 23054
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16592 22642 16620 24278
rect 16764 23792 16816 23798
rect 16764 23734 16816 23740
rect 16776 23050 16804 23734
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16948 22704 17000 22710
rect 16948 22646 17000 22652
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15856 21690 15884 21966
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15856 21010 15884 21626
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15948 21146 15976 21286
rect 16316 21146 16344 21490
rect 16960 21350 16988 22646
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15856 20602 15884 20946
rect 15844 20596 15896 20602
rect 17052 20584 17080 24754
rect 17236 22094 17264 31878
rect 17604 31822 17632 32234
rect 17788 32026 17816 32370
rect 17776 32020 17828 32026
rect 17776 31962 17828 31968
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17500 31748 17552 31754
rect 17500 31690 17552 31696
rect 17512 31414 17540 31690
rect 17604 31464 17632 31758
rect 19352 31754 19380 32778
rect 19536 32774 19564 33254
rect 19720 33114 19748 33526
rect 20536 33516 20588 33522
rect 20536 33458 20588 33464
rect 20548 33318 20576 33458
rect 20732 33454 20760 33798
rect 21652 33658 21680 34342
rect 21088 33652 21140 33658
rect 21088 33594 21140 33600
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 20720 33448 20772 33454
rect 20720 33390 20772 33396
rect 20536 33312 20588 33318
rect 20536 33254 20588 33260
rect 20996 33312 21048 33318
rect 20996 33254 21048 33260
rect 19708 33108 19760 33114
rect 19708 33050 19760 33056
rect 19524 32768 19576 32774
rect 19524 32710 19576 32716
rect 19616 32768 19668 32774
rect 19616 32710 19668 32716
rect 19536 32026 19564 32710
rect 19628 32570 19656 32710
rect 19616 32564 19668 32570
rect 19616 32506 19668 32512
rect 20548 32434 20576 33254
rect 21008 32910 21036 33254
rect 20996 32904 21048 32910
rect 20996 32846 21048 32852
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20720 32428 20772 32434
rect 20720 32370 20772 32376
rect 19984 32292 20036 32298
rect 19984 32234 20036 32240
rect 19524 32020 19576 32026
rect 19524 31962 19576 31968
rect 19996 31958 20024 32234
rect 20168 32224 20220 32230
rect 20168 32166 20220 32172
rect 20180 31958 20208 32166
rect 19984 31952 20036 31958
rect 19984 31894 20036 31900
rect 20168 31952 20220 31958
rect 20168 31894 20220 31900
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19708 31816 19760 31822
rect 19708 31758 19760 31764
rect 18880 31748 18932 31754
rect 18880 31690 18932 31696
rect 19260 31726 19380 31754
rect 17738 31580 18046 31589
rect 17738 31578 17744 31580
rect 17800 31578 17824 31580
rect 17880 31578 17904 31580
rect 17960 31578 17984 31580
rect 18040 31578 18046 31580
rect 17800 31526 17802 31578
rect 17982 31526 17984 31578
rect 17738 31524 17744 31526
rect 17800 31524 17824 31526
rect 17880 31524 17904 31526
rect 17960 31524 17984 31526
rect 18040 31524 18046 31526
rect 17738 31515 18046 31524
rect 17604 31436 17724 31464
rect 17500 31408 17552 31414
rect 17500 31350 17552 31356
rect 17512 30870 17540 31350
rect 17696 31346 17724 31436
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17684 31204 17736 31210
rect 17684 31146 17736 31152
rect 17696 30870 17724 31146
rect 17776 31136 17828 31142
rect 17776 31078 17828 31084
rect 17788 30870 17816 31078
rect 17880 30938 17908 31282
rect 18892 30938 18920 31690
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 18880 30932 18932 30938
rect 18880 30874 18932 30880
rect 17500 30864 17552 30870
rect 17500 30806 17552 30812
rect 17684 30864 17736 30870
rect 17684 30806 17736 30812
rect 17776 30864 17828 30870
rect 17776 30806 17828 30812
rect 17592 30796 17644 30802
rect 17592 30738 17644 30744
rect 17408 30660 17460 30666
rect 17408 30602 17460 30608
rect 17420 30190 17448 30602
rect 17408 30184 17460 30190
rect 17408 30126 17460 30132
rect 17420 29730 17448 30126
rect 17604 30054 17632 30738
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 17738 30492 18046 30501
rect 17738 30490 17744 30492
rect 17800 30490 17824 30492
rect 17880 30490 17904 30492
rect 17960 30490 17984 30492
rect 18040 30490 18046 30492
rect 17800 30438 17802 30490
rect 17982 30438 17984 30490
rect 17738 30436 17744 30438
rect 17800 30436 17824 30438
rect 17880 30436 17904 30438
rect 17960 30436 17984 30438
rect 18040 30436 18046 30438
rect 17738 30427 18046 30436
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 17420 29702 17540 29730
rect 17512 29646 17540 29702
rect 17604 29646 17632 29990
rect 18156 29850 18184 30670
rect 18144 29844 18196 29850
rect 18144 29786 18196 29792
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17500 29640 17552 29646
rect 17500 29582 17552 29588
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17420 29306 17448 29582
rect 18144 29572 18196 29578
rect 18144 29514 18196 29520
rect 17738 29404 18046 29413
rect 17738 29402 17744 29404
rect 17800 29402 17824 29404
rect 17880 29402 17904 29404
rect 17960 29402 17984 29404
rect 18040 29402 18046 29404
rect 17800 29350 17802 29402
rect 17982 29350 17984 29402
rect 17738 29348 17744 29350
rect 17800 29348 17824 29350
rect 17880 29348 17904 29350
rect 17960 29348 17984 29350
rect 18040 29348 18046 29350
rect 17738 29339 18046 29348
rect 18156 29306 18184 29514
rect 18604 29504 18656 29510
rect 18604 29446 18656 29452
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18616 29170 18644 29446
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18604 29164 18656 29170
rect 18604 29106 18656 29112
rect 18788 29164 18840 29170
rect 18788 29106 18840 29112
rect 17500 29096 17552 29102
rect 17500 29038 17552 29044
rect 17776 29096 17828 29102
rect 17828 29056 18000 29084
rect 17776 29038 17828 29044
rect 17512 28422 17540 29038
rect 17972 28762 18000 29056
rect 17960 28756 18012 28762
rect 17960 28698 18012 28704
rect 18524 28558 18552 29106
rect 18616 28626 18644 29106
rect 18604 28620 18656 28626
rect 18604 28562 18656 28568
rect 18800 28558 18828 29106
rect 18892 28966 18920 30874
rect 19260 29714 19288 31726
rect 19444 31482 19472 31758
rect 19616 31680 19668 31686
rect 19616 31622 19668 31628
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19628 31414 19656 31622
rect 19616 31408 19668 31414
rect 19616 31350 19668 31356
rect 19720 31346 19748 31758
rect 20180 31754 20208 31894
rect 20088 31726 20208 31754
rect 19708 31340 19760 31346
rect 19708 31282 19760 31288
rect 20088 31226 20116 31726
rect 20364 31482 20392 32370
rect 20548 31754 20576 32370
rect 20732 32298 20760 32370
rect 21008 32366 21036 32846
rect 21100 32366 21128 33594
rect 21836 33454 21864 34410
rect 21935 34300 22243 34309
rect 21935 34298 21941 34300
rect 21997 34298 22021 34300
rect 22077 34298 22101 34300
rect 22157 34298 22181 34300
rect 22237 34298 22243 34300
rect 21997 34246 21999 34298
rect 22179 34246 22181 34298
rect 21935 34244 21941 34246
rect 21997 34244 22021 34246
rect 22077 34244 22101 34246
rect 22157 34244 22181 34246
rect 22237 34244 22243 34246
rect 21935 34235 22243 34244
rect 22664 34202 22692 34478
rect 22652 34196 22704 34202
rect 22652 34138 22704 34144
rect 23124 33590 23152 34478
rect 24124 34400 24176 34406
rect 24124 34342 24176 34348
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23112 33584 23164 33590
rect 23032 33544 23112 33572
rect 21824 33448 21876 33454
rect 21824 33390 21876 33396
rect 22192 33448 22244 33454
rect 22244 33396 22324 33402
rect 22192 33390 22324 33396
rect 20996 32360 21048 32366
rect 20996 32302 21048 32308
rect 21088 32360 21140 32366
rect 21088 32302 21140 32308
rect 20720 32292 20772 32298
rect 20720 32234 20772 32240
rect 20628 32224 20680 32230
rect 20628 32166 20680 32172
rect 20640 32026 20668 32166
rect 20628 32020 20680 32026
rect 20628 31962 20680 31968
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 20352 31476 20404 31482
rect 20352 31418 20404 31424
rect 20088 31198 20208 31226
rect 20180 31142 20208 31198
rect 20168 31136 20220 31142
rect 20168 31078 20220 31084
rect 20180 30054 20208 31078
rect 20548 30802 20576 31690
rect 21008 31414 21036 32302
rect 21100 31414 21128 32302
rect 21836 31822 21864 33390
rect 22204 33374 22324 33390
rect 21935 33212 22243 33221
rect 21935 33210 21941 33212
rect 21997 33210 22021 33212
rect 22077 33210 22101 33212
rect 22157 33210 22181 33212
rect 22237 33210 22243 33212
rect 21997 33158 21999 33210
rect 22179 33158 22181 33210
rect 21935 33156 21941 33158
rect 21997 33156 22021 33158
rect 22077 33156 22101 33158
rect 22157 33156 22181 33158
rect 22237 33156 22243 33158
rect 21935 33147 22243 33156
rect 22296 33114 22324 33374
rect 23032 33114 23060 33544
rect 23112 33526 23164 33532
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 23020 33108 23072 33114
rect 23020 33050 23072 33056
rect 21935 32124 22243 32133
rect 21935 32122 21941 32124
rect 21997 32122 22021 32124
rect 22077 32122 22101 32124
rect 22157 32122 22181 32124
rect 22237 32122 22243 32124
rect 21997 32070 21999 32122
rect 22179 32070 22181 32122
rect 21935 32068 21941 32070
rect 21997 32068 22021 32070
rect 22077 32068 22101 32070
rect 22157 32068 22181 32070
rect 22237 32068 22243 32070
rect 21935 32059 22243 32068
rect 21824 31816 21876 31822
rect 21824 31758 21876 31764
rect 20996 31408 21048 31414
rect 20996 31350 21048 31356
rect 21088 31408 21140 31414
rect 21140 31356 21220 31362
rect 21088 31350 21220 31356
rect 20536 30796 20588 30802
rect 20536 30738 20588 30744
rect 21008 30410 21036 31350
rect 21100 31334 21220 31350
rect 21088 31272 21140 31278
rect 21088 31214 21140 31220
rect 21100 30938 21128 31214
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 21192 30870 21220 31334
rect 21364 31204 21416 31210
rect 21364 31146 21416 31152
rect 21376 30938 21404 31146
rect 21364 30932 21416 30938
rect 21364 30874 21416 30880
rect 21180 30864 21232 30870
rect 21180 30806 21232 30812
rect 21008 30382 21128 30410
rect 21100 30190 21128 30382
rect 21192 30190 21220 30806
rect 21836 30802 21864 31758
rect 23032 31754 23060 33050
rect 23400 32978 23428 34002
rect 24136 33998 24164 34342
rect 24228 34066 24256 34954
rect 26132 34844 26440 34853
rect 26132 34842 26138 34844
rect 26194 34842 26218 34844
rect 26274 34842 26298 34844
rect 26354 34842 26378 34844
rect 26434 34842 26440 34844
rect 26194 34790 26196 34842
rect 26376 34790 26378 34842
rect 26132 34788 26138 34790
rect 26194 34788 26218 34790
rect 26274 34788 26298 34790
rect 26354 34788 26378 34790
rect 26434 34788 26440 34790
rect 26132 34779 26440 34788
rect 27080 34746 27108 34954
rect 32680 34944 32732 34950
rect 32680 34886 32732 34892
rect 24308 34740 24360 34746
rect 24308 34682 24360 34688
rect 27068 34740 27120 34746
rect 27068 34682 27120 34688
rect 24320 34610 24348 34682
rect 32692 34678 32720 34886
rect 34526 34844 34834 34853
rect 34526 34842 34532 34844
rect 34588 34842 34612 34844
rect 34668 34842 34692 34844
rect 34748 34842 34772 34844
rect 34828 34842 34834 34844
rect 34588 34790 34590 34842
rect 34770 34790 34772 34842
rect 34526 34788 34532 34790
rect 34588 34788 34612 34790
rect 34668 34788 34692 34790
rect 34748 34788 34772 34790
rect 34828 34788 34834 34790
rect 34526 34779 34834 34788
rect 32680 34672 32732 34678
rect 31022 34640 31078 34649
rect 24308 34604 24360 34610
rect 32680 34614 32732 34620
rect 31022 34575 31078 34584
rect 24308 34546 24360 34552
rect 30329 34300 30637 34309
rect 30329 34298 30335 34300
rect 30391 34298 30415 34300
rect 30471 34298 30495 34300
rect 30551 34298 30575 34300
rect 30631 34298 30637 34300
rect 30391 34246 30393 34298
rect 30573 34246 30575 34298
rect 30329 34244 30335 34246
rect 30391 34244 30415 34246
rect 30471 34244 30495 34246
rect 30551 34244 30575 34246
rect 30631 34244 30637 34246
rect 30329 34235 30637 34244
rect 24216 34060 24268 34066
rect 24216 34002 24268 34008
rect 24124 33992 24176 33998
rect 24124 33934 24176 33940
rect 23756 33856 23808 33862
rect 23756 33798 23808 33804
rect 23940 33856 23992 33862
rect 23940 33798 23992 33804
rect 23768 33658 23796 33798
rect 23756 33652 23808 33658
rect 23756 33594 23808 33600
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23584 32978 23612 33254
rect 23388 32972 23440 32978
rect 23388 32914 23440 32920
rect 23572 32972 23624 32978
rect 23572 32914 23624 32920
rect 23400 32858 23428 32914
rect 23308 32830 23428 32858
rect 22284 31748 22336 31754
rect 22284 31690 22336 31696
rect 23020 31748 23072 31754
rect 23020 31690 23072 31696
rect 22296 31482 22324 31690
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 23308 31362 23336 32830
rect 23848 32496 23900 32502
rect 23848 32438 23900 32444
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23400 31482 23428 31962
rect 23768 31686 23796 32370
rect 23756 31680 23808 31686
rect 23756 31622 23808 31628
rect 23860 31482 23888 32438
rect 23952 32230 23980 33798
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 24124 32224 24176 32230
rect 24124 32166 24176 32172
rect 24136 31890 24164 32166
rect 24124 31884 24176 31890
rect 24124 31826 24176 31832
rect 23388 31476 23440 31482
rect 23388 31418 23440 31424
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23308 31334 23428 31362
rect 23400 31278 23428 31334
rect 23388 31272 23440 31278
rect 23388 31214 23440 31220
rect 21935 31036 22243 31045
rect 21935 31034 21941 31036
rect 21997 31034 22021 31036
rect 22077 31034 22101 31036
rect 22157 31034 22181 31036
rect 22237 31034 22243 31036
rect 21997 30982 21999 31034
rect 22179 30982 22181 31034
rect 21935 30980 21941 30982
rect 21997 30980 22021 30982
rect 22077 30980 22101 30982
rect 22157 30980 22181 30982
rect 22237 30980 22243 30982
rect 21935 30971 22243 30980
rect 21824 30796 21876 30802
rect 21824 30738 21876 30744
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 21284 30258 21312 30602
rect 21376 30394 21404 30670
rect 21364 30388 21416 30394
rect 21364 30330 21416 30336
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 21088 30184 21140 30190
rect 21088 30126 21140 30132
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 20168 30048 20220 30054
rect 20088 29996 20168 30002
rect 20088 29990 20220 29996
rect 20088 29974 20208 29990
rect 19248 29708 19300 29714
rect 19248 29650 19300 29656
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 18880 28960 18932 28966
rect 18880 28902 18932 28908
rect 18892 28762 18920 28902
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 19352 28558 19380 29582
rect 19904 29306 19932 29650
rect 20088 29646 20116 29974
rect 21008 29850 21036 30126
rect 20996 29844 21048 29850
rect 20996 29786 21048 29792
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 19892 29300 19944 29306
rect 19892 29242 19944 29248
rect 19708 29232 19760 29238
rect 19708 29174 19760 29180
rect 19720 29102 19748 29174
rect 19524 29096 19576 29102
rect 19524 29038 19576 29044
rect 19616 29096 19668 29102
rect 19616 29038 19668 29044
rect 19708 29096 19760 29102
rect 19708 29038 19760 29044
rect 19536 28762 19564 29038
rect 19628 28762 19656 29038
rect 20088 29034 20116 29582
rect 20812 29572 20864 29578
rect 20812 29514 20864 29520
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20364 29102 20392 29446
rect 20444 29164 20496 29170
rect 20444 29106 20496 29112
rect 20352 29096 20404 29102
rect 20352 29038 20404 29044
rect 20076 29028 20128 29034
rect 20076 28970 20128 28976
rect 19524 28756 19576 28762
rect 19524 28698 19576 28704
rect 19616 28756 19668 28762
rect 19616 28698 19668 28704
rect 20456 28558 20484 29106
rect 20720 29096 20772 29102
rect 20720 29038 20772 29044
rect 20732 28762 20760 29038
rect 20720 28756 20772 28762
rect 20720 28698 20772 28704
rect 20824 28558 20852 29514
rect 20996 29164 21048 29170
rect 20996 29106 21048 29112
rect 21008 28762 21036 29106
rect 21100 29034 21128 30126
rect 21192 29510 21220 30126
rect 21376 29578 21404 30330
rect 21836 30190 21864 30738
rect 23112 30320 23164 30326
rect 23164 30268 23336 30274
rect 23112 30262 23336 30268
rect 23124 30246 23336 30262
rect 23124 30190 23152 30246
rect 21824 30184 21876 30190
rect 21824 30126 21876 30132
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 23112 30184 23164 30190
rect 23112 30126 23164 30132
rect 21364 29572 21416 29578
rect 21364 29514 21416 29520
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 21192 29170 21220 29446
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21088 29028 21140 29034
rect 21088 28970 21140 28976
rect 21836 28762 21864 30126
rect 21935 29948 22243 29957
rect 21935 29946 21941 29948
rect 21997 29946 22021 29948
rect 22077 29946 22101 29948
rect 22157 29946 22181 29948
rect 22237 29946 22243 29948
rect 21997 29894 21999 29946
rect 22179 29894 22181 29946
rect 21935 29892 21941 29894
rect 21997 29892 22021 29894
rect 22077 29892 22101 29894
rect 22157 29892 22181 29894
rect 22237 29892 22243 29894
rect 21935 29883 22243 29892
rect 22388 29850 22416 30126
rect 22376 29844 22428 29850
rect 22376 29786 22428 29792
rect 23112 29232 23164 29238
rect 23112 29174 23164 29180
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 21935 28860 22243 28869
rect 21935 28858 21941 28860
rect 21997 28858 22021 28860
rect 22077 28858 22101 28860
rect 22157 28858 22181 28860
rect 22237 28858 22243 28860
rect 21997 28806 21999 28858
rect 22179 28806 22181 28858
rect 21935 28804 21941 28806
rect 21997 28804 22021 28806
rect 22077 28804 22101 28806
rect 22157 28804 22181 28806
rect 22237 28804 22243 28806
rect 21935 28795 22243 28804
rect 20996 28756 21048 28762
rect 20996 28698 21048 28704
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 18788 28552 18840 28558
rect 18788 28494 18840 28500
rect 18880 28552 18932 28558
rect 18880 28494 18932 28500
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17512 27470 17540 28358
rect 17738 28316 18046 28325
rect 17738 28314 17744 28316
rect 17800 28314 17824 28316
rect 17880 28314 17904 28316
rect 17960 28314 17984 28316
rect 18040 28314 18046 28316
rect 17800 28262 17802 28314
rect 17982 28262 17984 28314
rect 17738 28260 17744 28262
rect 17800 28260 17824 28262
rect 17880 28260 17904 28262
rect 17960 28260 17984 28262
rect 18040 28260 18046 28262
rect 17738 28251 18046 28260
rect 18892 27470 18920 28494
rect 20076 28484 20128 28490
rect 20076 28426 20128 28432
rect 20088 28150 20116 28426
rect 21836 28218 21864 28698
rect 22296 28490 22324 28902
rect 23124 28762 23152 29174
rect 23112 28756 23164 28762
rect 23112 28698 23164 28704
rect 23308 28490 23336 30246
rect 23400 29730 23428 31214
rect 24228 30258 24256 34002
rect 26792 33992 26844 33998
rect 26792 33934 26844 33940
rect 26516 33924 26568 33930
rect 26516 33866 26568 33872
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 25056 33658 25084 33798
rect 26132 33756 26440 33765
rect 26132 33754 26138 33756
rect 26194 33754 26218 33756
rect 26274 33754 26298 33756
rect 26354 33754 26378 33756
rect 26434 33754 26440 33756
rect 26194 33702 26196 33754
rect 26376 33702 26378 33754
rect 26132 33700 26138 33702
rect 26194 33700 26218 33702
rect 26274 33700 26298 33702
rect 26354 33700 26378 33702
rect 26434 33700 26440 33702
rect 26132 33691 26440 33700
rect 26528 33658 26556 33866
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 26516 33652 26568 33658
rect 26516 33594 26568 33600
rect 24584 33108 24636 33114
rect 24584 33050 24636 33056
rect 24308 32972 24360 32978
rect 24308 32914 24360 32920
rect 24320 32502 24348 32914
rect 24400 32836 24452 32842
rect 24400 32778 24452 32784
rect 24308 32496 24360 32502
rect 24308 32438 24360 32444
rect 24412 32434 24440 32778
rect 24596 32434 24624 33050
rect 24780 32910 24808 33594
rect 25964 33448 26016 33454
rect 25964 33390 26016 33396
rect 25976 33114 26004 33390
rect 25964 33108 26016 33114
rect 25964 33050 26016 33056
rect 24768 32904 24820 32910
rect 24768 32846 24820 32852
rect 24952 32836 25004 32842
rect 24872 32796 24952 32824
rect 24400 32428 24452 32434
rect 24400 32370 24452 32376
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24412 32314 24440 32370
rect 24412 32286 24716 32314
rect 24688 30326 24716 32286
rect 24872 31686 24900 32796
rect 24952 32778 25004 32784
rect 25044 32836 25096 32842
rect 25044 32778 25096 32784
rect 25056 32570 25084 32778
rect 26132 32668 26440 32677
rect 26132 32666 26138 32668
rect 26194 32666 26218 32668
rect 26274 32666 26298 32668
rect 26354 32666 26378 32668
rect 26434 32666 26440 32668
rect 26194 32614 26196 32666
rect 26376 32614 26378 32666
rect 26132 32612 26138 32614
rect 26194 32612 26218 32614
rect 26274 32612 26298 32614
rect 26354 32612 26378 32614
rect 26434 32612 26440 32614
rect 26132 32603 26440 32612
rect 25044 32564 25096 32570
rect 25044 32506 25096 32512
rect 26804 32434 26832 33934
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 26976 32904 27028 32910
rect 26976 32846 27028 32852
rect 26988 32502 27016 32846
rect 27172 32502 27200 33798
rect 30329 33212 30637 33221
rect 30329 33210 30335 33212
rect 30391 33210 30415 33212
rect 30471 33210 30495 33212
rect 30551 33210 30575 33212
rect 30631 33210 30637 33212
rect 30391 33158 30393 33210
rect 30573 33158 30575 33210
rect 30329 33156 30335 33158
rect 30391 33156 30415 33158
rect 30471 33156 30495 33158
rect 30551 33156 30575 33158
rect 30631 33156 30637 33158
rect 30329 33147 30637 33156
rect 28356 32768 28408 32774
rect 28356 32710 28408 32716
rect 26976 32496 27028 32502
rect 26976 32438 27028 32444
rect 27160 32496 27212 32502
rect 27160 32438 27212 32444
rect 26516 32428 26568 32434
rect 26516 32370 26568 32376
rect 26792 32428 26844 32434
rect 26792 32370 26844 32376
rect 25136 32360 25188 32366
rect 25136 32302 25188 32308
rect 25688 32360 25740 32366
rect 25688 32302 25740 32308
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24780 30938 24808 31078
rect 24768 30932 24820 30938
rect 24768 30874 24820 30880
rect 24676 30320 24728 30326
rect 24676 30262 24728 30268
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23860 29850 23888 29990
rect 23848 29844 23900 29850
rect 23848 29786 23900 29792
rect 23400 29714 23612 29730
rect 23400 29708 23624 29714
rect 23400 29702 23572 29708
rect 23400 29102 23428 29702
rect 23572 29650 23624 29656
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24504 29170 24532 29582
rect 24688 29170 24716 30262
rect 24768 30252 24820 30258
rect 24768 30194 24820 30200
rect 24780 29170 24808 30194
rect 24872 29714 24900 31622
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24964 30394 24992 31282
rect 25148 30666 25176 32302
rect 25700 32026 25728 32302
rect 26528 32026 26556 32370
rect 25688 32020 25740 32026
rect 25688 31962 25740 31968
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 26132 31580 26440 31589
rect 26132 31578 26138 31580
rect 26194 31578 26218 31580
rect 26274 31578 26298 31580
rect 26354 31578 26378 31580
rect 26434 31578 26440 31580
rect 26194 31526 26196 31578
rect 26376 31526 26378 31578
rect 26132 31524 26138 31526
rect 26194 31524 26218 31526
rect 26274 31524 26298 31526
rect 26354 31524 26378 31526
rect 26434 31524 26440 31526
rect 26132 31515 26440 31524
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25136 30660 25188 30666
rect 25056 30620 25136 30648
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 25056 29646 25084 30620
rect 25136 30602 25188 30608
rect 25596 30592 25648 30598
rect 25596 30534 25648 30540
rect 25608 30394 25636 30534
rect 25596 30388 25648 30394
rect 25596 30330 25648 30336
rect 25884 30258 25912 31078
rect 26516 30660 26568 30666
rect 26516 30602 26568 30608
rect 26132 30492 26440 30501
rect 26132 30490 26138 30492
rect 26194 30490 26218 30492
rect 26274 30490 26298 30492
rect 26354 30490 26378 30492
rect 26434 30490 26440 30492
rect 26194 30438 26196 30490
rect 26376 30438 26378 30490
rect 26132 30436 26138 30438
rect 26194 30436 26218 30438
rect 26274 30436 26298 30438
rect 26354 30436 26378 30438
rect 26434 30436 26440 30438
rect 26132 30427 26440 30436
rect 26528 30394 26556 30602
rect 26516 30388 26568 30394
rect 26516 30330 26568 30336
rect 26056 30320 26108 30326
rect 26056 30262 26108 30268
rect 25872 30252 25924 30258
rect 25872 30194 25924 30200
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25884 29850 25912 29990
rect 25872 29844 25924 29850
rect 25872 29786 25924 29792
rect 26068 29714 26096 30262
rect 26240 30252 26292 30258
rect 26292 30212 26556 30240
rect 26240 30194 26292 30200
rect 26056 29708 26108 29714
rect 26056 29650 26108 29656
rect 25044 29640 25096 29646
rect 25044 29582 25096 29588
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 24492 29164 24544 29170
rect 24492 29106 24544 29112
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 22284 28484 22336 28490
rect 22284 28426 22336 28432
rect 23296 28484 23348 28490
rect 23296 28426 23348 28432
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 18972 27940 19024 27946
rect 18972 27882 19024 27888
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 18880 27464 18932 27470
rect 18880 27406 18932 27412
rect 17512 26586 17540 27406
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17604 27130 17632 27270
rect 17738 27228 18046 27237
rect 17738 27226 17744 27228
rect 17800 27226 17824 27228
rect 17880 27226 17904 27228
rect 17960 27226 17984 27228
rect 18040 27226 18046 27228
rect 17800 27174 17802 27226
rect 17982 27174 17984 27226
rect 17738 27172 17744 27174
rect 17800 27172 17824 27174
rect 17880 27172 17904 27174
rect 17960 27172 17984 27174
rect 18040 27172 18046 27174
rect 17738 27163 18046 27172
rect 18892 27130 18920 27406
rect 17592 27124 17644 27130
rect 17592 27066 17644 27072
rect 18880 27124 18932 27130
rect 18880 27066 18932 27072
rect 18984 27062 19012 27882
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 21935 27772 22243 27781
rect 21935 27770 21941 27772
rect 21997 27770 22021 27772
rect 22077 27770 22101 27772
rect 22157 27770 22181 27772
rect 22237 27770 22243 27772
rect 21997 27718 21999 27770
rect 22179 27718 22181 27770
rect 21935 27716 21941 27718
rect 21997 27716 22021 27718
rect 22077 27716 22101 27718
rect 22157 27716 22181 27718
rect 22237 27716 22243 27718
rect 21935 27707 22243 27716
rect 19064 27464 19116 27470
rect 19064 27406 19116 27412
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 19076 26926 19104 27406
rect 19248 27328 19300 27334
rect 19248 27270 19300 27276
rect 19260 27130 19288 27270
rect 19248 27124 19300 27130
rect 19248 27066 19300 27072
rect 19064 26920 19116 26926
rect 19064 26862 19116 26868
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 19076 26450 19104 26862
rect 19444 26586 19472 27406
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20824 27130 20852 27338
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 20076 27056 20128 27062
rect 20076 26998 20128 27004
rect 19432 26580 19484 26586
rect 19432 26522 19484 26528
rect 19064 26444 19116 26450
rect 19064 26386 19116 26392
rect 19984 26444 20036 26450
rect 19984 26386 20036 26392
rect 17738 26140 18046 26149
rect 17738 26138 17744 26140
rect 17800 26138 17824 26140
rect 17880 26138 17904 26140
rect 17960 26138 17984 26140
rect 18040 26138 18046 26140
rect 17800 26086 17802 26138
rect 17982 26086 17984 26138
rect 17738 26084 17744 26086
rect 17800 26084 17824 26086
rect 17880 26084 17904 26086
rect 17960 26084 17984 26086
rect 18040 26084 18046 26086
rect 17738 26075 18046 26084
rect 19996 25906 20024 26386
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 20088 25242 20116 26998
rect 22296 26994 22324 27814
rect 22388 27674 22416 28086
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 22940 27130 22968 27406
rect 23308 27402 23336 28426
rect 23400 28150 23428 29038
rect 23584 28558 23612 29106
rect 24504 28626 24532 29106
rect 24492 28620 24544 28626
rect 24492 28562 24544 28568
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23388 28144 23440 28150
rect 23388 28086 23440 28092
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23492 27538 23520 27950
rect 23584 27946 23612 28494
rect 23848 28484 23900 28490
rect 23848 28426 23900 28432
rect 23572 27940 23624 27946
rect 23572 27882 23624 27888
rect 23860 27674 23888 28426
rect 24308 28416 24360 28422
rect 24308 28358 24360 28364
rect 23848 27668 23900 27674
rect 23848 27610 23900 27616
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23296 27396 23348 27402
rect 23296 27338 23348 27344
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 23308 26790 23336 27338
rect 23492 27130 23520 27474
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23860 26926 23888 27610
rect 23848 26920 23900 26926
rect 23848 26862 23900 26868
rect 20904 26784 20956 26790
rect 20904 26726 20956 26732
rect 23296 26784 23348 26790
rect 23296 26726 23348 26732
rect 20916 26450 20944 26726
rect 21935 26684 22243 26693
rect 21935 26682 21941 26684
rect 21997 26682 22021 26684
rect 22077 26682 22101 26684
rect 22157 26682 22181 26684
rect 22237 26682 22243 26684
rect 21997 26630 21999 26682
rect 22179 26630 22181 26682
rect 21935 26628 21941 26630
rect 21997 26628 22021 26630
rect 22077 26628 22101 26630
rect 22157 26628 22181 26630
rect 22237 26628 22243 26630
rect 21935 26619 22243 26628
rect 20904 26444 20956 26450
rect 20904 26386 20956 26392
rect 20996 26376 21048 26382
rect 20996 26318 21048 26324
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20732 25498 20760 26250
rect 21008 26042 21036 26318
rect 23308 26314 23336 26726
rect 23296 26308 23348 26314
rect 23296 26250 23348 26256
rect 23572 26308 23624 26314
rect 23572 26250 23624 26256
rect 23112 26240 23164 26246
rect 23112 26182 23164 26188
rect 23124 26042 23152 26182
rect 20996 26036 21048 26042
rect 20996 25978 21048 25984
rect 23112 26036 23164 26042
rect 23112 25978 23164 25984
rect 23308 25974 23336 26250
rect 23296 25968 23348 25974
rect 23296 25910 23348 25916
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 19996 25226 20116 25242
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19984 25220 20128 25226
rect 20036 25214 20076 25220
rect 19984 25162 20036 25168
rect 20076 25162 20128 25168
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 19064 25152 19116 25158
rect 19064 25094 19116 25100
rect 17738 25052 18046 25061
rect 17738 25050 17744 25052
rect 17800 25050 17824 25052
rect 17880 25050 17904 25052
rect 17960 25050 17984 25052
rect 18040 25050 18046 25052
rect 17800 24998 17802 25050
rect 17982 24998 17984 25050
rect 17738 24996 17744 24998
rect 17800 24996 17824 24998
rect 17880 24996 17904 24998
rect 17960 24996 17984 24998
rect 18040 24996 18046 24998
rect 17738 24987 18046 24996
rect 18248 24954 18276 25094
rect 18236 24948 18288 24954
rect 18236 24890 18288 24896
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18432 24410 18460 24754
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 19076 24342 19104 25094
rect 19536 24954 19564 25162
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19352 24410 19380 24754
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 17328 22982 17356 24006
rect 17316 22976 17368 22982
rect 17316 22918 17368 22924
rect 17328 22710 17356 22918
rect 17512 22778 17540 24142
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 17738 23964 18046 23973
rect 17738 23962 17744 23964
rect 17800 23962 17824 23964
rect 17880 23962 17904 23964
rect 17960 23962 17984 23964
rect 18040 23962 18046 23964
rect 17800 23910 17802 23962
rect 17982 23910 17984 23962
rect 17738 23908 17744 23910
rect 17800 23908 17824 23910
rect 17880 23908 17904 23910
rect 17960 23908 17984 23910
rect 18040 23908 18046 23910
rect 17738 23899 18046 23908
rect 18800 23186 18828 24074
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23866 19472 24006
rect 19536 23866 19564 24142
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19248 23724 19300 23730
rect 19248 23666 19300 23672
rect 19260 23322 19288 23666
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18236 23044 18288 23050
rect 18236 22986 18288 22992
rect 17738 22876 18046 22885
rect 17738 22874 17744 22876
rect 17800 22874 17824 22876
rect 17880 22874 17904 22876
rect 17960 22874 17984 22876
rect 18040 22874 18046 22876
rect 17800 22822 17802 22874
rect 17982 22822 17984 22874
rect 17738 22820 17744 22822
rect 17800 22820 17824 22822
rect 17880 22820 17904 22822
rect 17960 22820 17984 22822
rect 18040 22820 18046 22822
rect 17738 22811 18046 22820
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17316 22704 17368 22710
rect 17316 22646 17368 22652
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 17236 22066 17448 22094
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 15844 20538 15896 20544
rect 16960 20556 17080 20584
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15764 18426 15792 18702
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15488 17678 15516 18090
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15212 16114 15240 16526
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 14832 15496 14884 15502
rect 14830 15464 14832 15473
rect 14884 15464 14886 15473
rect 14830 15399 14886 15408
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15120 14618 15148 14758
rect 15212 14618 15240 15642
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 15304 13938 15332 16594
rect 15488 16590 15516 16934
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 16114 15424 16390
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 14414 15424 15846
rect 15488 15026 15516 16526
rect 15580 16522 15608 18022
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15580 16114 15608 16458
rect 15672 16454 15700 16934
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15764 16130 15792 16730
rect 15856 16590 15884 18090
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16316 17678 16344 18022
rect 16960 17814 16988 20556
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17052 19786 17080 20402
rect 17236 20058 17264 20470
rect 17328 20466 17356 20742
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17144 19310 17172 19654
rect 17236 19514 17264 19994
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17328 19378 17356 19654
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 16040 16794 16068 17478
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15672 16102 15792 16130
rect 15672 15178 15700 16102
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15580 15150 15700 15178
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15580 14906 15608 15150
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15488 14878 15608 14906
rect 15488 14414 15516 14878
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14414 15608 14758
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15396 14006 15424 14350
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15488 13326 15516 14350
rect 15672 13530 15700 14962
rect 15764 14414 15792 15982
rect 15856 15706 15884 16526
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 16040 15026 16068 15438
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15764 13938 15792 14350
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13541 10364 13849 10373
rect 13541 10362 13547 10364
rect 13603 10362 13627 10364
rect 13683 10362 13707 10364
rect 13763 10362 13787 10364
rect 13843 10362 13849 10364
rect 13603 10310 13605 10362
rect 13785 10310 13787 10362
rect 13541 10308 13547 10310
rect 13603 10308 13627 10310
rect 13683 10308 13707 10310
rect 13763 10308 13787 10310
rect 13843 10308 13849 10310
rect 13541 10299 13849 10308
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9761 13584 9998
rect 14108 9926 14136 12650
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13556 9586 13584 9687
rect 13726 9616 13782 9625
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13544 9580 13596 9586
rect 13726 9551 13728 9560
rect 13544 9522 13596 9528
rect 13780 9551 13782 9560
rect 13728 9522 13780 9528
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 13541 9276 13849 9285
rect 13541 9274 13547 9276
rect 13603 9274 13627 9276
rect 13683 9274 13707 9276
rect 13763 9274 13787 9276
rect 13843 9274 13849 9276
rect 13603 9222 13605 9274
rect 13785 9222 13787 9274
rect 13541 9220 13547 9222
rect 13603 9220 13627 9222
rect 13683 9220 13707 9222
rect 13763 9220 13787 9222
rect 13843 9220 13849 9222
rect 13541 9211 13849 9220
rect 14476 9178 14504 9318
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 12308 8928 12572 8956
rect 12256 8910 12308 8916
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 9344 8732 9652 8741
rect 9344 8730 9350 8732
rect 9406 8730 9430 8732
rect 9486 8730 9510 8732
rect 9566 8730 9590 8732
rect 9646 8730 9652 8732
rect 9406 8678 9408 8730
rect 9588 8678 9590 8730
rect 9344 8676 9350 8678
rect 9406 8676 9430 8678
rect 9486 8676 9510 8678
rect 9566 8676 9590 8678
rect 9646 8676 9652 8678
rect 9344 8667 9652 8676
rect 5147 8188 5455 8197
rect 5147 8186 5153 8188
rect 5209 8186 5233 8188
rect 5289 8186 5313 8188
rect 5369 8186 5393 8188
rect 5449 8186 5455 8188
rect 5209 8134 5211 8186
rect 5391 8134 5393 8186
rect 5147 8132 5153 8134
rect 5209 8132 5233 8134
rect 5289 8132 5313 8134
rect 5369 8132 5393 8134
rect 5449 8132 5455 8134
rect 5147 8123 5455 8132
rect 13541 8188 13849 8197
rect 13541 8186 13547 8188
rect 13603 8186 13627 8188
rect 13683 8186 13707 8188
rect 13763 8186 13787 8188
rect 13843 8186 13849 8188
rect 13603 8134 13605 8186
rect 13785 8134 13787 8186
rect 13541 8132 13547 8134
rect 13603 8132 13627 8134
rect 13683 8132 13707 8134
rect 13763 8132 13787 8134
rect 13843 8132 13849 8134
rect 13541 8123 13849 8132
rect 13924 8090 13952 8774
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 9344 7644 9652 7653
rect 9344 7642 9350 7644
rect 9406 7642 9430 7644
rect 9486 7642 9510 7644
rect 9566 7642 9590 7644
rect 9646 7642 9652 7644
rect 9406 7590 9408 7642
rect 9588 7590 9590 7642
rect 9344 7588 9350 7590
rect 9406 7588 9430 7590
rect 9486 7588 9510 7590
rect 9566 7588 9590 7590
rect 9646 7588 9652 7590
rect 9344 7579 9652 7588
rect 12176 7342 12204 7890
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 12452 7546 12480 7754
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 13924 7478 13952 7754
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 14568 7410 14596 11154
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14660 8906 14688 9590
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 8974 14780 9454
rect 15028 9450 15056 12650
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11218 15240 11494
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15488 9654 15516 12582
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15198 9480 15254 9489
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15108 9444 15160 9450
rect 15198 9415 15254 9424
rect 15108 9386 15160 9392
rect 15120 8974 15148 9386
rect 15212 9382 15240 9415
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 15108 8968 15160 8974
rect 15488 8956 15516 9590
rect 15672 9382 15700 13262
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12782 15792 13126
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15856 9654 15884 14350
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15948 13326 15976 14214
rect 16040 13938 16068 14418
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 16040 13326 16068 13738
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15752 9512 15804 9518
rect 15844 9512 15896 9518
rect 15752 9454 15804 9460
rect 15842 9480 15844 9489
rect 15896 9480 15898 9489
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15568 8968 15620 8974
rect 15488 8928 15568 8956
rect 15108 8910 15160 8916
rect 15568 8910 15620 8916
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 5147 7100 5455 7109
rect 5147 7098 5153 7100
rect 5209 7098 5233 7100
rect 5289 7098 5313 7100
rect 5369 7098 5393 7100
rect 5449 7098 5455 7100
rect 5209 7046 5211 7098
rect 5391 7046 5393 7098
rect 5147 7044 5153 7046
rect 5209 7044 5233 7046
rect 5289 7044 5313 7046
rect 5369 7044 5393 7046
rect 5449 7044 5455 7046
rect 5147 7035 5455 7044
rect 7944 7002 7972 7278
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1688 6458 1716 6666
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 2700 6322 2728 6734
rect 3252 6390 3280 6734
rect 9344 6556 9652 6565
rect 9344 6554 9350 6556
rect 9406 6554 9430 6556
rect 9486 6554 9510 6556
rect 9566 6554 9590 6556
rect 9646 6554 9652 6556
rect 9406 6502 9408 6554
rect 9588 6502 9590 6554
rect 9344 6500 9350 6502
rect 9406 6500 9430 6502
rect 9486 6500 9510 6502
rect 9566 6500 9590 6502
rect 9646 6500 9652 6502
rect 9344 6491 9652 6500
rect 10704 6458 10732 7278
rect 13280 6458 13308 7278
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13372 6390 13400 7278
rect 13541 7100 13849 7109
rect 13541 7098 13547 7100
rect 13603 7098 13627 7100
rect 13683 7098 13707 7100
rect 13763 7098 13787 7100
rect 13843 7098 13849 7100
rect 13603 7046 13605 7098
rect 13785 7046 13787 7098
rect 13541 7044 13547 7046
rect 13603 7044 13627 7046
rect 13683 7044 13707 7046
rect 13763 7044 13787 7046
rect 13843 7044 13849 7046
rect 13541 7035 13849 7044
rect 14568 6458 14596 7346
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 952 6225 980 6258
rect 7472 6248 7524 6254
rect 938 6216 994 6225
rect 7472 6190 7524 6196
rect 938 6151 994 6160
rect 5147 6012 5455 6021
rect 5147 6010 5153 6012
rect 5209 6010 5233 6012
rect 5289 6010 5313 6012
rect 5369 6010 5393 6012
rect 5449 6010 5455 6012
rect 5209 5958 5211 6010
rect 5391 5958 5393 6010
rect 5147 5956 5153 5958
rect 5209 5956 5233 5958
rect 5289 5956 5313 5958
rect 5369 5956 5393 5958
rect 5449 5956 5455 5958
rect 5147 5947 5455 5956
rect 5147 4924 5455 4933
rect 5147 4922 5153 4924
rect 5209 4922 5233 4924
rect 5289 4922 5313 4924
rect 5369 4922 5393 4924
rect 5449 4922 5455 4924
rect 5209 4870 5211 4922
rect 5391 4870 5393 4922
rect 5147 4868 5153 4870
rect 5209 4868 5233 4870
rect 5289 4868 5313 4870
rect 5369 4868 5393 4870
rect 5449 4868 5455 4870
rect 5147 4859 5455 4868
rect 5147 3836 5455 3845
rect 5147 3834 5153 3836
rect 5209 3834 5233 3836
rect 5289 3834 5313 3836
rect 5369 3834 5393 3836
rect 5449 3834 5455 3836
rect 5209 3782 5211 3834
rect 5391 3782 5393 3834
rect 5147 3780 5153 3782
rect 5209 3780 5233 3782
rect 5289 3780 5313 3782
rect 5369 3780 5393 3782
rect 5449 3780 5455 3782
rect 5147 3771 5455 3780
rect 5147 2748 5455 2757
rect 5147 2746 5153 2748
rect 5209 2746 5233 2748
rect 5289 2746 5313 2748
rect 5369 2746 5393 2748
rect 5449 2746 5455 2748
rect 5209 2694 5211 2746
rect 5391 2694 5393 2746
rect 5147 2692 5153 2694
rect 5209 2692 5233 2694
rect 5289 2692 5313 2694
rect 5369 2692 5393 2694
rect 5449 2692 5455 2694
rect 5147 2683 5455 2692
rect 7484 2650 7512 6190
rect 9344 5468 9652 5477
rect 9344 5466 9350 5468
rect 9406 5466 9430 5468
rect 9486 5466 9510 5468
rect 9566 5466 9590 5468
rect 9646 5466 9652 5468
rect 9406 5414 9408 5466
rect 9588 5414 9590 5466
rect 9344 5412 9350 5414
rect 9406 5412 9430 5414
rect 9486 5412 9510 5414
rect 9566 5412 9590 5414
rect 9646 5412 9652 5414
rect 9344 5403 9652 5412
rect 9344 4380 9652 4389
rect 9344 4378 9350 4380
rect 9406 4378 9430 4380
rect 9486 4378 9510 4380
rect 9566 4378 9590 4380
rect 9646 4378 9652 4380
rect 9406 4326 9408 4378
rect 9588 4326 9590 4378
rect 9344 4324 9350 4326
rect 9406 4324 9430 4326
rect 9486 4324 9510 4326
rect 9566 4324 9590 4326
rect 9646 4324 9652 4326
rect 9344 4315 9652 4324
rect 9344 3292 9652 3301
rect 9344 3290 9350 3292
rect 9406 3290 9430 3292
rect 9486 3290 9510 3292
rect 9566 3290 9590 3292
rect 9646 3290 9652 3292
rect 9406 3238 9408 3290
rect 9588 3238 9590 3290
rect 9344 3236 9350 3238
rect 9406 3236 9430 3238
rect 9486 3236 9510 3238
rect 9566 3236 9590 3238
rect 9646 3236 9652 3238
rect 9344 3227 9652 3236
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 32 800 60 2382
rect 5920 1306 5948 2382
rect 11808 2310 11836 6326
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 12820 5234 12848 6190
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13280 5914 13308 6054
rect 13541 6012 13849 6021
rect 13541 6010 13547 6012
rect 13603 6010 13627 6012
rect 13683 6010 13707 6012
rect 13763 6010 13787 6012
rect 13843 6010 13849 6012
rect 13603 5958 13605 6010
rect 13785 5958 13787 6010
rect 13541 5956 13547 5958
rect 13603 5956 13627 5958
rect 13683 5956 13707 5958
rect 13763 5956 13787 5958
rect 13843 5956 13849 5958
rect 13541 5947 13849 5956
rect 14108 5914 14136 6190
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12820 4282 12848 5170
rect 14660 5166 14688 8842
rect 14752 5166 14780 8910
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14844 6322 14872 7414
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15212 6458 15240 6666
rect 15580 6662 15608 8910
rect 15672 8838 15700 9318
rect 15764 9178 15792 9454
rect 15842 9415 15898 9424
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15764 8634 15792 8910
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15764 7290 15792 8570
rect 15856 8090 15884 8842
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15844 7540 15896 7546
rect 15948 7528 15976 10950
rect 15896 7500 15976 7528
rect 15844 7482 15896 7488
rect 15764 7262 15976 7290
rect 15948 6798 15976 7262
rect 16040 7206 16068 13262
rect 16132 12986 16160 16526
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16224 12918 16252 16050
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16316 15026 16344 15574
rect 16408 15570 16436 17750
rect 16960 17678 16988 17750
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17420 17218 17448 22066
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17512 21622 17540 21898
rect 17738 21788 18046 21797
rect 17738 21786 17744 21788
rect 17800 21786 17824 21788
rect 17880 21786 17904 21788
rect 17960 21786 17984 21788
rect 18040 21786 18046 21788
rect 17800 21734 17802 21786
rect 17982 21734 17984 21786
rect 17738 21732 17744 21734
rect 17800 21732 17824 21734
rect 17880 21732 17904 21734
rect 17960 21732 17984 21734
rect 18040 21732 18046 21734
rect 17738 21723 18046 21732
rect 18156 21622 18184 22578
rect 18248 22574 18276 22986
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 18800 22094 18828 23122
rect 18880 23044 18932 23050
rect 18880 22986 18932 22992
rect 18892 22778 18920 22986
rect 19260 22778 19288 23258
rect 19720 22982 19748 24074
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 18972 22500 19024 22506
rect 18972 22442 19024 22448
rect 18524 22066 18828 22094
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18248 21622 18276 21966
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18236 21616 18288 21622
rect 18236 21558 18288 21564
rect 17880 21350 17908 21558
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17512 20602 17540 20878
rect 17880 20874 17908 21286
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 17972 20806 18000 21422
rect 18064 21146 18092 21422
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17604 20482 17632 20742
rect 17738 20700 18046 20709
rect 17738 20698 17744 20700
rect 17800 20698 17824 20700
rect 17880 20698 17904 20700
rect 17960 20698 17984 20700
rect 18040 20698 18046 20700
rect 17800 20646 17802 20698
rect 17982 20646 17984 20698
rect 17738 20644 17744 20646
rect 17800 20644 17824 20646
rect 17880 20644 17904 20646
rect 17960 20644 17984 20646
rect 18040 20644 18046 20646
rect 17738 20635 18046 20644
rect 18156 20602 18184 21558
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 17512 20454 17632 20482
rect 17868 20460 17920 20466
rect 17512 19718 17540 20454
rect 17868 20402 17920 20408
rect 17880 20262 17908 20402
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 18248 20058 18276 20878
rect 18524 20806 18552 22066
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18616 21622 18644 21830
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18524 19854 18552 20742
rect 18800 20534 18828 20810
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17512 18426 17540 19654
rect 17604 19514 17632 19722
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 17738 19612 18046 19621
rect 17738 19610 17744 19612
rect 17800 19610 17824 19612
rect 17880 19610 17904 19612
rect 17960 19610 17984 19612
rect 18040 19610 18046 19612
rect 17800 19558 17802 19610
rect 17982 19558 17984 19610
rect 17738 19556 17744 19558
rect 17800 19556 17824 19558
rect 17880 19556 17904 19558
rect 17960 19556 17984 19558
rect 18040 19556 18046 19558
rect 17738 19547 18046 19556
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17592 19236 17644 19242
rect 17592 19178 17644 19184
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17512 17338 17540 18362
rect 17604 18272 17632 19178
rect 18156 18834 18184 19654
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 17738 18524 18046 18533
rect 17738 18522 17744 18524
rect 17800 18522 17824 18524
rect 17880 18522 17904 18524
rect 17960 18522 17984 18524
rect 18040 18522 18046 18524
rect 17800 18470 17802 18522
rect 17982 18470 17984 18522
rect 17738 18468 17744 18470
rect 17800 18468 17824 18470
rect 17880 18468 17904 18470
rect 17960 18468 17984 18470
rect 18040 18468 18046 18470
rect 17738 18459 18046 18468
rect 18524 18358 18552 19790
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18708 18426 18736 18702
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18892 18426 18920 18566
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 17684 18284 17736 18290
rect 17604 18244 17684 18272
rect 17684 18226 17736 18232
rect 17696 17814 17724 18226
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 17684 17808 17736 17814
rect 17684 17750 17736 17756
rect 18064 17678 18092 18158
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17328 17190 17448 17218
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16408 14940 16436 15506
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 15094 16528 15302
rect 16488 15088 16540 15094
rect 16488 15030 16540 15036
rect 16580 14952 16632 14958
rect 16408 14912 16580 14940
rect 16580 14894 16632 14900
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16316 14414 16344 14826
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16684 14074 16712 15438
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16868 14618 16896 14962
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17144 14618 17172 14894
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16132 9042 16160 9318
rect 16224 9178 16252 9318
rect 16316 9178 16344 13806
rect 16868 12434 16896 14418
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16868 12406 16988 12434
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 11898 16528 12038
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16132 7342 16160 7822
rect 16224 7410 16252 7822
rect 16408 7818 16436 9114
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16500 8634 16528 8910
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16408 7546 16436 7754
rect 16684 7546 16712 8842
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 16132 6866 16160 7278
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14844 5234 14872 6258
rect 15948 5914 15976 6734
rect 16224 6730 16252 7346
rect 16408 7002 16436 7482
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16212 6724 16264 6730
rect 16212 6666 16264 6672
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 15764 5166 15792 5238
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 13188 4826 13216 5102
rect 13541 4924 13849 4933
rect 13541 4922 13547 4924
rect 13603 4922 13627 4924
rect 13683 4922 13707 4924
rect 13763 4922 13787 4924
rect 13843 4922 13849 4924
rect 13603 4870 13605 4922
rect 13785 4870 13787 4922
rect 13541 4868 13547 4870
rect 13603 4868 13627 4870
rect 13683 4868 13707 4870
rect 13763 4868 13787 4870
rect 13843 4868 13849 4870
rect 13541 4859 13849 4868
rect 16224 4826 16252 5102
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12820 4078 12848 4218
rect 13832 4078 13860 4558
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14384 4214 14412 4422
rect 14660 4282 14688 4558
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 16500 4078 16528 5170
rect 16776 4486 16804 11698
rect 16868 11694 16896 12174
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 12176 2650 12204 4014
rect 13541 3836 13849 3845
rect 13541 3834 13547 3836
rect 13603 3834 13627 3836
rect 13683 3834 13707 3836
rect 13763 3834 13787 3836
rect 13843 3834 13849 3836
rect 13603 3782 13605 3834
rect 13785 3782 13787 3834
rect 13541 3780 13547 3782
rect 13603 3780 13627 3782
rect 13683 3780 13707 3782
rect 13763 3780 13787 3782
rect 13843 3780 13849 3782
rect 13541 3771 13849 3780
rect 13541 2748 13849 2757
rect 13541 2746 13547 2748
rect 13603 2746 13627 2748
rect 13683 2746 13707 2748
rect 13763 2746 13787 2748
rect 13843 2746 13849 2748
rect 13603 2694 13605 2746
rect 13785 2694 13787 2746
rect 13541 2692 13547 2694
rect 13603 2692 13627 2694
rect 13683 2692 13707 2694
rect 13763 2692 13787 2694
rect 13843 2692 13849 2694
rect 13541 2683 13849 2692
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 15672 2514 15700 4014
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 16960 2446 16988 12406
rect 17144 12238 17172 12786
rect 17328 12434 17356 17190
rect 17512 12832 17540 17274
rect 17604 17270 17632 17546
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 17738 17436 18046 17445
rect 17738 17434 17744 17436
rect 17800 17434 17824 17436
rect 17880 17434 17904 17436
rect 17960 17434 17984 17436
rect 18040 17434 18046 17436
rect 17800 17382 17802 17434
rect 17982 17382 17984 17434
rect 17738 17380 17744 17382
rect 17800 17380 17824 17382
rect 17880 17380 17904 17382
rect 17960 17380 17984 17382
rect 18040 17380 18046 17382
rect 17738 17371 18046 17380
rect 18156 17338 18184 17478
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 17592 17264 17644 17270
rect 17592 17206 17644 17212
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 18156 16590 18184 16934
rect 18248 16590 18276 18158
rect 18524 18086 18552 18294
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18524 17202 18552 18022
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18708 17202 18736 17478
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18328 17128 18380 17134
rect 18380 17088 18460 17116
rect 18328 17070 18380 17076
rect 18432 16998 18460 17088
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 17738 16348 18046 16357
rect 17738 16346 17744 16348
rect 17800 16346 17824 16348
rect 17880 16346 17904 16348
rect 17960 16346 17984 16348
rect 18040 16346 18046 16348
rect 17800 16294 17802 16346
rect 17982 16294 17984 16346
rect 17738 16292 17744 16294
rect 17800 16292 17824 16294
rect 17880 16292 17904 16294
rect 17960 16292 17984 16294
rect 18040 16292 18046 16294
rect 17738 16283 18046 16292
rect 18248 16046 18276 16526
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 16250 18460 16390
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17738 15260 18046 15269
rect 17738 15258 17744 15260
rect 17800 15258 17824 15260
rect 17880 15258 17904 15260
rect 17960 15258 17984 15260
rect 18040 15258 18046 15260
rect 17800 15206 17802 15258
rect 17982 15206 17984 15258
rect 17738 15204 17744 15206
rect 17800 15204 17824 15206
rect 17880 15204 17904 15206
rect 17960 15204 17984 15206
rect 18040 15204 18046 15206
rect 17738 15195 18046 15204
rect 18156 15026 18184 15302
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17604 14346 17632 14826
rect 18156 14414 18184 14962
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17738 14172 18046 14181
rect 17738 14170 17744 14172
rect 17800 14170 17824 14172
rect 17880 14170 17904 14172
rect 17960 14170 17984 14172
rect 18040 14170 18046 14172
rect 17800 14118 17802 14170
rect 17982 14118 17984 14170
rect 17738 14116 17744 14118
rect 17800 14116 17824 14118
rect 17880 14116 17904 14118
rect 17960 14116 17984 14118
rect 18040 14116 18046 14118
rect 17738 14107 18046 14116
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 17738 13084 18046 13093
rect 17738 13082 17744 13084
rect 17800 13082 17824 13084
rect 17880 13082 17904 13084
rect 17960 13082 17984 13084
rect 18040 13082 18046 13084
rect 17800 13030 17802 13082
rect 17982 13030 17984 13082
rect 17738 13028 17744 13030
rect 17800 13028 17824 13030
rect 17880 13028 17904 13030
rect 17960 13028 17984 13030
rect 18040 13028 18046 13030
rect 17738 13019 18046 13028
rect 17236 12406 17356 12434
rect 17420 12804 17540 12832
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 17052 11898 17080 12106
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17236 11762 17264 12406
rect 17420 12102 17448 12804
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17512 12306 17540 12582
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17604 12102 17632 12378
rect 18156 12306 18184 13942
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 17408 12096 17460 12102
rect 17592 12096 17644 12102
rect 17460 12056 17540 12084
rect 17408 12038 17460 12044
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 17052 11286 17080 11630
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 17420 10674 17448 11766
rect 17512 10810 17540 12056
rect 17592 12038 17644 12044
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 17604 11286 17632 12038
rect 17738 11996 18046 12005
rect 17738 11994 17744 11996
rect 17800 11994 17824 11996
rect 17880 11994 17904 11996
rect 17960 11994 17984 11996
rect 18040 11994 18046 11996
rect 17800 11942 17802 11994
rect 17982 11942 17984 11994
rect 17738 11940 17744 11942
rect 17800 11940 17824 11942
rect 17880 11940 17904 11942
rect 17960 11940 17984 11942
rect 18040 11940 18046 11942
rect 17738 11931 18046 11940
rect 18156 11898 18184 12038
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18248 11830 18276 15982
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18340 14618 18368 14962
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18432 14362 18460 14826
rect 18340 14334 18460 14362
rect 18340 13938 18368 14334
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 13938 18460 14214
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18340 12170 18368 12786
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18432 11898 18460 12378
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18432 11558 18460 11834
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 17972 11354 18000 11494
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18524 11286 18552 17138
rect 18708 12442 18736 17138
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18800 12238 18828 17206
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18616 11694 18644 12038
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 17592 11280 17644 11286
rect 17592 11222 17644 11228
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17420 10266 17448 10610
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17236 8090 17264 9658
rect 17328 9654 17356 9862
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17328 8634 17356 9590
rect 17420 9518 17448 9930
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17420 9178 17448 9454
rect 17512 9382 17540 10746
rect 17604 10674 17632 11222
rect 17738 10908 18046 10917
rect 17738 10906 17744 10908
rect 17800 10906 17824 10908
rect 17880 10906 17904 10908
rect 17960 10906 17984 10908
rect 18040 10906 18046 10908
rect 17800 10854 17802 10906
rect 17982 10854 17984 10906
rect 17738 10852 17744 10854
rect 17800 10852 17824 10854
rect 17880 10852 17904 10854
rect 17960 10852 17984 10854
rect 18040 10852 18046 10854
rect 17738 10843 18046 10852
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17604 9722 17632 10610
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 17880 10266 17908 10542
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 17738 9820 18046 9829
rect 17738 9818 17744 9820
rect 17800 9818 17824 9820
rect 17880 9818 17904 9820
rect 17960 9818 17984 9820
rect 18040 9818 18046 9820
rect 17800 9766 17802 9818
rect 17982 9766 17984 9818
rect 17738 9764 17744 9766
rect 17800 9764 17824 9766
rect 17880 9764 17904 9766
rect 17960 9764 17984 9766
rect 18040 9764 18046 9766
rect 17738 9755 18046 9764
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 18156 9654 18184 10202
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18156 9466 18184 9590
rect 18432 9586 18460 10542
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18064 9438 18184 9466
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17328 7954 17356 8570
rect 17408 8016 17460 8022
rect 17408 7958 17460 7964
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17420 7546 17448 7958
rect 17512 7886 17540 9318
rect 18064 8906 18092 9438
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 9178 18184 9318
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17604 8634 17632 8774
rect 17738 8732 18046 8741
rect 17738 8730 17744 8732
rect 17800 8730 17824 8732
rect 17880 8730 17904 8732
rect 17960 8730 17984 8732
rect 18040 8730 18046 8732
rect 17800 8678 17802 8730
rect 17982 8678 17984 8730
rect 17738 8676 17744 8678
rect 17800 8676 17824 8678
rect 17880 8676 17904 8678
rect 17960 8676 17984 8678
rect 18040 8676 18046 8678
rect 17738 8667 18046 8676
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 18156 8514 18184 8774
rect 18064 8486 18184 8514
rect 18236 8492 18288 8498
rect 18064 8430 18092 8486
rect 18236 8434 18288 8440
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17500 7744 17552 7750
rect 17604 7732 17632 8026
rect 18064 7818 18092 8366
rect 18248 8022 18276 8434
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 18052 7812 18104 7818
rect 18052 7754 18104 7760
rect 17552 7704 17632 7732
rect 17500 7686 17552 7692
rect 17738 7644 18046 7653
rect 17738 7642 17744 7644
rect 17800 7642 17824 7644
rect 17880 7642 17904 7644
rect 17960 7642 17984 7644
rect 18040 7642 18046 7644
rect 17800 7590 17802 7642
rect 17982 7590 17984 7642
rect 17738 7588 17744 7590
rect 17800 7588 17824 7590
rect 17880 7588 17904 7590
rect 17960 7588 17984 7590
rect 18040 7588 18046 7590
rect 17738 7579 18046 7588
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 18432 7410 18460 9522
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18708 9178 18736 9454
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18984 8566 19012 22442
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19720 21554 19748 21830
rect 19904 21690 19932 23054
rect 20088 22982 20116 25162
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 24206 20208 24754
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19260 20874 19288 21422
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19514 19380 19654
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19628 18970 19656 19858
rect 19720 19854 19748 21490
rect 20180 20942 20208 24142
rect 20732 23866 20760 25434
rect 21008 24750 21036 25842
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 22928 25832 22980 25838
rect 22928 25774 22980 25780
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 21284 24410 21312 24754
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21560 24410 21588 24550
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21548 24404 21600 24410
rect 21548 24346 21600 24352
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20640 23050 20668 23122
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20640 21894 20668 22986
rect 20732 22642 20760 23802
rect 21652 23322 21680 25774
rect 21935 25596 22243 25605
rect 21935 25594 21941 25596
rect 21997 25594 22021 25596
rect 22077 25594 22101 25596
rect 22157 25594 22181 25596
rect 22237 25594 22243 25596
rect 21997 25542 21999 25594
rect 22179 25542 22181 25594
rect 21935 25540 21941 25542
rect 21997 25540 22021 25542
rect 22077 25540 22101 25542
rect 22157 25540 22181 25542
rect 22237 25540 22243 25542
rect 21935 25531 22243 25540
rect 21935 24508 22243 24517
rect 21935 24506 21941 24508
rect 21997 24506 22021 24508
rect 22077 24506 22101 24508
rect 22157 24506 22181 24508
rect 22237 24506 22243 24508
rect 21997 24454 21999 24506
rect 22179 24454 22181 24506
rect 21935 24452 21941 24454
rect 21997 24452 22021 24454
rect 22077 24452 22101 24454
rect 22157 24452 22181 24454
rect 22237 24452 22243 24454
rect 21935 24443 22243 24452
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 21935 23420 22243 23429
rect 21935 23418 21941 23420
rect 21997 23418 22021 23420
rect 22077 23418 22101 23420
rect 22157 23418 22181 23420
rect 22237 23418 22243 23420
rect 21997 23366 21999 23418
rect 22179 23366 22181 23418
rect 21935 23364 21941 23366
rect 21997 23364 22021 23366
rect 22077 23364 22101 23366
rect 22157 23364 22181 23366
rect 22237 23364 22243 23366
rect 21935 23355 22243 23364
rect 22296 23322 22324 23666
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 22284 23316 22336 23322
rect 22284 23258 22336 23264
rect 21652 22710 21680 23258
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20732 21554 20760 22578
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20812 21412 20864 21418
rect 20812 21354 20864 21360
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20640 21146 20668 21286
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20732 21026 20760 21286
rect 20824 21146 20852 21354
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20916 21146 20944 21286
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 21008 21026 21036 22578
rect 21180 22500 21232 22506
rect 21180 22442 21232 22448
rect 21192 21622 21220 22442
rect 21652 21622 21680 22646
rect 21935 22332 22243 22341
rect 21935 22330 21941 22332
rect 21997 22330 22021 22332
rect 22077 22330 22101 22332
rect 22157 22330 22181 22332
rect 22237 22330 22243 22332
rect 21997 22278 21999 22330
rect 22179 22278 22181 22330
rect 21935 22276 21941 22278
rect 21997 22276 22021 22278
rect 22077 22276 22101 22278
rect 22157 22276 22181 22278
rect 22237 22276 22243 22278
rect 21935 22267 22243 22276
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21652 21434 21680 21558
rect 21652 21406 21772 21434
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 20732 20998 21036 21026
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 20272 18902 20300 19314
rect 20364 19310 20392 20742
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20260 18896 20312 18902
rect 20260 18838 20312 18844
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 19524 18352 19576 18358
rect 19628 18306 19656 18634
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 19576 18300 19656 18306
rect 19524 18294 19656 18300
rect 19536 18278 19656 18294
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19352 17134 19380 17818
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19628 16114 19656 18278
rect 20260 18148 20312 18154
rect 20260 18090 20312 18096
rect 19892 17808 19944 17814
rect 19892 17750 19944 17756
rect 19904 16658 19932 17750
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19892 16652 19944 16658
rect 19720 16612 19892 16640
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19260 15162 19288 15370
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19156 14884 19208 14890
rect 19156 14826 19208 14832
rect 19168 14346 19196 14826
rect 19352 14618 19380 14894
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19444 14414 19472 15506
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19536 15094 19564 15302
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19168 13938 19196 14282
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19444 13870 19472 14350
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19628 11762 19656 16050
rect 19720 15026 19748 16612
rect 19892 16594 19944 16600
rect 19996 16250 20024 17070
rect 20180 16726 20208 17614
rect 20272 17610 20300 18090
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 20180 15502 20208 16662
rect 20456 16590 20484 18566
rect 20640 17882 20668 19314
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20272 15910 20300 16526
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 19984 15496 20036 15502
rect 19982 15464 19984 15473
rect 20168 15496 20220 15502
rect 20036 15464 20038 15473
rect 20168 15438 20220 15444
rect 19982 15399 20038 15408
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19720 14414 19748 14962
rect 19996 14618 20024 15302
rect 20180 15162 20208 15438
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 19720 12170 19748 12310
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19720 11898 19748 12106
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19076 9518 19104 10202
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19904 9450 19932 14214
rect 20088 11762 20116 14826
rect 20272 14346 20300 15846
rect 20456 15434 20484 16526
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20444 15428 20496 15434
rect 20444 15370 20496 15376
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20364 15162 20392 15302
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20364 13938 20392 14350
rect 20548 14278 20576 14962
rect 20640 14482 20668 15438
rect 20732 14890 20760 20998
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21560 20602 21588 20878
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21652 20534 21680 21286
rect 21744 21146 21772 21406
rect 21935 21244 22243 21253
rect 21935 21242 21941 21244
rect 21997 21242 22021 21244
rect 22077 21242 22101 21244
rect 22157 21242 22181 21244
rect 22237 21242 22243 21244
rect 21997 21190 21999 21242
rect 22179 21190 22181 21242
rect 21935 21188 21941 21190
rect 21997 21188 22021 21190
rect 22077 21188 22101 21190
rect 22157 21188 22181 21190
rect 22237 21188 22243 21190
rect 21935 21179 22243 21188
rect 22480 21146 22508 24074
rect 22940 23186 22968 25774
rect 23124 24614 23152 25842
rect 23308 24750 23336 25910
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23124 24274 23152 24550
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 23124 23882 23152 24210
rect 23032 23866 23152 23882
rect 23308 23866 23336 24686
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23400 24070 23428 24550
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23020 23860 23152 23866
rect 23072 23854 23152 23860
rect 23296 23860 23348 23866
rect 23020 23802 23072 23808
rect 23296 23802 23348 23808
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 22664 21554 22692 23054
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 22940 21690 22968 22918
rect 23032 22030 23060 23802
rect 23308 23186 23336 23802
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23124 22098 23152 23122
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 22928 21684 22980 21690
rect 22928 21626 22980 21632
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21640 20528 21692 20534
rect 21546 20496 21602 20505
rect 21640 20470 21692 20476
rect 21546 20431 21602 20440
rect 21732 20460 21784 20466
rect 21560 20330 21588 20431
rect 21732 20402 21784 20408
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21192 19990 21220 20198
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20916 17678 20944 19246
rect 21744 18358 21772 20402
rect 21836 18902 21864 20878
rect 22376 20868 22428 20874
rect 22376 20810 22428 20816
rect 22388 20262 22416 20810
rect 22664 20806 22692 21490
rect 22940 20942 22968 21626
rect 23032 21486 23060 21966
rect 23020 21480 23072 21486
rect 23020 21422 23072 21428
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 21935 20156 22243 20165
rect 21935 20154 21941 20156
rect 21997 20154 22021 20156
rect 22077 20154 22101 20156
rect 22157 20154 22181 20156
rect 22237 20154 22243 20156
rect 21997 20102 21999 20154
rect 22179 20102 22181 20154
rect 21935 20100 21941 20102
rect 21997 20100 22021 20102
rect 22077 20100 22101 20102
rect 22157 20100 22181 20102
rect 22237 20100 22243 20102
rect 21935 20091 22243 20100
rect 22480 20058 22508 20402
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 21935 19068 22243 19077
rect 21935 19066 21941 19068
rect 21997 19066 22021 19068
rect 22077 19066 22101 19068
rect 22157 19066 22181 19068
rect 22237 19066 22243 19068
rect 21997 19014 21999 19066
rect 22179 19014 22181 19066
rect 21935 19012 21941 19014
rect 21997 19012 22021 19014
rect 22077 19012 22101 19014
rect 22157 19012 22181 19014
rect 22237 19012 22243 19014
rect 21935 19003 22243 19012
rect 21824 18896 21876 18902
rect 22296 18850 22324 19654
rect 22572 19446 22600 19790
rect 22560 19440 22612 19446
rect 22560 19382 22612 19388
rect 21824 18838 21876 18844
rect 22204 18822 22324 18850
rect 22468 18896 22520 18902
rect 22468 18838 22520 18844
rect 22204 18766 22232 18822
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22284 18692 22336 18698
rect 22284 18634 22336 18640
rect 21732 18352 21784 18358
rect 21732 18294 21784 18300
rect 22296 18154 22324 18634
rect 22480 18442 22508 18838
rect 22572 18766 22600 19382
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22480 18414 22600 18442
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 21935 17980 22243 17989
rect 21935 17978 21941 17980
rect 21997 17978 22021 17980
rect 22077 17978 22101 17980
rect 22157 17978 22181 17980
rect 22237 17978 22243 17980
rect 21997 17926 21999 17978
rect 22179 17926 22181 17978
rect 21935 17924 21941 17926
rect 21997 17924 22021 17926
rect 22077 17924 22101 17926
rect 22157 17924 22181 17926
rect 22237 17924 22243 17926
rect 21935 17915 22243 17924
rect 22296 17882 22324 18090
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 20916 15706 20944 17614
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21008 17202 21036 17478
rect 21652 17202 21680 17614
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21192 16794 21220 16934
rect 21935 16892 22243 16901
rect 21935 16890 21941 16892
rect 21997 16890 22021 16892
rect 22077 16890 22101 16892
rect 22157 16890 22181 16892
rect 22237 16890 22243 16892
rect 21997 16838 21999 16890
rect 22179 16838 22181 16890
rect 21935 16836 21941 16838
rect 21997 16836 22021 16838
rect 22077 16836 22101 16838
rect 22157 16836 22181 16838
rect 22237 16836 22243 16838
rect 21935 16827 22243 16836
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21652 15706 21680 16526
rect 22296 16250 22324 17070
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 21935 15804 22243 15813
rect 21935 15802 21941 15804
rect 21997 15802 22021 15804
rect 22077 15802 22101 15804
rect 22157 15802 22181 15804
rect 22237 15802 22243 15804
rect 21997 15750 21999 15802
rect 22179 15750 22181 15802
rect 21935 15748 21941 15750
rect 21997 15748 22021 15750
rect 22077 15748 22101 15750
rect 22157 15748 22181 15750
rect 22237 15748 22243 15750
rect 21935 15739 22243 15748
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20824 14278 20852 14962
rect 20916 14498 20944 15642
rect 22296 15570 22324 15982
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 21008 15026 21036 15370
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 21100 14618 21128 14962
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21180 14544 21232 14550
rect 20916 14492 21180 14498
rect 20916 14486 21232 14492
rect 20916 14470 21220 14486
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20548 13938 20576 14214
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20364 13462 20392 13874
rect 20548 13530 20576 13874
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20352 13456 20404 13462
rect 20352 13398 20404 13404
rect 20548 13258 20576 13466
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20364 12986 20392 13126
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20364 12434 20392 12922
rect 20272 12406 20392 12434
rect 20444 12436 20496 12442
rect 20272 12238 20300 12406
rect 20444 12378 20496 12384
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11762 20208 12038
rect 20456 11762 20484 12378
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 19996 10674 20024 11698
rect 20088 11082 20116 11698
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 20180 10810 20208 11562
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19996 9926 20024 10610
rect 20180 9994 20208 10746
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19996 9586 20024 9862
rect 20166 9616 20222 9625
rect 19984 9580 20036 9586
rect 20166 9551 20222 9560
rect 19984 9522 20036 9528
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 18984 7886 19012 8502
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 7002 17448 7142
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17738 6556 18046 6565
rect 17738 6554 17744 6556
rect 17800 6554 17824 6556
rect 17880 6554 17904 6556
rect 17960 6554 17984 6556
rect 18040 6554 18046 6556
rect 17800 6502 17802 6554
rect 17982 6502 17984 6554
rect 17738 6500 17744 6502
rect 17800 6500 17824 6502
rect 17880 6500 17904 6502
rect 17960 6500 17984 6502
rect 18040 6500 18046 6502
rect 17738 6491 18046 6500
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 17144 5302 17172 5578
rect 17738 5468 18046 5477
rect 17738 5466 17744 5468
rect 17800 5466 17824 5468
rect 17880 5466 17904 5468
rect 17960 5466 17984 5468
rect 18040 5466 18046 5468
rect 17800 5414 17802 5466
rect 17982 5414 17984 5466
rect 17738 5412 17744 5414
rect 17800 5412 17824 5414
rect 17880 5412 17904 5414
rect 17960 5412 17984 5414
rect 18040 5412 18046 5414
rect 17738 5403 18046 5412
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17144 4214 17172 5238
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 17738 4380 18046 4389
rect 17738 4378 17744 4380
rect 17800 4378 17824 4380
rect 17880 4378 17904 4380
rect 17960 4378 17984 4380
rect 18040 4378 18046 4380
rect 17800 4326 17802 4378
rect 17982 4326 17984 4378
rect 17738 4324 17744 4326
rect 17800 4324 17824 4326
rect 17880 4324 17904 4326
rect 17960 4324 17984 4326
rect 18040 4324 18046 4326
rect 17738 4315 18046 4324
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17144 3534 17172 4150
rect 18156 3738 18184 4558
rect 18248 4078 18276 7346
rect 18432 7002 18460 7346
rect 18800 7002 18828 7754
rect 18984 7562 19012 7822
rect 18984 7546 19104 7562
rect 18972 7540 19104 7546
rect 19024 7534 19104 7540
rect 18972 7482 19024 7488
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18984 6390 19012 7346
rect 19076 6390 19104 7534
rect 19260 7478 19288 8230
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19708 8016 19760 8022
rect 19708 7958 19760 7964
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19168 6458 19196 6666
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 18972 6384 19024 6390
rect 18972 6326 19024 6332
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19260 5778 19288 7278
rect 19628 7274 19656 7890
rect 19720 7546 19748 7958
rect 19904 7750 19932 8026
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19616 7268 19668 7274
rect 19616 7210 19668 7216
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19536 6798 19564 7142
rect 19812 6934 19840 7686
rect 19800 6928 19852 6934
rect 19800 6870 19852 6876
rect 19904 6798 19932 7686
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19996 6730 20024 9522
rect 20180 9518 20208 9551
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20732 9466 20760 14010
rect 20824 13938 20852 14214
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 21468 13802 21496 14350
rect 21456 13796 21508 13802
rect 21456 13738 21508 13744
rect 21468 13326 21496 13738
rect 21560 13394 21588 14894
rect 21652 14346 21680 15438
rect 21744 15162 21772 15438
rect 22008 15428 22060 15434
rect 22284 15428 22336 15434
rect 22060 15388 22284 15416
rect 22008 15370 22060 15376
rect 22284 15370 22336 15376
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21935 14716 22243 14725
rect 21935 14714 21941 14716
rect 21997 14714 22021 14716
rect 22077 14714 22101 14716
rect 22157 14714 22181 14716
rect 22237 14714 22243 14716
rect 21997 14662 21999 14714
rect 22179 14662 22181 14714
rect 21935 14660 21941 14662
rect 21997 14660 22021 14662
rect 22077 14660 22101 14662
rect 22157 14660 22181 14662
rect 22237 14660 22243 14662
rect 21935 14651 22243 14660
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12764 21128 13126
rect 21100 12736 21312 12764
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20916 11354 20944 11630
rect 21008 11354 21036 12038
rect 21100 11898 21128 12038
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20548 8906 20576 9454
rect 20732 9438 21036 9466
rect 21008 9382 21036 9438
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20640 8974 20668 9318
rect 20916 9178 20944 9318
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20536 8900 20588 8906
rect 20536 8842 20588 8848
rect 21008 8498 21036 9318
rect 21192 9178 21220 9522
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21284 8974 21312 12736
rect 21560 12442 21588 13330
rect 21652 13326 21680 13398
rect 21744 13326 21772 13806
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21560 11898 21588 12174
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21468 11354 21496 11494
rect 21560 11354 21588 11698
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21652 9654 21680 11630
rect 21744 9654 21772 11766
rect 21836 9692 21864 14418
rect 21935 13628 22243 13637
rect 21935 13626 21941 13628
rect 21997 13626 22021 13628
rect 22077 13626 22101 13628
rect 22157 13626 22181 13628
rect 22237 13626 22243 13628
rect 21997 13574 21999 13626
rect 22179 13574 22181 13626
rect 21935 13572 21941 13574
rect 21997 13572 22021 13574
rect 22077 13572 22101 13574
rect 22157 13572 22181 13574
rect 22237 13572 22243 13574
rect 21935 13563 22243 13572
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 21928 12986 21956 13194
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 22296 12918 22324 13126
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 21935 12540 22243 12549
rect 21935 12538 21941 12540
rect 21997 12538 22021 12540
rect 22077 12538 22101 12540
rect 22157 12538 22181 12540
rect 22237 12538 22243 12540
rect 21997 12486 21999 12538
rect 22179 12486 22181 12538
rect 21935 12484 21941 12486
rect 21997 12484 22021 12486
rect 22077 12484 22101 12486
rect 22157 12484 22181 12486
rect 22237 12484 22243 12486
rect 21935 12475 22243 12484
rect 22296 12238 22324 12582
rect 22388 12442 22416 18226
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22388 11898 22416 12106
rect 22480 11898 22508 18226
rect 22572 17882 22600 18414
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22572 15450 22600 17478
rect 22664 15978 22692 20742
rect 22756 20482 22784 20878
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22756 20454 22876 20482
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22756 18766 22784 19790
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22848 18612 22876 20454
rect 22940 20262 22968 20742
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 23032 19922 23060 21422
rect 23124 21162 23152 22034
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23216 21350 23244 21830
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 23124 21134 23244 21162
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 23124 20534 23152 21014
rect 23112 20528 23164 20534
rect 23112 20470 23164 20476
rect 23216 19922 23244 21134
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23308 19854 23336 21830
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23492 19394 23520 25162
rect 23584 22438 23612 26250
rect 23664 25968 23716 25974
rect 23664 25910 23716 25916
rect 23676 24954 23704 25910
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 24124 23588 24176 23594
rect 24124 23530 24176 23536
rect 24136 23118 24164 23530
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 23572 22432 23624 22438
rect 23572 22374 23624 22380
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23676 22030 23704 22374
rect 24320 22234 24348 28358
rect 24504 27690 24532 28562
rect 24688 28558 24716 29106
rect 25056 28994 25084 29582
rect 26528 29578 26556 30212
rect 26804 29714 26832 32370
rect 27172 32230 27200 32438
rect 26976 32224 27028 32230
rect 26976 32166 27028 32172
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 27988 32224 28040 32230
rect 27988 32166 28040 32172
rect 26988 31890 27016 32166
rect 26976 31884 27028 31890
rect 26976 31826 27028 31832
rect 27160 31884 27212 31890
rect 27160 31826 27212 31832
rect 27172 31754 27200 31826
rect 27172 31726 27384 31754
rect 26976 31680 27028 31686
rect 26976 31622 27028 31628
rect 26988 31482 27016 31622
rect 26976 31476 27028 31482
rect 26976 31418 27028 31424
rect 27356 29850 27384 31726
rect 27804 31748 27856 31754
rect 27804 31690 27856 31696
rect 27620 31272 27672 31278
rect 27620 31214 27672 31220
rect 27632 30938 27660 31214
rect 27620 30932 27672 30938
rect 27620 30874 27672 30880
rect 27816 30598 27844 31690
rect 28000 30666 28028 32166
rect 28080 32020 28132 32026
rect 28080 31962 28132 31968
rect 28092 31822 28120 31962
rect 28368 31822 28396 32710
rect 28540 32496 28592 32502
rect 28540 32438 28592 32444
rect 28816 32496 28868 32502
rect 28816 32438 28868 32444
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 28092 30682 28120 31758
rect 28448 31748 28500 31754
rect 28448 31690 28500 31696
rect 28356 31680 28408 31686
rect 28356 31622 28408 31628
rect 27988 30660 28040 30666
rect 28092 30654 28212 30682
rect 27988 30602 28040 30608
rect 27804 30592 27856 30598
rect 27804 30534 27856 30540
rect 28080 30592 28132 30598
rect 28080 30534 28132 30540
rect 28092 30054 28120 30534
rect 28184 30394 28212 30654
rect 28172 30388 28224 30394
rect 28172 30330 28224 30336
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 27344 29844 27396 29850
rect 27344 29786 27396 29792
rect 26792 29708 26844 29714
rect 26792 29650 26844 29656
rect 26056 29572 26108 29578
rect 26056 29514 26108 29520
rect 26516 29572 26568 29578
rect 26516 29514 26568 29520
rect 26068 29306 26096 29514
rect 26132 29404 26440 29413
rect 26132 29402 26138 29404
rect 26194 29402 26218 29404
rect 26274 29402 26298 29404
rect 26354 29402 26378 29404
rect 26434 29402 26440 29404
rect 26194 29350 26196 29402
rect 26376 29350 26378 29402
rect 26132 29348 26138 29350
rect 26194 29348 26218 29350
rect 26274 29348 26298 29350
rect 26354 29348 26378 29350
rect 26434 29348 26440 29350
rect 26132 29339 26440 29348
rect 26528 29306 26556 29514
rect 26056 29300 26108 29306
rect 26056 29242 26108 29248
rect 26516 29300 26568 29306
rect 26516 29242 26568 29248
rect 26804 29170 26832 29650
rect 26792 29164 26844 29170
rect 26792 29106 26844 29112
rect 24964 28966 25084 28994
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24964 28014 24992 28966
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 26700 28552 26752 28558
rect 26700 28494 26752 28500
rect 24952 28008 25004 28014
rect 24952 27950 25004 27956
rect 25148 27878 25176 28494
rect 25780 28484 25832 28490
rect 25780 28426 25832 28432
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 24504 27662 24900 27690
rect 24872 26926 24900 27662
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24688 25226 24716 25842
rect 24872 25820 24900 26862
rect 25042 26480 25098 26489
rect 25042 26415 25098 26424
rect 25056 26382 25084 26415
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 25044 25832 25096 25838
rect 24872 25792 25044 25820
rect 25044 25774 25096 25780
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24872 24954 24900 25638
rect 24860 24948 24912 24954
rect 24860 24890 24912 24896
rect 24400 24744 24452 24750
rect 24400 24686 24452 24692
rect 24412 22642 24440 24686
rect 24872 24682 24900 24890
rect 25056 24886 25084 25774
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 24860 24676 24912 24682
rect 24860 24618 24912 24624
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24676 23656 24728 23662
rect 24676 23598 24728 23604
rect 24688 23118 24716 23598
rect 24872 23322 24900 24074
rect 25148 23610 25176 27814
rect 25608 26994 25636 28018
rect 25792 28014 25820 28426
rect 26132 28316 26440 28325
rect 26132 28314 26138 28316
rect 26194 28314 26218 28316
rect 26274 28314 26298 28316
rect 26354 28314 26378 28316
rect 26434 28314 26440 28316
rect 26194 28262 26196 28314
rect 26376 28262 26378 28314
rect 26132 28260 26138 28262
rect 26194 28260 26218 28262
rect 26274 28260 26298 28262
rect 26354 28260 26378 28262
rect 26434 28260 26440 28262
rect 26132 28251 26440 28260
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25884 27130 25912 27338
rect 26132 27228 26440 27237
rect 26132 27226 26138 27228
rect 26194 27226 26218 27228
rect 26274 27226 26298 27228
rect 26354 27226 26378 27228
rect 26434 27226 26440 27228
rect 26194 27174 26196 27226
rect 26376 27174 26378 27226
rect 26132 27172 26138 27174
rect 26194 27172 26218 27174
rect 26274 27172 26298 27174
rect 26354 27172 26378 27174
rect 26434 27172 26440 27174
rect 26132 27163 26440 27172
rect 26712 27130 26740 28494
rect 26804 28082 26832 29106
rect 27160 29028 27212 29034
rect 27160 28970 27212 28976
rect 26976 28416 27028 28422
rect 26976 28358 27028 28364
rect 26988 28218 27016 28358
rect 26976 28212 27028 28218
rect 26976 28154 27028 28160
rect 26792 28076 26844 28082
rect 26792 28018 26844 28024
rect 26804 27690 26832 28018
rect 26804 27662 26924 27690
rect 26896 27538 26924 27662
rect 26884 27532 26936 27538
rect 26884 27474 26936 27480
rect 27172 27402 27200 28970
rect 27160 27396 27212 27402
rect 27160 27338 27212 27344
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 26700 27124 26752 27130
rect 26700 27066 26752 27072
rect 27356 26994 27384 29786
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27724 28218 27752 28494
rect 27712 28212 27764 28218
rect 27712 28154 27764 28160
rect 27896 28008 27948 28014
rect 27896 27950 27948 27956
rect 27620 27872 27672 27878
rect 27620 27814 27672 27820
rect 27632 27674 27660 27814
rect 27620 27668 27672 27674
rect 27620 27610 27672 27616
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 27712 27396 27764 27402
rect 27764 27356 27844 27384
rect 27712 27338 27764 27344
rect 25228 26988 25280 26994
rect 25228 26930 25280 26936
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 25240 26586 25268 26930
rect 25228 26580 25280 26586
rect 25228 26522 25280 26528
rect 25332 25702 25360 26930
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 25320 25696 25372 25702
rect 25320 25638 25372 25644
rect 25424 25226 25452 26182
rect 25516 26042 25544 26250
rect 25504 26036 25556 26042
rect 25504 25978 25556 25984
rect 25608 25906 25636 26930
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 27252 26920 27304 26926
rect 27252 26862 27304 26868
rect 25688 26852 25740 26858
rect 25688 26794 25740 26800
rect 25596 25900 25648 25906
rect 25596 25842 25648 25848
rect 25700 25770 25728 26794
rect 26132 26140 26440 26149
rect 26132 26138 26138 26140
rect 26194 26138 26218 26140
rect 26274 26138 26298 26140
rect 26354 26138 26378 26140
rect 26434 26138 26440 26140
rect 26194 26086 26196 26138
rect 26376 26086 26378 26138
rect 26132 26084 26138 26086
rect 26194 26084 26218 26086
rect 26274 26084 26298 26086
rect 26354 26084 26378 26086
rect 26434 26084 26440 26086
rect 26132 26075 26440 26084
rect 26528 25906 26556 26862
rect 27160 26852 27212 26858
rect 27160 26794 27212 26800
rect 27172 25906 27200 26794
rect 27264 25906 27292 26862
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 26608 25900 26660 25906
rect 26608 25842 26660 25848
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 25688 25764 25740 25770
rect 25688 25706 25740 25712
rect 26528 25498 26556 25842
rect 26516 25492 26568 25498
rect 26516 25434 26568 25440
rect 26620 25294 26648 25842
rect 27160 25764 27212 25770
rect 27160 25706 27212 25712
rect 26608 25288 26660 25294
rect 26608 25230 26660 25236
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25424 24274 25452 25162
rect 26976 25152 27028 25158
rect 26976 25094 27028 25100
rect 26132 25052 26440 25061
rect 26132 25050 26138 25052
rect 26194 25050 26218 25052
rect 26274 25050 26298 25052
rect 26354 25050 26378 25052
rect 26434 25050 26440 25052
rect 26194 24998 26196 25050
rect 26376 24998 26378 25050
rect 26132 24996 26138 24998
rect 26194 24996 26218 24998
rect 26274 24996 26298 24998
rect 26354 24996 26378 24998
rect 26434 24996 26440 24998
rect 26132 24987 26440 24996
rect 26988 24818 27016 25094
rect 27172 24818 27200 25706
rect 26976 24812 27028 24818
rect 26976 24754 27028 24760
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 26516 24744 26568 24750
rect 26516 24686 26568 24692
rect 27068 24744 27120 24750
rect 27068 24686 27120 24692
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25872 24200 25924 24206
rect 26148 24200 26200 24206
rect 25872 24142 25924 24148
rect 25976 24148 26148 24154
rect 25976 24142 26200 24148
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 25228 23792 25280 23798
rect 25332 23746 25360 24074
rect 25280 23740 25360 23746
rect 25228 23734 25360 23740
rect 25240 23718 25360 23734
rect 25148 23582 25268 23610
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 25148 23118 25176 23462
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 25136 23112 25188 23118
rect 25136 23054 25188 23060
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24952 22568 25004 22574
rect 24952 22510 25004 22516
rect 24964 22234 24992 22510
rect 24308 22228 24360 22234
rect 24308 22170 24360 22176
rect 24952 22228 25004 22234
rect 24952 22170 25004 22176
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23860 21486 23888 21830
rect 24596 21486 24624 21966
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 24584 21480 24636 21486
rect 24584 21422 24636 21428
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 24412 20505 24440 20742
rect 24398 20496 24454 20505
rect 24872 20466 24900 22034
rect 24964 21690 24992 22170
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 25136 21616 25188 21622
rect 25136 21558 25188 21564
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24398 20431 24454 20440
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 23756 19984 23808 19990
rect 23808 19944 23980 19972
rect 23756 19926 23808 19932
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23400 19366 23520 19394
rect 23400 19242 23428 19366
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23388 19236 23440 19242
rect 23388 19178 23440 19184
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 22756 18584 22876 18612
rect 22928 18624 22980 18630
rect 22756 16794 22784 18584
rect 22928 18566 22980 18572
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 22940 18290 22968 18566
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 23032 18222 23060 18566
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 23124 18154 23152 18566
rect 23112 18148 23164 18154
rect 23112 18090 23164 18096
rect 23216 17882 23244 18906
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 23308 18426 23336 18566
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 22928 17604 22980 17610
rect 22848 17564 22928 17592
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22744 16176 22796 16182
rect 22848 16164 22876 17564
rect 22928 17546 22980 17552
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22796 16136 22876 16164
rect 22744 16118 22796 16124
rect 22940 16114 22968 16526
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22652 15972 22704 15978
rect 22652 15914 22704 15920
rect 22756 15638 22784 15982
rect 22940 15706 22968 16050
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 22744 15632 22796 15638
rect 22744 15574 22796 15580
rect 22650 15464 22706 15473
rect 22572 15422 22650 15450
rect 22650 15399 22706 15408
rect 22756 15094 22784 15574
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22756 14414 22784 15030
rect 22848 15026 22876 15370
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22940 14958 22968 15302
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22940 14414 22968 14894
rect 23032 14482 23060 14962
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22744 14408 22796 14414
rect 22928 14408 22980 14414
rect 22744 14350 22796 14356
rect 22848 14368 22928 14396
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22572 12306 22600 14214
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22652 13456 22704 13462
rect 22652 13398 22704 13404
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22572 11762 22600 12242
rect 22664 11830 22692 13398
rect 22652 11824 22704 11830
rect 22652 11766 22704 11772
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 21935 11452 22243 11461
rect 21935 11450 21941 11452
rect 21997 11450 22021 11452
rect 22077 11450 22101 11452
rect 22157 11450 22181 11452
rect 22237 11450 22243 11452
rect 21997 11398 21999 11450
rect 22179 11398 22181 11450
rect 21935 11396 21941 11398
rect 21997 11396 22021 11398
rect 22077 11396 22101 11398
rect 22157 11396 22181 11398
rect 22237 11396 22243 11398
rect 21935 11387 22243 11396
rect 22664 11150 22692 11766
rect 22756 11762 22784 13466
rect 22848 13462 22876 14368
rect 22928 14350 22980 14356
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22940 13326 22968 13738
rect 23124 13530 23152 16050
rect 23216 15434 23244 16186
rect 23296 16108 23348 16114
rect 23296 16050 23348 16056
rect 23308 15910 23336 16050
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23308 15570 23336 15846
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23294 15464 23350 15473
rect 23204 15428 23256 15434
rect 23294 15399 23296 15408
rect 23204 15370 23256 15376
rect 23348 15399 23350 15408
rect 23296 15370 23348 15376
rect 23216 15042 23244 15370
rect 23216 15026 23336 15042
rect 23216 15020 23348 15026
rect 23216 15014 23296 15020
rect 23296 14962 23348 14968
rect 23308 14414 23336 14962
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22940 12850 22968 13262
rect 23308 13190 23336 14350
rect 23400 13326 23428 19178
rect 23492 18290 23520 19246
rect 23676 18290 23704 19654
rect 23768 19446 23796 19790
rect 23756 19440 23808 19446
rect 23756 19382 23808 19388
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23492 17814 23520 18022
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23480 17808 23532 17814
rect 23480 17750 23532 17756
rect 23492 17678 23520 17750
rect 23584 17678 23612 17818
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23492 15978 23520 17478
rect 23676 16794 23704 17546
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23768 16250 23796 19382
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23860 17678 23888 18022
rect 23952 17882 23980 19944
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24412 19310 24440 19654
rect 25056 19446 25084 21490
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24952 19236 25004 19242
rect 24952 19178 25004 19184
rect 24964 18902 24992 19178
rect 25148 19174 25176 21558
rect 25240 21486 25268 23582
rect 25332 21894 25360 23718
rect 25884 23186 25912 24142
rect 25976 24126 26188 24142
rect 25976 23798 26004 24126
rect 26132 23964 26440 23973
rect 26132 23962 26138 23964
rect 26194 23962 26218 23964
rect 26274 23962 26298 23964
rect 26354 23962 26378 23964
rect 26434 23962 26440 23964
rect 26194 23910 26196 23962
rect 26376 23910 26378 23962
rect 26132 23908 26138 23910
rect 26194 23908 26218 23910
rect 26274 23908 26298 23910
rect 26354 23908 26378 23910
rect 26434 23908 26440 23910
rect 26132 23899 26440 23908
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 25872 23180 25924 23186
rect 25872 23122 25924 23128
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25332 21554 25360 21830
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25424 20534 25452 20742
rect 25412 20528 25464 20534
rect 25412 20470 25464 20476
rect 25608 20058 25636 20878
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25700 19854 25728 20198
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 24952 18896 25004 18902
rect 24952 18838 25004 18844
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 24136 16522 24164 18158
rect 24412 17882 24440 18702
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18426 24624 18566
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24964 18358 24992 18838
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24780 16794 24808 17750
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24780 16538 24808 16730
rect 24872 16658 24900 17478
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24688 16510 24808 16538
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 24136 16114 24164 16458
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24412 16250 24440 16390
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23492 15638 23520 15914
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 24136 15570 24164 16050
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24136 14074 24164 15506
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23676 13530 23704 13874
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 24136 13394 24164 14010
rect 24688 13394 24716 16510
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24780 16250 24808 16390
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 25596 16040 25648 16046
rect 25596 15982 25648 15988
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24964 15162 24992 15302
rect 25516 15162 25544 15438
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25608 14006 25636 15982
rect 25976 14958 26004 23734
rect 26528 23730 26556 24686
rect 27080 24274 27108 24686
rect 27068 24268 27120 24274
rect 27068 24210 27120 24216
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 26608 24064 26660 24070
rect 26608 24006 26660 24012
rect 26620 23866 26648 24006
rect 27172 23866 27200 24142
rect 26608 23860 26660 23866
rect 26608 23802 26660 23808
rect 27160 23860 27212 23866
rect 27160 23802 27212 23808
rect 26516 23724 26568 23730
rect 26516 23666 26568 23672
rect 26132 22876 26440 22885
rect 26132 22874 26138 22876
rect 26194 22874 26218 22876
rect 26274 22874 26298 22876
rect 26354 22874 26378 22876
rect 26434 22874 26440 22876
rect 26194 22822 26196 22874
rect 26376 22822 26378 22874
rect 26132 22820 26138 22822
rect 26194 22820 26218 22822
rect 26274 22820 26298 22822
rect 26354 22820 26378 22822
rect 26434 22820 26440 22822
rect 26132 22811 26440 22820
rect 26132 21788 26440 21797
rect 26132 21786 26138 21788
rect 26194 21786 26218 21788
rect 26274 21786 26298 21788
rect 26354 21786 26378 21788
rect 26434 21786 26440 21788
rect 26194 21734 26196 21786
rect 26376 21734 26378 21786
rect 26132 21732 26138 21734
rect 26194 21732 26218 21734
rect 26274 21732 26298 21734
rect 26354 21732 26378 21734
rect 26434 21732 26440 21734
rect 26132 21723 26440 21732
rect 26528 21350 26556 23666
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 27264 23186 27292 23462
rect 27252 23180 27304 23186
rect 27252 23122 27304 23128
rect 27540 22094 27568 27338
rect 27816 25514 27844 27356
rect 27908 27062 27936 27950
rect 28184 27554 28212 30330
rect 28264 30320 28316 30326
rect 28264 30262 28316 30268
rect 28276 29306 28304 30262
rect 28368 30190 28396 31622
rect 28460 31482 28488 31690
rect 28448 31476 28500 31482
rect 28448 31418 28500 31424
rect 28552 30326 28580 32438
rect 28828 32230 28856 32438
rect 28908 32360 28960 32366
rect 28908 32302 28960 32308
rect 28816 32224 28868 32230
rect 28816 32166 28868 32172
rect 28920 32026 28948 32302
rect 30329 32124 30637 32133
rect 30329 32122 30335 32124
rect 30391 32122 30415 32124
rect 30471 32122 30495 32124
rect 30551 32122 30575 32124
rect 30631 32122 30637 32124
rect 30391 32070 30393 32122
rect 30573 32070 30575 32122
rect 30329 32068 30335 32070
rect 30391 32068 30415 32070
rect 30471 32068 30495 32070
rect 30551 32068 30575 32070
rect 30631 32068 30637 32070
rect 30329 32059 30637 32068
rect 28908 32020 28960 32026
rect 28908 31962 28960 31968
rect 29736 31272 29788 31278
rect 29736 31214 29788 31220
rect 28908 30660 28960 30666
rect 28908 30602 28960 30608
rect 28540 30320 28592 30326
rect 28540 30262 28592 30268
rect 28920 30240 28948 30602
rect 29748 30394 29776 31214
rect 30329 31036 30637 31045
rect 30329 31034 30335 31036
rect 30391 31034 30415 31036
rect 30471 31034 30495 31036
rect 30551 31034 30575 31036
rect 30631 31034 30637 31036
rect 30391 30982 30393 31034
rect 30573 30982 30575 31034
rect 30329 30980 30335 30982
rect 30391 30980 30415 30982
rect 30471 30980 30495 30982
rect 30551 30980 30575 30982
rect 30631 30980 30637 30982
rect 30329 30971 30637 30980
rect 29736 30388 29788 30394
rect 29736 30330 29788 30336
rect 29276 30252 29328 30258
rect 28920 30212 29276 30240
rect 28356 30184 28408 30190
rect 28356 30126 28408 30132
rect 28264 29300 28316 29306
rect 28264 29242 28316 29248
rect 28092 27538 28212 27554
rect 28276 27538 28304 29242
rect 29196 29238 29224 30212
rect 29276 30194 29328 30200
rect 30329 29948 30637 29957
rect 30329 29946 30335 29948
rect 30391 29946 30415 29948
rect 30471 29946 30495 29948
rect 30551 29946 30575 29948
rect 30631 29946 30637 29948
rect 30391 29894 30393 29946
rect 30573 29894 30575 29946
rect 30329 29892 30335 29894
rect 30391 29892 30415 29894
rect 30471 29892 30495 29894
rect 30551 29892 30575 29894
rect 30631 29892 30637 29894
rect 30329 29883 30637 29892
rect 29460 29640 29512 29646
rect 29460 29582 29512 29588
rect 30840 29640 30892 29646
rect 30840 29582 30892 29588
rect 29368 29504 29420 29510
rect 29368 29446 29420 29452
rect 29184 29232 29236 29238
rect 29184 29174 29236 29180
rect 29196 28966 29224 29174
rect 29380 29034 29408 29446
rect 29472 29238 29500 29582
rect 29552 29504 29604 29510
rect 29552 29446 29604 29452
rect 29460 29232 29512 29238
rect 29460 29174 29512 29180
rect 29564 29170 29592 29446
rect 29552 29164 29604 29170
rect 29552 29106 29604 29112
rect 29368 29028 29420 29034
rect 29368 28970 29420 28976
rect 29184 28960 29236 28966
rect 28460 28886 28948 28914
rect 29184 28902 29236 28908
rect 28460 28762 28488 28886
rect 28448 28756 28500 28762
rect 28448 28698 28500 28704
rect 28540 28756 28592 28762
rect 28540 28698 28592 28704
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28552 28370 28580 28698
rect 28816 28688 28868 28694
rect 28644 28636 28816 28642
rect 28644 28630 28868 28636
rect 28920 28642 28948 28886
rect 28644 28614 28856 28630
rect 28920 28626 28994 28642
rect 28920 28620 29006 28626
rect 28920 28614 28954 28620
rect 28644 28558 28672 28614
rect 28954 28562 29006 28568
rect 28632 28552 28684 28558
rect 28632 28494 28684 28500
rect 28954 28484 29006 28490
rect 28828 28444 28954 28472
rect 28828 28370 28856 28444
rect 28954 28426 29006 28432
rect 29092 28416 29144 28422
rect 28368 28014 28396 28358
rect 28552 28342 28856 28370
rect 28920 28364 29092 28370
rect 28920 28358 29144 28364
rect 28920 28342 29132 28358
rect 28356 28008 28408 28014
rect 28356 27950 28408 27956
rect 28080 27532 28212 27538
rect 28132 27526 28212 27532
rect 28264 27532 28316 27538
rect 28080 27474 28132 27480
rect 28264 27474 28316 27480
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 27896 27056 27948 27062
rect 27896 26998 27948 27004
rect 27908 26586 27936 26998
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 27896 26580 27948 26586
rect 27896 26522 27948 26528
rect 28000 26314 28028 26930
rect 28080 26784 28132 26790
rect 28080 26726 28132 26732
rect 28092 26382 28120 26726
rect 28080 26376 28132 26382
rect 28080 26318 28132 26324
rect 27988 26308 28040 26314
rect 27988 26250 28040 26256
rect 27724 25486 27844 25514
rect 27724 23866 27752 25486
rect 27804 25424 27856 25430
rect 27804 25366 27856 25372
rect 27712 23860 27764 23866
rect 27712 23802 27764 23808
rect 27356 22066 27568 22094
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 26620 21690 26648 21830
rect 26608 21684 26660 21690
rect 26608 21626 26660 21632
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26620 21146 26648 21490
rect 26884 21344 26936 21350
rect 26884 21286 26936 21292
rect 26608 21140 26660 21146
rect 26608 21082 26660 21088
rect 26896 21010 26924 21286
rect 26884 21004 26936 21010
rect 26884 20946 26936 20952
rect 26132 20700 26440 20709
rect 26132 20698 26138 20700
rect 26194 20698 26218 20700
rect 26274 20698 26298 20700
rect 26354 20698 26378 20700
rect 26434 20698 26440 20700
rect 26194 20646 26196 20698
rect 26376 20646 26378 20698
rect 26132 20644 26138 20646
rect 26194 20644 26218 20646
rect 26274 20644 26298 20646
rect 26354 20644 26378 20646
rect 26434 20644 26440 20646
rect 26132 20635 26440 20644
rect 26896 19922 26924 20946
rect 26988 20602 27016 21490
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26132 19612 26440 19621
rect 26132 19610 26138 19612
rect 26194 19610 26218 19612
rect 26274 19610 26298 19612
rect 26354 19610 26378 19612
rect 26434 19610 26440 19612
rect 26194 19558 26196 19610
rect 26376 19558 26378 19610
rect 26132 19556 26138 19558
rect 26194 19556 26218 19558
rect 26274 19556 26298 19558
rect 26354 19556 26378 19558
rect 26434 19556 26440 19558
rect 26132 19547 26440 19556
rect 26804 19446 26832 19790
rect 26792 19440 26844 19446
rect 26792 19382 26844 19388
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26528 18970 26556 19314
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 26132 18524 26440 18533
rect 26132 18522 26138 18524
rect 26194 18522 26218 18524
rect 26274 18522 26298 18524
rect 26354 18522 26378 18524
rect 26434 18522 26440 18524
rect 26194 18470 26196 18522
rect 26376 18470 26378 18522
rect 26132 18468 26138 18470
rect 26194 18468 26218 18470
rect 26274 18468 26298 18470
rect 26354 18468 26378 18470
rect 26434 18468 26440 18470
rect 26132 18459 26440 18468
rect 26804 18426 26832 19110
rect 26896 18834 26924 19858
rect 26988 19378 27016 20538
rect 27356 19446 27384 22066
rect 27712 21616 27764 21622
rect 27712 21558 27764 21564
rect 27724 20534 27752 21558
rect 27712 20528 27764 20534
rect 27712 20470 27764 20476
rect 27724 20262 27752 20470
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27816 19922 27844 25366
rect 27896 24064 27948 24070
rect 27896 24006 27948 24012
rect 27908 23866 27936 24006
rect 27896 23860 27948 23866
rect 27896 23802 27948 23808
rect 28000 23186 28028 26250
rect 28184 25906 28212 27406
rect 28276 26994 28304 27474
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 28172 25900 28224 25906
rect 28172 25842 28224 25848
rect 28276 24818 28304 26930
rect 28368 25684 28396 27950
rect 28920 27606 28948 28342
rect 28908 27600 28960 27606
rect 28908 27542 28960 27548
rect 29092 27396 29144 27402
rect 29092 27338 29144 27344
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28460 26382 28488 27270
rect 28540 26920 28592 26926
rect 28540 26862 28592 26868
rect 28632 26920 28684 26926
rect 28632 26862 28684 26868
rect 28552 26586 28580 26862
rect 28540 26580 28592 26586
rect 28540 26522 28592 26528
rect 28644 26466 28672 26862
rect 28552 26438 28672 26466
rect 28908 26512 28960 26518
rect 28908 26454 28960 26460
rect 28552 26382 28580 26438
rect 28448 26376 28500 26382
rect 28448 26318 28500 26324
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28448 25696 28500 25702
rect 28368 25656 28448 25684
rect 28448 25638 28500 25644
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28356 23724 28408 23730
rect 28356 23666 28408 23672
rect 28368 23322 28396 23666
rect 28356 23316 28408 23322
rect 28356 23258 28408 23264
rect 27988 23180 28040 23186
rect 27988 23122 28040 23128
rect 28000 20482 28028 23122
rect 28460 23100 28488 25638
rect 28552 24342 28580 26318
rect 28632 26308 28684 26314
rect 28632 26250 28684 26256
rect 28644 24750 28672 26250
rect 28816 25492 28868 25498
rect 28816 25434 28868 25440
rect 28828 24750 28856 25434
rect 28632 24744 28684 24750
rect 28632 24686 28684 24692
rect 28816 24744 28868 24750
rect 28816 24686 28868 24692
rect 28540 24336 28592 24342
rect 28540 24278 28592 24284
rect 28644 23798 28672 24686
rect 28632 23792 28684 23798
rect 28632 23734 28684 23740
rect 28540 23656 28592 23662
rect 28540 23598 28592 23604
rect 28552 23254 28580 23598
rect 28540 23248 28592 23254
rect 28540 23190 28592 23196
rect 28920 23186 28948 26454
rect 29104 26382 29132 27338
rect 29196 27130 29224 28902
rect 29380 28762 29408 28970
rect 29368 28756 29420 28762
rect 29368 28698 29420 28704
rect 29564 28626 29592 29106
rect 29644 28960 29696 28966
rect 29644 28902 29696 28908
rect 29656 28626 29684 28902
rect 30329 28860 30637 28869
rect 30329 28858 30335 28860
rect 30391 28858 30415 28860
rect 30471 28858 30495 28860
rect 30551 28858 30575 28860
rect 30631 28858 30637 28860
rect 30391 28806 30393 28858
rect 30573 28806 30575 28858
rect 30329 28804 30335 28806
rect 30391 28804 30415 28806
rect 30471 28804 30495 28806
rect 30551 28804 30575 28806
rect 30631 28804 30637 28806
rect 30329 28795 30637 28804
rect 30852 28762 30880 29582
rect 30840 28756 30892 28762
rect 30840 28698 30892 28704
rect 29552 28620 29604 28626
rect 29552 28562 29604 28568
rect 29644 28620 29696 28626
rect 29644 28562 29696 28568
rect 30564 28552 30616 28558
rect 30564 28494 30616 28500
rect 30576 28218 30604 28494
rect 30656 28416 30708 28422
rect 30656 28358 30708 28364
rect 30564 28212 30616 28218
rect 30564 28154 30616 28160
rect 30329 27772 30637 27781
rect 30329 27770 30335 27772
rect 30391 27770 30415 27772
rect 30471 27770 30495 27772
rect 30551 27770 30575 27772
rect 30631 27770 30637 27772
rect 30391 27718 30393 27770
rect 30573 27718 30575 27770
rect 30329 27716 30335 27718
rect 30391 27716 30415 27718
rect 30471 27716 30495 27718
rect 30551 27716 30575 27718
rect 30631 27716 30637 27718
rect 30329 27707 30637 27716
rect 30668 27402 30696 28358
rect 30748 28144 30800 28150
rect 30748 28086 30800 28092
rect 30760 27674 30788 28086
rect 30932 27940 30984 27946
rect 30932 27882 30984 27888
rect 30944 27674 30972 27882
rect 30748 27668 30800 27674
rect 30748 27610 30800 27616
rect 30932 27668 30984 27674
rect 30932 27610 30984 27616
rect 30656 27396 30708 27402
rect 30656 27338 30708 27344
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 30668 26994 30696 27338
rect 30656 26988 30708 26994
rect 30656 26930 30708 26936
rect 29920 26784 29972 26790
rect 29920 26726 29972 26732
rect 29092 26376 29144 26382
rect 29092 26318 29144 26324
rect 29828 26376 29880 26382
rect 29828 26318 29880 26324
rect 29000 25968 29052 25974
rect 29000 25910 29052 25916
rect 29012 24886 29040 25910
rect 29840 25498 29868 26318
rect 29828 25492 29880 25498
rect 29828 25434 29880 25440
rect 29840 25226 29868 25434
rect 29184 25220 29236 25226
rect 29184 25162 29236 25168
rect 29828 25220 29880 25226
rect 29828 25162 29880 25168
rect 29000 24880 29052 24886
rect 29000 24822 29052 24828
rect 29196 24682 29224 25162
rect 29460 24812 29512 24818
rect 29460 24754 29512 24760
rect 29184 24676 29236 24682
rect 29184 24618 29236 24624
rect 29472 24206 29500 24754
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 29828 24132 29880 24138
rect 29828 24074 29880 24080
rect 29736 23724 29788 23730
rect 29736 23666 29788 23672
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 28460 23072 28580 23100
rect 28172 20800 28224 20806
rect 28172 20742 28224 20748
rect 28080 20528 28132 20534
rect 28000 20476 28080 20482
rect 28000 20470 28132 20476
rect 28000 20454 28120 20470
rect 28000 20262 28028 20454
rect 28184 20262 28212 20742
rect 27988 20256 28040 20262
rect 27988 20198 28040 20204
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 27804 19916 27856 19922
rect 27804 19858 27856 19864
rect 28448 19916 28500 19922
rect 28448 19858 28500 19864
rect 28172 19780 28224 19786
rect 28172 19722 28224 19728
rect 27344 19440 27396 19446
rect 27344 19382 27396 19388
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 26884 18828 26936 18834
rect 26884 18770 26936 18776
rect 26792 18420 26844 18426
rect 26792 18362 26844 18368
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26620 17542 26648 17614
rect 26608 17536 26660 17542
rect 26608 17478 26660 17484
rect 26700 17536 26752 17542
rect 26700 17478 26752 17484
rect 26132 17436 26440 17445
rect 26132 17434 26138 17436
rect 26194 17434 26218 17436
rect 26274 17434 26298 17436
rect 26354 17434 26378 17436
rect 26434 17434 26440 17436
rect 26194 17382 26196 17434
rect 26376 17382 26378 17434
rect 26132 17380 26138 17382
rect 26194 17380 26218 17382
rect 26274 17380 26298 17382
rect 26354 17380 26378 17382
rect 26434 17380 26440 17382
rect 26132 17371 26440 17380
rect 26712 16794 26740 17478
rect 26700 16788 26752 16794
rect 26700 16730 26752 16736
rect 26804 16522 26832 18362
rect 26896 17814 26924 18770
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 26884 17808 26936 17814
rect 26884 17750 26936 17756
rect 27816 17746 27844 18022
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 28184 17678 28212 19722
rect 28264 18692 28316 18698
rect 28264 18634 28316 18640
rect 28276 18086 28304 18634
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28276 17678 28304 18022
rect 27988 17672 28040 17678
rect 28172 17672 28224 17678
rect 27988 17614 28040 17620
rect 28092 17632 28172 17660
rect 27620 17604 27672 17610
rect 27620 17546 27672 17552
rect 27896 17604 27948 17610
rect 27896 17546 27948 17552
rect 27632 17066 27660 17546
rect 27620 17060 27672 17066
rect 27620 17002 27672 17008
rect 27632 16794 27660 17002
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26792 16516 26844 16522
rect 26712 16476 26792 16504
rect 26132 16348 26440 16357
rect 26132 16346 26138 16348
rect 26194 16346 26218 16348
rect 26274 16346 26298 16348
rect 26354 16346 26378 16348
rect 26434 16346 26440 16348
rect 26194 16294 26196 16346
rect 26376 16294 26378 16346
rect 26132 16292 26138 16294
rect 26194 16292 26218 16294
rect 26274 16292 26298 16294
rect 26354 16292 26378 16294
rect 26434 16292 26440 16294
rect 26132 16283 26440 16292
rect 26712 16182 26740 16476
rect 26792 16458 26844 16464
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26700 16176 26752 16182
rect 26700 16118 26752 16124
rect 26804 15706 26832 16186
rect 26896 16114 26924 16594
rect 27712 16448 27764 16454
rect 27712 16390 27764 16396
rect 27724 16250 27752 16390
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 26884 16108 26936 16114
rect 26884 16050 26936 16056
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26132 15260 26440 15269
rect 26132 15258 26138 15260
rect 26194 15258 26218 15260
rect 26274 15258 26298 15260
rect 26354 15258 26378 15260
rect 26434 15258 26440 15260
rect 26194 15206 26196 15258
rect 26376 15206 26378 15258
rect 26132 15204 26138 15206
rect 26194 15204 26218 15206
rect 26274 15204 26298 15206
rect 26354 15204 26378 15206
rect 26434 15204 26440 15206
rect 26132 15195 26440 15204
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25976 14482 26004 14894
rect 26896 14550 26924 16050
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27448 15434 27476 15982
rect 27908 15638 27936 17546
rect 28000 17338 28028 17614
rect 27988 17332 28040 17338
rect 27988 17274 28040 17280
rect 28092 15638 28120 17632
rect 28172 17614 28224 17620
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28368 17354 28396 18226
rect 28460 17678 28488 19858
rect 28552 17882 28580 23072
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28644 21894 28672 22578
rect 28632 21888 28684 21894
rect 28632 21830 28684 21836
rect 28816 21344 28868 21350
rect 28816 21286 28868 21292
rect 28828 21146 28856 21286
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28736 20058 28764 20878
rect 28724 20052 28776 20058
rect 28724 19994 28776 20000
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 28736 18834 28764 19246
rect 28920 18850 28948 23122
rect 29092 23112 29144 23118
rect 29092 23054 29144 23060
rect 29104 22574 29132 23054
rect 29748 22778 29776 23666
rect 29736 22772 29788 22778
rect 29736 22714 29788 22720
rect 29840 22658 29868 24074
rect 29932 23730 29960 26726
rect 30329 26684 30637 26693
rect 30329 26682 30335 26684
rect 30391 26682 30415 26684
rect 30471 26682 30495 26684
rect 30551 26682 30575 26684
rect 30631 26682 30637 26684
rect 30391 26630 30393 26682
rect 30573 26630 30575 26682
rect 30329 26628 30335 26630
rect 30391 26628 30415 26630
rect 30471 26628 30495 26630
rect 30551 26628 30575 26630
rect 30631 26628 30637 26630
rect 30329 26619 30637 26628
rect 30472 26240 30524 26246
rect 30472 26182 30524 26188
rect 30484 26042 30512 26182
rect 30472 26036 30524 26042
rect 30472 25978 30524 25984
rect 30012 25900 30064 25906
rect 30012 25842 30064 25848
rect 30024 25498 30052 25842
rect 30656 25832 30708 25838
rect 30656 25774 30708 25780
rect 30329 25596 30637 25605
rect 30329 25594 30335 25596
rect 30391 25594 30415 25596
rect 30471 25594 30495 25596
rect 30551 25594 30575 25596
rect 30631 25594 30637 25596
rect 30391 25542 30393 25594
rect 30573 25542 30575 25594
rect 30329 25540 30335 25542
rect 30391 25540 30415 25542
rect 30471 25540 30495 25542
rect 30551 25540 30575 25542
rect 30631 25540 30637 25542
rect 30329 25531 30637 25540
rect 30012 25492 30064 25498
rect 30012 25434 30064 25440
rect 30196 25152 30248 25158
rect 30196 25094 30248 25100
rect 30208 24886 30236 25094
rect 30668 24954 30696 25774
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30656 24948 30708 24954
rect 30656 24890 30708 24896
rect 30196 24880 30248 24886
rect 30196 24822 30248 24828
rect 30012 24676 30064 24682
rect 30012 24618 30064 24624
rect 30024 23730 30052 24618
rect 30208 24324 30236 24822
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 30329 24508 30637 24517
rect 30329 24506 30335 24508
rect 30391 24506 30415 24508
rect 30471 24506 30495 24508
rect 30551 24506 30575 24508
rect 30631 24506 30637 24508
rect 30391 24454 30393 24506
rect 30573 24454 30575 24506
rect 30329 24452 30335 24454
rect 30391 24452 30415 24454
rect 30471 24452 30495 24454
rect 30551 24452 30575 24454
rect 30631 24452 30637 24454
rect 30329 24443 30637 24452
rect 30208 24296 30328 24324
rect 30104 24064 30156 24070
rect 30104 24006 30156 24012
rect 30116 23730 30144 24006
rect 30300 23730 30328 24296
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 30012 23724 30064 23730
rect 30012 23666 30064 23672
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 29932 23254 29960 23666
rect 30329 23420 30637 23429
rect 30329 23418 30335 23420
rect 30391 23418 30415 23420
rect 30471 23418 30495 23420
rect 30551 23418 30575 23420
rect 30631 23418 30637 23420
rect 30391 23366 30393 23418
rect 30573 23366 30575 23418
rect 30329 23364 30335 23366
rect 30391 23364 30415 23366
rect 30471 23364 30495 23366
rect 30551 23364 30575 23366
rect 30631 23364 30637 23366
rect 30329 23355 30637 23364
rect 30668 23322 30696 24550
rect 30656 23316 30708 23322
rect 30656 23258 30708 23264
rect 29920 23248 29972 23254
rect 30852 23202 30880 25094
rect 29920 23190 29972 23196
rect 29932 22778 29960 23190
rect 30668 23174 30880 23202
rect 30012 22976 30064 22982
rect 30012 22918 30064 22924
rect 29920 22772 29972 22778
rect 29920 22714 29972 22720
rect 29748 22630 29868 22658
rect 29092 22568 29144 22574
rect 29092 22510 29144 22516
rect 29748 22438 29776 22630
rect 30024 22574 30052 22918
rect 30012 22568 30064 22574
rect 30012 22510 30064 22516
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 29748 20602 29776 22374
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 29828 21344 29880 21350
rect 29828 21286 29880 21292
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29368 19848 29420 19854
rect 29368 19790 29420 19796
rect 29380 18970 29408 19790
rect 29368 18964 29420 18970
rect 29368 18906 29420 18912
rect 28724 18828 28776 18834
rect 28920 18822 29040 18850
rect 28724 18770 28776 18776
rect 29012 18766 29040 18822
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 28644 17882 28672 18702
rect 28540 17876 28592 17882
rect 28540 17818 28592 17824
rect 28632 17876 28684 17882
rect 28632 17818 28684 17824
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28184 17326 28396 17354
rect 28184 16182 28212 17326
rect 28552 17218 28580 17818
rect 29012 17338 29040 18702
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29380 18086 29408 18566
rect 29748 18290 29776 20538
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 29368 18080 29420 18086
rect 29368 18022 29420 18028
rect 29552 17536 29604 17542
rect 29552 17478 29604 17484
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 28368 17202 28856 17218
rect 28368 17196 28868 17202
rect 28368 17190 28816 17196
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28172 16176 28224 16182
rect 28172 16118 28224 16124
rect 28184 16046 28212 16118
rect 28172 16040 28224 16046
rect 28172 15982 28224 15988
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 27896 15632 27948 15638
rect 27896 15574 27948 15580
rect 28080 15632 28132 15638
rect 28080 15574 28132 15580
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 26884 14544 26936 14550
rect 26884 14486 26936 14492
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 25700 14074 25728 14350
rect 26528 14334 26740 14362
rect 26528 14278 26556 14334
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 25596 14000 25648 14006
rect 25596 13942 25648 13948
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12986 23336 13126
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 22928 12844 22980 12850
rect 22848 12804 22928 12832
rect 22848 12306 22876 12804
rect 22928 12786 22980 12792
rect 23308 12374 23336 12922
rect 23400 12918 23428 13262
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23572 13184 23624 13190
rect 23572 13126 23624 13132
rect 23388 12912 23440 12918
rect 23388 12854 23440 12860
rect 23584 12782 23612 13126
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23492 12442 23520 12718
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23584 12306 23612 12718
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23676 12170 23704 13194
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22756 11150 22784 11698
rect 22836 11620 22888 11626
rect 22836 11562 22888 11568
rect 22928 11620 22980 11626
rect 22928 11562 22980 11568
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22572 10962 22600 11018
rect 22848 10962 22876 11562
rect 22940 11218 22968 11562
rect 22928 11212 22980 11218
rect 22928 11154 22980 11160
rect 22572 10934 22876 10962
rect 21935 10364 22243 10373
rect 21935 10362 21941 10364
rect 21997 10362 22021 10364
rect 22077 10362 22101 10364
rect 22157 10362 22181 10364
rect 22237 10362 22243 10364
rect 21997 10310 21999 10362
rect 22179 10310 22181 10362
rect 21935 10308 21941 10310
rect 21997 10308 22021 10310
rect 22077 10308 22101 10310
rect 22157 10308 22181 10310
rect 22237 10308 22243 10310
rect 21935 10299 22243 10308
rect 21824 9686 21876 9692
rect 21640 9648 21692 9654
rect 21640 9590 21692 9596
rect 21732 9648 21784 9654
rect 22572 9654 22600 10934
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22940 10266 22968 10406
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 23124 9722 23152 10610
rect 23480 10124 23532 10130
rect 23480 10066 23532 10072
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 22560 9648 22612 9654
rect 21876 9634 22416 9636
rect 21824 9628 22416 9634
rect 21836 9608 22416 9628
rect 21732 9590 21784 9596
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21376 8634 21404 9522
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22020 9364 22048 9454
rect 21836 9336 22048 9364
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20456 7886 20484 8230
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20456 7546 20484 7822
rect 21468 7750 21496 8434
rect 21652 7750 21680 8978
rect 21732 8900 21784 8906
rect 21732 8842 21784 8848
rect 21744 8362 21772 8842
rect 21836 8566 21864 9336
rect 21935 9276 22243 9285
rect 21935 9274 21941 9276
rect 21997 9274 22021 9276
rect 22077 9274 22101 9276
rect 22157 9274 22181 9276
rect 22237 9274 22243 9276
rect 21997 9222 21999 9274
rect 22179 9222 22181 9274
rect 21935 9220 21941 9222
rect 21997 9220 22021 9222
rect 22077 9220 22101 9222
rect 22157 9220 22181 9222
rect 22237 9220 22243 9222
rect 21935 9211 22243 9220
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21928 8634 21956 8978
rect 21916 8628 21968 8634
rect 21916 8570 21968 8576
rect 21824 8560 21876 8566
rect 21824 8502 21876 8508
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21836 8242 21864 8502
rect 21744 8214 21864 8242
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6458 19380 6598
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19536 5778 19564 6054
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19260 5522 19288 5714
rect 19996 5642 20024 6666
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 19260 5494 19380 5522
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 19352 3602 19380 5494
rect 19996 5370 20024 5578
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4078 19472 4422
rect 19904 4146 19932 5102
rect 19996 4214 20024 5306
rect 20272 5302 20300 6054
rect 20548 5914 20576 6258
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 21468 5642 21496 7686
rect 21652 7546 21680 7686
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 21468 5302 21496 5578
rect 21744 5556 21772 8214
rect 21935 8188 22243 8197
rect 21935 8186 21941 8188
rect 21997 8186 22021 8188
rect 22077 8186 22101 8188
rect 22157 8186 22181 8188
rect 22237 8186 22243 8188
rect 21997 8134 21999 8186
rect 22179 8134 22181 8186
rect 21935 8132 21941 8134
rect 21997 8132 22021 8134
rect 22077 8132 22101 8134
rect 22157 8132 22181 8134
rect 22237 8132 22243 8134
rect 21935 8123 22243 8132
rect 22296 7954 22324 9454
rect 22388 9042 22416 9608
rect 22558 9616 22560 9625
rect 22612 9616 22614 9625
rect 22558 9551 22614 9560
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22100 7472 22152 7478
rect 22152 7420 22232 7426
rect 22100 7414 22232 7420
rect 22112 7398 22232 7414
rect 22204 7342 22232 7398
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 21935 7100 22243 7109
rect 21935 7098 21941 7100
rect 21997 7098 22021 7100
rect 22077 7098 22101 7100
rect 22157 7098 22181 7100
rect 22237 7098 22243 7100
rect 21997 7046 21999 7098
rect 22179 7046 22181 7098
rect 21935 7044 21941 7046
rect 21997 7044 22021 7046
rect 22077 7044 22101 7046
rect 22157 7044 22181 7046
rect 22237 7044 22243 7046
rect 21935 7035 22243 7044
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21836 5914 21864 6054
rect 21935 6012 22243 6021
rect 21935 6010 21941 6012
rect 21997 6010 22021 6012
rect 22077 6010 22101 6012
rect 22157 6010 22181 6012
rect 22237 6010 22243 6012
rect 21997 5958 21999 6010
rect 22179 5958 22181 6010
rect 21935 5956 21941 5958
rect 21997 5956 22021 5958
rect 22077 5956 22101 5958
rect 22157 5956 22181 5958
rect 22237 5956 22243 5958
rect 21935 5947 22243 5956
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 22296 5778 22324 7142
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 21824 5568 21876 5574
rect 21744 5528 21824 5556
rect 21824 5510 21876 5516
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21192 4690 21220 5102
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21836 4622 21864 4966
rect 21935 4924 22243 4933
rect 21935 4922 21941 4924
rect 21997 4922 22021 4924
rect 22077 4922 22101 4924
rect 22157 4922 22181 4924
rect 22237 4922 22243 4924
rect 21997 4870 21999 4922
rect 22179 4870 22181 4922
rect 21935 4868 21941 4870
rect 21997 4868 22021 4870
rect 22077 4868 22101 4870
rect 22157 4868 22181 4870
rect 22237 4868 22243 4870
rect 21935 4859 22243 4868
rect 22296 4690 22324 5714
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 22388 4078 22416 8298
rect 22480 6458 22508 8910
rect 22572 8498 22600 9386
rect 23492 8498 23520 10066
rect 23768 9178 23796 12174
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11898 24072 12038
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 24136 10674 24164 13330
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24124 10668 24176 10674
rect 24124 10610 24176 10616
rect 24136 10130 24164 10610
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22480 5370 22508 6258
rect 22664 6254 22692 7890
rect 22940 7546 22968 8230
rect 23124 8090 23152 8434
rect 23768 8430 23796 8774
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23492 7954 23520 8298
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23768 7546 23796 7822
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 24228 7410 24256 12718
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24688 12170 24716 12582
rect 24676 12164 24728 12170
rect 24676 12106 24728 12112
rect 24872 11898 24900 12786
rect 24964 12186 24992 13330
rect 25516 12918 25544 13874
rect 25504 12912 25556 12918
rect 25504 12854 25556 12860
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 25056 12442 25084 12786
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 25608 12220 25636 13942
rect 26068 13326 26096 14214
rect 26132 14172 26440 14181
rect 26132 14170 26138 14172
rect 26194 14170 26218 14172
rect 26274 14170 26298 14172
rect 26354 14170 26378 14172
rect 26434 14170 26440 14172
rect 26194 14118 26196 14170
rect 26376 14118 26378 14170
rect 26132 14116 26138 14118
rect 26194 14116 26218 14118
rect 26274 14116 26298 14118
rect 26354 14116 26378 14118
rect 26434 14116 26440 14118
rect 26132 14107 26440 14116
rect 26620 14074 26648 14214
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26516 14000 26568 14006
rect 26516 13942 26568 13948
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 26132 13084 26440 13093
rect 26132 13082 26138 13084
rect 26194 13082 26218 13084
rect 26274 13082 26298 13084
rect 26354 13082 26378 13084
rect 26434 13082 26440 13084
rect 26194 13030 26196 13082
rect 26376 13030 26378 13082
rect 26132 13028 26138 13030
rect 26194 13028 26218 13030
rect 26274 13028 26298 13030
rect 26354 13028 26378 13030
rect 26434 13028 26440 13030
rect 26132 13019 26440 13028
rect 26528 12306 26556 13942
rect 26712 13870 26740 14334
rect 26896 14006 26924 14486
rect 26884 14000 26936 14006
rect 26884 13942 26936 13948
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26712 13530 26740 13806
rect 27252 13728 27304 13734
rect 27252 13670 27304 13676
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 27264 13394 27292 13670
rect 27252 13388 27304 13394
rect 27252 13330 27304 13336
rect 27356 12850 27384 14894
rect 27448 13258 27476 15370
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27540 15162 27568 15302
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27908 14532 27936 15574
rect 28092 15094 28120 15574
rect 28184 15570 28212 15846
rect 28276 15706 28304 16526
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 28080 15088 28132 15094
rect 28132 15036 28304 15042
rect 28080 15030 28304 15036
rect 28092 15014 28304 15030
rect 27908 14504 28028 14532
rect 27620 14476 27672 14482
rect 27620 14418 27672 14424
rect 27528 14340 27580 14346
rect 27528 14282 27580 14288
rect 27540 14074 27568 14282
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27632 13394 27660 14418
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27908 14074 27936 14282
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 28000 13802 28028 14504
rect 27988 13796 28040 13802
rect 27988 13738 28040 13744
rect 27620 13388 27672 13394
rect 27620 13330 27672 13336
rect 28172 13320 28224 13326
rect 28172 13262 28224 13268
rect 27436 13252 27488 13258
rect 27436 13194 27488 13200
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 26988 12434 27016 12582
rect 26804 12406 27016 12434
rect 26804 12306 26832 12406
rect 27448 12306 27476 13194
rect 27896 13184 27948 13190
rect 27896 13126 27948 13132
rect 27908 12850 27936 13126
rect 27896 12844 27948 12850
rect 27896 12786 27948 12792
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27988 12776 28040 12782
rect 27988 12718 28040 12724
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26792 12300 26844 12306
rect 26792 12242 26844 12248
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 25688 12232 25740 12238
rect 25608 12192 25688 12220
rect 24964 12158 25084 12186
rect 25688 12174 25740 12180
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24964 11898 24992 12038
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 25056 11694 25084 12158
rect 26132 11996 26440 12005
rect 26132 11994 26138 11996
rect 26194 11994 26218 11996
rect 26274 11994 26298 11996
rect 26354 11994 26378 11996
rect 26434 11994 26440 11996
rect 26194 11942 26196 11994
rect 26376 11942 26378 11994
rect 26132 11940 26138 11942
rect 26194 11940 26218 11942
rect 26274 11940 26298 11942
rect 26354 11940 26378 11942
rect 26434 11940 26440 11942
rect 26132 11931 26440 11940
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24320 10130 24348 11630
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24504 10266 24532 10610
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24400 10192 24452 10198
rect 24400 10134 24452 10140
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24412 9586 24440 10134
rect 25056 9994 25084 11630
rect 27540 11558 27568 12718
rect 28000 11830 28028 12718
rect 28184 12102 28212 13262
rect 28172 12096 28224 12102
rect 28172 12038 28224 12044
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 27528 11552 27580 11558
rect 27528 11494 27580 11500
rect 26516 11280 26568 11286
rect 26516 11222 26568 11228
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25700 10810 25728 11018
rect 26132 10908 26440 10917
rect 26132 10906 26138 10908
rect 26194 10906 26218 10908
rect 26274 10906 26298 10908
rect 26354 10906 26378 10908
rect 26434 10906 26440 10908
rect 26194 10854 26196 10906
rect 26376 10854 26378 10906
rect 26132 10852 26138 10854
rect 26194 10852 26218 10854
rect 26274 10852 26298 10854
rect 26354 10852 26378 10854
rect 26434 10852 26440 10854
rect 26132 10843 26440 10852
rect 25688 10804 25740 10810
rect 25688 10746 25740 10752
rect 25136 10736 25188 10742
rect 25136 10678 25188 10684
rect 25148 10062 25176 10678
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25044 9988 25096 9994
rect 25044 9930 25096 9936
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 25056 9518 25084 9930
rect 26132 9820 26440 9829
rect 26132 9818 26138 9820
rect 26194 9818 26218 9820
rect 26274 9818 26298 9820
rect 26354 9818 26378 9820
rect 26434 9818 26440 9820
rect 26194 9766 26196 9818
rect 26376 9766 26378 9818
rect 26132 9764 26138 9766
rect 26194 9764 26218 9766
rect 26274 9764 26298 9766
rect 26354 9764 26378 9766
rect 26434 9764 26440 9766
rect 26132 9755 26440 9764
rect 26528 9654 26556 11222
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26712 10810 26740 11086
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 27540 10606 27568 11494
rect 27620 11212 27672 11218
rect 28000 11200 28028 11766
rect 27672 11172 28028 11200
rect 27620 11154 27672 11160
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26620 10130 26648 10406
rect 26608 10124 26660 10130
rect 26608 10066 26660 10072
rect 26516 9648 26568 9654
rect 26516 9590 26568 9596
rect 27540 9518 27568 10542
rect 27632 10266 27660 11154
rect 28172 10532 28224 10538
rect 28172 10474 28224 10480
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26344 9042 26372 9318
rect 26332 9036 26384 9042
rect 26332 8978 26384 8984
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25608 8634 25636 8774
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 26068 8498 26096 8910
rect 26132 8732 26440 8741
rect 26132 8730 26138 8732
rect 26194 8730 26218 8732
rect 26274 8730 26298 8732
rect 26354 8730 26378 8732
rect 26434 8730 26440 8732
rect 26194 8678 26196 8730
rect 26376 8678 26378 8730
rect 26132 8676 26138 8678
rect 26194 8676 26218 8678
rect 26274 8676 26298 8678
rect 26354 8676 26378 8678
rect 26434 8676 26440 8678
rect 26132 8667 26440 8676
rect 26528 8498 26556 9318
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 26620 8566 26648 8842
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24412 7546 24440 7686
rect 24780 7546 24808 7686
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 22652 6248 22704 6254
rect 22572 6208 22652 6236
rect 22572 5914 22600 6208
rect 22652 6190 22704 6196
rect 23400 5914 23428 6598
rect 23584 6458 23612 6734
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22572 5166 22600 5850
rect 23768 5642 23796 7346
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 23756 5636 23808 5642
rect 23756 5578 23808 5584
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23492 5370 23520 5510
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 22560 5160 22612 5166
rect 22560 5102 22612 5108
rect 23676 4826 23704 5170
rect 23768 5098 23796 5578
rect 24136 5574 24164 6054
rect 24228 5778 24256 7346
rect 24872 7206 24900 8434
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24964 7954 24992 8366
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 26068 6866 26096 8434
rect 26132 7644 26440 7653
rect 26132 7642 26138 7644
rect 26194 7642 26218 7644
rect 26274 7642 26298 7644
rect 26354 7642 26378 7644
rect 26434 7642 26440 7644
rect 26194 7590 26196 7642
rect 26376 7590 26378 7642
rect 26132 7588 26138 7590
rect 26194 7588 26218 7590
rect 26274 7588 26298 7590
rect 26354 7588 26378 7590
rect 26434 7588 26440 7590
rect 26132 7579 26440 7588
rect 26056 6860 26108 6866
rect 26056 6802 26108 6808
rect 26620 6730 26648 8502
rect 27068 8288 27120 8294
rect 27068 8230 27120 8236
rect 27080 7954 27108 8230
rect 27172 7954 27200 9454
rect 27344 8832 27396 8838
rect 27396 8780 27568 8786
rect 27344 8774 27568 8780
rect 27356 8758 27568 8774
rect 27068 7948 27120 7954
rect 27068 7890 27120 7896
rect 27160 7948 27212 7954
rect 27160 7890 27212 7896
rect 26976 7744 27028 7750
rect 26976 7686 27028 7692
rect 27068 7744 27120 7750
rect 27068 7686 27120 7692
rect 26988 7546 27016 7686
rect 26976 7540 27028 7546
rect 26976 7482 27028 7488
rect 27080 7002 27108 7686
rect 27068 6996 27120 7002
rect 27068 6938 27120 6944
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 26608 6724 26660 6730
rect 26608 6666 26660 6672
rect 26132 6556 26440 6565
rect 26132 6554 26138 6556
rect 26194 6554 26218 6556
rect 26274 6554 26298 6556
rect 26354 6554 26378 6556
rect 26434 6554 26440 6556
rect 26194 6502 26196 6554
rect 26376 6502 26378 6554
rect 26132 6500 26138 6502
rect 26194 6500 26218 6502
rect 26274 6500 26298 6502
rect 26354 6500 26378 6502
rect 26434 6500 26440 6502
rect 26132 6491 26440 6500
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 24768 5840 24820 5846
rect 24768 5782 24820 5788
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 23756 5092 23808 5098
rect 23756 5034 23808 5040
rect 23664 4820 23716 4826
rect 23664 4762 23716 4768
rect 23768 4622 23796 5034
rect 23756 4616 23808 4622
rect 23756 4558 23808 4564
rect 23480 4548 23532 4554
rect 23480 4490 23532 4496
rect 23492 4282 23520 4490
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 24228 4146 24256 5714
rect 24780 5216 24808 5782
rect 24872 5370 24900 6054
rect 24964 5370 24992 6190
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 25332 5778 25360 6054
rect 25320 5772 25372 5778
rect 25320 5714 25372 5720
rect 25884 5370 25912 6190
rect 26620 5778 26648 6666
rect 26792 6180 26844 6186
rect 26792 6122 26844 6128
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26608 5772 26660 5778
rect 26608 5714 26660 5720
rect 26132 5468 26440 5477
rect 26132 5466 26138 5468
rect 26194 5466 26218 5468
rect 26274 5466 26298 5468
rect 26354 5466 26378 5468
rect 26434 5466 26440 5468
rect 26194 5414 26196 5466
rect 26376 5414 26378 5466
rect 26132 5412 26138 5414
rect 26194 5412 26218 5414
rect 26274 5412 26298 5414
rect 26354 5412 26378 5414
rect 26434 5412 26440 5414
rect 26132 5403 26440 5412
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 25872 5364 25924 5370
rect 25872 5306 25924 5312
rect 24860 5228 24912 5234
rect 24780 5188 24860 5216
rect 24860 5170 24912 5176
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 25056 4826 25084 5170
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25240 4758 25268 5170
rect 25228 4752 25280 4758
rect 25228 4694 25280 4700
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24412 4282 24440 4422
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 24504 4214 24532 4558
rect 25964 4480 26016 4486
rect 25964 4422 26016 4428
rect 25976 4282 26004 4422
rect 26132 4380 26440 4389
rect 26132 4378 26138 4380
rect 26194 4378 26218 4380
rect 26274 4378 26298 4380
rect 26354 4378 26378 4380
rect 26434 4378 26440 4380
rect 26194 4326 26196 4378
rect 26376 4326 26378 4378
rect 26132 4324 26138 4326
rect 26194 4324 26218 4326
rect 26274 4324 26298 4326
rect 26354 4324 26378 4326
rect 26434 4324 26440 4326
rect 26132 4315 26440 4324
rect 25964 4276 26016 4282
rect 25964 4218 26016 4224
rect 26620 4214 26648 5714
rect 26712 5642 26740 5850
rect 26700 5636 26752 5642
rect 26700 5578 26752 5584
rect 26804 5370 26832 6122
rect 26884 5568 26936 5574
rect 26884 5510 26936 5516
rect 26896 5370 26924 5510
rect 26792 5364 26844 5370
rect 26792 5306 26844 5312
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 26792 5092 26844 5098
rect 26792 5034 26844 5040
rect 26804 4214 26832 5034
rect 24492 4208 24544 4214
rect 24492 4150 24544 4156
rect 26608 4208 26660 4214
rect 26608 4150 26660 4156
rect 26792 4208 26844 4214
rect 26792 4150 26844 4156
rect 26988 4146 27016 6802
rect 27172 5234 27200 7890
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 27264 7546 27292 7822
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 27540 6866 27568 8758
rect 27632 8430 27660 10202
rect 28184 9994 28212 10474
rect 28276 10062 28304 15014
rect 28368 13938 28396 17190
rect 28816 17138 28868 17144
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 28920 16454 28948 17138
rect 28908 16448 28960 16454
rect 28908 16390 28960 16396
rect 28920 15910 28948 16390
rect 29012 16114 29040 17274
rect 29564 17270 29592 17478
rect 29552 17264 29604 17270
rect 29552 17206 29604 17212
rect 29276 17196 29328 17202
rect 29276 17138 29328 17144
rect 29288 16794 29316 17138
rect 29276 16788 29328 16794
rect 29276 16730 29328 16736
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29368 16108 29420 16114
rect 29368 16050 29420 16056
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 29012 15366 29040 16050
rect 29380 15484 29408 16050
rect 29460 15904 29512 15910
rect 29460 15846 29512 15852
rect 29472 15706 29500 15846
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 29552 15496 29604 15502
rect 29380 15456 29552 15484
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 29380 15026 29408 15456
rect 29748 15484 29776 15642
rect 29604 15456 29776 15484
rect 29552 15438 29604 15444
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 28632 14816 28684 14822
rect 28632 14758 28684 14764
rect 28644 13938 28672 14758
rect 29380 14618 29408 14962
rect 29368 14612 29420 14618
rect 29368 14554 29420 14560
rect 29368 14340 29420 14346
rect 29368 14282 29420 14288
rect 28356 13932 28408 13938
rect 28356 13874 28408 13880
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 28172 9988 28224 9994
rect 28172 9930 28224 9936
rect 27896 9716 27948 9722
rect 27896 9658 27948 9664
rect 27804 9580 27856 9586
rect 27804 9522 27856 9528
rect 27816 9178 27844 9522
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27908 8974 27936 9658
rect 28276 9042 28304 9998
rect 28368 9926 28396 13874
rect 28816 13796 28868 13802
rect 28816 13738 28868 13744
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28552 10470 28580 11086
rect 28724 11008 28776 11014
rect 28724 10950 28776 10956
rect 28736 10674 28764 10950
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28540 10464 28592 10470
rect 28540 10406 28592 10412
rect 28828 10062 28856 13738
rect 29380 12434 29408 14282
rect 29552 13252 29604 13258
rect 29552 13194 29604 13200
rect 29012 12406 29408 12434
rect 29012 12306 29040 12406
rect 29000 12300 29052 12306
rect 29000 12242 29052 12248
rect 29012 11762 29040 12242
rect 29564 12238 29592 13194
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29012 11218 29040 11698
rect 29564 11694 29592 12174
rect 29748 12170 29776 12378
rect 29736 12164 29788 12170
rect 29736 12106 29788 12112
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 29000 11212 29052 11218
rect 29000 11154 29052 11160
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 28356 9920 28408 9926
rect 28356 9862 28408 9868
rect 28264 9036 28316 9042
rect 28264 8978 28316 8984
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 27724 7886 27752 8298
rect 27908 7954 27936 8910
rect 28368 8838 28396 9862
rect 28828 9722 28856 9998
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 28356 8832 28408 8838
rect 28724 8832 28776 8838
rect 28408 8780 28488 8786
rect 28356 8774 28488 8780
rect 28724 8774 28776 8780
rect 28368 8758 28488 8774
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28368 8090 28396 8366
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28460 7954 28488 8758
rect 27896 7948 27948 7954
rect 27896 7890 27948 7896
rect 28448 7948 28500 7954
rect 28448 7890 28500 7896
rect 28736 7886 28764 8774
rect 29012 8634 29040 11154
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 27804 7812 27856 7818
rect 27804 7754 27856 7760
rect 27816 7002 27844 7754
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 27528 6860 27580 6866
rect 27528 6802 27580 6808
rect 27344 6452 27396 6458
rect 27540 6440 27568 6802
rect 27396 6412 27568 6440
rect 27344 6394 27396 6400
rect 27540 6322 27568 6412
rect 27816 6390 27844 6938
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27344 6248 27396 6254
rect 27396 6196 27660 6202
rect 27344 6190 27660 6196
rect 27356 6174 27660 6190
rect 27632 5778 27660 6174
rect 27896 6180 27948 6186
rect 27896 6122 27948 6128
rect 27804 6112 27856 6118
rect 27804 6054 27856 6060
rect 27620 5772 27672 5778
rect 27620 5714 27672 5720
rect 27816 5574 27844 6054
rect 27908 5642 27936 6122
rect 27896 5636 27948 5642
rect 27896 5578 27948 5584
rect 27804 5568 27856 5574
rect 27804 5510 27856 5516
rect 28552 5370 28580 7822
rect 28816 6724 28868 6730
rect 28816 6666 28868 6672
rect 28828 5778 28856 6666
rect 29564 6458 29592 9522
rect 29840 9382 29868 21286
rect 29932 21146 29960 21490
rect 29920 21140 29972 21146
rect 29920 21082 29972 21088
rect 30024 20482 30052 22510
rect 30329 22332 30637 22341
rect 30329 22330 30335 22332
rect 30391 22330 30415 22332
rect 30471 22330 30495 22332
rect 30551 22330 30575 22332
rect 30631 22330 30637 22332
rect 30391 22278 30393 22330
rect 30573 22278 30575 22330
rect 30329 22276 30335 22278
rect 30391 22276 30415 22278
rect 30471 22276 30495 22278
rect 30551 22276 30575 22278
rect 30631 22276 30637 22278
rect 30329 22267 30637 22276
rect 30668 22094 30696 23174
rect 30840 23044 30892 23050
rect 30840 22986 30892 22992
rect 30748 22976 30800 22982
rect 30748 22918 30800 22924
rect 30760 22778 30788 22918
rect 30748 22772 30800 22778
rect 30748 22714 30800 22720
rect 30576 22066 30696 22094
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 30300 21350 30328 21966
rect 30576 21350 30604 22066
rect 30656 21684 30708 21690
rect 30656 21626 30708 21632
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 30288 21344 30340 21350
rect 30288 21286 30340 21292
rect 30564 21344 30616 21350
rect 30564 21286 30616 21292
rect 30116 21078 30144 21286
rect 30329 21244 30637 21253
rect 30329 21242 30335 21244
rect 30391 21242 30415 21244
rect 30471 21242 30495 21244
rect 30551 21242 30575 21244
rect 30631 21242 30637 21244
rect 30391 21190 30393 21242
rect 30573 21190 30575 21242
rect 30329 21188 30335 21190
rect 30391 21188 30415 21190
rect 30471 21188 30495 21190
rect 30551 21188 30575 21190
rect 30631 21188 30637 21190
rect 30329 21179 30637 21188
rect 30104 21072 30156 21078
rect 30104 21014 30156 21020
rect 30668 21010 30696 21626
rect 30748 21480 30800 21486
rect 30748 21422 30800 21428
rect 30760 21146 30788 21422
rect 30852 21350 30880 22986
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30944 21146 30972 21490
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 30840 21140 30892 21146
rect 30840 21082 30892 21088
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 30656 21004 30708 21010
rect 30656 20946 30708 20952
rect 30748 20528 30800 20534
rect 30024 20454 30144 20482
rect 30748 20470 30800 20476
rect 30012 20324 30064 20330
rect 30012 20266 30064 20272
rect 29920 20256 29972 20262
rect 29920 20198 29972 20204
rect 29932 20058 29960 20198
rect 30024 20058 30052 20266
rect 29920 20052 29972 20058
rect 29920 19994 29972 20000
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 30012 17808 30064 17814
rect 30012 17750 30064 17756
rect 30024 16250 30052 17750
rect 30012 16244 30064 16250
rect 30012 16186 30064 16192
rect 30116 15094 30144 20454
rect 30329 20156 30637 20165
rect 30329 20154 30335 20156
rect 30391 20154 30415 20156
rect 30471 20154 30495 20156
rect 30551 20154 30575 20156
rect 30631 20154 30637 20156
rect 30391 20102 30393 20154
rect 30573 20102 30575 20154
rect 30329 20100 30335 20102
rect 30391 20100 30415 20102
rect 30471 20100 30495 20102
rect 30551 20100 30575 20102
rect 30631 20100 30637 20102
rect 30329 20091 30637 20100
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 30392 19446 30420 19654
rect 30380 19440 30432 19446
rect 30380 19382 30432 19388
rect 30656 19236 30708 19242
rect 30656 19178 30708 19184
rect 30196 19168 30248 19174
rect 30196 19110 30248 19116
rect 30208 18698 30236 19110
rect 30329 19068 30637 19077
rect 30329 19066 30335 19068
rect 30391 19066 30415 19068
rect 30471 19066 30495 19068
rect 30551 19066 30575 19068
rect 30631 19066 30637 19068
rect 30391 19014 30393 19066
rect 30573 19014 30575 19066
rect 30329 19012 30335 19014
rect 30391 19012 30415 19014
rect 30471 19012 30495 19014
rect 30551 19012 30575 19014
rect 30631 19012 30637 19014
rect 30329 19003 30637 19012
rect 30668 18766 30696 19178
rect 30564 18760 30616 18766
rect 30564 18702 30616 18708
rect 30656 18760 30708 18766
rect 30656 18702 30708 18708
rect 30196 18692 30248 18698
rect 30196 18634 30248 18640
rect 30576 18170 30604 18702
rect 30576 18142 30696 18170
rect 30329 17980 30637 17989
rect 30329 17978 30335 17980
rect 30391 17978 30415 17980
rect 30471 17978 30495 17980
rect 30551 17978 30575 17980
rect 30631 17978 30637 17980
rect 30391 17926 30393 17978
rect 30573 17926 30575 17978
rect 30329 17924 30335 17926
rect 30391 17924 30415 17926
rect 30471 17924 30495 17926
rect 30551 17924 30575 17926
rect 30631 17924 30637 17926
rect 30329 17915 30637 17924
rect 30668 17814 30696 18142
rect 30656 17808 30708 17814
rect 30656 17750 30708 17756
rect 30656 16992 30708 16998
rect 30656 16934 30708 16940
rect 30329 16892 30637 16901
rect 30329 16890 30335 16892
rect 30391 16890 30415 16892
rect 30471 16890 30495 16892
rect 30551 16890 30575 16892
rect 30631 16890 30637 16892
rect 30391 16838 30393 16890
rect 30573 16838 30575 16890
rect 30329 16836 30335 16838
rect 30391 16836 30415 16838
rect 30471 16836 30495 16838
rect 30551 16836 30575 16838
rect 30631 16836 30637 16838
rect 30329 16827 30637 16836
rect 30668 16658 30696 16934
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30329 15804 30637 15813
rect 30329 15802 30335 15804
rect 30391 15802 30415 15804
rect 30471 15802 30495 15804
rect 30551 15802 30575 15804
rect 30631 15802 30637 15804
rect 30391 15750 30393 15802
rect 30573 15750 30575 15802
rect 30329 15748 30335 15750
rect 30391 15748 30415 15750
rect 30471 15748 30495 15750
rect 30551 15748 30575 15750
rect 30631 15748 30637 15750
rect 30329 15739 30637 15748
rect 30104 15088 30156 15094
rect 30104 15030 30156 15036
rect 30760 14958 30788 20470
rect 30852 18970 30880 21082
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 30944 20602 30972 20810
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 31036 19446 31064 34575
rect 32404 34536 32456 34542
rect 32404 34478 32456 34484
rect 32416 32978 32444 34478
rect 32956 34400 33008 34406
rect 32956 34342 33008 34348
rect 33876 34400 33928 34406
rect 33876 34342 33928 34348
rect 32968 33930 32996 34342
rect 33888 34066 33916 34342
rect 33876 34060 33928 34066
rect 33876 34002 33928 34008
rect 32956 33924 33008 33930
rect 32956 33866 33008 33872
rect 32404 32972 32456 32978
rect 32404 32914 32456 32920
rect 32416 32434 32444 32914
rect 32968 32910 32996 33866
rect 34336 33856 34388 33862
rect 34336 33798 34388 33804
rect 32956 32904 33008 32910
rect 32956 32846 33008 32852
rect 32588 32768 32640 32774
rect 32588 32710 32640 32716
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 31116 29776 31168 29782
rect 31116 29718 31168 29724
rect 31128 29238 31156 29718
rect 31116 29232 31168 29238
rect 31116 29174 31168 29180
rect 32600 28218 32628 32710
rect 32588 28212 32640 28218
rect 32588 28154 32640 28160
rect 32968 27470 32996 32846
rect 34348 32842 34376 33798
rect 34526 33756 34834 33765
rect 34526 33754 34532 33756
rect 34588 33754 34612 33756
rect 34668 33754 34692 33756
rect 34748 33754 34772 33756
rect 34828 33754 34834 33756
rect 34588 33702 34590 33754
rect 34770 33702 34772 33754
rect 34526 33700 34532 33702
rect 34588 33700 34612 33702
rect 34668 33700 34692 33702
rect 34748 33700 34772 33702
rect 34828 33700 34834 33702
rect 34526 33691 34834 33700
rect 34336 32836 34388 32842
rect 34336 32778 34388 32784
rect 34526 32668 34834 32677
rect 34526 32666 34532 32668
rect 34588 32666 34612 32668
rect 34668 32666 34692 32668
rect 34748 32666 34772 32668
rect 34828 32666 34834 32668
rect 34588 32614 34590 32666
rect 34770 32614 34772 32666
rect 34526 32612 34532 32614
rect 34588 32612 34612 32614
rect 34668 32612 34692 32614
rect 34748 32612 34772 32614
rect 34828 32612 34834 32614
rect 34526 32603 34834 32612
rect 34526 31580 34834 31589
rect 34526 31578 34532 31580
rect 34588 31578 34612 31580
rect 34668 31578 34692 31580
rect 34748 31578 34772 31580
rect 34828 31578 34834 31580
rect 34588 31526 34590 31578
rect 34770 31526 34772 31578
rect 34526 31524 34532 31526
rect 34588 31524 34612 31526
rect 34668 31524 34692 31526
rect 34748 31524 34772 31526
rect 34828 31524 34834 31526
rect 34526 31515 34834 31524
rect 34526 30492 34834 30501
rect 34526 30490 34532 30492
rect 34588 30490 34612 30492
rect 34668 30490 34692 30492
rect 34748 30490 34772 30492
rect 34828 30490 34834 30492
rect 34588 30438 34590 30490
rect 34770 30438 34772 30490
rect 34526 30436 34532 30438
rect 34588 30436 34612 30438
rect 34668 30436 34692 30438
rect 34748 30436 34772 30438
rect 34828 30436 34834 30438
rect 34526 30427 34834 30436
rect 34526 29404 34834 29413
rect 34526 29402 34532 29404
rect 34588 29402 34612 29404
rect 34668 29402 34692 29404
rect 34748 29402 34772 29404
rect 34828 29402 34834 29404
rect 34588 29350 34590 29402
rect 34770 29350 34772 29402
rect 34526 29348 34532 29350
rect 34588 29348 34612 29350
rect 34668 29348 34692 29350
rect 34748 29348 34772 29350
rect 34828 29348 34834 29350
rect 34526 29339 34834 29348
rect 34526 28316 34834 28325
rect 34526 28314 34532 28316
rect 34588 28314 34612 28316
rect 34668 28314 34692 28316
rect 34748 28314 34772 28316
rect 34828 28314 34834 28316
rect 34588 28262 34590 28314
rect 34770 28262 34772 28314
rect 34526 28260 34532 28262
rect 34588 28260 34612 28262
rect 34668 28260 34692 28262
rect 34748 28260 34772 28262
rect 34828 28260 34834 28262
rect 34526 28251 34834 28260
rect 34796 28008 34848 28014
rect 34794 27976 34796 27985
rect 34848 27976 34850 27985
rect 34794 27911 34850 27920
rect 33600 27532 33652 27538
rect 33600 27474 33652 27480
rect 32956 27464 33008 27470
rect 32956 27406 33008 27412
rect 31760 27396 31812 27402
rect 31760 27338 31812 27344
rect 32772 27396 32824 27402
rect 32772 27338 32824 27344
rect 31772 27062 31800 27338
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32784 27282 32812 27338
rect 31760 27056 31812 27062
rect 31760 26998 31812 27004
rect 32496 26988 32548 26994
rect 32496 26930 32548 26936
rect 31576 26784 31628 26790
rect 31576 26726 31628 26732
rect 31588 26382 31616 26726
rect 31576 26376 31628 26382
rect 31576 26318 31628 26324
rect 31392 26308 31444 26314
rect 31392 26250 31444 26256
rect 31404 26194 31432 26250
rect 31404 26166 31524 26194
rect 31392 25356 31444 25362
rect 31392 25298 31444 25304
rect 31404 24818 31432 25298
rect 31300 24812 31352 24818
rect 31300 24754 31352 24760
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 31312 24070 31340 24754
rect 31300 24064 31352 24070
rect 31300 24006 31352 24012
rect 31300 23520 31352 23526
rect 31300 23462 31352 23468
rect 31312 23118 31340 23462
rect 31116 23112 31168 23118
rect 31300 23112 31352 23118
rect 31168 23060 31248 23066
rect 31116 23054 31248 23060
rect 31300 23054 31352 23060
rect 31128 23038 31248 23054
rect 31116 22976 31168 22982
rect 31116 22918 31168 22924
rect 31128 22778 31156 22918
rect 31116 22772 31168 22778
rect 31116 22714 31168 22720
rect 31220 21690 31248 23038
rect 31208 21684 31260 21690
rect 31208 21626 31260 21632
rect 31404 21622 31432 24754
rect 31496 23798 31524 26166
rect 31588 24698 31616 26318
rect 32312 26240 32364 26246
rect 32312 26182 32364 26188
rect 32324 25906 32352 26182
rect 32508 25906 32536 26930
rect 32600 26489 32628 27270
rect 32784 27254 32904 27282
rect 32586 26480 32642 26489
rect 32586 26415 32642 26424
rect 32876 26314 32904 27254
rect 33612 26586 33640 27474
rect 34526 27228 34834 27237
rect 34526 27226 34532 27228
rect 34588 27226 34612 27228
rect 34668 27226 34692 27228
rect 34748 27226 34772 27228
rect 34828 27226 34834 27228
rect 34588 27174 34590 27226
rect 34770 27174 34772 27226
rect 34526 27172 34532 27174
rect 34588 27172 34612 27174
rect 34668 27172 34692 27174
rect 34748 27172 34772 27174
rect 34828 27172 34834 27174
rect 34526 27163 34834 27172
rect 33600 26580 33652 26586
rect 33600 26522 33652 26528
rect 32864 26308 32916 26314
rect 32864 26250 32916 26256
rect 33048 26308 33100 26314
rect 33048 26250 33100 26256
rect 32876 26194 32904 26250
rect 32876 26166 32996 26194
rect 32312 25900 32364 25906
rect 32312 25842 32364 25848
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 31852 25288 31904 25294
rect 31852 25230 31904 25236
rect 31864 24954 31892 25230
rect 31852 24948 31904 24954
rect 31852 24890 31904 24896
rect 31588 24670 31708 24698
rect 31576 24608 31628 24614
rect 31576 24550 31628 24556
rect 31588 24410 31616 24550
rect 31576 24404 31628 24410
rect 31576 24346 31628 24352
rect 31484 23792 31536 23798
rect 31484 23734 31536 23740
rect 31496 21962 31524 23734
rect 31680 23526 31708 24670
rect 32128 24336 32180 24342
rect 32128 24278 32180 24284
rect 32140 23730 32168 24278
rect 32508 23746 32536 25842
rect 32600 25498 32628 25842
rect 32588 25492 32640 25498
rect 32588 25434 32640 25440
rect 32588 25220 32640 25226
rect 32588 25162 32640 25168
rect 32600 24410 32628 25162
rect 32588 24404 32640 24410
rect 32588 24346 32640 24352
rect 32968 24206 32996 26166
rect 33060 26042 33088 26250
rect 34526 26140 34834 26149
rect 34526 26138 34532 26140
rect 34588 26138 34612 26140
rect 34668 26138 34692 26140
rect 34748 26138 34772 26140
rect 34828 26138 34834 26140
rect 34588 26086 34590 26138
rect 34770 26086 34772 26138
rect 34526 26084 34532 26086
rect 34588 26084 34612 26086
rect 34668 26084 34692 26086
rect 34748 26084 34772 26086
rect 34828 26084 34834 26086
rect 34526 26075 34834 26084
rect 33048 26036 33100 26042
rect 33048 25978 33100 25984
rect 33416 25356 33468 25362
rect 33416 25298 33468 25304
rect 32956 24200 33008 24206
rect 32956 24142 33008 24148
rect 32508 23730 32628 23746
rect 32128 23724 32180 23730
rect 32508 23724 32640 23730
rect 32508 23718 32588 23724
rect 32128 23666 32180 23672
rect 32588 23666 32640 23672
rect 32772 23724 32824 23730
rect 32772 23666 32824 23672
rect 31668 23520 31720 23526
rect 31668 23462 31720 23468
rect 31680 22030 31708 23462
rect 32220 22568 32272 22574
rect 32220 22510 32272 22516
rect 32128 22500 32180 22506
rect 32128 22442 32180 22448
rect 32140 22094 32168 22442
rect 32232 22234 32260 22510
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 32508 22098 32536 22374
rect 32140 22066 32260 22094
rect 31668 22024 31720 22030
rect 31668 21966 31720 21972
rect 31484 21956 31536 21962
rect 31484 21898 31536 21904
rect 31392 21616 31444 21622
rect 31392 21558 31444 21564
rect 31116 21480 31168 21486
rect 31496 21434 31524 21898
rect 31116 21422 31168 21428
rect 31128 21146 31156 21422
rect 31220 21406 31524 21434
rect 31116 21140 31168 21146
rect 31116 21082 31168 21088
rect 31128 20534 31156 21082
rect 31116 20528 31168 20534
rect 31116 20470 31168 20476
rect 31024 19440 31076 19446
rect 31024 19382 31076 19388
rect 30840 18964 30892 18970
rect 30840 18906 30892 18912
rect 31220 18850 31248 21406
rect 31300 21344 31352 21350
rect 31300 21286 31352 21292
rect 31484 21344 31536 21350
rect 31484 21286 31536 21292
rect 30852 18822 31248 18850
rect 30852 15484 30880 18822
rect 31312 17762 31340 21286
rect 31392 20596 31444 20602
rect 31392 20538 31444 20544
rect 31404 19514 31432 20538
rect 31392 19508 31444 19514
rect 31392 19450 31444 19456
rect 31392 19304 31444 19310
rect 31392 19246 31444 19252
rect 31404 18630 31432 19246
rect 31392 18624 31444 18630
rect 31392 18566 31444 18572
rect 31496 17882 31524 21286
rect 32036 20936 32088 20942
rect 32036 20878 32088 20884
rect 31576 19168 31628 19174
rect 31576 19110 31628 19116
rect 31588 18766 31616 19110
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31576 18624 31628 18630
rect 31576 18566 31628 18572
rect 31588 18358 31616 18566
rect 31576 18352 31628 18358
rect 31576 18294 31628 18300
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 31116 17740 31168 17746
rect 31312 17734 31524 17762
rect 31588 17746 31616 18294
rect 31116 17682 31168 17688
rect 30932 17536 30984 17542
rect 30932 17478 30984 17484
rect 30944 17270 30972 17478
rect 30932 17264 30984 17270
rect 30932 17206 30984 17212
rect 31128 17202 31156 17682
rect 31024 17196 31076 17202
rect 31024 17138 31076 17144
rect 31116 17196 31168 17202
rect 31116 17138 31168 17144
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 30932 17060 30984 17066
rect 30932 17002 30984 17008
rect 30944 16590 30972 17002
rect 31036 16794 31064 17138
rect 31220 16794 31248 17138
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 31208 16788 31260 16794
rect 31208 16730 31260 16736
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 31024 16584 31076 16590
rect 31024 16526 31076 16532
rect 31036 16114 31064 16526
rect 31024 16108 31076 16114
rect 31024 16050 31076 16056
rect 31036 15978 31064 16050
rect 31024 15972 31076 15978
rect 31024 15914 31076 15920
rect 31036 15638 31064 15914
rect 31024 15632 31076 15638
rect 31024 15574 31076 15580
rect 30852 15456 31064 15484
rect 30932 15088 30984 15094
rect 30932 15030 30984 15036
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 30329 14716 30637 14725
rect 30329 14714 30335 14716
rect 30391 14714 30415 14716
rect 30471 14714 30495 14716
rect 30551 14714 30575 14716
rect 30631 14714 30637 14716
rect 30391 14662 30393 14714
rect 30573 14662 30575 14714
rect 30329 14660 30335 14662
rect 30391 14660 30415 14662
rect 30471 14660 30495 14662
rect 30551 14660 30575 14662
rect 30631 14660 30637 14662
rect 30329 14651 30637 14660
rect 30656 13932 30708 13938
rect 30656 13874 30708 13880
rect 30196 13728 30248 13734
rect 30196 13670 30248 13676
rect 30208 13258 30236 13670
rect 30329 13628 30637 13637
rect 30329 13626 30335 13628
rect 30391 13626 30415 13628
rect 30471 13626 30495 13628
rect 30551 13626 30575 13628
rect 30631 13626 30637 13628
rect 30391 13574 30393 13626
rect 30573 13574 30575 13626
rect 30329 13572 30335 13574
rect 30391 13572 30415 13574
rect 30471 13572 30495 13574
rect 30551 13572 30575 13574
rect 30631 13572 30637 13574
rect 30329 13563 30637 13572
rect 30668 13530 30696 13874
rect 30656 13524 30708 13530
rect 30656 13466 30708 13472
rect 30668 13258 30696 13466
rect 30196 13252 30248 13258
rect 30196 13194 30248 13200
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30329 12540 30637 12549
rect 30329 12538 30335 12540
rect 30391 12538 30415 12540
rect 30471 12538 30495 12540
rect 30551 12538 30575 12540
rect 30631 12538 30637 12540
rect 30391 12486 30393 12538
rect 30573 12486 30575 12538
rect 30329 12484 30335 12486
rect 30391 12484 30415 12486
rect 30471 12484 30495 12486
rect 30551 12484 30575 12486
rect 30631 12484 30637 12486
rect 30329 12475 30637 12484
rect 30944 12442 30972 15030
rect 30932 12436 30984 12442
rect 30932 12378 30984 12384
rect 31036 12374 31064 15456
rect 31312 15144 31340 16730
rect 31392 16448 31444 16454
rect 31392 16390 31444 16396
rect 31404 16114 31432 16390
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31404 15706 31432 16050
rect 31392 15700 31444 15706
rect 31392 15642 31444 15648
rect 31128 15116 31340 15144
rect 31128 14346 31156 15116
rect 31208 15020 31260 15026
rect 31208 14962 31260 14968
rect 31116 14340 31168 14346
rect 31116 14282 31168 14288
rect 31128 14074 31156 14282
rect 31116 14068 31168 14074
rect 31116 14010 31168 14016
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 31128 13394 31156 13874
rect 31116 13388 31168 13394
rect 31116 13330 31168 13336
rect 31220 12434 31248 14962
rect 31496 14822 31524 17734
rect 31576 17740 31628 17746
rect 31576 17682 31628 17688
rect 31680 17338 31708 18702
rect 31852 18624 31904 18630
rect 31852 18566 31904 18572
rect 31864 18290 31892 18566
rect 31852 18284 31904 18290
rect 31852 18226 31904 18232
rect 31852 17672 31904 17678
rect 31852 17614 31904 17620
rect 31668 17332 31720 17338
rect 31668 17274 31720 17280
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31588 15094 31616 17138
rect 31864 16454 31892 17614
rect 31852 16448 31904 16454
rect 31852 16390 31904 16396
rect 31576 15088 31628 15094
rect 31576 15030 31628 15036
rect 31668 15020 31720 15026
rect 31668 14962 31720 14968
rect 31300 14816 31352 14822
rect 31300 14758 31352 14764
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31312 13530 31340 14758
rect 31392 14408 31444 14414
rect 31444 14356 31524 14362
rect 31392 14350 31524 14356
rect 31404 14334 31524 14350
rect 31496 13938 31524 14334
rect 31576 14272 31628 14278
rect 31576 14214 31628 14220
rect 31588 13938 31616 14214
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 31576 13932 31628 13938
rect 31576 13874 31628 13880
rect 31496 13530 31524 13874
rect 31680 13682 31708 14962
rect 31864 14958 31892 16390
rect 31944 15360 31996 15366
rect 31944 15302 31996 15308
rect 31852 14952 31904 14958
rect 31852 14894 31904 14900
rect 31852 14816 31904 14822
rect 31852 14758 31904 14764
rect 31864 14464 31892 14758
rect 31956 14550 31984 15302
rect 31944 14544 31996 14550
rect 31944 14486 31996 14492
rect 31588 13654 31708 13682
rect 31772 14436 31892 14464
rect 31300 13524 31352 13530
rect 31300 13466 31352 13472
rect 31484 13524 31536 13530
rect 31484 13466 31536 13472
rect 31300 12980 31352 12986
rect 31300 12922 31352 12928
rect 31128 12406 31248 12434
rect 31024 12368 31076 12374
rect 31024 12310 31076 12316
rect 30012 12232 30064 12238
rect 30012 12174 30064 12180
rect 30024 11558 30052 12174
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 30564 12096 30616 12102
rect 30564 12038 30616 12044
rect 30208 11830 30236 12038
rect 30576 11898 30604 12038
rect 30564 11892 30616 11898
rect 30564 11834 30616 11840
rect 30196 11824 30248 11830
rect 30196 11766 30248 11772
rect 30012 11552 30064 11558
rect 30012 11494 30064 11500
rect 30024 11286 30052 11494
rect 30329 11452 30637 11461
rect 30329 11450 30335 11452
rect 30391 11450 30415 11452
rect 30471 11450 30495 11452
rect 30551 11450 30575 11452
rect 30631 11450 30637 11452
rect 30391 11398 30393 11450
rect 30573 11398 30575 11450
rect 30329 11396 30335 11398
rect 30391 11396 30415 11398
rect 30471 11396 30495 11398
rect 30551 11396 30575 11398
rect 30631 11396 30637 11398
rect 30329 11387 30637 11396
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30012 11280 30064 11286
rect 30012 11222 30064 11228
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30300 10742 30328 11086
rect 30288 10736 30340 10742
rect 30288 10678 30340 10684
rect 30668 10538 30696 11290
rect 30932 11212 30984 11218
rect 30932 11154 30984 11160
rect 30944 10742 30972 11154
rect 30932 10736 30984 10742
rect 30932 10678 30984 10684
rect 30656 10532 30708 10538
rect 30656 10474 30708 10480
rect 30329 10364 30637 10373
rect 30329 10362 30335 10364
rect 30391 10362 30415 10364
rect 30471 10362 30495 10364
rect 30551 10362 30575 10364
rect 30631 10362 30637 10364
rect 30391 10310 30393 10362
rect 30573 10310 30575 10362
rect 30329 10308 30335 10310
rect 30391 10308 30415 10310
rect 30471 10308 30495 10310
rect 30551 10308 30575 10310
rect 30631 10308 30637 10310
rect 30329 10299 30637 10308
rect 31036 10198 31064 12310
rect 31024 10192 31076 10198
rect 31024 10134 31076 10140
rect 30840 9580 30892 9586
rect 30840 9522 30892 9528
rect 29920 9512 29972 9518
rect 29920 9454 29972 9460
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29828 8900 29880 8906
rect 29828 8842 29880 8848
rect 29840 8634 29868 8842
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 29736 7812 29788 7818
rect 29736 7754 29788 7760
rect 29644 6656 29696 6662
rect 29644 6598 29696 6604
rect 29552 6452 29604 6458
rect 29552 6394 29604 6400
rect 29368 6180 29420 6186
rect 29368 6122 29420 6128
rect 29380 5914 29408 6122
rect 29656 5914 29684 6598
rect 29748 6458 29776 7754
rect 29840 7206 29868 8570
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 29932 6866 29960 9454
rect 30329 9276 30637 9285
rect 30329 9274 30335 9276
rect 30391 9274 30415 9276
rect 30471 9274 30495 9276
rect 30551 9274 30575 9276
rect 30631 9274 30637 9276
rect 30391 9222 30393 9274
rect 30573 9222 30575 9274
rect 30329 9220 30335 9222
rect 30391 9220 30415 9222
rect 30471 9220 30495 9222
rect 30551 9220 30575 9222
rect 30631 9220 30637 9222
rect 30329 9211 30637 9220
rect 30852 9178 30880 9522
rect 31036 9330 31064 10134
rect 31128 9450 31156 12406
rect 31312 12322 31340 12922
rect 31484 12844 31536 12850
rect 31484 12786 31536 12792
rect 31392 12436 31444 12442
rect 31392 12378 31444 12384
rect 31220 12294 31340 12322
rect 31220 12238 31248 12294
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 31312 11830 31340 12174
rect 31300 11824 31352 11830
rect 31300 11766 31352 11772
rect 31208 11552 31260 11558
rect 31208 11494 31260 11500
rect 31220 11014 31248 11494
rect 31312 11354 31340 11766
rect 31404 11626 31432 12378
rect 31496 12288 31524 12786
rect 31588 12442 31616 13654
rect 31668 13524 31720 13530
rect 31668 13466 31720 13472
rect 31576 12436 31628 12442
rect 31576 12378 31628 12384
rect 31496 12260 31616 12288
rect 31484 12164 31536 12170
rect 31484 12106 31536 12112
rect 31392 11620 31444 11626
rect 31392 11562 31444 11568
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31312 11150 31340 11290
rect 31300 11144 31352 11150
rect 31300 11086 31352 11092
rect 31208 11008 31260 11014
rect 31208 10950 31260 10956
rect 31220 10470 31248 10950
rect 31300 10532 31352 10538
rect 31300 10474 31352 10480
rect 31208 10464 31260 10470
rect 31208 10406 31260 10412
rect 31116 9444 31168 9450
rect 31116 9386 31168 9392
rect 31220 9382 31248 10406
rect 31312 10266 31340 10474
rect 31300 10260 31352 10266
rect 31300 10202 31352 10208
rect 31300 9512 31352 9518
rect 31300 9454 31352 9460
rect 31208 9376 31260 9382
rect 31036 9302 31156 9330
rect 31208 9318 31260 9324
rect 30840 9172 30892 9178
rect 30840 9114 30892 9120
rect 30852 8498 30880 9114
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 30329 8188 30637 8197
rect 30329 8186 30335 8188
rect 30391 8186 30415 8188
rect 30471 8186 30495 8188
rect 30551 8186 30575 8188
rect 30631 8186 30637 8188
rect 30391 8134 30393 8186
rect 30573 8134 30575 8186
rect 30329 8132 30335 8134
rect 30391 8132 30415 8134
rect 30471 8132 30495 8134
rect 30551 8132 30575 8134
rect 30631 8132 30637 8134
rect 30329 8123 30637 8132
rect 30840 7744 30892 7750
rect 30840 7686 30892 7692
rect 30852 7478 30880 7686
rect 30840 7472 30892 7478
rect 30840 7414 30892 7420
rect 30329 7100 30637 7109
rect 30329 7098 30335 7100
rect 30391 7098 30415 7100
rect 30471 7098 30495 7100
rect 30551 7098 30575 7100
rect 30631 7098 30637 7100
rect 30391 7046 30393 7098
rect 30573 7046 30575 7098
rect 30329 7044 30335 7046
rect 30391 7044 30415 7046
rect 30471 7044 30495 7046
rect 30551 7044 30575 7046
rect 30631 7044 30637 7046
rect 30329 7035 30637 7044
rect 29920 6860 29972 6866
rect 29920 6802 29972 6808
rect 30852 6798 30880 7414
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30196 6724 30248 6730
rect 30196 6666 30248 6672
rect 29736 6452 29788 6458
rect 29736 6394 29788 6400
rect 30208 6322 30236 6666
rect 30760 6458 30788 6734
rect 30944 6730 30972 7142
rect 31036 7002 31064 8366
rect 31024 6996 31076 7002
rect 31024 6938 31076 6944
rect 30932 6724 30984 6730
rect 30932 6666 30984 6672
rect 30748 6452 30800 6458
rect 30748 6394 30800 6400
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 30196 6316 30248 6322
rect 30380 6316 30432 6322
rect 30196 6258 30248 6264
rect 30300 6276 30380 6304
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29840 5914 29868 6190
rect 29368 5908 29420 5914
rect 29368 5850 29420 5856
rect 29644 5908 29696 5914
rect 29644 5850 29696 5856
rect 29828 5908 29880 5914
rect 29828 5850 29880 5856
rect 28816 5772 28868 5778
rect 28816 5714 28868 5720
rect 28540 5364 28592 5370
rect 28540 5306 28592 5312
rect 27160 5228 27212 5234
rect 27160 5170 27212 5176
rect 27172 4758 27200 5170
rect 28828 5166 28856 5714
rect 28908 5228 28960 5234
rect 28908 5170 28960 5176
rect 28816 5160 28868 5166
rect 28816 5102 28868 5108
rect 27344 5092 27396 5098
rect 27344 5034 27396 5040
rect 27356 4826 27384 5034
rect 28920 4826 28948 5170
rect 29368 5160 29420 5166
rect 29368 5102 29420 5108
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 28908 4820 28960 4826
rect 28908 4762 28960 4768
rect 27160 4752 27212 4758
rect 27160 4694 27212 4700
rect 28920 4282 28948 4762
rect 29380 4758 29408 5102
rect 29932 5098 29960 6258
rect 30104 6248 30156 6254
rect 30104 6190 30156 6196
rect 29920 5092 29972 5098
rect 29920 5034 29972 5040
rect 30116 4826 30144 6190
rect 30300 6168 30328 6276
rect 30380 6258 30432 6264
rect 30208 6140 30328 6168
rect 30208 5914 30236 6140
rect 30329 6012 30637 6021
rect 30329 6010 30335 6012
rect 30391 6010 30415 6012
rect 30471 6010 30495 6012
rect 30551 6010 30575 6012
rect 30631 6010 30637 6012
rect 30391 5958 30393 6010
rect 30573 5958 30575 6010
rect 30329 5956 30335 5958
rect 30391 5956 30415 5958
rect 30471 5956 30495 5958
rect 30551 5956 30575 5958
rect 30631 5956 30637 5958
rect 30329 5947 30637 5956
rect 30196 5908 30248 5914
rect 30196 5850 30248 5856
rect 30208 5166 30236 5850
rect 31128 5574 31156 9302
rect 31312 7818 31340 9454
rect 31496 9450 31524 12106
rect 31588 11354 31616 12260
rect 31680 12238 31708 13466
rect 31772 13308 31800 14436
rect 31852 14340 31904 14346
rect 31852 14282 31904 14288
rect 31944 14340 31996 14346
rect 31944 14282 31996 14288
rect 31864 13734 31892 14282
rect 31956 14074 31984 14282
rect 31944 14068 31996 14074
rect 31944 14010 31996 14016
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 31852 13728 31904 13734
rect 31852 13670 31904 13676
rect 31772 13280 31892 13308
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31772 12442 31800 12786
rect 31760 12436 31812 12442
rect 31760 12378 31812 12384
rect 31772 12238 31800 12378
rect 31668 12232 31720 12238
rect 31668 12174 31720 12180
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31668 11552 31720 11558
rect 31668 11494 31720 11500
rect 31576 11348 31628 11354
rect 31576 11290 31628 11296
rect 31680 11150 31708 11494
rect 31760 11280 31812 11286
rect 31760 11222 31812 11228
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31772 10674 31800 11222
rect 31576 10668 31628 10674
rect 31576 10610 31628 10616
rect 31760 10668 31812 10674
rect 31760 10610 31812 10616
rect 31588 10198 31616 10610
rect 31772 10470 31800 10610
rect 31760 10464 31812 10470
rect 31760 10406 31812 10412
rect 31576 10192 31628 10198
rect 31576 10134 31628 10140
rect 31668 9580 31720 9586
rect 31668 9522 31720 9528
rect 31484 9444 31536 9450
rect 31484 9386 31536 9392
rect 31576 9104 31628 9110
rect 31576 9046 31628 9052
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 31404 8498 31432 8774
rect 31496 8566 31524 8842
rect 31484 8560 31536 8566
rect 31484 8502 31536 8508
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 31404 8090 31432 8434
rect 31496 8294 31524 8502
rect 31588 8430 31616 9046
rect 31680 9042 31708 9522
rect 31760 9172 31812 9178
rect 31760 9114 31812 9120
rect 31668 9036 31720 9042
rect 31668 8978 31720 8984
rect 31772 8838 31800 9114
rect 31760 8832 31812 8838
rect 31760 8774 31812 8780
rect 31576 8424 31628 8430
rect 31576 8366 31628 8372
rect 31484 8288 31536 8294
rect 31484 8230 31536 8236
rect 31392 8084 31444 8090
rect 31392 8026 31444 8032
rect 31300 7812 31352 7818
rect 31300 7754 31352 7760
rect 31496 7410 31524 8230
rect 31484 7404 31536 7410
rect 31484 7346 31536 7352
rect 31576 7336 31628 7342
rect 31576 7278 31628 7284
rect 31484 7200 31536 7206
rect 31484 7142 31536 7148
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 31116 5568 31168 5574
rect 31116 5510 31168 5516
rect 30392 5370 30420 5510
rect 31496 5370 31524 7142
rect 31588 6798 31616 7278
rect 31576 6792 31628 6798
rect 31576 6734 31628 6740
rect 31772 6458 31800 8774
rect 31864 7546 31892 13280
rect 31956 12986 31984 13874
rect 31944 12980 31996 12986
rect 31944 12922 31996 12928
rect 32048 12866 32076 20878
rect 32128 19236 32180 19242
rect 32128 19178 32180 19184
rect 32140 17678 32168 19178
rect 32232 18766 32260 22066
rect 32496 22092 32548 22098
rect 32496 22034 32548 22040
rect 32600 21894 32628 23666
rect 32680 22024 32732 22030
rect 32680 21966 32732 21972
rect 32588 21888 32640 21894
rect 32588 21830 32640 21836
rect 32600 20942 32628 21830
rect 32588 20936 32640 20942
rect 32588 20878 32640 20884
rect 32692 20602 32720 21966
rect 32784 21894 32812 23666
rect 32968 22642 32996 24142
rect 32956 22636 33008 22642
rect 32956 22578 33008 22584
rect 32772 21888 32824 21894
rect 32772 21830 32824 21836
rect 32968 20942 32996 22578
rect 33428 22166 33456 25298
rect 34526 25052 34834 25061
rect 34526 25050 34532 25052
rect 34588 25050 34612 25052
rect 34668 25050 34692 25052
rect 34748 25050 34772 25052
rect 34828 25050 34834 25052
rect 34588 24998 34590 25050
rect 34770 24998 34772 25050
rect 34526 24996 34532 24998
rect 34588 24996 34612 24998
rect 34668 24996 34692 24998
rect 34748 24996 34772 24998
rect 34828 24996 34834 24998
rect 34526 24987 34834 24996
rect 34336 24200 34388 24206
rect 34336 24142 34388 24148
rect 34060 24132 34112 24138
rect 34060 24074 34112 24080
rect 34072 23866 34100 24074
rect 34060 23860 34112 23866
rect 34060 23802 34112 23808
rect 34348 22438 34376 24142
rect 34526 23964 34834 23973
rect 34526 23962 34532 23964
rect 34588 23962 34612 23964
rect 34668 23962 34692 23964
rect 34748 23962 34772 23964
rect 34828 23962 34834 23964
rect 34588 23910 34590 23962
rect 34770 23910 34772 23962
rect 34526 23908 34532 23910
rect 34588 23908 34612 23910
rect 34668 23908 34692 23910
rect 34748 23908 34772 23910
rect 34828 23908 34834 23910
rect 34526 23899 34834 23908
rect 34526 22876 34834 22885
rect 34526 22874 34532 22876
rect 34588 22874 34612 22876
rect 34668 22874 34692 22876
rect 34748 22874 34772 22876
rect 34828 22874 34834 22876
rect 34588 22822 34590 22874
rect 34770 22822 34772 22874
rect 34526 22820 34532 22822
rect 34588 22820 34612 22822
rect 34668 22820 34692 22822
rect 34748 22820 34772 22822
rect 34828 22820 34834 22822
rect 34526 22811 34834 22820
rect 34336 22432 34388 22438
rect 34336 22374 34388 22380
rect 33416 22160 33468 22166
rect 33416 22102 33468 22108
rect 33232 21888 33284 21894
rect 33232 21830 33284 21836
rect 33244 21690 33272 21830
rect 33232 21684 33284 21690
rect 33232 21626 33284 21632
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 32680 20596 32732 20602
rect 32680 20538 32732 20544
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 33060 19514 33088 20402
rect 33428 20398 33456 22102
rect 34348 21010 34376 22374
rect 34526 21788 34834 21797
rect 34526 21786 34532 21788
rect 34588 21786 34612 21788
rect 34668 21786 34692 21788
rect 34748 21786 34772 21788
rect 34828 21786 34834 21788
rect 34588 21734 34590 21786
rect 34770 21734 34772 21786
rect 34526 21732 34532 21734
rect 34588 21732 34612 21734
rect 34668 21732 34692 21734
rect 34748 21732 34772 21734
rect 34828 21732 34834 21734
rect 34526 21723 34834 21732
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34808 21185 34836 21490
rect 34794 21176 34850 21185
rect 34794 21111 34850 21120
rect 34336 21004 34388 21010
rect 34336 20946 34388 20952
rect 34526 20700 34834 20709
rect 34526 20698 34532 20700
rect 34588 20698 34612 20700
rect 34668 20698 34692 20700
rect 34748 20698 34772 20700
rect 34828 20698 34834 20700
rect 34588 20646 34590 20698
rect 34770 20646 34772 20698
rect 34526 20644 34532 20646
rect 34588 20644 34612 20646
rect 34668 20644 34692 20646
rect 34748 20644 34772 20646
rect 34828 20644 34834 20646
rect 34526 20635 34834 20644
rect 33416 20392 33468 20398
rect 33416 20334 33468 20340
rect 33048 19508 33100 19514
rect 33048 19450 33100 19456
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 32312 18896 32364 18902
rect 32508 18850 32536 19314
rect 32680 19304 32732 19310
rect 32680 19246 32732 19252
rect 32692 18970 32720 19246
rect 32680 18964 32732 18970
rect 32680 18906 32732 18912
rect 32364 18844 32536 18850
rect 32312 18838 32536 18844
rect 32324 18822 32536 18838
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32232 18086 32260 18702
rect 32220 18080 32272 18086
rect 32220 18022 32272 18028
rect 32508 17678 32536 18822
rect 32956 18760 33008 18766
rect 32956 18702 33008 18708
rect 32680 18692 32732 18698
rect 32680 18634 32732 18640
rect 32588 18284 32640 18290
rect 32588 18226 32640 18232
rect 32600 17882 32628 18226
rect 32588 17876 32640 17882
rect 32588 17818 32640 17824
rect 32128 17672 32180 17678
rect 32128 17614 32180 17620
rect 32496 17672 32548 17678
rect 32496 17614 32548 17620
rect 32220 17536 32272 17542
rect 32220 17478 32272 17484
rect 32232 16114 32260 17478
rect 32692 17338 32720 18634
rect 32864 18624 32916 18630
rect 32864 18566 32916 18572
rect 32876 18426 32904 18566
rect 32864 18420 32916 18426
rect 32864 18362 32916 18368
rect 32968 18358 32996 18702
rect 32956 18352 33008 18358
rect 32956 18294 33008 18300
rect 32864 18080 32916 18086
rect 32864 18022 32916 18028
rect 32772 17604 32824 17610
rect 32772 17546 32824 17552
rect 32680 17332 32732 17338
rect 32680 17274 32732 17280
rect 32784 17202 32812 17546
rect 32772 17196 32824 17202
rect 32772 17138 32824 17144
rect 32772 16516 32824 16522
rect 32772 16458 32824 16464
rect 32588 16448 32640 16454
rect 32588 16390 32640 16396
rect 32600 16250 32628 16390
rect 32588 16244 32640 16250
rect 32588 16186 32640 16192
rect 32220 16108 32272 16114
rect 32220 16050 32272 16056
rect 32232 14618 32260 16050
rect 32784 15978 32812 16458
rect 32876 16182 32904 18022
rect 33428 17338 33456 20334
rect 34526 19612 34834 19621
rect 34526 19610 34532 19612
rect 34588 19610 34612 19612
rect 34668 19610 34692 19612
rect 34748 19610 34772 19612
rect 34828 19610 34834 19612
rect 34588 19558 34590 19610
rect 34770 19558 34772 19610
rect 34526 19556 34532 19558
rect 34588 19556 34612 19558
rect 34668 19556 34692 19558
rect 34748 19556 34772 19558
rect 34828 19556 34834 19558
rect 34526 19547 34834 19556
rect 34526 18524 34834 18533
rect 34526 18522 34532 18524
rect 34588 18522 34612 18524
rect 34668 18522 34692 18524
rect 34748 18522 34772 18524
rect 34828 18522 34834 18524
rect 34588 18470 34590 18522
rect 34770 18470 34772 18522
rect 34526 18468 34532 18470
rect 34588 18468 34612 18470
rect 34668 18468 34692 18470
rect 34748 18468 34772 18470
rect 34828 18468 34834 18470
rect 34526 18459 34834 18468
rect 33508 17536 33560 17542
rect 33508 17478 33560 17484
rect 33416 17332 33468 17338
rect 33416 17274 33468 17280
rect 32956 17196 33008 17202
rect 32956 17138 33008 17144
rect 33140 17196 33192 17202
rect 33140 17138 33192 17144
rect 32968 16454 32996 17138
rect 33152 16794 33180 17138
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 33152 16590 33180 16730
rect 33140 16584 33192 16590
rect 33140 16526 33192 16532
rect 32956 16448 33008 16454
rect 32956 16390 33008 16396
rect 32864 16176 32916 16182
rect 32864 16118 32916 16124
rect 32772 15972 32824 15978
rect 32772 15914 32824 15920
rect 32876 15026 32904 16118
rect 32968 15910 32996 16390
rect 32956 15904 33008 15910
rect 32956 15846 33008 15852
rect 33428 15366 33456 17274
rect 33520 16794 33548 17478
rect 34526 17436 34834 17445
rect 34526 17434 34532 17436
rect 34588 17434 34612 17436
rect 34668 17434 34692 17436
rect 34748 17434 34772 17436
rect 34828 17434 34834 17436
rect 34588 17382 34590 17434
rect 34770 17382 34772 17434
rect 34526 17380 34532 17382
rect 34588 17380 34612 17382
rect 34668 17380 34692 17382
rect 34748 17380 34772 17382
rect 34828 17380 34834 17382
rect 34526 17371 34834 17380
rect 33692 17196 33744 17202
rect 33692 17138 33744 17144
rect 33704 16794 33732 17138
rect 33508 16788 33560 16794
rect 33508 16730 33560 16736
rect 33692 16788 33744 16794
rect 33692 16730 33744 16736
rect 34526 16348 34834 16357
rect 34526 16346 34532 16348
rect 34588 16346 34612 16348
rect 34668 16346 34692 16348
rect 34748 16346 34772 16348
rect 34828 16346 34834 16348
rect 34588 16294 34590 16346
rect 34770 16294 34772 16346
rect 34526 16292 34532 16294
rect 34588 16292 34612 16294
rect 34668 16292 34692 16294
rect 34748 16292 34772 16294
rect 34828 16292 34834 16294
rect 34526 16283 34834 16292
rect 33416 15360 33468 15366
rect 33416 15302 33468 15308
rect 33428 15094 33456 15302
rect 34526 15260 34834 15269
rect 34526 15258 34532 15260
rect 34588 15258 34612 15260
rect 34668 15258 34692 15260
rect 34748 15258 34772 15260
rect 34828 15258 34834 15260
rect 34588 15206 34590 15258
rect 34770 15206 34772 15258
rect 34526 15204 34532 15206
rect 34588 15204 34612 15206
rect 34668 15204 34692 15206
rect 34748 15204 34772 15206
rect 34828 15204 34834 15206
rect 34526 15195 34834 15204
rect 33416 15088 33468 15094
rect 33416 15030 33468 15036
rect 32864 15020 32916 15026
rect 32864 14962 32916 14968
rect 32220 14612 32272 14618
rect 32220 14554 32272 14560
rect 32876 14414 32904 14962
rect 32864 14408 32916 14414
rect 32864 14350 32916 14356
rect 32220 14272 32272 14278
rect 32220 14214 32272 14220
rect 32312 14272 32364 14278
rect 32312 14214 32364 14220
rect 32232 13938 32260 14214
rect 32324 14006 32352 14214
rect 32312 14000 32364 14006
rect 32312 13942 32364 13948
rect 32220 13932 32272 13938
rect 32220 13874 32272 13880
rect 32680 13184 32732 13190
rect 32680 13126 32732 13132
rect 31956 12838 32076 12866
rect 32692 12850 32720 13126
rect 32680 12844 32732 12850
rect 31956 11626 31984 12838
rect 32680 12786 32732 12792
rect 33428 12782 33456 15030
rect 34152 14816 34204 14822
rect 34152 14758 34204 14764
rect 34164 14414 34192 14758
rect 34704 14544 34756 14550
rect 34704 14486 34756 14492
rect 34152 14408 34204 14414
rect 34716 14385 34744 14486
rect 34152 14350 34204 14356
rect 34702 14376 34758 14385
rect 34702 14311 34758 14320
rect 34526 14172 34834 14181
rect 34526 14170 34532 14172
rect 34588 14170 34612 14172
rect 34668 14170 34692 14172
rect 34748 14170 34772 14172
rect 34828 14170 34834 14172
rect 34588 14118 34590 14170
rect 34770 14118 34772 14170
rect 34526 14116 34532 14118
rect 34588 14116 34612 14118
rect 34668 14116 34692 14118
rect 34748 14116 34772 14118
rect 34828 14116 34834 14118
rect 34526 14107 34834 14116
rect 34526 13084 34834 13093
rect 34526 13082 34532 13084
rect 34588 13082 34612 13084
rect 34668 13082 34692 13084
rect 34748 13082 34772 13084
rect 34828 13082 34834 13084
rect 34588 13030 34590 13082
rect 34770 13030 34772 13082
rect 34526 13028 34532 13030
rect 34588 13028 34612 13030
rect 34668 13028 34692 13030
rect 34748 13028 34772 13030
rect 34828 13028 34834 13030
rect 34526 13019 34834 13028
rect 33876 12844 33928 12850
rect 33876 12786 33928 12792
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 34152 12844 34204 12850
rect 34152 12786 34204 12792
rect 33416 12776 33468 12782
rect 33416 12718 33468 12724
rect 33692 12776 33744 12782
rect 33692 12718 33744 12724
rect 32036 12640 32088 12646
rect 32036 12582 32088 12588
rect 32048 12170 32076 12582
rect 33704 12434 33732 12718
rect 33888 12442 33916 12786
rect 33876 12436 33928 12442
rect 33704 12406 33824 12434
rect 32036 12164 32088 12170
rect 32036 12106 32088 12112
rect 31944 11620 31996 11626
rect 31944 11562 31996 11568
rect 32496 11552 32548 11558
rect 32496 11494 32548 11500
rect 32036 11212 32088 11218
rect 32036 11154 32088 11160
rect 31944 10464 31996 10470
rect 31944 10406 31996 10412
rect 31852 7540 31904 7546
rect 31852 7482 31904 7488
rect 31956 6914 31984 10406
rect 32048 9178 32076 11154
rect 32508 10674 32536 11494
rect 33048 11008 33100 11014
rect 33048 10950 33100 10956
rect 33060 10810 33088 10950
rect 33048 10804 33100 10810
rect 33048 10746 33100 10752
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 33048 10668 33100 10674
rect 33048 10610 33100 10616
rect 32220 10600 32272 10606
rect 32220 10542 32272 10548
rect 32128 10464 32180 10470
rect 32128 10406 32180 10412
rect 32140 10266 32168 10406
rect 32128 10260 32180 10266
rect 32128 10202 32180 10208
rect 32232 10198 32260 10542
rect 32220 10192 32272 10198
rect 32220 10134 32272 10140
rect 32220 9988 32272 9994
rect 32220 9930 32272 9936
rect 32232 9178 32260 9930
rect 32036 9172 32088 9178
rect 32036 9114 32088 9120
rect 32220 9172 32272 9178
rect 32220 9114 32272 9120
rect 32404 9036 32456 9042
rect 32404 8978 32456 8984
rect 31864 6886 31984 6914
rect 31760 6452 31812 6458
rect 31760 6394 31812 6400
rect 31772 5914 31800 6394
rect 31760 5908 31812 5914
rect 31760 5850 31812 5856
rect 31864 5710 31892 6886
rect 32416 6866 32444 8978
rect 32404 6860 32456 6866
rect 32404 6802 32456 6808
rect 32508 6390 32536 10610
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 32968 8566 32996 9862
rect 33060 9042 33088 10610
rect 33796 10606 33824 12406
rect 33876 12378 33928 12384
rect 33784 10600 33836 10606
rect 33784 10542 33836 10548
rect 33888 10538 33916 12378
rect 33980 12102 34008 12786
rect 34164 12442 34192 12786
rect 34152 12436 34204 12442
rect 34152 12378 34204 12384
rect 33968 12096 34020 12102
rect 33968 12038 34020 12044
rect 34526 11996 34834 12005
rect 34526 11994 34532 11996
rect 34588 11994 34612 11996
rect 34668 11994 34692 11996
rect 34748 11994 34772 11996
rect 34828 11994 34834 11996
rect 34588 11942 34590 11994
rect 34770 11942 34772 11994
rect 34526 11940 34532 11942
rect 34588 11940 34612 11942
rect 34668 11940 34692 11942
rect 34748 11940 34772 11942
rect 34828 11940 34834 11942
rect 34526 11931 34834 11940
rect 34526 10908 34834 10917
rect 34526 10906 34532 10908
rect 34588 10906 34612 10908
rect 34668 10906 34692 10908
rect 34748 10906 34772 10908
rect 34828 10906 34834 10908
rect 34588 10854 34590 10906
rect 34770 10854 34772 10906
rect 34526 10852 34532 10854
rect 34588 10852 34612 10854
rect 34668 10852 34692 10854
rect 34748 10852 34772 10854
rect 34828 10852 34834 10854
rect 34526 10843 34834 10852
rect 33876 10532 33928 10538
rect 33876 10474 33928 10480
rect 33888 10266 33916 10474
rect 33876 10260 33928 10266
rect 33876 10202 33928 10208
rect 34336 10056 34388 10062
rect 34336 9998 34388 10004
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33060 8634 33088 8774
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 32956 8560 33008 8566
rect 32956 8502 33008 8508
rect 32968 7886 32996 8502
rect 34060 8288 34112 8294
rect 34060 8230 34112 8236
rect 34072 7954 34100 8230
rect 34060 7948 34112 7954
rect 34060 7890 34112 7896
rect 34348 7886 34376 9998
rect 34526 9820 34834 9829
rect 34526 9818 34532 9820
rect 34588 9818 34612 9820
rect 34668 9818 34692 9820
rect 34748 9818 34772 9820
rect 34828 9818 34834 9820
rect 34588 9766 34590 9818
rect 34770 9766 34772 9818
rect 34526 9764 34532 9766
rect 34588 9764 34612 9766
rect 34668 9764 34692 9766
rect 34748 9764 34772 9766
rect 34828 9764 34834 9766
rect 34526 9755 34834 9764
rect 34526 8732 34834 8741
rect 34526 8730 34532 8732
rect 34588 8730 34612 8732
rect 34668 8730 34692 8732
rect 34748 8730 34772 8732
rect 34828 8730 34834 8732
rect 34588 8678 34590 8730
rect 34770 8678 34772 8730
rect 34526 8676 34532 8678
rect 34588 8676 34612 8678
rect 34668 8676 34692 8678
rect 34748 8676 34772 8678
rect 34828 8676 34834 8678
rect 34526 8667 34834 8676
rect 34796 8356 34848 8362
rect 34796 8298 34848 8304
rect 34808 8265 34836 8298
rect 34794 8256 34850 8265
rect 34794 8191 34850 8200
rect 32956 7880 33008 7886
rect 32956 7822 33008 7828
rect 34336 7880 34388 7886
rect 34336 7822 34388 7828
rect 32588 7268 32640 7274
rect 32588 7210 32640 7216
rect 32600 6866 32628 7210
rect 32588 6860 32640 6866
rect 32588 6802 32640 6808
rect 32496 6384 32548 6390
rect 32496 6326 32548 6332
rect 32128 6316 32180 6322
rect 32128 6258 32180 6264
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 31484 5364 31536 5370
rect 31484 5306 31536 5312
rect 30656 5228 30708 5234
rect 30656 5170 30708 5176
rect 30196 5160 30248 5166
rect 30196 5102 30248 5108
rect 30196 5024 30248 5030
rect 30196 4966 30248 4972
rect 30104 4820 30156 4826
rect 30104 4762 30156 4768
rect 29368 4752 29420 4758
rect 29368 4694 29420 4700
rect 30208 4282 30236 4966
rect 30329 4924 30637 4933
rect 30329 4922 30335 4924
rect 30391 4922 30415 4924
rect 30471 4922 30495 4924
rect 30551 4922 30575 4924
rect 30631 4922 30637 4924
rect 30391 4870 30393 4922
rect 30573 4870 30575 4922
rect 30329 4868 30335 4870
rect 30391 4868 30415 4870
rect 30471 4868 30495 4870
rect 30551 4868 30575 4870
rect 30631 4868 30637 4870
rect 30329 4859 30637 4868
rect 30668 4826 30696 5170
rect 30656 4820 30708 4826
rect 30656 4762 30708 4768
rect 28908 4276 28960 4282
rect 28908 4218 28960 4224
rect 30196 4276 30248 4282
rect 30196 4218 30248 4224
rect 32140 4214 32168 6258
rect 32508 5710 32536 6326
rect 32968 6322 32996 7822
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 32956 6316 33008 6322
rect 32956 6258 33008 6264
rect 33060 5710 33088 6598
rect 34348 6322 34376 7822
rect 34526 7644 34834 7653
rect 34526 7642 34532 7644
rect 34588 7642 34612 7644
rect 34668 7642 34692 7644
rect 34748 7642 34772 7644
rect 34828 7642 34834 7644
rect 34588 7590 34590 7642
rect 34770 7590 34772 7642
rect 34526 7588 34532 7590
rect 34588 7588 34612 7590
rect 34668 7588 34692 7590
rect 34748 7588 34772 7590
rect 34828 7588 34834 7590
rect 34526 7579 34834 7588
rect 34526 6556 34834 6565
rect 34526 6554 34532 6556
rect 34588 6554 34612 6556
rect 34668 6554 34692 6556
rect 34748 6554 34772 6556
rect 34828 6554 34834 6556
rect 34588 6502 34590 6554
rect 34770 6502 34772 6554
rect 34526 6500 34532 6502
rect 34588 6500 34612 6502
rect 34668 6500 34692 6502
rect 34748 6500 34772 6502
rect 34828 6500 34834 6502
rect 34526 6491 34834 6500
rect 34336 6316 34388 6322
rect 34336 6258 34388 6264
rect 34060 6248 34112 6254
rect 34060 6190 34112 6196
rect 34072 5914 34100 6190
rect 34060 5908 34112 5914
rect 34060 5850 34112 5856
rect 32496 5704 32548 5710
rect 32496 5646 32548 5652
rect 33048 5704 33100 5710
rect 33048 5646 33100 5652
rect 32128 4208 32180 4214
rect 32128 4150 32180 4156
rect 34348 4146 34376 6258
rect 34526 5468 34834 5477
rect 34526 5466 34532 5468
rect 34588 5466 34612 5468
rect 34668 5466 34692 5468
rect 34748 5466 34772 5468
rect 34828 5466 34834 5468
rect 34588 5414 34590 5466
rect 34770 5414 34772 5466
rect 34526 5412 34532 5414
rect 34588 5412 34612 5414
rect 34668 5412 34692 5414
rect 34748 5412 34772 5414
rect 34828 5412 34834 5414
rect 34526 5403 34834 5412
rect 34526 4380 34834 4389
rect 34526 4378 34532 4380
rect 34588 4378 34612 4380
rect 34668 4378 34692 4380
rect 34748 4378 34772 4380
rect 34828 4378 34834 4380
rect 34588 4326 34590 4378
rect 34770 4326 34772 4378
rect 34526 4324 34532 4326
rect 34588 4324 34612 4326
rect 34668 4324 34692 4326
rect 34748 4324 34772 4326
rect 34828 4324 34834 4326
rect 34526 4315 34834 4324
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 34336 4140 34388 4146
rect 34336 4082 34388 4088
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 31668 4072 31720 4078
rect 31668 4014 31720 4020
rect 21935 3836 22243 3845
rect 21935 3834 21941 3836
rect 21997 3834 22021 3836
rect 22077 3834 22101 3836
rect 22157 3834 22181 3836
rect 22237 3834 22243 3836
rect 21997 3782 21999 3834
rect 22179 3782 22181 3834
rect 21935 3780 21941 3782
rect 21997 3780 22021 3782
rect 22077 3780 22101 3782
rect 22157 3780 22181 3782
rect 22237 3780 22243 3782
rect 21935 3771 22243 3780
rect 30329 3836 30637 3845
rect 30329 3834 30335 3836
rect 30391 3834 30415 3836
rect 30471 3834 30495 3836
rect 30551 3834 30575 3836
rect 30631 3834 30637 3836
rect 30391 3782 30393 3834
rect 30573 3782 30575 3834
rect 30329 3780 30335 3782
rect 30391 3780 30415 3782
rect 30471 3780 30495 3782
rect 30551 3780 30575 3782
rect 30631 3780 30637 3782
rect 30329 3771 30637 3780
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 24584 3460 24636 3466
rect 24584 3402 24636 3408
rect 17738 3292 18046 3301
rect 17738 3290 17744 3292
rect 17800 3290 17824 3292
rect 17880 3290 17904 3292
rect 17960 3290 17984 3292
rect 18040 3290 18046 3292
rect 17800 3238 17802 3290
rect 17982 3238 17984 3290
rect 17738 3236 17744 3238
rect 17800 3236 17824 3238
rect 17880 3236 17904 3238
rect 17960 3236 17984 3238
rect 18040 3236 18046 3238
rect 17738 3227 18046 3236
rect 21935 2748 22243 2757
rect 21935 2746 21941 2748
rect 21997 2746 22021 2748
rect 22077 2746 22101 2748
rect 22157 2746 22181 2748
rect 22237 2746 22243 2748
rect 21997 2694 21999 2746
rect 22179 2694 22181 2746
rect 21935 2692 21941 2694
rect 21997 2692 22021 2694
rect 22077 2692 22101 2694
rect 22157 2692 22181 2694
rect 22237 2692 22243 2694
rect 21935 2683 22243 2692
rect 24596 2650 24624 3402
rect 26132 3292 26440 3301
rect 26132 3290 26138 3292
rect 26194 3290 26218 3292
rect 26274 3290 26298 3292
rect 26354 3290 26378 3292
rect 26434 3290 26440 3292
rect 26194 3238 26196 3290
rect 26376 3238 26378 3290
rect 26132 3236 26138 3238
rect 26194 3236 26218 3238
rect 26274 3236 26298 3238
rect 26354 3236 26378 3238
rect 26434 3236 26440 3238
rect 26132 3227 26440 3236
rect 30329 2748 30637 2757
rect 30329 2746 30335 2748
rect 30391 2746 30415 2748
rect 30471 2746 30495 2748
rect 30551 2746 30575 2748
rect 30631 2746 30637 2748
rect 30391 2694 30393 2746
rect 30573 2694 30575 2746
rect 30329 2692 30335 2694
rect 30391 2692 30415 2694
rect 30471 2692 30495 2694
rect 30551 2692 30575 2694
rect 30631 2692 30637 2694
rect 30329 2683 30637 2692
rect 31680 2650 31708 4014
rect 34526 3292 34834 3301
rect 34526 3290 34532 3292
rect 34588 3290 34612 3292
rect 34668 3290 34692 3292
rect 34748 3290 34772 3292
rect 34828 3290 34834 3292
rect 34588 3238 34590 3290
rect 34770 3238 34772 3290
rect 34526 3236 34532 3238
rect 34588 3236 34612 3238
rect 34668 3236 34692 3238
rect 34748 3236 34772 3238
rect 34828 3236 34834 3238
rect 34526 3227 34834 3236
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 9344 2204 9652 2213
rect 9344 2202 9350 2204
rect 9406 2202 9430 2204
rect 9486 2202 9510 2204
rect 9566 2202 9590 2204
rect 9646 2202 9652 2204
rect 9406 2150 9408 2202
rect 9588 2150 9590 2202
rect 9344 2148 9350 2150
rect 9406 2148 9430 2150
rect 9486 2148 9510 2150
rect 9566 2148 9590 2150
rect 9646 2148 9652 2150
rect 9344 2139 9652 2148
rect 5828 1278 5948 1306
rect 5828 800 5856 1278
rect 12268 800 12296 2382
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 17738 2204 18046 2213
rect 17738 2202 17744 2204
rect 17800 2202 17824 2204
rect 17880 2202 17904 2204
rect 17960 2202 17984 2204
rect 18040 2202 18046 2204
rect 17800 2150 17802 2202
rect 17982 2150 17984 2202
rect 17738 2148 17744 2150
rect 17800 2148 17824 2150
rect 17880 2148 17904 2150
rect 17960 2148 17984 2150
rect 18040 2148 18046 2150
rect 17738 2139 18046 2148
rect 18708 870 18828 898
rect 18708 800 18736 870
rect 18 0 74 800
rect 5814 0 5870 800
rect 12254 0 12310 800
rect 18694 0 18750 800
rect 18800 762 18828 870
rect 19076 762 19104 2246
rect 24504 800 24532 2382
rect 26132 2204 26440 2213
rect 26132 2202 26138 2204
rect 26194 2202 26218 2204
rect 26274 2202 26298 2204
rect 26354 2202 26378 2204
rect 26434 2202 26440 2204
rect 26194 2150 26196 2202
rect 26376 2150 26378 2202
rect 26132 2148 26138 2150
rect 26194 2148 26218 2150
rect 26274 2148 26298 2150
rect 26354 2148 26378 2150
rect 26434 2148 26440 2150
rect 26132 2139 26440 2148
rect 31036 1306 31064 2382
rect 34428 2304 34480 2310
rect 34428 2246 34480 2252
rect 34440 1442 34468 2246
rect 34526 2204 34834 2213
rect 34526 2202 34532 2204
rect 34588 2202 34612 2204
rect 34668 2202 34692 2204
rect 34748 2202 34772 2204
rect 34828 2202 34834 2204
rect 34588 2150 34590 2202
rect 34770 2150 34772 2202
rect 34526 2148 34532 2150
rect 34588 2148 34612 2150
rect 34668 2148 34692 2150
rect 34748 2148 34772 2150
rect 34828 2148 34834 2150
rect 34526 2139 34834 2148
rect 34518 1456 34574 1465
rect 34440 1414 34518 1442
rect 34518 1391 34574 1400
rect 30944 1278 31064 1306
rect 30944 800 30972 1278
rect 18800 734 19104 762
rect 24490 0 24546 800
rect 30930 0 30986 800
<< via2 >>
rect 5153 35386 5209 35388
rect 5233 35386 5289 35388
rect 5313 35386 5369 35388
rect 5393 35386 5449 35388
rect 5153 35334 5199 35386
rect 5199 35334 5209 35386
rect 5233 35334 5263 35386
rect 5263 35334 5275 35386
rect 5275 35334 5289 35386
rect 5313 35334 5327 35386
rect 5327 35334 5339 35386
rect 5339 35334 5369 35386
rect 5393 35334 5403 35386
rect 5403 35334 5449 35386
rect 5153 35332 5209 35334
rect 5233 35332 5289 35334
rect 5313 35332 5369 35334
rect 5393 35332 5449 35334
rect 13547 35386 13603 35388
rect 13627 35386 13683 35388
rect 13707 35386 13763 35388
rect 13787 35386 13843 35388
rect 13547 35334 13593 35386
rect 13593 35334 13603 35386
rect 13627 35334 13657 35386
rect 13657 35334 13669 35386
rect 13669 35334 13683 35386
rect 13707 35334 13721 35386
rect 13721 35334 13733 35386
rect 13733 35334 13763 35386
rect 13787 35334 13797 35386
rect 13797 35334 13843 35386
rect 13547 35332 13603 35334
rect 13627 35332 13683 35334
rect 13707 35332 13763 35334
rect 13787 35332 13843 35334
rect 938 32680 994 32736
rect 1398 26152 1454 26208
rect 938 19796 940 19816
rect 940 19796 992 19816
rect 992 19796 994 19816
rect 938 19760 994 19796
rect 5153 34298 5209 34300
rect 5233 34298 5289 34300
rect 5313 34298 5369 34300
rect 5393 34298 5449 34300
rect 5153 34246 5199 34298
rect 5199 34246 5209 34298
rect 5233 34246 5263 34298
rect 5263 34246 5275 34298
rect 5275 34246 5289 34298
rect 5313 34246 5327 34298
rect 5327 34246 5339 34298
rect 5339 34246 5369 34298
rect 5393 34246 5403 34298
rect 5403 34246 5449 34298
rect 5153 34244 5209 34246
rect 5233 34244 5289 34246
rect 5313 34244 5369 34246
rect 5393 34244 5449 34246
rect 5153 33210 5209 33212
rect 5233 33210 5289 33212
rect 5313 33210 5369 33212
rect 5393 33210 5449 33212
rect 5153 33158 5199 33210
rect 5199 33158 5209 33210
rect 5233 33158 5263 33210
rect 5263 33158 5275 33210
rect 5275 33158 5289 33210
rect 5313 33158 5327 33210
rect 5327 33158 5339 33210
rect 5339 33158 5369 33210
rect 5393 33158 5403 33210
rect 5403 33158 5449 33210
rect 5153 33156 5209 33158
rect 5233 33156 5289 33158
rect 5313 33156 5369 33158
rect 5393 33156 5449 33158
rect 5153 32122 5209 32124
rect 5233 32122 5289 32124
rect 5313 32122 5369 32124
rect 5393 32122 5449 32124
rect 5153 32070 5199 32122
rect 5199 32070 5209 32122
rect 5233 32070 5263 32122
rect 5263 32070 5275 32122
rect 5275 32070 5289 32122
rect 5313 32070 5327 32122
rect 5327 32070 5339 32122
rect 5339 32070 5369 32122
rect 5393 32070 5403 32122
rect 5403 32070 5449 32122
rect 5153 32068 5209 32070
rect 5233 32068 5289 32070
rect 5313 32068 5369 32070
rect 5393 32068 5449 32070
rect 9350 34842 9406 34844
rect 9430 34842 9486 34844
rect 9510 34842 9566 34844
rect 9590 34842 9646 34844
rect 9350 34790 9396 34842
rect 9396 34790 9406 34842
rect 9430 34790 9460 34842
rect 9460 34790 9472 34842
rect 9472 34790 9486 34842
rect 9510 34790 9524 34842
rect 9524 34790 9536 34842
rect 9536 34790 9566 34842
rect 9590 34790 9600 34842
rect 9600 34790 9646 34842
rect 9350 34788 9406 34790
rect 9430 34788 9486 34790
rect 9510 34788 9566 34790
rect 9590 34788 9646 34790
rect 5153 31034 5209 31036
rect 5233 31034 5289 31036
rect 5313 31034 5369 31036
rect 5393 31034 5449 31036
rect 5153 30982 5199 31034
rect 5199 30982 5209 31034
rect 5233 30982 5263 31034
rect 5263 30982 5275 31034
rect 5275 30982 5289 31034
rect 5313 30982 5327 31034
rect 5327 30982 5339 31034
rect 5339 30982 5369 31034
rect 5393 30982 5403 31034
rect 5403 30982 5449 31034
rect 5153 30980 5209 30982
rect 5233 30980 5289 30982
rect 5313 30980 5369 30982
rect 5393 30980 5449 30982
rect 5153 29946 5209 29948
rect 5233 29946 5289 29948
rect 5313 29946 5369 29948
rect 5393 29946 5449 29948
rect 5153 29894 5199 29946
rect 5199 29894 5209 29946
rect 5233 29894 5263 29946
rect 5263 29894 5275 29946
rect 5275 29894 5289 29946
rect 5313 29894 5327 29946
rect 5327 29894 5339 29946
rect 5339 29894 5369 29946
rect 5393 29894 5403 29946
rect 5403 29894 5449 29946
rect 5153 29892 5209 29894
rect 5233 29892 5289 29894
rect 5313 29892 5369 29894
rect 5393 29892 5449 29894
rect 5153 28858 5209 28860
rect 5233 28858 5289 28860
rect 5313 28858 5369 28860
rect 5393 28858 5449 28860
rect 5153 28806 5199 28858
rect 5199 28806 5209 28858
rect 5233 28806 5263 28858
rect 5263 28806 5275 28858
rect 5275 28806 5289 28858
rect 5313 28806 5327 28858
rect 5327 28806 5339 28858
rect 5339 28806 5369 28858
rect 5393 28806 5403 28858
rect 5403 28806 5449 28858
rect 5153 28804 5209 28806
rect 5233 28804 5289 28806
rect 5313 28804 5369 28806
rect 5393 28804 5449 28806
rect 5153 27770 5209 27772
rect 5233 27770 5289 27772
rect 5313 27770 5369 27772
rect 5393 27770 5449 27772
rect 5153 27718 5199 27770
rect 5199 27718 5209 27770
rect 5233 27718 5263 27770
rect 5263 27718 5275 27770
rect 5275 27718 5289 27770
rect 5313 27718 5327 27770
rect 5327 27718 5339 27770
rect 5339 27718 5369 27770
rect 5393 27718 5403 27770
rect 5403 27718 5449 27770
rect 5153 27716 5209 27718
rect 5233 27716 5289 27718
rect 5313 27716 5369 27718
rect 5393 27716 5449 27718
rect 9350 33754 9406 33756
rect 9430 33754 9486 33756
rect 9510 33754 9566 33756
rect 9590 33754 9646 33756
rect 9350 33702 9396 33754
rect 9396 33702 9406 33754
rect 9430 33702 9460 33754
rect 9460 33702 9472 33754
rect 9472 33702 9486 33754
rect 9510 33702 9524 33754
rect 9524 33702 9536 33754
rect 9536 33702 9566 33754
rect 9590 33702 9600 33754
rect 9600 33702 9646 33754
rect 9350 33700 9406 33702
rect 9430 33700 9486 33702
rect 9510 33700 9566 33702
rect 9590 33700 9646 33702
rect 9350 32666 9406 32668
rect 9430 32666 9486 32668
rect 9510 32666 9566 32668
rect 9590 32666 9646 32668
rect 9350 32614 9396 32666
rect 9396 32614 9406 32666
rect 9430 32614 9460 32666
rect 9460 32614 9472 32666
rect 9472 32614 9486 32666
rect 9510 32614 9524 32666
rect 9524 32614 9536 32666
rect 9536 32614 9566 32666
rect 9590 32614 9600 32666
rect 9600 32614 9646 32666
rect 9350 32612 9406 32614
rect 9430 32612 9486 32614
rect 9510 32612 9566 32614
rect 9590 32612 9646 32614
rect 9350 31578 9406 31580
rect 9430 31578 9486 31580
rect 9510 31578 9566 31580
rect 9590 31578 9646 31580
rect 9350 31526 9396 31578
rect 9396 31526 9406 31578
rect 9430 31526 9460 31578
rect 9460 31526 9472 31578
rect 9472 31526 9486 31578
rect 9510 31526 9524 31578
rect 9524 31526 9536 31578
rect 9536 31526 9566 31578
rect 9590 31526 9600 31578
rect 9600 31526 9646 31578
rect 9350 31524 9406 31526
rect 9430 31524 9486 31526
rect 9510 31524 9566 31526
rect 9590 31524 9646 31526
rect 5153 26682 5209 26684
rect 5233 26682 5289 26684
rect 5313 26682 5369 26684
rect 5393 26682 5449 26684
rect 5153 26630 5199 26682
rect 5199 26630 5209 26682
rect 5233 26630 5263 26682
rect 5263 26630 5275 26682
rect 5275 26630 5289 26682
rect 5313 26630 5327 26682
rect 5327 26630 5339 26682
rect 5339 26630 5369 26682
rect 5393 26630 5403 26682
rect 5403 26630 5449 26682
rect 5153 26628 5209 26630
rect 5233 26628 5289 26630
rect 5313 26628 5369 26630
rect 5393 26628 5449 26630
rect 5153 25594 5209 25596
rect 5233 25594 5289 25596
rect 5313 25594 5369 25596
rect 5393 25594 5449 25596
rect 5153 25542 5199 25594
rect 5199 25542 5209 25594
rect 5233 25542 5263 25594
rect 5263 25542 5275 25594
rect 5275 25542 5289 25594
rect 5313 25542 5327 25594
rect 5327 25542 5339 25594
rect 5339 25542 5369 25594
rect 5393 25542 5403 25594
rect 5403 25542 5449 25594
rect 5153 25540 5209 25542
rect 5233 25540 5289 25542
rect 5313 25540 5369 25542
rect 5393 25540 5449 25542
rect 9350 30490 9406 30492
rect 9430 30490 9486 30492
rect 9510 30490 9566 30492
rect 9590 30490 9646 30492
rect 9350 30438 9396 30490
rect 9396 30438 9406 30490
rect 9430 30438 9460 30490
rect 9460 30438 9472 30490
rect 9472 30438 9486 30490
rect 9510 30438 9524 30490
rect 9524 30438 9536 30490
rect 9536 30438 9566 30490
rect 9590 30438 9600 30490
rect 9600 30438 9646 30490
rect 9350 30436 9406 30438
rect 9430 30436 9486 30438
rect 9510 30436 9566 30438
rect 9590 30436 9646 30438
rect 9126 29572 9182 29608
rect 9126 29552 9128 29572
rect 9128 29552 9180 29572
rect 9180 29552 9182 29572
rect 5153 24506 5209 24508
rect 5233 24506 5289 24508
rect 5313 24506 5369 24508
rect 5393 24506 5449 24508
rect 5153 24454 5199 24506
rect 5199 24454 5209 24506
rect 5233 24454 5263 24506
rect 5263 24454 5275 24506
rect 5275 24454 5289 24506
rect 5313 24454 5327 24506
rect 5327 24454 5339 24506
rect 5339 24454 5369 24506
rect 5393 24454 5403 24506
rect 5403 24454 5449 24506
rect 5153 24452 5209 24454
rect 5233 24452 5289 24454
rect 5313 24452 5369 24454
rect 5393 24452 5449 24454
rect 5153 23418 5209 23420
rect 5233 23418 5289 23420
rect 5313 23418 5369 23420
rect 5393 23418 5449 23420
rect 5153 23366 5199 23418
rect 5199 23366 5209 23418
rect 5233 23366 5263 23418
rect 5263 23366 5275 23418
rect 5275 23366 5289 23418
rect 5313 23366 5327 23418
rect 5327 23366 5339 23418
rect 5339 23366 5369 23418
rect 5393 23366 5403 23418
rect 5403 23366 5449 23418
rect 5153 23364 5209 23366
rect 5233 23364 5289 23366
rect 5313 23364 5369 23366
rect 5393 23364 5449 23366
rect 9350 29402 9406 29404
rect 9430 29402 9486 29404
rect 9510 29402 9566 29404
rect 9590 29402 9646 29404
rect 9350 29350 9396 29402
rect 9396 29350 9406 29402
rect 9430 29350 9460 29402
rect 9460 29350 9472 29402
rect 9472 29350 9486 29402
rect 9510 29350 9524 29402
rect 9524 29350 9536 29402
rect 9536 29350 9566 29402
rect 9590 29350 9600 29402
rect 9600 29350 9646 29402
rect 9350 29348 9406 29350
rect 9430 29348 9486 29350
rect 9510 29348 9566 29350
rect 9590 29348 9646 29350
rect 938 12960 994 13016
rect 3146 19352 3202 19408
rect 5153 22330 5209 22332
rect 5233 22330 5289 22332
rect 5313 22330 5369 22332
rect 5393 22330 5449 22332
rect 5153 22278 5199 22330
rect 5199 22278 5209 22330
rect 5233 22278 5263 22330
rect 5263 22278 5275 22330
rect 5275 22278 5289 22330
rect 5313 22278 5327 22330
rect 5327 22278 5339 22330
rect 5339 22278 5369 22330
rect 5393 22278 5403 22330
rect 5403 22278 5449 22330
rect 5153 22276 5209 22278
rect 5233 22276 5289 22278
rect 5313 22276 5369 22278
rect 5393 22276 5449 22278
rect 5153 21242 5209 21244
rect 5233 21242 5289 21244
rect 5313 21242 5369 21244
rect 5393 21242 5449 21244
rect 5153 21190 5199 21242
rect 5199 21190 5209 21242
rect 5233 21190 5263 21242
rect 5263 21190 5275 21242
rect 5275 21190 5289 21242
rect 5313 21190 5327 21242
rect 5327 21190 5339 21242
rect 5339 21190 5369 21242
rect 5393 21190 5403 21242
rect 5403 21190 5449 21242
rect 5153 21188 5209 21190
rect 5233 21188 5289 21190
rect 5313 21188 5369 21190
rect 5393 21188 5449 21190
rect 5153 20154 5209 20156
rect 5233 20154 5289 20156
rect 5313 20154 5369 20156
rect 5393 20154 5449 20156
rect 5153 20102 5199 20154
rect 5199 20102 5209 20154
rect 5233 20102 5263 20154
rect 5263 20102 5275 20154
rect 5275 20102 5289 20154
rect 5313 20102 5327 20154
rect 5327 20102 5339 20154
rect 5339 20102 5369 20154
rect 5393 20102 5403 20154
rect 5403 20102 5449 20154
rect 5153 20100 5209 20102
rect 5233 20100 5289 20102
rect 5313 20100 5369 20102
rect 5393 20100 5449 20102
rect 4618 18808 4674 18864
rect 3606 17196 3662 17232
rect 3606 17176 3608 17196
rect 3608 17176 3660 17196
rect 3660 17176 3662 17196
rect 4434 16632 4490 16688
rect 4250 13912 4306 13968
rect 5722 20304 5778 20360
rect 5153 19066 5209 19068
rect 5233 19066 5289 19068
rect 5313 19066 5369 19068
rect 5393 19066 5449 19068
rect 5153 19014 5199 19066
rect 5199 19014 5209 19066
rect 5233 19014 5263 19066
rect 5263 19014 5275 19066
rect 5275 19014 5289 19066
rect 5313 19014 5327 19066
rect 5327 19014 5339 19066
rect 5339 19014 5369 19066
rect 5393 19014 5403 19066
rect 5403 19014 5449 19066
rect 5153 19012 5209 19014
rect 5233 19012 5289 19014
rect 5313 19012 5369 19014
rect 5393 19012 5449 19014
rect 5153 17978 5209 17980
rect 5233 17978 5289 17980
rect 5313 17978 5369 17980
rect 5393 17978 5449 17980
rect 5153 17926 5199 17978
rect 5199 17926 5209 17978
rect 5233 17926 5263 17978
rect 5263 17926 5275 17978
rect 5275 17926 5289 17978
rect 5313 17926 5327 17978
rect 5327 17926 5339 17978
rect 5339 17926 5369 17978
rect 5393 17926 5403 17978
rect 5403 17926 5449 17978
rect 5153 17924 5209 17926
rect 5233 17924 5289 17926
rect 5313 17924 5369 17926
rect 5393 17924 5449 17926
rect 4618 13932 4674 13968
rect 4618 13912 4620 13932
rect 4620 13912 4672 13932
rect 4672 13912 4674 13932
rect 5153 16890 5209 16892
rect 5233 16890 5289 16892
rect 5313 16890 5369 16892
rect 5393 16890 5449 16892
rect 5153 16838 5199 16890
rect 5199 16838 5209 16890
rect 5233 16838 5263 16890
rect 5263 16838 5275 16890
rect 5275 16838 5289 16890
rect 5313 16838 5327 16890
rect 5327 16838 5339 16890
rect 5339 16838 5369 16890
rect 5393 16838 5403 16890
rect 5403 16838 5449 16890
rect 5153 16836 5209 16838
rect 5233 16836 5289 16838
rect 5313 16836 5369 16838
rect 5393 16836 5449 16838
rect 5998 19780 6054 19816
rect 5998 19760 6000 19780
rect 6000 19760 6052 19780
rect 6052 19760 6054 19780
rect 5153 15802 5209 15804
rect 5233 15802 5289 15804
rect 5313 15802 5369 15804
rect 5393 15802 5449 15804
rect 5153 15750 5199 15802
rect 5199 15750 5209 15802
rect 5233 15750 5263 15802
rect 5263 15750 5275 15802
rect 5275 15750 5289 15802
rect 5313 15750 5327 15802
rect 5327 15750 5339 15802
rect 5339 15750 5369 15802
rect 5393 15750 5403 15802
rect 5403 15750 5449 15802
rect 5153 15748 5209 15750
rect 5233 15748 5289 15750
rect 5313 15748 5369 15750
rect 5393 15748 5449 15750
rect 7102 17720 7158 17776
rect 6826 16532 6828 16552
rect 6828 16532 6880 16552
rect 6880 16532 6882 16552
rect 6826 16496 6882 16532
rect 5814 15156 5870 15192
rect 5814 15136 5816 15156
rect 5816 15136 5868 15156
rect 5868 15136 5870 15156
rect 5153 14714 5209 14716
rect 5233 14714 5289 14716
rect 5313 14714 5369 14716
rect 5393 14714 5449 14716
rect 5153 14662 5199 14714
rect 5199 14662 5209 14714
rect 5233 14662 5263 14714
rect 5263 14662 5275 14714
rect 5275 14662 5289 14714
rect 5313 14662 5327 14714
rect 5327 14662 5339 14714
rect 5339 14662 5369 14714
rect 5393 14662 5403 14714
rect 5403 14662 5449 14714
rect 5153 14660 5209 14662
rect 5233 14660 5289 14662
rect 5313 14660 5369 14662
rect 5393 14660 5449 14662
rect 5153 13626 5209 13628
rect 5233 13626 5289 13628
rect 5313 13626 5369 13628
rect 5393 13626 5449 13628
rect 5153 13574 5199 13626
rect 5199 13574 5209 13626
rect 5233 13574 5263 13626
rect 5263 13574 5275 13626
rect 5275 13574 5289 13626
rect 5313 13574 5327 13626
rect 5327 13574 5339 13626
rect 5339 13574 5369 13626
rect 5393 13574 5403 13626
rect 5403 13574 5449 13626
rect 5153 13572 5209 13574
rect 5233 13572 5289 13574
rect 5313 13572 5369 13574
rect 5393 13572 5449 13574
rect 5153 12538 5209 12540
rect 5233 12538 5289 12540
rect 5313 12538 5369 12540
rect 5393 12538 5449 12540
rect 5153 12486 5199 12538
rect 5199 12486 5209 12538
rect 5233 12486 5263 12538
rect 5263 12486 5275 12538
rect 5275 12486 5289 12538
rect 5313 12486 5327 12538
rect 5327 12486 5339 12538
rect 5339 12486 5369 12538
rect 5393 12486 5403 12538
rect 5403 12486 5449 12538
rect 5153 12484 5209 12486
rect 5233 12484 5289 12486
rect 5313 12484 5369 12486
rect 5393 12484 5449 12486
rect 5446 12164 5502 12200
rect 5446 12144 5448 12164
rect 5448 12144 5500 12164
rect 5500 12144 5502 12164
rect 5078 11756 5134 11792
rect 5078 11736 5080 11756
rect 5080 11736 5132 11756
rect 5132 11736 5134 11756
rect 5153 11450 5209 11452
rect 5233 11450 5289 11452
rect 5313 11450 5369 11452
rect 5393 11450 5449 11452
rect 5153 11398 5199 11450
rect 5199 11398 5209 11450
rect 5233 11398 5263 11450
rect 5263 11398 5275 11450
rect 5275 11398 5289 11450
rect 5313 11398 5327 11450
rect 5327 11398 5339 11450
rect 5339 11398 5369 11450
rect 5393 11398 5403 11450
rect 5403 11398 5449 11450
rect 5153 11396 5209 11398
rect 5233 11396 5289 11398
rect 5313 11396 5369 11398
rect 5393 11396 5449 11398
rect 6918 15408 6974 15464
rect 7010 14864 7066 14920
rect 7378 17196 7434 17232
rect 7378 17176 7380 17196
rect 7380 17176 7432 17196
rect 7432 17176 7434 17196
rect 7930 16768 7986 16824
rect 7746 16632 7802 16688
rect 8114 16224 8170 16280
rect 8298 16360 8354 16416
rect 6274 10920 6330 10976
rect 5153 10362 5209 10364
rect 5233 10362 5289 10364
rect 5313 10362 5369 10364
rect 5393 10362 5449 10364
rect 5153 10310 5199 10362
rect 5199 10310 5209 10362
rect 5233 10310 5263 10362
rect 5263 10310 5275 10362
rect 5275 10310 5289 10362
rect 5313 10310 5327 10362
rect 5327 10310 5339 10362
rect 5339 10310 5369 10362
rect 5393 10310 5403 10362
rect 5403 10310 5449 10362
rect 5153 10308 5209 10310
rect 5233 10308 5289 10310
rect 5313 10308 5369 10310
rect 5393 10308 5449 10310
rect 6826 11056 6882 11112
rect 7470 12416 7526 12472
rect 7930 15136 7986 15192
rect 8482 19352 8538 19408
rect 8298 13368 8354 13424
rect 8758 18828 8814 18864
rect 8758 18808 8760 18828
rect 8760 18808 8812 18828
rect 8812 18808 8814 18828
rect 9350 28314 9406 28316
rect 9430 28314 9486 28316
rect 9510 28314 9566 28316
rect 9590 28314 9646 28316
rect 9350 28262 9396 28314
rect 9396 28262 9406 28314
rect 9430 28262 9460 28314
rect 9460 28262 9472 28314
rect 9472 28262 9486 28314
rect 9510 28262 9524 28314
rect 9524 28262 9536 28314
rect 9536 28262 9566 28314
rect 9590 28262 9600 28314
rect 9600 28262 9646 28314
rect 9350 28260 9406 28262
rect 9430 28260 9486 28262
rect 9510 28260 9566 28262
rect 9590 28260 9646 28262
rect 9350 27226 9406 27228
rect 9430 27226 9486 27228
rect 9510 27226 9566 27228
rect 9590 27226 9646 27228
rect 9350 27174 9396 27226
rect 9396 27174 9406 27226
rect 9430 27174 9460 27226
rect 9460 27174 9472 27226
rect 9472 27174 9486 27226
rect 9510 27174 9524 27226
rect 9524 27174 9536 27226
rect 9536 27174 9566 27226
rect 9590 27174 9600 27226
rect 9600 27174 9646 27226
rect 9350 27172 9406 27174
rect 9430 27172 9486 27174
rect 9510 27172 9566 27174
rect 9590 27172 9646 27174
rect 10230 29552 10286 29608
rect 13547 34298 13603 34300
rect 13627 34298 13683 34300
rect 13707 34298 13763 34300
rect 13787 34298 13843 34300
rect 13547 34246 13593 34298
rect 13593 34246 13603 34298
rect 13627 34246 13657 34298
rect 13657 34246 13669 34298
rect 13669 34246 13683 34298
rect 13707 34246 13721 34298
rect 13721 34246 13733 34298
rect 13733 34246 13763 34298
rect 13787 34246 13797 34298
rect 13797 34246 13843 34298
rect 13547 34244 13603 34246
rect 13627 34244 13683 34246
rect 13707 34244 13763 34246
rect 13787 34244 13843 34246
rect 13547 33210 13603 33212
rect 13627 33210 13683 33212
rect 13707 33210 13763 33212
rect 13787 33210 13843 33212
rect 13547 33158 13593 33210
rect 13593 33158 13603 33210
rect 13627 33158 13657 33210
rect 13657 33158 13669 33210
rect 13669 33158 13683 33210
rect 13707 33158 13721 33210
rect 13721 33158 13733 33210
rect 13733 33158 13763 33210
rect 13787 33158 13797 33210
rect 13797 33158 13843 33210
rect 13547 33156 13603 33158
rect 13627 33156 13683 33158
rect 13707 33156 13763 33158
rect 13787 33156 13843 33158
rect 21941 35386 21997 35388
rect 22021 35386 22077 35388
rect 22101 35386 22157 35388
rect 22181 35386 22237 35388
rect 21941 35334 21987 35386
rect 21987 35334 21997 35386
rect 22021 35334 22051 35386
rect 22051 35334 22063 35386
rect 22063 35334 22077 35386
rect 22101 35334 22115 35386
rect 22115 35334 22127 35386
rect 22127 35334 22157 35386
rect 22181 35334 22191 35386
rect 22191 35334 22237 35386
rect 21941 35332 21997 35334
rect 22021 35332 22077 35334
rect 22101 35332 22157 35334
rect 22181 35332 22237 35334
rect 30335 35386 30391 35388
rect 30415 35386 30471 35388
rect 30495 35386 30551 35388
rect 30575 35386 30631 35388
rect 30335 35334 30381 35386
rect 30381 35334 30391 35386
rect 30415 35334 30445 35386
rect 30445 35334 30457 35386
rect 30457 35334 30471 35386
rect 30495 35334 30509 35386
rect 30509 35334 30521 35386
rect 30521 35334 30551 35386
rect 30575 35334 30585 35386
rect 30585 35334 30631 35386
rect 30335 35332 30391 35334
rect 30415 35332 30471 35334
rect 30495 35332 30551 35334
rect 30575 35332 30631 35334
rect 9350 26138 9406 26140
rect 9430 26138 9486 26140
rect 9510 26138 9566 26140
rect 9590 26138 9646 26140
rect 9350 26086 9396 26138
rect 9396 26086 9406 26138
rect 9430 26086 9460 26138
rect 9460 26086 9472 26138
rect 9472 26086 9486 26138
rect 9510 26086 9524 26138
rect 9524 26086 9536 26138
rect 9536 26086 9566 26138
rect 9590 26086 9600 26138
rect 9600 26086 9646 26138
rect 9350 26084 9406 26086
rect 9430 26084 9486 26086
rect 9510 26084 9566 26086
rect 9590 26084 9646 26086
rect 9350 25050 9406 25052
rect 9430 25050 9486 25052
rect 9510 25050 9566 25052
rect 9590 25050 9646 25052
rect 9350 24998 9396 25050
rect 9396 24998 9406 25050
rect 9430 24998 9460 25050
rect 9460 24998 9472 25050
rect 9472 24998 9486 25050
rect 9510 24998 9524 25050
rect 9524 24998 9536 25050
rect 9536 24998 9566 25050
rect 9590 24998 9600 25050
rect 9600 24998 9646 25050
rect 9350 24996 9406 24998
rect 9430 24996 9486 24998
rect 9510 24996 9566 24998
rect 9590 24996 9646 24998
rect 9350 23962 9406 23964
rect 9430 23962 9486 23964
rect 9510 23962 9566 23964
rect 9590 23962 9646 23964
rect 9350 23910 9396 23962
rect 9396 23910 9406 23962
rect 9430 23910 9460 23962
rect 9460 23910 9472 23962
rect 9472 23910 9486 23962
rect 9510 23910 9524 23962
rect 9524 23910 9536 23962
rect 9536 23910 9566 23962
rect 9590 23910 9600 23962
rect 9600 23910 9646 23962
rect 9350 23908 9406 23910
rect 9430 23908 9486 23910
rect 9510 23908 9566 23910
rect 9590 23908 9646 23910
rect 13547 32122 13603 32124
rect 13627 32122 13683 32124
rect 13707 32122 13763 32124
rect 13787 32122 13843 32124
rect 13547 32070 13593 32122
rect 13593 32070 13603 32122
rect 13627 32070 13657 32122
rect 13657 32070 13669 32122
rect 13669 32070 13683 32122
rect 13707 32070 13721 32122
rect 13721 32070 13733 32122
rect 13733 32070 13763 32122
rect 13787 32070 13797 32122
rect 13797 32070 13843 32122
rect 13547 32068 13603 32070
rect 13627 32068 13683 32070
rect 13707 32068 13763 32070
rect 13787 32068 13843 32070
rect 13547 31034 13603 31036
rect 13627 31034 13683 31036
rect 13707 31034 13763 31036
rect 13787 31034 13843 31036
rect 13547 30982 13593 31034
rect 13593 30982 13603 31034
rect 13627 30982 13657 31034
rect 13657 30982 13669 31034
rect 13669 30982 13683 31034
rect 13707 30982 13721 31034
rect 13721 30982 13733 31034
rect 13733 30982 13763 31034
rect 13787 30982 13797 31034
rect 13797 30982 13843 31034
rect 13547 30980 13603 30982
rect 13627 30980 13683 30982
rect 13707 30980 13763 30982
rect 13787 30980 13843 30982
rect 17744 34842 17800 34844
rect 17824 34842 17880 34844
rect 17904 34842 17960 34844
rect 17984 34842 18040 34844
rect 17744 34790 17790 34842
rect 17790 34790 17800 34842
rect 17824 34790 17854 34842
rect 17854 34790 17866 34842
rect 17866 34790 17880 34842
rect 17904 34790 17918 34842
rect 17918 34790 17930 34842
rect 17930 34790 17960 34842
rect 17984 34790 17994 34842
rect 17994 34790 18040 34842
rect 17744 34788 17800 34790
rect 17824 34788 17880 34790
rect 17904 34788 17960 34790
rect 17984 34788 18040 34790
rect 17744 33754 17800 33756
rect 17824 33754 17880 33756
rect 17904 33754 17960 33756
rect 17984 33754 18040 33756
rect 17744 33702 17790 33754
rect 17790 33702 17800 33754
rect 17824 33702 17854 33754
rect 17854 33702 17866 33754
rect 17866 33702 17880 33754
rect 17904 33702 17918 33754
rect 17918 33702 17930 33754
rect 17930 33702 17960 33754
rect 17984 33702 17994 33754
rect 17994 33702 18040 33754
rect 17744 33700 17800 33702
rect 17824 33700 17880 33702
rect 17904 33700 17960 33702
rect 17984 33700 18040 33702
rect 17744 32666 17800 32668
rect 17824 32666 17880 32668
rect 17904 32666 17960 32668
rect 17984 32666 18040 32668
rect 17744 32614 17790 32666
rect 17790 32614 17800 32666
rect 17824 32614 17854 32666
rect 17854 32614 17866 32666
rect 17866 32614 17880 32666
rect 17904 32614 17918 32666
rect 17918 32614 17930 32666
rect 17930 32614 17960 32666
rect 17984 32614 17994 32666
rect 17994 32614 18040 32666
rect 17744 32612 17800 32614
rect 17824 32612 17880 32614
rect 17904 32612 17960 32614
rect 17984 32612 18040 32614
rect 9350 22874 9406 22876
rect 9430 22874 9486 22876
rect 9510 22874 9566 22876
rect 9590 22874 9646 22876
rect 9350 22822 9396 22874
rect 9396 22822 9406 22874
rect 9430 22822 9460 22874
rect 9460 22822 9472 22874
rect 9472 22822 9486 22874
rect 9510 22822 9524 22874
rect 9524 22822 9536 22874
rect 9536 22822 9566 22874
rect 9590 22822 9600 22874
rect 9600 22822 9646 22874
rect 9350 22820 9406 22822
rect 9430 22820 9486 22822
rect 9510 22820 9566 22822
rect 9590 22820 9646 22822
rect 9350 21786 9406 21788
rect 9430 21786 9486 21788
rect 9510 21786 9566 21788
rect 9590 21786 9646 21788
rect 9350 21734 9396 21786
rect 9396 21734 9406 21786
rect 9430 21734 9460 21786
rect 9460 21734 9472 21786
rect 9472 21734 9486 21786
rect 9510 21734 9524 21786
rect 9524 21734 9536 21786
rect 9536 21734 9566 21786
rect 9590 21734 9600 21786
rect 9600 21734 9646 21786
rect 9350 21732 9406 21734
rect 9430 21732 9486 21734
rect 9510 21732 9566 21734
rect 9590 21732 9646 21734
rect 9350 20698 9406 20700
rect 9430 20698 9486 20700
rect 9510 20698 9566 20700
rect 9590 20698 9646 20700
rect 9350 20646 9396 20698
rect 9396 20646 9406 20698
rect 9430 20646 9460 20698
rect 9460 20646 9472 20698
rect 9472 20646 9486 20698
rect 9510 20646 9524 20698
rect 9524 20646 9536 20698
rect 9536 20646 9566 20698
rect 9590 20646 9600 20698
rect 9600 20646 9646 20698
rect 9350 20644 9406 20646
rect 9430 20644 9486 20646
rect 9510 20644 9566 20646
rect 9590 20644 9646 20646
rect 9350 19610 9406 19612
rect 9430 19610 9486 19612
rect 9510 19610 9566 19612
rect 9590 19610 9646 19612
rect 9350 19558 9396 19610
rect 9396 19558 9406 19610
rect 9430 19558 9460 19610
rect 9460 19558 9472 19610
rect 9472 19558 9486 19610
rect 9510 19558 9524 19610
rect 9524 19558 9536 19610
rect 9536 19558 9566 19610
rect 9590 19558 9600 19610
rect 9600 19558 9646 19610
rect 9350 19556 9406 19558
rect 9430 19556 9486 19558
rect 9510 19556 9566 19558
rect 9590 19556 9646 19558
rect 9678 18708 9680 18728
rect 9680 18708 9732 18728
rect 9732 18708 9734 18728
rect 9678 18672 9734 18708
rect 9350 18522 9406 18524
rect 9430 18522 9486 18524
rect 9510 18522 9566 18524
rect 9590 18522 9646 18524
rect 9350 18470 9396 18522
rect 9396 18470 9406 18522
rect 9430 18470 9460 18522
rect 9460 18470 9472 18522
rect 9472 18470 9486 18522
rect 9510 18470 9524 18522
rect 9524 18470 9536 18522
rect 9536 18470 9566 18522
rect 9590 18470 9600 18522
rect 9600 18470 9646 18522
rect 9350 18468 9406 18470
rect 9430 18468 9486 18470
rect 9510 18468 9566 18470
rect 9590 18468 9646 18470
rect 8942 17756 8944 17776
rect 8944 17756 8996 17776
rect 8996 17756 8998 17776
rect 8942 17720 8998 17756
rect 9310 17720 9366 17776
rect 8850 16632 8906 16688
rect 8758 16360 8814 16416
rect 8758 16224 8814 16280
rect 8574 16088 8630 16144
rect 8574 14728 8630 14784
rect 8390 11600 8446 11656
rect 8390 11500 8392 11520
rect 8392 11500 8444 11520
rect 8444 11500 8446 11520
rect 8390 11464 8446 11500
rect 8574 10920 8630 10976
rect 9350 17434 9406 17436
rect 9430 17434 9486 17436
rect 9510 17434 9566 17436
rect 9590 17434 9646 17436
rect 9350 17382 9396 17434
rect 9396 17382 9406 17434
rect 9430 17382 9460 17434
rect 9460 17382 9472 17434
rect 9472 17382 9486 17434
rect 9510 17382 9524 17434
rect 9524 17382 9536 17434
rect 9536 17382 9566 17434
rect 9590 17382 9600 17434
rect 9600 17382 9646 17434
rect 9350 17380 9406 17382
rect 9430 17380 9486 17382
rect 9510 17380 9566 17382
rect 9590 17380 9646 17382
rect 9310 16768 9366 16824
rect 9402 16532 9404 16552
rect 9404 16532 9456 16552
rect 9456 16532 9458 16552
rect 9402 16496 9458 16532
rect 9350 16346 9406 16348
rect 9430 16346 9486 16348
rect 9510 16346 9566 16348
rect 9590 16346 9646 16348
rect 9350 16294 9396 16346
rect 9396 16294 9406 16346
rect 9430 16294 9460 16346
rect 9460 16294 9472 16346
rect 9472 16294 9486 16346
rect 9510 16294 9524 16346
rect 9524 16294 9536 16346
rect 9536 16294 9566 16346
rect 9590 16294 9600 16346
rect 9600 16294 9646 16346
rect 9350 16292 9406 16294
rect 9430 16292 9486 16294
rect 9510 16292 9566 16294
rect 9590 16292 9646 16294
rect 9218 15952 9274 16008
rect 9678 15544 9734 15600
rect 9770 15272 9826 15328
rect 9350 15258 9406 15260
rect 9430 15258 9486 15260
rect 9510 15258 9566 15260
rect 9590 15258 9646 15260
rect 9350 15206 9396 15258
rect 9396 15206 9406 15258
rect 9430 15206 9460 15258
rect 9460 15206 9472 15258
rect 9472 15206 9486 15258
rect 9510 15206 9524 15258
rect 9524 15206 9536 15258
rect 9536 15206 9566 15258
rect 9590 15206 9600 15258
rect 9600 15206 9646 15258
rect 9350 15204 9406 15206
rect 9430 15204 9486 15206
rect 9510 15204 9566 15206
rect 9590 15204 9646 15206
rect 9350 14170 9406 14172
rect 9430 14170 9486 14172
rect 9510 14170 9566 14172
rect 9590 14170 9646 14172
rect 9350 14118 9396 14170
rect 9396 14118 9406 14170
rect 9430 14118 9460 14170
rect 9460 14118 9472 14170
rect 9472 14118 9486 14170
rect 9510 14118 9524 14170
rect 9524 14118 9536 14170
rect 9536 14118 9566 14170
rect 9590 14118 9600 14170
rect 9600 14118 9646 14170
rect 9350 14116 9406 14118
rect 9430 14116 9486 14118
rect 9510 14116 9566 14118
rect 9590 14116 9646 14118
rect 9350 13082 9406 13084
rect 9430 13082 9486 13084
rect 9510 13082 9566 13084
rect 9590 13082 9646 13084
rect 9350 13030 9396 13082
rect 9396 13030 9406 13082
rect 9430 13030 9460 13082
rect 9460 13030 9472 13082
rect 9472 13030 9486 13082
rect 9510 13030 9524 13082
rect 9524 13030 9536 13082
rect 9536 13030 9566 13082
rect 9590 13030 9600 13082
rect 9600 13030 9646 13082
rect 9350 13028 9406 13030
rect 9430 13028 9486 13030
rect 9510 13028 9566 13030
rect 9590 13028 9646 13030
rect 9310 12416 9366 12472
rect 9350 11994 9406 11996
rect 9430 11994 9486 11996
rect 9510 11994 9566 11996
rect 9590 11994 9646 11996
rect 9350 11942 9396 11994
rect 9396 11942 9406 11994
rect 9430 11942 9460 11994
rect 9460 11942 9472 11994
rect 9472 11942 9486 11994
rect 9510 11942 9524 11994
rect 9524 11942 9536 11994
rect 9536 11942 9566 11994
rect 9590 11942 9600 11994
rect 9600 11942 9646 11994
rect 9350 11940 9406 11942
rect 9430 11940 9486 11942
rect 9510 11940 9566 11942
rect 9590 11940 9646 11942
rect 9402 11600 9458 11656
rect 9770 11464 9826 11520
rect 9126 11328 9182 11384
rect 5153 9274 5209 9276
rect 5233 9274 5289 9276
rect 5313 9274 5369 9276
rect 5393 9274 5449 9276
rect 5153 9222 5199 9274
rect 5199 9222 5209 9274
rect 5233 9222 5263 9274
rect 5263 9222 5275 9274
rect 5275 9222 5289 9274
rect 5313 9222 5327 9274
rect 5327 9222 5339 9274
rect 5339 9222 5369 9274
rect 5393 9222 5403 9274
rect 5403 9222 5449 9274
rect 5153 9220 5209 9222
rect 5233 9220 5289 9222
rect 5313 9220 5369 9222
rect 5393 9220 5449 9222
rect 9350 10906 9406 10908
rect 9430 10906 9486 10908
rect 9510 10906 9566 10908
rect 9590 10906 9646 10908
rect 9350 10854 9396 10906
rect 9396 10854 9406 10906
rect 9430 10854 9460 10906
rect 9460 10854 9472 10906
rect 9472 10854 9486 10906
rect 9510 10854 9524 10906
rect 9524 10854 9536 10906
rect 9536 10854 9566 10906
rect 9590 10854 9600 10906
rect 9600 10854 9646 10906
rect 9350 10852 9406 10854
rect 9430 10852 9486 10854
rect 9510 10852 9566 10854
rect 9590 10852 9646 10854
rect 9350 9818 9406 9820
rect 9430 9818 9486 9820
rect 9510 9818 9566 9820
rect 9590 9818 9646 9820
rect 9350 9766 9396 9818
rect 9396 9766 9406 9818
rect 9430 9766 9460 9818
rect 9460 9766 9472 9818
rect 9472 9766 9486 9818
rect 9510 9766 9524 9818
rect 9524 9766 9536 9818
rect 9536 9766 9566 9818
rect 9590 9766 9600 9818
rect 9600 9766 9646 9818
rect 9350 9764 9406 9766
rect 9430 9764 9486 9766
rect 9510 9764 9566 9766
rect 9590 9764 9646 9766
rect 10322 11872 10378 11928
rect 10414 11772 10416 11792
rect 10416 11772 10468 11792
rect 10468 11772 10470 11792
rect 10414 11736 10470 11772
rect 10046 11328 10102 11384
rect 12254 20304 12310 20360
rect 11978 19760 12034 19816
rect 11702 19372 11758 19408
rect 11702 19352 11704 19372
rect 11704 19352 11756 19372
rect 11756 19352 11758 19372
rect 11518 15580 11520 15600
rect 11520 15580 11572 15600
rect 11572 15580 11574 15600
rect 11518 15544 11574 15580
rect 11242 13912 11298 13968
rect 11242 13368 11298 13424
rect 12070 18692 12126 18728
rect 12070 18672 12072 18692
rect 12072 18672 12124 18692
rect 12124 18672 12126 18692
rect 11794 16088 11850 16144
rect 10874 9696 10930 9752
rect 11886 15020 11942 15056
rect 13547 29946 13603 29948
rect 13627 29946 13683 29948
rect 13707 29946 13763 29948
rect 13787 29946 13843 29948
rect 13547 29894 13593 29946
rect 13593 29894 13603 29946
rect 13627 29894 13657 29946
rect 13657 29894 13669 29946
rect 13669 29894 13683 29946
rect 13707 29894 13721 29946
rect 13721 29894 13733 29946
rect 13733 29894 13763 29946
rect 13787 29894 13797 29946
rect 13797 29894 13843 29946
rect 13547 29892 13603 29894
rect 13627 29892 13683 29894
rect 13707 29892 13763 29894
rect 13787 29892 13843 29894
rect 13547 28858 13603 28860
rect 13627 28858 13683 28860
rect 13707 28858 13763 28860
rect 13787 28858 13843 28860
rect 13547 28806 13593 28858
rect 13593 28806 13603 28858
rect 13627 28806 13657 28858
rect 13657 28806 13669 28858
rect 13669 28806 13683 28858
rect 13707 28806 13721 28858
rect 13721 28806 13733 28858
rect 13733 28806 13763 28858
rect 13787 28806 13797 28858
rect 13797 28806 13843 28858
rect 13547 28804 13603 28806
rect 13627 28804 13683 28806
rect 13707 28804 13763 28806
rect 13787 28804 13843 28806
rect 13547 27770 13603 27772
rect 13627 27770 13683 27772
rect 13707 27770 13763 27772
rect 13787 27770 13843 27772
rect 13547 27718 13593 27770
rect 13593 27718 13603 27770
rect 13627 27718 13657 27770
rect 13657 27718 13669 27770
rect 13669 27718 13683 27770
rect 13707 27718 13721 27770
rect 13721 27718 13733 27770
rect 13733 27718 13763 27770
rect 13787 27718 13797 27770
rect 13797 27718 13843 27770
rect 13547 27716 13603 27718
rect 13627 27716 13683 27718
rect 13707 27716 13763 27718
rect 13787 27716 13843 27718
rect 13547 26682 13603 26684
rect 13627 26682 13683 26684
rect 13707 26682 13763 26684
rect 13787 26682 13843 26684
rect 13547 26630 13593 26682
rect 13593 26630 13603 26682
rect 13627 26630 13657 26682
rect 13657 26630 13669 26682
rect 13669 26630 13683 26682
rect 13707 26630 13721 26682
rect 13721 26630 13733 26682
rect 13733 26630 13763 26682
rect 13787 26630 13797 26682
rect 13797 26630 13843 26682
rect 13547 26628 13603 26630
rect 13627 26628 13683 26630
rect 13707 26628 13763 26630
rect 13787 26628 13843 26630
rect 13547 25594 13603 25596
rect 13627 25594 13683 25596
rect 13707 25594 13763 25596
rect 13787 25594 13843 25596
rect 13547 25542 13593 25594
rect 13593 25542 13603 25594
rect 13627 25542 13657 25594
rect 13657 25542 13669 25594
rect 13669 25542 13683 25594
rect 13707 25542 13721 25594
rect 13721 25542 13733 25594
rect 13733 25542 13763 25594
rect 13787 25542 13797 25594
rect 13797 25542 13843 25594
rect 13547 25540 13603 25542
rect 13627 25540 13683 25542
rect 13707 25540 13763 25542
rect 13787 25540 13843 25542
rect 13547 24506 13603 24508
rect 13627 24506 13683 24508
rect 13707 24506 13763 24508
rect 13787 24506 13843 24508
rect 13547 24454 13593 24506
rect 13593 24454 13603 24506
rect 13627 24454 13657 24506
rect 13657 24454 13669 24506
rect 13669 24454 13683 24506
rect 13707 24454 13721 24506
rect 13721 24454 13733 24506
rect 13733 24454 13763 24506
rect 13787 24454 13797 24506
rect 13797 24454 13843 24506
rect 13547 24452 13603 24454
rect 13627 24452 13683 24454
rect 13707 24452 13763 24454
rect 13787 24452 13843 24454
rect 13547 23418 13603 23420
rect 13627 23418 13683 23420
rect 13707 23418 13763 23420
rect 13787 23418 13843 23420
rect 13547 23366 13593 23418
rect 13593 23366 13603 23418
rect 13627 23366 13657 23418
rect 13657 23366 13669 23418
rect 13669 23366 13683 23418
rect 13707 23366 13721 23418
rect 13721 23366 13733 23418
rect 13733 23366 13763 23418
rect 13787 23366 13797 23418
rect 13797 23366 13843 23418
rect 13547 23364 13603 23366
rect 13627 23364 13683 23366
rect 13707 23364 13763 23366
rect 13787 23364 13843 23366
rect 13547 22330 13603 22332
rect 13627 22330 13683 22332
rect 13707 22330 13763 22332
rect 13787 22330 13843 22332
rect 13547 22278 13593 22330
rect 13593 22278 13603 22330
rect 13627 22278 13657 22330
rect 13657 22278 13669 22330
rect 13669 22278 13683 22330
rect 13707 22278 13721 22330
rect 13721 22278 13733 22330
rect 13733 22278 13763 22330
rect 13787 22278 13797 22330
rect 13797 22278 13843 22330
rect 13547 22276 13603 22278
rect 13627 22276 13683 22278
rect 13707 22276 13763 22278
rect 13787 22276 13843 22278
rect 13547 21242 13603 21244
rect 13627 21242 13683 21244
rect 13707 21242 13763 21244
rect 13787 21242 13843 21244
rect 13547 21190 13593 21242
rect 13593 21190 13603 21242
rect 13627 21190 13657 21242
rect 13657 21190 13669 21242
rect 13669 21190 13683 21242
rect 13707 21190 13721 21242
rect 13721 21190 13733 21242
rect 13733 21190 13763 21242
rect 13787 21190 13797 21242
rect 13797 21190 13843 21242
rect 13547 21188 13603 21190
rect 13627 21188 13683 21190
rect 13707 21188 13763 21190
rect 13787 21188 13843 21190
rect 12898 19352 12954 19408
rect 13547 20154 13603 20156
rect 13627 20154 13683 20156
rect 13707 20154 13763 20156
rect 13787 20154 13843 20156
rect 13547 20102 13593 20154
rect 13593 20102 13603 20154
rect 13627 20102 13657 20154
rect 13657 20102 13669 20154
rect 13669 20102 13683 20154
rect 13707 20102 13721 20154
rect 13721 20102 13733 20154
rect 13733 20102 13763 20154
rect 13787 20102 13797 20154
rect 13797 20102 13843 20154
rect 13547 20100 13603 20102
rect 13627 20100 13683 20102
rect 13707 20100 13763 20102
rect 13787 20100 13843 20102
rect 12162 15272 12218 15328
rect 11886 15000 11888 15020
rect 11888 15000 11940 15020
rect 11940 15000 11942 15020
rect 13547 19066 13603 19068
rect 13627 19066 13683 19068
rect 13707 19066 13763 19068
rect 13787 19066 13843 19068
rect 13547 19014 13593 19066
rect 13593 19014 13603 19066
rect 13627 19014 13657 19066
rect 13657 19014 13669 19066
rect 13669 19014 13683 19066
rect 13707 19014 13721 19066
rect 13721 19014 13733 19066
rect 13733 19014 13763 19066
rect 13787 19014 13797 19066
rect 13797 19014 13843 19066
rect 13547 19012 13603 19014
rect 13627 19012 13683 19014
rect 13707 19012 13763 19014
rect 13787 19012 13843 19014
rect 12806 14864 12862 14920
rect 11886 11892 11942 11928
rect 11886 11872 11888 11892
rect 11888 11872 11940 11892
rect 11940 11872 11942 11892
rect 11886 11756 11942 11792
rect 11886 11736 11888 11756
rect 11888 11736 11940 11756
rect 11940 11736 11942 11756
rect 12162 9560 12218 9616
rect 13547 17978 13603 17980
rect 13627 17978 13683 17980
rect 13707 17978 13763 17980
rect 13787 17978 13843 17980
rect 13547 17926 13593 17978
rect 13593 17926 13603 17978
rect 13627 17926 13657 17978
rect 13657 17926 13669 17978
rect 13669 17926 13683 17978
rect 13707 17926 13721 17978
rect 13721 17926 13733 17978
rect 13733 17926 13763 17978
rect 13787 17926 13797 17978
rect 13797 17926 13843 17978
rect 13547 17924 13603 17926
rect 13627 17924 13683 17926
rect 13707 17924 13763 17926
rect 13787 17924 13843 17926
rect 13547 16890 13603 16892
rect 13627 16890 13683 16892
rect 13707 16890 13763 16892
rect 13787 16890 13843 16892
rect 13547 16838 13593 16890
rect 13593 16838 13603 16890
rect 13627 16838 13657 16890
rect 13657 16838 13669 16890
rect 13669 16838 13683 16890
rect 13707 16838 13721 16890
rect 13721 16838 13733 16890
rect 13733 16838 13763 16890
rect 13787 16838 13797 16890
rect 13797 16838 13843 16890
rect 13547 16836 13603 16838
rect 13627 16836 13683 16838
rect 13707 16836 13763 16838
rect 13787 16836 13843 16838
rect 13547 15802 13603 15804
rect 13627 15802 13683 15804
rect 13707 15802 13763 15804
rect 13787 15802 13843 15804
rect 13547 15750 13593 15802
rect 13593 15750 13603 15802
rect 13627 15750 13657 15802
rect 13657 15750 13669 15802
rect 13669 15750 13683 15802
rect 13707 15750 13721 15802
rect 13721 15750 13733 15802
rect 13733 15750 13763 15802
rect 13787 15750 13797 15802
rect 13797 15750 13843 15802
rect 13547 15748 13603 15750
rect 13627 15748 13683 15750
rect 13707 15748 13763 15750
rect 13787 15748 13843 15750
rect 12714 12180 12716 12200
rect 12716 12180 12768 12200
rect 12768 12180 12770 12200
rect 12714 12144 12770 12180
rect 12530 11092 12532 11112
rect 12532 11092 12584 11112
rect 12584 11092 12586 11112
rect 12530 11056 12586 11092
rect 13174 11872 13230 11928
rect 13450 15020 13506 15056
rect 13450 15000 13452 15020
rect 13452 15000 13504 15020
rect 13504 15000 13506 15020
rect 13547 14714 13603 14716
rect 13627 14714 13683 14716
rect 13707 14714 13763 14716
rect 13787 14714 13843 14716
rect 13547 14662 13593 14714
rect 13593 14662 13603 14714
rect 13627 14662 13657 14714
rect 13657 14662 13669 14714
rect 13669 14662 13683 14714
rect 13707 14662 13721 14714
rect 13721 14662 13733 14714
rect 13733 14662 13763 14714
rect 13787 14662 13797 14714
rect 13797 14662 13843 14714
rect 13547 14660 13603 14662
rect 13627 14660 13683 14662
rect 13707 14660 13763 14662
rect 13787 14660 13843 14662
rect 13358 13948 13360 13968
rect 13360 13948 13412 13968
rect 13412 13948 13414 13968
rect 13358 13912 13414 13948
rect 13547 13626 13603 13628
rect 13627 13626 13683 13628
rect 13707 13626 13763 13628
rect 13787 13626 13843 13628
rect 13547 13574 13593 13626
rect 13593 13574 13603 13626
rect 13627 13574 13657 13626
rect 13657 13574 13669 13626
rect 13669 13574 13683 13626
rect 13707 13574 13721 13626
rect 13721 13574 13733 13626
rect 13733 13574 13763 13626
rect 13787 13574 13797 13626
rect 13797 13574 13843 13626
rect 13547 13572 13603 13574
rect 13627 13572 13683 13574
rect 13707 13572 13763 13574
rect 13787 13572 13843 13574
rect 13547 12538 13603 12540
rect 13627 12538 13683 12540
rect 13707 12538 13763 12540
rect 13787 12538 13843 12540
rect 13547 12486 13593 12538
rect 13593 12486 13603 12538
rect 13627 12486 13657 12538
rect 13657 12486 13669 12538
rect 13669 12486 13683 12538
rect 13707 12486 13721 12538
rect 13721 12486 13733 12538
rect 13733 12486 13763 12538
rect 13787 12486 13797 12538
rect 13797 12486 13843 12538
rect 13547 12484 13603 12486
rect 13627 12484 13683 12486
rect 13707 12484 13763 12486
rect 13787 12484 13843 12486
rect 12438 9696 12494 9752
rect 13726 11872 13782 11928
rect 13547 11450 13603 11452
rect 13627 11450 13683 11452
rect 13707 11450 13763 11452
rect 13787 11450 13843 11452
rect 13547 11398 13593 11450
rect 13593 11398 13603 11450
rect 13627 11398 13657 11450
rect 13657 11398 13669 11450
rect 13669 11398 13683 11450
rect 13707 11398 13721 11450
rect 13721 11398 13733 11450
rect 13733 11398 13763 11450
rect 13787 11398 13797 11450
rect 13797 11398 13843 11450
rect 13547 11396 13603 11398
rect 13627 11396 13683 11398
rect 13707 11396 13763 11398
rect 13787 11396 13843 11398
rect 17744 31578 17800 31580
rect 17824 31578 17880 31580
rect 17904 31578 17960 31580
rect 17984 31578 18040 31580
rect 17744 31526 17790 31578
rect 17790 31526 17800 31578
rect 17824 31526 17854 31578
rect 17854 31526 17866 31578
rect 17866 31526 17880 31578
rect 17904 31526 17918 31578
rect 17918 31526 17930 31578
rect 17930 31526 17960 31578
rect 17984 31526 17994 31578
rect 17994 31526 18040 31578
rect 17744 31524 17800 31526
rect 17824 31524 17880 31526
rect 17904 31524 17960 31526
rect 17984 31524 18040 31526
rect 17744 30490 17800 30492
rect 17824 30490 17880 30492
rect 17904 30490 17960 30492
rect 17984 30490 18040 30492
rect 17744 30438 17790 30490
rect 17790 30438 17800 30490
rect 17824 30438 17854 30490
rect 17854 30438 17866 30490
rect 17866 30438 17880 30490
rect 17904 30438 17918 30490
rect 17918 30438 17930 30490
rect 17930 30438 17960 30490
rect 17984 30438 17994 30490
rect 17994 30438 18040 30490
rect 17744 30436 17800 30438
rect 17824 30436 17880 30438
rect 17904 30436 17960 30438
rect 17984 30436 18040 30438
rect 17744 29402 17800 29404
rect 17824 29402 17880 29404
rect 17904 29402 17960 29404
rect 17984 29402 18040 29404
rect 17744 29350 17790 29402
rect 17790 29350 17800 29402
rect 17824 29350 17854 29402
rect 17854 29350 17866 29402
rect 17866 29350 17880 29402
rect 17904 29350 17918 29402
rect 17918 29350 17930 29402
rect 17930 29350 17960 29402
rect 17984 29350 17994 29402
rect 17994 29350 18040 29402
rect 17744 29348 17800 29350
rect 17824 29348 17880 29350
rect 17904 29348 17960 29350
rect 17984 29348 18040 29350
rect 21941 34298 21997 34300
rect 22021 34298 22077 34300
rect 22101 34298 22157 34300
rect 22181 34298 22237 34300
rect 21941 34246 21987 34298
rect 21987 34246 21997 34298
rect 22021 34246 22051 34298
rect 22051 34246 22063 34298
rect 22063 34246 22077 34298
rect 22101 34246 22115 34298
rect 22115 34246 22127 34298
rect 22127 34246 22157 34298
rect 22181 34246 22191 34298
rect 22191 34246 22237 34298
rect 21941 34244 21997 34246
rect 22021 34244 22077 34246
rect 22101 34244 22157 34246
rect 22181 34244 22237 34246
rect 21941 33210 21997 33212
rect 22021 33210 22077 33212
rect 22101 33210 22157 33212
rect 22181 33210 22237 33212
rect 21941 33158 21987 33210
rect 21987 33158 21997 33210
rect 22021 33158 22051 33210
rect 22051 33158 22063 33210
rect 22063 33158 22077 33210
rect 22101 33158 22115 33210
rect 22115 33158 22127 33210
rect 22127 33158 22157 33210
rect 22181 33158 22191 33210
rect 22191 33158 22237 33210
rect 21941 33156 21997 33158
rect 22021 33156 22077 33158
rect 22101 33156 22157 33158
rect 22181 33156 22237 33158
rect 21941 32122 21997 32124
rect 22021 32122 22077 32124
rect 22101 32122 22157 32124
rect 22181 32122 22237 32124
rect 21941 32070 21987 32122
rect 21987 32070 21997 32122
rect 22021 32070 22051 32122
rect 22051 32070 22063 32122
rect 22063 32070 22077 32122
rect 22101 32070 22115 32122
rect 22115 32070 22127 32122
rect 22127 32070 22157 32122
rect 22181 32070 22191 32122
rect 22191 32070 22237 32122
rect 21941 32068 21997 32070
rect 22021 32068 22077 32070
rect 22101 32068 22157 32070
rect 22181 32068 22237 32070
rect 26138 34842 26194 34844
rect 26218 34842 26274 34844
rect 26298 34842 26354 34844
rect 26378 34842 26434 34844
rect 26138 34790 26184 34842
rect 26184 34790 26194 34842
rect 26218 34790 26248 34842
rect 26248 34790 26260 34842
rect 26260 34790 26274 34842
rect 26298 34790 26312 34842
rect 26312 34790 26324 34842
rect 26324 34790 26354 34842
rect 26378 34790 26388 34842
rect 26388 34790 26434 34842
rect 26138 34788 26194 34790
rect 26218 34788 26274 34790
rect 26298 34788 26354 34790
rect 26378 34788 26434 34790
rect 34532 34842 34588 34844
rect 34612 34842 34668 34844
rect 34692 34842 34748 34844
rect 34772 34842 34828 34844
rect 34532 34790 34578 34842
rect 34578 34790 34588 34842
rect 34612 34790 34642 34842
rect 34642 34790 34654 34842
rect 34654 34790 34668 34842
rect 34692 34790 34706 34842
rect 34706 34790 34718 34842
rect 34718 34790 34748 34842
rect 34772 34790 34782 34842
rect 34782 34790 34828 34842
rect 34532 34788 34588 34790
rect 34612 34788 34668 34790
rect 34692 34788 34748 34790
rect 34772 34788 34828 34790
rect 31022 34584 31078 34640
rect 30335 34298 30391 34300
rect 30415 34298 30471 34300
rect 30495 34298 30551 34300
rect 30575 34298 30631 34300
rect 30335 34246 30381 34298
rect 30381 34246 30391 34298
rect 30415 34246 30445 34298
rect 30445 34246 30457 34298
rect 30457 34246 30471 34298
rect 30495 34246 30509 34298
rect 30509 34246 30521 34298
rect 30521 34246 30551 34298
rect 30575 34246 30585 34298
rect 30585 34246 30631 34298
rect 30335 34244 30391 34246
rect 30415 34244 30471 34246
rect 30495 34244 30551 34246
rect 30575 34244 30631 34246
rect 21941 31034 21997 31036
rect 22021 31034 22077 31036
rect 22101 31034 22157 31036
rect 22181 31034 22237 31036
rect 21941 30982 21987 31034
rect 21987 30982 21997 31034
rect 22021 30982 22051 31034
rect 22051 30982 22063 31034
rect 22063 30982 22077 31034
rect 22101 30982 22115 31034
rect 22115 30982 22127 31034
rect 22127 30982 22157 31034
rect 22181 30982 22191 31034
rect 22191 30982 22237 31034
rect 21941 30980 21997 30982
rect 22021 30980 22077 30982
rect 22101 30980 22157 30982
rect 22181 30980 22237 30982
rect 21941 29946 21997 29948
rect 22021 29946 22077 29948
rect 22101 29946 22157 29948
rect 22181 29946 22237 29948
rect 21941 29894 21987 29946
rect 21987 29894 21997 29946
rect 22021 29894 22051 29946
rect 22051 29894 22063 29946
rect 22063 29894 22077 29946
rect 22101 29894 22115 29946
rect 22115 29894 22127 29946
rect 22127 29894 22157 29946
rect 22181 29894 22191 29946
rect 22191 29894 22237 29946
rect 21941 29892 21997 29894
rect 22021 29892 22077 29894
rect 22101 29892 22157 29894
rect 22181 29892 22237 29894
rect 21941 28858 21997 28860
rect 22021 28858 22077 28860
rect 22101 28858 22157 28860
rect 22181 28858 22237 28860
rect 21941 28806 21987 28858
rect 21987 28806 21997 28858
rect 22021 28806 22051 28858
rect 22051 28806 22063 28858
rect 22063 28806 22077 28858
rect 22101 28806 22115 28858
rect 22115 28806 22127 28858
rect 22127 28806 22157 28858
rect 22181 28806 22191 28858
rect 22191 28806 22237 28858
rect 21941 28804 21997 28806
rect 22021 28804 22077 28806
rect 22101 28804 22157 28806
rect 22181 28804 22237 28806
rect 17744 28314 17800 28316
rect 17824 28314 17880 28316
rect 17904 28314 17960 28316
rect 17984 28314 18040 28316
rect 17744 28262 17790 28314
rect 17790 28262 17800 28314
rect 17824 28262 17854 28314
rect 17854 28262 17866 28314
rect 17866 28262 17880 28314
rect 17904 28262 17918 28314
rect 17918 28262 17930 28314
rect 17930 28262 17960 28314
rect 17984 28262 17994 28314
rect 17994 28262 18040 28314
rect 17744 28260 17800 28262
rect 17824 28260 17880 28262
rect 17904 28260 17960 28262
rect 17984 28260 18040 28262
rect 26138 33754 26194 33756
rect 26218 33754 26274 33756
rect 26298 33754 26354 33756
rect 26378 33754 26434 33756
rect 26138 33702 26184 33754
rect 26184 33702 26194 33754
rect 26218 33702 26248 33754
rect 26248 33702 26260 33754
rect 26260 33702 26274 33754
rect 26298 33702 26312 33754
rect 26312 33702 26324 33754
rect 26324 33702 26354 33754
rect 26378 33702 26388 33754
rect 26388 33702 26434 33754
rect 26138 33700 26194 33702
rect 26218 33700 26274 33702
rect 26298 33700 26354 33702
rect 26378 33700 26434 33702
rect 26138 32666 26194 32668
rect 26218 32666 26274 32668
rect 26298 32666 26354 32668
rect 26378 32666 26434 32668
rect 26138 32614 26184 32666
rect 26184 32614 26194 32666
rect 26218 32614 26248 32666
rect 26248 32614 26260 32666
rect 26260 32614 26274 32666
rect 26298 32614 26312 32666
rect 26312 32614 26324 32666
rect 26324 32614 26354 32666
rect 26378 32614 26388 32666
rect 26388 32614 26434 32666
rect 26138 32612 26194 32614
rect 26218 32612 26274 32614
rect 26298 32612 26354 32614
rect 26378 32612 26434 32614
rect 30335 33210 30391 33212
rect 30415 33210 30471 33212
rect 30495 33210 30551 33212
rect 30575 33210 30631 33212
rect 30335 33158 30381 33210
rect 30381 33158 30391 33210
rect 30415 33158 30445 33210
rect 30445 33158 30457 33210
rect 30457 33158 30471 33210
rect 30495 33158 30509 33210
rect 30509 33158 30521 33210
rect 30521 33158 30551 33210
rect 30575 33158 30585 33210
rect 30585 33158 30631 33210
rect 30335 33156 30391 33158
rect 30415 33156 30471 33158
rect 30495 33156 30551 33158
rect 30575 33156 30631 33158
rect 26138 31578 26194 31580
rect 26218 31578 26274 31580
rect 26298 31578 26354 31580
rect 26378 31578 26434 31580
rect 26138 31526 26184 31578
rect 26184 31526 26194 31578
rect 26218 31526 26248 31578
rect 26248 31526 26260 31578
rect 26260 31526 26274 31578
rect 26298 31526 26312 31578
rect 26312 31526 26324 31578
rect 26324 31526 26354 31578
rect 26378 31526 26388 31578
rect 26388 31526 26434 31578
rect 26138 31524 26194 31526
rect 26218 31524 26274 31526
rect 26298 31524 26354 31526
rect 26378 31524 26434 31526
rect 26138 30490 26194 30492
rect 26218 30490 26274 30492
rect 26298 30490 26354 30492
rect 26378 30490 26434 30492
rect 26138 30438 26184 30490
rect 26184 30438 26194 30490
rect 26218 30438 26248 30490
rect 26248 30438 26260 30490
rect 26260 30438 26274 30490
rect 26298 30438 26312 30490
rect 26312 30438 26324 30490
rect 26324 30438 26354 30490
rect 26378 30438 26388 30490
rect 26388 30438 26434 30490
rect 26138 30436 26194 30438
rect 26218 30436 26274 30438
rect 26298 30436 26354 30438
rect 26378 30436 26434 30438
rect 17744 27226 17800 27228
rect 17824 27226 17880 27228
rect 17904 27226 17960 27228
rect 17984 27226 18040 27228
rect 17744 27174 17790 27226
rect 17790 27174 17800 27226
rect 17824 27174 17854 27226
rect 17854 27174 17866 27226
rect 17866 27174 17880 27226
rect 17904 27174 17918 27226
rect 17918 27174 17930 27226
rect 17930 27174 17960 27226
rect 17984 27174 17994 27226
rect 17994 27174 18040 27226
rect 17744 27172 17800 27174
rect 17824 27172 17880 27174
rect 17904 27172 17960 27174
rect 17984 27172 18040 27174
rect 21941 27770 21997 27772
rect 22021 27770 22077 27772
rect 22101 27770 22157 27772
rect 22181 27770 22237 27772
rect 21941 27718 21987 27770
rect 21987 27718 21997 27770
rect 22021 27718 22051 27770
rect 22051 27718 22063 27770
rect 22063 27718 22077 27770
rect 22101 27718 22115 27770
rect 22115 27718 22127 27770
rect 22127 27718 22157 27770
rect 22181 27718 22191 27770
rect 22191 27718 22237 27770
rect 21941 27716 21997 27718
rect 22021 27716 22077 27718
rect 22101 27716 22157 27718
rect 22181 27716 22237 27718
rect 17744 26138 17800 26140
rect 17824 26138 17880 26140
rect 17904 26138 17960 26140
rect 17984 26138 18040 26140
rect 17744 26086 17790 26138
rect 17790 26086 17800 26138
rect 17824 26086 17854 26138
rect 17854 26086 17866 26138
rect 17866 26086 17880 26138
rect 17904 26086 17918 26138
rect 17918 26086 17930 26138
rect 17930 26086 17960 26138
rect 17984 26086 17994 26138
rect 17994 26086 18040 26138
rect 17744 26084 17800 26086
rect 17824 26084 17880 26086
rect 17904 26084 17960 26086
rect 17984 26084 18040 26086
rect 21941 26682 21997 26684
rect 22021 26682 22077 26684
rect 22101 26682 22157 26684
rect 22181 26682 22237 26684
rect 21941 26630 21987 26682
rect 21987 26630 21997 26682
rect 22021 26630 22051 26682
rect 22051 26630 22063 26682
rect 22063 26630 22077 26682
rect 22101 26630 22115 26682
rect 22115 26630 22127 26682
rect 22127 26630 22157 26682
rect 22181 26630 22191 26682
rect 22191 26630 22237 26682
rect 21941 26628 21997 26630
rect 22021 26628 22077 26630
rect 22101 26628 22157 26630
rect 22181 26628 22237 26630
rect 17744 25050 17800 25052
rect 17824 25050 17880 25052
rect 17904 25050 17960 25052
rect 17984 25050 18040 25052
rect 17744 24998 17790 25050
rect 17790 24998 17800 25050
rect 17824 24998 17854 25050
rect 17854 24998 17866 25050
rect 17866 24998 17880 25050
rect 17904 24998 17918 25050
rect 17918 24998 17930 25050
rect 17930 24998 17960 25050
rect 17984 24998 17994 25050
rect 17994 24998 18040 25050
rect 17744 24996 17800 24998
rect 17824 24996 17880 24998
rect 17904 24996 17960 24998
rect 17984 24996 18040 24998
rect 17744 23962 17800 23964
rect 17824 23962 17880 23964
rect 17904 23962 17960 23964
rect 17984 23962 18040 23964
rect 17744 23910 17790 23962
rect 17790 23910 17800 23962
rect 17824 23910 17854 23962
rect 17854 23910 17866 23962
rect 17866 23910 17880 23962
rect 17904 23910 17918 23962
rect 17918 23910 17930 23962
rect 17930 23910 17960 23962
rect 17984 23910 17994 23962
rect 17994 23910 18040 23962
rect 17744 23908 17800 23910
rect 17824 23908 17880 23910
rect 17904 23908 17960 23910
rect 17984 23908 18040 23910
rect 17744 22874 17800 22876
rect 17824 22874 17880 22876
rect 17904 22874 17960 22876
rect 17984 22874 18040 22876
rect 17744 22822 17790 22874
rect 17790 22822 17800 22874
rect 17824 22822 17854 22874
rect 17854 22822 17866 22874
rect 17866 22822 17880 22874
rect 17904 22822 17918 22874
rect 17918 22822 17930 22874
rect 17930 22822 17960 22874
rect 17984 22822 17994 22874
rect 17994 22822 18040 22874
rect 17744 22820 17800 22822
rect 17824 22820 17880 22822
rect 17904 22820 17960 22822
rect 17984 22820 18040 22822
rect 14830 15444 14832 15464
rect 14832 15444 14884 15464
rect 14884 15444 14886 15464
rect 14830 15408 14886 15444
rect 13547 10362 13603 10364
rect 13627 10362 13683 10364
rect 13707 10362 13763 10364
rect 13787 10362 13843 10364
rect 13547 10310 13593 10362
rect 13593 10310 13603 10362
rect 13627 10310 13657 10362
rect 13657 10310 13669 10362
rect 13669 10310 13683 10362
rect 13707 10310 13721 10362
rect 13721 10310 13733 10362
rect 13733 10310 13763 10362
rect 13787 10310 13797 10362
rect 13797 10310 13843 10362
rect 13547 10308 13603 10310
rect 13627 10308 13683 10310
rect 13707 10308 13763 10310
rect 13787 10308 13843 10310
rect 13542 9696 13598 9752
rect 13726 9580 13782 9616
rect 13726 9560 13728 9580
rect 13728 9560 13780 9580
rect 13780 9560 13782 9580
rect 13547 9274 13603 9276
rect 13627 9274 13683 9276
rect 13707 9274 13763 9276
rect 13787 9274 13843 9276
rect 13547 9222 13593 9274
rect 13593 9222 13603 9274
rect 13627 9222 13657 9274
rect 13657 9222 13669 9274
rect 13669 9222 13683 9274
rect 13707 9222 13721 9274
rect 13721 9222 13733 9274
rect 13733 9222 13763 9274
rect 13787 9222 13797 9274
rect 13797 9222 13843 9274
rect 13547 9220 13603 9222
rect 13627 9220 13683 9222
rect 13707 9220 13763 9222
rect 13787 9220 13843 9222
rect 9350 8730 9406 8732
rect 9430 8730 9486 8732
rect 9510 8730 9566 8732
rect 9590 8730 9646 8732
rect 9350 8678 9396 8730
rect 9396 8678 9406 8730
rect 9430 8678 9460 8730
rect 9460 8678 9472 8730
rect 9472 8678 9486 8730
rect 9510 8678 9524 8730
rect 9524 8678 9536 8730
rect 9536 8678 9566 8730
rect 9590 8678 9600 8730
rect 9600 8678 9646 8730
rect 9350 8676 9406 8678
rect 9430 8676 9486 8678
rect 9510 8676 9566 8678
rect 9590 8676 9646 8678
rect 5153 8186 5209 8188
rect 5233 8186 5289 8188
rect 5313 8186 5369 8188
rect 5393 8186 5449 8188
rect 5153 8134 5199 8186
rect 5199 8134 5209 8186
rect 5233 8134 5263 8186
rect 5263 8134 5275 8186
rect 5275 8134 5289 8186
rect 5313 8134 5327 8186
rect 5327 8134 5339 8186
rect 5339 8134 5369 8186
rect 5393 8134 5403 8186
rect 5403 8134 5449 8186
rect 5153 8132 5209 8134
rect 5233 8132 5289 8134
rect 5313 8132 5369 8134
rect 5393 8132 5449 8134
rect 13547 8186 13603 8188
rect 13627 8186 13683 8188
rect 13707 8186 13763 8188
rect 13787 8186 13843 8188
rect 13547 8134 13593 8186
rect 13593 8134 13603 8186
rect 13627 8134 13657 8186
rect 13657 8134 13669 8186
rect 13669 8134 13683 8186
rect 13707 8134 13721 8186
rect 13721 8134 13733 8186
rect 13733 8134 13763 8186
rect 13787 8134 13797 8186
rect 13797 8134 13843 8186
rect 13547 8132 13603 8134
rect 13627 8132 13683 8134
rect 13707 8132 13763 8134
rect 13787 8132 13843 8134
rect 9350 7642 9406 7644
rect 9430 7642 9486 7644
rect 9510 7642 9566 7644
rect 9590 7642 9646 7644
rect 9350 7590 9396 7642
rect 9396 7590 9406 7642
rect 9430 7590 9460 7642
rect 9460 7590 9472 7642
rect 9472 7590 9486 7642
rect 9510 7590 9524 7642
rect 9524 7590 9536 7642
rect 9536 7590 9566 7642
rect 9590 7590 9600 7642
rect 9600 7590 9646 7642
rect 9350 7588 9406 7590
rect 9430 7588 9486 7590
rect 9510 7588 9566 7590
rect 9590 7588 9646 7590
rect 15198 9424 15254 9480
rect 15842 9460 15844 9480
rect 15844 9460 15896 9480
rect 15896 9460 15898 9480
rect 5153 7098 5209 7100
rect 5233 7098 5289 7100
rect 5313 7098 5369 7100
rect 5393 7098 5449 7100
rect 5153 7046 5199 7098
rect 5199 7046 5209 7098
rect 5233 7046 5263 7098
rect 5263 7046 5275 7098
rect 5275 7046 5289 7098
rect 5313 7046 5327 7098
rect 5327 7046 5339 7098
rect 5339 7046 5369 7098
rect 5393 7046 5403 7098
rect 5403 7046 5449 7098
rect 5153 7044 5209 7046
rect 5233 7044 5289 7046
rect 5313 7044 5369 7046
rect 5393 7044 5449 7046
rect 9350 6554 9406 6556
rect 9430 6554 9486 6556
rect 9510 6554 9566 6556
rect 9590 6554 9646 6556
rect 9350 6502 9396 6554
rect 9396 6502 9406 6554
rect 9430 6502 9460 6554
rect 9460 6502 9472 6554
rect 9472 6502 9486 6554
rect 9510 6502 9524 6554
rect 9524 6502 9536 6554
rect 9536 6502 9566 6554
rect 9590 6502 9600 6554
rect 9600 6502 9646 6554
rect 9350 6500 9406 6502
rect 9430 6500 9486 6502
rect 9510 6500 9566 6502
rect 9590 6500 9646 6502
rect 13547 7098 13603 7100
rect 13627 7098 13683 7100
rect 13707 7098 13763 7100
rect 13787 7098 13843 7100
rect 13547 7046 13593 7098
rect 13593 7046 13603 7098
rect 13627 7046 13657 7098
rect 13657 7046 13669 7098
rect 13669 7046 13683 7098
rect 13707 7046 13721 7098
rect 13721 7046 13733 7098
rect 13733 7046 13763 7098
rect 13787 7046 13797 7098
rect 13797 7046 13843 7098
rect 13547 7044 13603 7046
rect 13627 7044 13683 7046
rect 13707 7044 13763 7046
rect 13787 7044 13843 7046
rect 938 6160 994 6216
rect 5153 6010 5209 6012
rect 5233 6010 5289 6012
rect 5313 6010 5369 6012
rect 5393 6010 5449 6012
rect 5153 5958 5199 6010
rect 5199 5958 5209 6010
rect 5233 5958 5263 6010
rect 5263 5958 5275 6010
rect 5275 5958 5289 6010
rect 5313 5958 5327 6010
rect 5327 5958 5339 6010
rect 5339 5958 5369 6010
rect 5393 5958 5403 6010
rect 5403 5958 5449 6010
rect 5153 5956 5209 5958
rect 5233 5956 5289 5958
rect 5313 5956 5369 5958
rect 5393 5956 5449 5958
rect 5153 4922 5209 4924
rect 5233 4922 5289 4924
rect 5313 4922 5369 4924
rect 5393 4922 5449 4924
rect 5153 4870 5199 4922
rect 5199 4870 5209 4922
rect 5233 4870 5263 4922
rect 5263 4870 5275 4922
rect 5275 4870 5289 4922
rect 5313 4870 5327 4922
rect 5327 4870 5339 4922
rect 5339 4870 5369 4922
rect 5393 4870 5403 4922
rect 5403 4870 5449 4922
rect 5153 4868 5209 4870
rect 5233 4868 5289 4870
rect 5313 4868 5369 4870
rect 5393 4868 5449 4870
rect 5153 3834 5209 3836
rect 5233 3834 5289 3836
rect 5313 3834 5369 3836
rect 5393 3834 5449 3836
rect 5153 3782 5199 3834
rect 5199 3782 5209 3834
rect 5233 3782 5263 3834
rect 5263 3782 5275 3834
rect 5275 3782 5289 3834
rect 5313 3782 5327 3834
rect 5327 3782 5339 3834
rect 5339 3782 5369 3834
rect 5393 3782 5403 3834
rect 5403 3782 5449 3834
rect 5153 3780 5209 3782
rect 5233 3780 5289 3782
rect 5313 3780 5369 3782
rect 5393 3780 5449 3782
rect 5153 2746 5209 2748
rect 5233 2746 5289 2748
rect 5313 2746 5369 2748
rect 5393 2746 5449 2748
rect 5153 2694 5199 2746
rect 5199 2694 5209 2746
rect 5233 2694 5263 2746
rect 5263 2694 5275 2746
rect 5275 2694 5289 2746
rect 5313 2694 5327 2746
rect 5327 2694 5339 2746
rect 5339 2694 5369 2746
rect 5393 2694 5403 2746
rect 5403 2694 5449 2746
rect 5153 2692 5209 2694
rect 5233 2692 5289 2694
rect 5313 2692 5369 2694
rect 5393 2692 5449 2694
rect 9350 5466 9406 5468
rect 9430 5466 9486 5468
rect 9510 5466 9566 5468
rect 9590 5466 9646 5468
rect 9350 5414 9396 5466
rect 9396 5414 9406 5466
rect 9430 5414 9460 5466
rect 9460 5414 9472 5466
rect 9472 5414 9486 5466
rect 9510 5414 9524 5466
rect 9524 5414 9536 5466
rect 9536 5414 9566 5466
rect 9590 5414 9600 5466
rect 9600 5414 9646 5466
rect 9350 5412 9406 5414
rect 9430 5412 9486 5414
rect 9510 5412 9566 5414
rect 9590 5412 9646 5414
rect 9350 4378 9406 4380
rect 9430 4378 9486 4380
rect 9510 4378 9566 4380
rect 9590 4378 9646 4380
rect 9350 4326 9396 4378
rect 9396 4326 9406 4378
rect 9430 4326 9460 4378
rect 9460 4326 9472 4378
rect 9472 4326 9486 4378
rect 9510 4326 9524 4378
rect 9524 4326 9536 4378
rect 9536 4326 9566 4378
rect 9590 4326 9600 4378
rect 9600 4326 9646 4378
rect 9350 4324 9406 4326
rect 9430 4324 9486 4326
rect 9510 4324 9566 4326
rect 9590 4324 9646 4326
rect 9350 3290 9406 3292
rect 9430 3290 9486 3292
rect 9510 3290 9566 3292
rect 9590 3290 9646 3292
rect 9350 3238 9396 3290
rect 9396 3238 9406 3290
rect 9430 3238 9460 3290
rect 9460 3238 9472 3290
rect 9472 3238 9486 3290
rect 9510 3238 9524 3290
rect 9524 3238 9536 3290
rect 9536 3238 9566 3290
rect 9590 3238 9600 3290
rect 9600 3238 9646 3290
rect 9350 3236 9406 3238
rect 9430 3236 9486 3238
rect 9510 3236 9566 3238
rect 9590 3236 9646 3238
rect 13547 6010 13603 6012
rect 13627 6010 13683 6012
rect 13707 6010 13763 6012
rect 13787 6010 13843 6012
rect 13547 5958 13593 6010
rect 13593 5958 13603 6010
rect 13627 5958 13657 6010
rect 13657 5958 13669 6010
rect 13669 5958 13683 6010
rect 13707 5958 13721 6010
rect 13721 5958 13733 6010
rect 13733 5958 13763 6010
rect 13787 5958 13797 6010
rect 13797 5958 13843 6010
rect 13547 5956 13603 5958
rect 13627 5956 13683 5958
rect 13707 5956 13763 5958
rect 13787 5956 13843 5958
rect 15842 9424 15898 9460
rect 17744 21786 17800 21788
rect 17824 21786 17880 21788
rect 17904 21786 17960 21788
rect 17984 21786 18040 21788
rect 17744 21734 17790 21786
rect 17790 21734 17800 21786
rect 17824 21734 17854 21786
rect 17854 21734 17866 21786
rect 17866 21734 17880 21786
rect 17904 21734 17918 21786
rect 17918 21734 17930 21786
rect 17930 21734 17960 21786
rect 17984 21734 17994 21786
rect 17994 21734 18040 21786
rect 17744 21732 17800 21734
rect 17824 21732 17880 21734
rect 17904 21732 17960 21734
rect 17984 21732 18040 21734
rect 17744 20698 17800 20700
rect 17824 20698 17880 20700
rect 17904 20698 17960 20700
rect 17984 20698 18040 20700
rect 17744 20646 17790 20698
rect 17790 20646 17800 20698
rect 17824 20646 17854 20698
rect 17854 20646 17866 20698
rect 17866 20646 17880 20698
rect 17904 20646 17918 20698
rect 17918 20646 17930 20698
rect 17930 20646 17960 20698
rect 17984 20646 17994 20698
rect 17994 20646 18040 20698
rect 17744 20644 17800 20646
rect 17824 20644 17880 20646
rect 17904 20644 17960 20646
rect 17984 20644 18040 20646
rect 17744 19610 17800 19612
rect 17824 19610 17880 19612
rect 17904 19610 17960 19612
rect 17984 19610 18040 19612
rect 17744 19558 17790 19610
rect 17790 19558 17800 19610
rect 17824 19558 17854 19610
rect 17854 19558 17866 19610
rect 17866 19558 17880 19610
rect 17904 19558 17918 19610
rect 17918 19558 17930 19610
rect 17930 19558 17960 19610
rect 17984 19558 17994 19610
rect 17994 19558 18040 19610
rect 17744 19556 17800 19558
rect 17824 19556 17880 19558
rect 17904 19556 17960 19558
rect 17984 19556 18040 19558
rect 17744 18522 17800 18524
rect 17824 18522 17880 18524
rect 17904 18522 17960 18524
rect 17984 18522 18040 18524
rect 17744 18470 17790 18522
rect 17790 18470 17800 18522
rect 17824 18470 17854 18522
rect 17854 18470 17866 18522
rect 17866 18470 17880 18522
rect 17904 18470 17918 18522
rect 17918 18470 17930 18522
rect 17930 18470 17960 18522
rect 17984 18470 17994 18522
rect 17994 18470 18040 18522
rect 17744 18468 17800 18470
rect 17824 18468 17880 18470
rect 17904 18468 17960 18470
rect 17984 18468 18040 18470
rect 13547 4922 13603 4924
rect 13627 4922 13683 4924
rect 13707 4922 13763 4924
rect 13787 4922 13843 4924
rect 13547 4870 13593 4922
rect 13593 4870 13603 4922
rect 13627 4870 13657 4922
rect 13657 4870 13669 4922
rect 13669 4870 13683 4922
rect 13707 4870 13721 4922
rect 13721 4870 13733 4922
rect 13733 4870 13763 4922
rect 13787 4870 13797 4922
rect 13797 4870 13843 4922
rect 13547 4868 13603 4870
rect 13627 4868 13683 4870
rect 13707 4868 13763 4870
rect 13787 4868 13843 4870
rect 13547 3834 13603 3836
rect 13627 3834 13683 3836
rect 13707 3834 13763 3836
rect 13787 3834 13843 3836
rect 13547 3782 13593 3834
rect 13593 3782 13603 3834
rect 13627 3782 13657 3834
rect 13657 3782 13669 3834
rect 13669 3782 13683 3834
rect 13707 3782 13721 3834
rect 13721 3782 13733 3834
rect 13733 3782 13763 3834
rect 13787 3782 13797 3834
rect 13797 3782 13843 3834
rect 13547 3780 13603 3782
rect 13627 3780 13683 3782
rect 13707 3780 13763 3782
rect 13787 3780 13843 3782
rect 13547 2746 13603 2748
rect 13627 2746 13683 2748
rect 13707 2746 13763 2748
rect 13787 2746 13843 2748
rect 13547 2694 13593 2746
rect 13593 2694 13603 2746
rect 13627 2694 13657 2746
rect 13657 2694 13669 2746
rect 13669 2694 13683 2746
rect 13707 2694 13721 2746
rect 13721 2694 13733 2746
rect 13733 2694 13763 2746
rect 13787 2694 13797 2746
rect 13797 2694 13843 2746
rect 13547 2692 13603 2694
rect 13627 2692 13683 2694
rect 13707 2692 13763 2694
rect 13787 2692 13843 2694
rect 17744 17434 17800 17436
rect 17824 17434 17880 17436
rect 17904 17434 17960 17436
rect 17984 17434 18040 17436
rect 17744 17382 17790 17434
rect 17790 17382 17800 17434
rect 17824 17382 17854 17434
rect 17854 17382 17866 17434
rect 17866 17382 17880 17434
rect 17904 17382 17918 17434
rect 17918 17382 17930 17434
rect 17930 17382 17960 17434
rect 17984 17382 17994 17434
rect 17994 17382 18040 17434
rect 17744 17380 17800 17382
rect 17824 17380 17880 17382
rect 17904 17380 17960 17382
rect 17984 17380 18040 17382
rect 17744 16346 17800 16348
rect 17824 16346 17880 16348
rect 17904 16346 17960 16348
rect 17984 16346 18040 16348
rect 17744 16294 17790 16346
rect 17790 16294 17800 16346
rect 17824 16294 17854 16346
rect 17854 16294 17866 16346
rect 17866 16294 17880 16346
rect 17904 16294 17918 16346
rect 17918 16294 17930 16346
rect 17930 16294 17960 16346
rect 17984 16294 17994 16346
rect 17994 16294 18040 16346
rect 17744 16292 17800 16294
rect 17824 16292 17880 16294
rect 17904 16292 17960 16294
rect 17984 16292 18040 16294
rect 17744 15258 17800 15260
rect 17824 15258 17880 15260
rect 17904 15258 17960 15260
rect 17984 15258 18040 15260
rect 17744 15206 17790 15258
rect 17790 15206 17800 15258
rect 17824 15206 17854 15258
rect 17854 15206 17866 15258
rect 17866 15206 17880 15258
rect 17904 15206 17918 15258
rect 17918 15206 17930 15258
rect 17930 15206 17960 15258
rect 17984 15206 17994 15258
rect 17994 15206 18040 15258
rect 17744 15204 17800 15206
rect 17824 15204 17880 15206
rect 17904 15204 17960 15206
rect 17984 15204 18040 15206
rect 17744 14170 17800 14172
rect 17824 14170 17880 14172
rect 17904 14170 17960 14172
rect 17984 14170 18040 14172
rect 17744 14118 17790 14170
rect 17790 14118 17800 14170
rect 17824 14118 17854 14170
rect 17854 14118 17866 14170
rect 17866 14118 17880 14170
rect 17904 14118 17918 14170
rect 17918 14118 17930 14170
rect 17930 14118 17960 14170
rect 17984 14118 17994 14170
rect 17994 14118 18040 14170
rect 17744 14116 17800 14118
rect 17824 14116 17880 14118
rect 17904 14116 17960 14118
rect 17984 14116 18040 14118
rect 17744 13082 17800 13084
rect 17824 13082 17880 13084
rect 17904 13082 17960 13084
rect 17984 13082 18040 13084
rect 17744 13030 17790 13082
rect 17790 13030 17800 13082
rect 17824 13030 17854 13082
rect 17854 13030 17866 13082
rect 17866 13030 17880 13082
rect 17904 13030 17918 13082
rect 17918 13030 17930 13082
rect 17930 13030 17960 13082
rect 17984 13030 17994 13082
rect 17994 13030 18040 13082
rect 17744 13028 17800 13030
rect 17824 13028 17880 13030
rect 17904 13028 17960 13030
rect 17984 13028 18040 13030
rect 17744 11994 17800 11996
rect 17824 11994 17880 11996
rect 17904 11994 17960 11996
rect 17984 11994 18040 11996
rect 17744 11942 17790 11994
rect 17790 11942 17800 11994
rect 17824 11942 17854 11994
rect 17854 11942 17866 11994
rect 17866 11942 17880 11994
rect 17904 11942 17918 11994
rect 17918 11942 17930 11994
rect 17930 11942 17960 11994
rect 17984 11942 17994 11994
rect 17994 11942 18040 11994
rect 17744 11940 17800 11942
rect 17824 11940 17880 11942
rect 17904 11940 17960 11942
rect 17984 11940 18040 11942
rect 17744 10906 17800 10908
rect 17824 10906 17880 10908
rect 17904 10906 17960 10908
rect 17984 10906 18040 10908
rect 17744 10854 17790 10906
rect 17790 10854 17800 10906
rect 17824 10854 17854 10906
rect 17854 10854 17866 10906
rect 17866 10854 17880 10906
rect 17904 10854 17918 10906
rect 17918 10854 17930 10906
rect 17930 10854 17960 10906
rect 17984 10854 17994 10906
rect 17994 10854 18040 10906
rect 17744 10852 17800 10854
rect 17824 10852 17880 10854
rect 17904 10852 17960 10854
rect 17984 10852 18040 10854
rect 17744 9818 17800 9820
rect 17824 9818 17880 9820
rect 17904 9818 17960 9820
rect 17984 9818 18040 9820
rect 17744 9766 17790 9818
rect 17790 9766 17800 9818
rect 17824 9766 17854 9818
rect 17854 9766 17866 9818
rect 17866 9766 17880 9818
rect 17904 9766 17918 9818
rect 17918 9766 17930 9818
rect 17930 9766 17960 9818
rect 17984 9766 17994 9818
rect 17994 9766 18040 9818
rect 17744 9764 17800 9766
rect 17824 9764 17880 9766
rect 17904 9764 17960 9766
rect 17984 9764 18040 9766
rect 17744 8730 17800 8732
rect 17824 8730 17880 8732
rect 17904 8730 17960 8732
rect 17984 8730 18040 8732
rect 17744 8678 17790 8730
rect 17790 8678 17800 8730
rect 17824 8678 17854 8730
rect 17854 8678 17866 8730
rect 17866 8678 17880 8730
rect 17904 8678 17918 8730
rect 17918 8678 17930 8730
rect 17930 8678 17960 8730
rect 17984 8678 17994 8730
rect 17994 8678 18040 8730
rect 17744 8676 17800 8678
rect 17824 8676 17880 8678
rect 17904 8676 17960 8678
rect 17984 8676 18040 8678
rect 17744 7642 17800 7644
rect 17824 7642 17880 7644
rect 17904 7642 17960 7644
rect 17984 7642 18040 7644
rect 17744 7590 17790 7642
rect 17790 7590 17800 7642
rect 17824 7590 17854 7642
rect 17854 7590 17866 7642
rect 17866 7590 17880 7642
rect 17904 7590 17918 7642
rect 17918 7590 17930 7642
rect 17930 7590 17960 7642
rect 17984 7590 17994 7642
rect 17994 7590 18040 7642
rect 17744 7588 17800 7590
rect 17824 7588 17880 7590
rect 17904 7588 17960 7590
rect 17984 7588 18040 7590
rect 21941 25594 21997 25596
rect 22021 25594 22077 25596
rect 22101 25594 22157 25596
rect 22181 25594 22237 25596
rect 21941 25542 21987 25594
rect 21987 25542 21997 25594
rect 22021 25542 22051 25594
rect 22051 25542 22063 25594
rect 22063 25542 22077 25594
rect 22101 25542 22115 25594
rect 22115 25542 22127 25594
rect 22127 25542 22157 25594
rect 22181 25542 22191 25594
rect 22191 25542 22237 25594
rect 21941 25540 21997 25542
rect 22021 25540 22077 25542
rect 22101 25540 22157 25542
rect 22181 25540 22237 25542
rect 21941 24506 21997 24508
rect 22021 24506 22077 24508
rect 22101 24506 22157 24508
rect 22181 24506 22237 24508
rect 21941 24454 21987 24506
rect 21987 24454 21997 24506
rect 22021 24454 22051 24506
rect 22051 24454 22063 24506
rect 22063 24454 22077 24506
rect 22101 24454 22115 24506
rect 22115 24454 22127 24506
rect 22127 24454 22157 24506
rect 22181 24454 22191 24506
rect 22191 24454 22237 24506
rect 21941 24452 21997 24454
rect 22021 24452 22077 24454
rect 22101 24452 22157 24454
rect 22181 24452 22237 24454
rect 21941 23418 21997 23420
rect 22021 23418 22077 23420
rect 22101 23418 22157 23420
rect 22181 23418 22237 23420
rect 21941 23366 21987 23418
rect 21987 23366 21997 23418
rect 22021 23366 22051 23418
rect 22051 23366 22063 23418
rect 22063 23366 22077 23418
rect 22101 23366 22115 23418
rect 22115 23366 22127 23418
rect 22127 23366 22157 23418
rect 22181 23366 22191 23418
rect 22191 23366 22237 23418
rect 21941 23364 21997 23366
rect 22021 23364 22077 23366
rect 22101 23364 22157 23366
rect 22181 23364 22237 23366
rect 21941 22330 21997 22332
rect 22021 22330 22077 22332
rect 22101 22330 22157 22332
rect 22181 22330 22237 22332
rect 21941 22278 21987 22330
rect 21987 22278 21997 22330
rect 22021 22278 22051 22330
rect 22051 22278 22063 22330
rect 22063 22278 22077 22330
rect 22101 22278 22115 22330
rect 22115 22278 22127 22330
rect 22127 22278 22157 22330
rect 22181 22278 22191 22330
rect 22191 22278 22237 22330
rect 21941 22276 21997 22278
rect 22021 22276 22077 22278
rect 22101 22276 22157 22278
rect 22181 22276 22237 22278
rect 19982 15444 19984 15464
rect 19984 15444 20036 15464
rect 20036 15444 20038 15464
rect 19982 15408 20038 15444
rect 21941 21242 21997 21244
rect 22021 21242 22077 21244
rect 22101 21242 22157 21244
rect 22181 21242 22237 21244
rect 21941 21190 21987 21242
rect 21987 21190 21997 21242
rect 22021 21190 22051 21242
rect 22051 21190 22063 21242
rect 22063 21190 22077 21242
rect 22101 21190 22115 21242
rect 22115 21190 22127 21242
rect 22127 21190 22157 21242
rect 22181 21190 22191 21242
rect 22191 21190 22237 21242
rect 21941 21188 21997 21190
rect 22021 21188 22077 21190
rect 22101 21188 22157 21190
rect 22181 21188 22237 21190
rect 21546 20440 21602 20496
rect 21941 20154 21997 20156
rect 22021 20154 22077 20156
rect 22101 20154 22157 20156
rect 22181 20154 22237 20156
rect 21941 20102 21987 20154
rect 21987 20102 21997 20154
rect 22021 20102 22051 20154
rect 22051 20102 22063 20154
rect 22063 20102 22077 20154
rect 22101 20102 22115 20154
rect 22115 20102 22127 20154
rect 22127 20102 22157 20154
rect 22181 20102 22191 20154
rect 22191 20102 22237 20154
rect 21941 20100 21997 20102
rect 22021 20100 22077 20102
rect 22101 20100 22157 20102
rect 22181 20100 22237 20102
rect 21941 19066 21997 19068
rect 22021 19066 22077 19068
rect 22101 19066 22157 19068
rect 22181 19066 22237 19068
rect 21941 19014 21987 19066
rect 21987 19014 21997 19066
rect 22021 19014 22051 19066
rect 22051 19014 22063 19066
rect 22063 19014 22077 19066
rect 22101 19014 22115 19066
rect 22115 19014 22127 19066
rect 22127 19014 22157 19066
rect 22181 19014 22191 19066
rect 22191 19014 22237 19066
rect 21941 19012 21997 19014
rect 22021 19012 22077 19014
rect 22101 19012 22157 19014
rect 22181 19012 22237 19014
rect 21941 17978 21997 17980
rect 22021 17978 22077 17980
rect 22101 17978 22157 17980
rect 22181 17978 22237 17980
rect 21941 17926 21987 17978
rect 21987 17926 21997 17978
rect 22021 17926 22051 17978
rect 22051 17926 22063 17978
rect 22063 17926 22077 17978
rect 22101 17926 22115 17978
rect 22115 17926 22127 17978
rect 22127 17926 22157 17978
rect 22181 17926 22191 17978
rect 22191 17926 22237 17978
rect 21941 17924 21997 17926
rect 22021 17924 22077 17926
rect 22101 17924 22157 17926
rect 22181 17924 22237 17926
rect 21941 16890 21997 16892
rect 22021 16890 22077 16892
rect 22101 16890 22157 16892
rect 22181 16890 22237 16892
rect 21941 16838 21987 16890
rect 21987 16838 21997 16890
rect 22021 16838 22051 16890
rect 22051 16838 22063 16890
rect 22063 16838 22077 16890
rect 22101 16838 22115 16890
rect 22115 16838 22127 16890
rect 22127 16838 22157 16890
rect 22181 16838 22191 16890
rect 22191 16838 22237 16890
rect 21941 16836 21997 16838
rect 22021 16836 22077 16838
rect 22101 16836 22157 16838
rect 22181 16836 22237 16838
rect 21941 15802 21997 15804
rect 22021 15802 22077 15804
rect 22101 15802 22157 15804
rect 22181 15802 22237 15804
rect 21941 15750 21987 15802
rect 21987 15750 21997 15802
rect 22021 15750 22051 15802
rect 22051 15750 22063 15802
rect 22063 15750 22077 15802
rect 22101 15750 22115 15802
rect 22115 15750 22127 15802
rect 22127 15750 22157 15802
rect 22181 15750 22191 15802
rect 22191 15750 22237 15802
rect 21941 15748 21997 15750
rect 22021 15748 22077 15750
rect 22101 15748 22157 15750
rect 22181 15748 22237 15750
rect 20166 9560 20222 9616
rect 17744 6554 17800 6556
rect 17824 6554 17880 6556
rect 17904 6554 17960 6556
rect 17984 6554 18040 6556
rect 17744 6502 17790 6554
rect 17790 6502 17800 6554
rect 17824 6502 17854 6554
rect 17854 6502 17866 6554
rect 17866 6502 17880 6554
rect 17904 6502 17918 6554
rect 17918 6502 17930 6554
rect 17930 6502 17960 6554
rect 17984 6502 17994 6554
rect 17994 6502 18040 6554
rect 17744 6500 17800 6502
rect 17824 6500 17880 6502
rect 17904 6500 17960 6502
rect 17984 6500 18040 6502
rect 17744 5466 17800 5468
rect 17824 5466 17880 5468
rect 17904 5466 17960 5468
rect 17984 5466 18040 5468
rect 17744 5414 17790 5466
rect 17790 5414 17800 5466
rect 17824 5414 17854 5466
rect 17854 5414 17866 5466
rect 17866 5414 17880 5466
rect 17904 5414 17918 5466
rect 17918 5414 17930 5466
rect 17930 5414 17960 5466
rect 17984 5414 17994 5466
rect 17994 5414 18040 5466
rect 17744 5412 17800 5414
rect 17824 5412 17880 5414
rect 17904 5412 17960 5414
rect 17984 5412 18040 5414
rect 17744 4378 17800 4380
rect 17824 4378 17880 4380
rect 17904 4378 17960 4380
rect 17984 4378 18040 4380
rect 17744 4326 17790 4378
rect 17790 4326 17800 4378
rect 17824 4326 17854 4378
rect 17854 4326 17866 4378
rect 17866 4326 17880 4378
rect 17904 4326 17918 4378
rect 17918 4326 17930 4378
rect 17930 4326 17960 4378
rect 17984 4326 17994 4378
rect 17994 4326 18040 4378
rect 17744 4324 17800 4326
rect 17824 4324 17880 4326
rect 17904 4324 17960 4326
rect 17984 4324 18040 4326
rect 21941 14714 21997 14716
rect 22021 14714 22077 14716
rect 22101 14714 22157 14716
rect 22181 14714 22237 14716
rect 21941 14662 21987 14714
rect 21987 14662 21997 14714
rect 22021 14662 22051 14714
rect 22051 14662 22063 14714
rect 22063 14662 22077 14714
rect 22101 14662 22115 14714
rect 22115 14662 22127 14714
rect 22127 14662 22157 14714
rect 22181 14662 22191 14714
rect 22191 14662 22237 14714
rect 21941 14660 21997 14662
rect 22021 14660 22077 14662
rect 22101 14660 22157 14662
rect 22181 14660 22237 14662
rect 21941 13626 21997 13628
rect 22021 13626 22077 13628
rect 22101 13626 22157 13628
rect 22181 13626 22237 13628
rect 21941 13574 21987 13626
rect 21987 13574 21997 13626
rect 22021 13574 22051 13626
rect 22051 13574 22063 13626
rect 22063 13574 22077 13626
rect 22101 13574 22115 13626
rect 22115 13574 22127 13626
rect 22127 13574 22157 13626
rect 22181 13574 22191 13626
rect 22191 13574 22237 13626
rect 21941 13572 21997 13574
rect 22021 13572 22077 13574
rect 22101 13572 22157 13574
rect 22181 13572 22237 13574
rect 21941 12538 21997 12540
rect 22021 12538 22077 12540
rect 22101 12538 22157 12540
rect 22181 12538 22237 12540
rect 21941 12486 21987 12538
rect 21987 12486 21997 12538
rect 22021 12486 22051 12538
rect 22051 12486 22063 12538
rect 22063 12486 22077 12538
rect 22101 12486 22115 12538
rect 22115 12486 22127 12538
rect 22127 12486 22157 12538
rect 22181 12486 22191 12538
rect 22191 12486 22237 12538
rect 21941 12484 21997 12486
rect 22021 12484 22077 12486
rect 22101 12484 22157 12486
rect 22181 12484 22237 12486
rect 26138 29402 26194 29404
rect 26218 29402 26274 29404
rect 26298 29402 26354 29404
rect 26378 29402 26434 29404
rect 26138 29350 26184 29402
rect 26184 29350 26194 29402
rect 26218 29350 26248 29402
rect 26248 29350 26260 29402
rect 26260 29350 26274 29402
rect 26298 29350 26312 29402
rect 26312 29350 26324 29402
rect 26324 29350 26354 29402
rect 26378 29350 26388 29402
rect 26388 29350 26434 29402
rect 26138 29348 26194 29350
rect 26218 29348 26274 29350
rect 26298 29348 26354 29350
rect 26378 29348 26434 29350
rect 25042 26424 25098 26480
rect 26138 28314 26194 28316
rect 26218 28314 26274 28316
rect 26298 28314 26354 28316
rect 26378 28314 26434 28316
rect 26138 28262 26184 28314
rect 26184 28262 26194 28314
rect 26218 28262 26248 28314
rect 26248 28262 26260 28314
rect 26260 28262 26274 28314
rect 26298 28262 26312 28314
rect 26312 28262 26324 28314
rect 26324 28262 26354 28314
rect 26378 28262 26388 28314
rect 26388 28262 26434 28314
rect 26138 28260 26194 28262
rect 26218 28260 26274 28262
rect 26298 28260 26354 28262
rect 26378 28260 26434 28262
rect 26138 27226 26194 27228
rect 26218 27226 26274 27228
rect 26298 27226 26354 27228
rect 26378 27226 26434 27228
rect 26138 27174 26184 27226
rect 26184 27174 26194 27226
rect 26218 27174 26248 27226
rect 26248 27174 26260 27226
rect 26260 27174 26274 27226
rect 26298 27174 26312 27226
rect 26312 27174 26324 27226
rect 26324 27174 26354 27226
rect 26378 27174 26388 27226
rect 26388 27174 26434 27226
rect 26138 27172 26194 27174
rect 26218 27172 26274 27174
rect 26298 27172 26354 27174
rect 26378 27172 26434 27174
rect 26138 26138 26194 26140
rect 26218 26138 26274 26140
rect 26298 26138 26354 26140
rect 26378 26138 26434 26140
rect 26138 26086 26184 26138
rect 26184 26086 26194 26138
rect 26218 26086 26248 26138
rect 26248 26086 26260 26138
rect 26260 26086 26274 26138
rect 26298 26086 26312 26138
rect 26312 26086 26324 26138
rect 26324 26086 26354 26138
rect 26378 26086 26388 26138
rect 26388 26086 26434 26138
rect 26138 26084 26194 26086
rect 26218 26084 26274 26086
rect 26298 26084 26354 26086
rect 26378 26084 26434 26086
rect 26138 25050 26194 25052
rect 26218 25050 26274 25052
rect 26298 25050 26354 25052
rect 26378 25050 26434 25052
rect 26138 24998 26184 25050
rect 26184 24998 26194 25050
rect 26218 24998 26248 25050
rect 26248 24998 26260 25050
rect 26260 24998 26274 25050
rect 26298 24998 26312 25050
rect 26312 24998 26324 25050
rect 26324 24998 26354 25050
rect 26378 24998 26388 25050
rect 26388 24998 26434 25050
rect 26138 24996 26194 24998
rect 26218 24996 26274 24998
rect 26298 24996 26354 24998
rect 26378 24996 26434 24998
rect 24398 20440 24454 20496
rect 22650 15408 22706 15464
rect 21941 11450 21997 11452
rect 22021 11450 22077 11452
rect 22101 11450 22157 11452
rect 22181 11450 22237 11452
rect 21941 11398 21987 11450
rect 21987 11398 21997 11450
rect 22021 11398 22051 11450
rect 22051 11398 22063 11450
rect 22063 11398 22077 11450
rect 22101 11398 22115 11450
rect 22115 11398 22127 11450
rect 22127 11398 22157 11450
rect 22181 11398 22191 11450
rect 22191 11398 22237 11450
rect 21941 11396 21997 11398
rect 22021 11396 22077 11398
rect 22101 11396 22157 11398
rect 22181 11396 22237 11398
rect 23294 15428 23350 15464
rect 23294 15408 23296 15428
rect 23296 15408 23348 15428
rect 23348 15408 23350 15428
rect 26138 23962 26194 23964
rect 26218 23962 26274 23964
rect 26298 23962 26354 23964
rect 26378 23962 26434 23964
rect 26138 23910 26184 23962
rect 26184 23910 26194 23962
rect 26218 23910 26248 23962
rect 26248 23910 26260 23962
rect 26260 23910 26274 23962
rect 26298 23910 26312 23962
rect 26312 23910 26324 23962
rect 26324 23910 26354 23962
rect 26378 23910 26388 23962
rect 26388 23910 26434 23962
rect 26138 23908 26194 23910
rect 26218 23908 26274 23910
rect 26298 23908 26354 23910
rect 26378 23908 26434 23910
rect 26138 22874 26194 22876
rect 26218 22874 26274 22876
rect 26298 22874 26354 22876
rect 26378 22874 26434 22876
rect 26138 22822 26184 22874
rect 26184 22822 26194 22874
rect 26218 22822 26248 22874
rect 26248 22822 26260 22874
rect 26260 22822 26274 22874
rect 26298 22822 26312 22874
rect 26312 22822 26324 22874
rect 26324 22822 26354 22874
rect 26378 22822 26388 22874
rect 26388 22822 26434 22874
rect 26138 22820 26194 22822
rect 26218 22820 26274 22822
rect 26298 22820 26354 22822
rect 26378 22820 26434 22822
rect 26138 21786 26194 21788
rect 26218 21786 26274 21788
rect 26298 21786 26354 21788
rect 26378 21786 26434 21788
rect 26138 21734 26184 21786
rect 26184 21734 26194 21786
rect 26218 21734 26248 21786
rect 26248 21734 26260 21786
rect 26260 21734 26274 21786
rect 26298 21734 26312 21786
rect 26312 21734 26324 21786
rect 26324 21734 26354 21786
rect 26378 21734 26388 21786
rect 26388 21734 26434 21786
rect 26138 21732 26194 21734
rect 26218 21732 26274 21734
rect 26298 21732 26354 21734
rect 26378 21732 26434 21734
rect 30335 32122 30391 32124
rect 30415 32122 30471 32124
rect 30495 32122 30551 32124
rect 30575 32122 30631 32124
rect 30335 32070 30381 32122
rect 30381 32070 30391 32122
rect 30415 32070 30445 32122
rect 30445 32070 30457 32122
rect 30457 32070 30471 32122
rect 30495 32070 30509 32122
rect 30509 32070 30521 32122
rect 30521 32070 30551 32122
rect 30575 32070 30585 32122
rect 30585 32070 30631 32122
rect 30335 32068 30391 32070
rect 30415 32068 30471 32070
rect 30495 32068 30551 32070
rect 30575 32068 30631 32070
rect 30335 31034 30391 31036
rect 30415 31034 30471 31036
rect 30495 31034 30551 31036
rect 30575 31034 30631 31036
rect 30335 30982 30381 31034
rect 30381 30982 30391 31034
rect 30415 30982 30445 31034
rect 30445 30982 30457 31034
rect 30457 30982 30471 31034
rect 30495 30982 30509 31034
rect 30509 30982 30521 31034
rect 30521 30982 30551 31034
rect 30575 30982 30585 31034
rect 30585 30982 30631 31034
rect 30335 30980 30391 30982
rect 30415 30980 30471 30982
rect 30495 30980 30551 30982
rect 30575 30980 30631 30982
rect 30335 29946 30391 29948
rect 30415 29946 30471 29948
rect 30495 29946 30551 29948
rect 30575 29946 30631 29948
rect 30335 29894 30381 29946
rect 30381 29894 30391 29946
rect 30415 29894 30445 29946
rect 30445 29894 30457 29946
rect 30457 29894 30471 29946
rect 30495 29894 30509 29946
rect 30509 29894 30521 29946
rect 30521 29894 30551 29946
rect 30575 29894 30585 29946
rect 30585 29894 30631 29946
rect 30335 29892 30391 29894
rect 30415 29892 30471 29894
rect 30495 29892 30551 29894
rect 30575 29892 30631 29894
rect 26138 20698 26194 20700
rect 26218 20698 26274 20700
rect 26298 20698 26354 20700
rect 26378 20698 26434 20700
rect 26138 20646 26184 20698
rect 26184 20646 26194 20698
rect 26218 20646 26248 20698
rect 26248 20646 26260 20698
rect 26260 20646 26274 20698
rect 26298 20646 26312 20698
rect 26312 20646 26324 20698
rect 26324 20646 26354 20698
rect 26378 20646 26388 20698
rect 26388 20646 26434 20698
rect 26138 20644 26194 20646
rect 26218 20644 26274 20646
rect 26298 20644 26354 20646
rect 26378 20644 26434 20646
rect 26138 19610 26194 19612
rect 26218 19610 26274 19612
rect 26298 19610 26354 19612
rect 26378 19610 26434 19612
rect 26138 19558 26184 19610
rect 26184 19558 26194 19610
rect 26218 19558 26248 19610
rect 26248 19558 26260 19610
rect 26260 19558 26274 19610
rect 26298 19558 26312 19610
rect 26312 19558 26324 19610
rect 26324 19558 26354 19610
rect 26378 19558 26388 19610
rect 26388 19558 26434 19610
rect 26138 19556 26194 19558
rect 26218 19556 26274 19558
rect 26298 19556 26354 19558
rect 26378 19556 26434 19558
rect 26138 18522 26194 18524
rect 26218 18522 26274 18524
rect 26298 18522 26354 18524
rect 26378 18522 26434 18524
rect 26138 18470 26184 18522
rect 26184 18470 26194 18522
rect 26218 18470 26248 18522
rect 26248 18470 26260 18522
rect 26260 18470 26274 18522
rect 26298 18470 26312 18522
rect 26312 18470 26324 18522
rect 26324 18470 26354 18522
rect 26378 18470 26388 18522
rect 26388 18470 26434 18522
rect 26138 18468 26194 18470
rect 26218 18468 26274 18470
rect 26298 18468 26354 18470
rect 26378 18468 26434 18470
rect 30335 28858 30391 28860
rect 30415 28858 30471 28860
rect 30495 28858 30551 28860
rect 30575 28858 30631 28860
rect 30335 28806 30381 28858
rect 30381 28806 30391 28858
rect 30415 28806 30445 28858
rect 30445 28806 30457 28858
rect 30457 28806 30471 28858
rect 30495 28806 30509 28858
rect 30509 28806 30521 28858
rect 30521 28806 30551 28858
rect 30575 28806 30585 28858
rect 30585 28806 30631 28858
rect 30335 28804 30391 28806
rect 30415 28804 30471 28806
rect 30495 28804 30551 28806
rect 30575 28804 30631 28806
rect 30335 27770 30391 27772
rect 30415 27770 30471 27772
rect 30495 27770 30551 27772
rect 30575 27770 30631 27772
rect 30335 27718 30381 27770
rect 30381 27718 30391 27770
rect 30415 27718 30445 27770
rect 30445 27718 30457 27770
rect 30457 27718 30471 27770
rect 30495 27718 30509 27770
rect 30509 27718 30521 27770
rect 30521 27718 30551 27770
rect 30575 27718 30585 27770
rect 30585 27718 30631 27770
rect 30335 27716 30391 27718
rect 30415 27716 30471 27718
rect 30495 27716 30551 27718
rect 30575 27716 30631 27718
rect 26138 17434 26194 17436
rect 26218 17434 26274 17436
rect 26298 17434 26354 17436
rect 26378 17434 26434 17436
rect 26138 17382 26184 17434
rect 26184 17382 26194 17434
rect 26218 17382 26248 17434
rect 26248 17382 26260 17434
rect 26260 17382 26274 17434
rect 26298 17382 26312 17434
rect 26312 17382 26324 17434
rect 26324 17382 26354 17434
rect 26378 17382 26388 17434
rect 26388 17382 26434 17434
rect 26138 17380 26194 17382
rect 26218 17380 26274 17382
rect 26298 17380 26354 17382
rect 26378 17380 26434 17382
rect 26138 16346 26194 16348
rect 26218 16346 26274 16348
rect 26298 16346 26354 16348
rect 26378 16346 26434 16348
rect 26138 16294 26184 16346
rect 26184 16294 26194 16346
rect 26218 16294 26248 16346
rect 26248 16294 26260 16346
rect 26260 16294 26274 16346
rect 26298 16294 26312 16346
rect 26312 16294 26324 16346
rect 26324 16294 26354 16346
rect 26378 16294 26388 16346
rect 26388 16294 26434 16346
rect 26138 16292 26194 16294
rect 26218 16292 26274 16294
rect 26298 16292 26354 16294
rect 26378 16292 26434 16294
rect 26138 15258 26194 15260
rect 26218 15258 26274 15260
rect 26298 15258 26354 15260
rect 26378 15258 26434 15260
rect 26138 15206 26184 15258
rect 26184 15206 26194 15258
rect 26218 15206 26248 15258
rect 26248 15206 26260 15258
rect 26260 15206 26274 15258
rect 26298 15206 26312 15258
rect 26312 15206 26324 15258
rect 26324 15206 26354 15258
rect 26378 15206 26388 15258
rect 26388 15206 26434 15258
rect 26138 15204 26194 15206
rect 26218 15204 26274 15206
rect 26298 15204 26354 15206
rect 26378 15204 26434 15206
rect 30335 26682 30391 26684
rect 30415 26682 30471 26684
rect 30495 26682 30551 26684
rect 30575 26682 30631 26684
rect 30335 26630 30381 26682
rect 30381 26630 30391 26682
rect 30415 26630 30445 26682
rect 30445 26630 30457 26682
rect 30457 26630 30471 26682
rect 30495 26630 30509 26682
rect 30509 26630 30521 26682
rect 30521 26630 30551 26682
rect 30575 26630 30585 26682
rect 30585 26630 30631 26682
rect 30335 26628 30391 26630
rect 30415 26628 30471 26630
rect 30495 26628 30551 26630
rect 30575 26628 30631 26630
rect 30335 25594 30391 25596
rect 30415 25594 30471 25596
rect 30495 25594 30551 25596
rect 30575 25594 30631 25596
rect 30335 25542 30381 25594
rect 30381 25542 30391 25594
rect 30415 25542 30445 25594
rect 30445 25542 30457 25594
rect 30457 25542 30471 25594
rect 30495 25542 30509 25594
rect 30509 25542 30521 25594
rect 30521 25542 30551 25594
rect 30575 25542 30585 25594
rect 30585 25542 30631 25594
rect 30335 25540 30391 25542
rect 30415 25540 30471 25542
rect 30495 25540 30551 25542
rect 30575 25540 30631 25542
rect 30335 24506 30391 24508
rect 30415 24506 30471 24508
rect 30495 24506 30551 24508
rect 30575 24506 30631 24508
rect 30335 24454 30381 24506
rect 30381 24454 30391 24506
rect 30415 24454 30445 24506
rect 30445 24454 30457 24506
rect 30457 24454 30471 24506
rect 30495 24454 30509 24506
rect 30509 24454 30521 24506
rect 30521 24454 30551 24506
rect 30575 24454 30585 24506
rect 30585 24454 30631 24506
rect 30335 24452 30391 24454
rect 30415 24452 30471 24454
rect 30495 24452 30551 24454
rect 30575 24452 30631 24454
rect 30335 23418 30391 23420
rect 30415 23418 30471 23420
rect 30495 23418 30551 23420
rect 30575 23418 30631 23420
rect 30335 23366 30381 23418
rect 30381 23366 30391 23418
rect 30415 23366 30445 23418
rect 30445 23366 30457 23418
rect 30457 23366 30471 23418
rect 30495 23366 30509 23418
rect 30509 23366 30521 23418
rect 30521 23366 30551 23418
rect 30575 23366 30585 23418
rect 30585 23366 30631 23418
rect 30335 23364 30391 23366
rect 30415 23364 30471 23366
rect 30495 23364 30551 23366
rect 30575 23364 30631 23366
rect 21941 10362 21997 10364
rect 22021 10362 22077 10364
rect 22101 10362 22157 10364
rect 22181 10362 22237 10364
rect 21941 10310 21987 10362
rect 21987 10310 21997 10362
rect 22021 10310 22051 10362
rect 22051 10310 22063 10362
rect 22063 10310 22077 10362
rect 22101 10310 22115 10362
rect 22115 10310 22127 10362
rect 22127 10310 22157 10362
rect 22181 10310 22191 10362
rect 22191 10310 22237 10362
rect 21941 10308 21997 10310
rect 22021 10308 22077 10310
rect 22101 10308 22157 10310
rect 22181 10308 22237 10310
rect 21941 9274 21997 9276
rect 22021 9274 22077 9276
rect 22101 9274 22157 9276
rect 22181 9274 22237 9276
rect 21941 9222 21987 9274
rect 21987 9222 21997 9274
rect 22021 9222 22051 9274
rect 22051 9222 22063 9274
rect 22063 9222 22077 9274
rect 22101 9222 22115 9274
rect 22115 9222 22127 9274
rect 22127 9222 22157 9274
rect 22181 9222 22191 9274
rect 22191 9222 22237 9274
rect 21941 9220 21997 9222
rect 22021 9220 22077 9222
rect 22101 9220 22157 9222
rect 22181 9220 22237 9222
rect 21941 8186 21997 8188
rect 22021 8186 22077 8188
rect 22101 8186 22157 8188
rect 22181 8186 22237 8188
rect 21941 8134 21987 8186
rect 21987 8134 21997 8186
rect 22021 8134 22051 8186
rect 22051 8134 22063 8186
rect 22063 8134 22077 8186
rect 22101 8134 22115 8186
rect 22115 8134 22127 8186
rect 22127 8134 22157 8186
rect 22181 8134 22191 8186
rect 22191 8134 22237 8186
rect 21941 8132 21997 8134
rect 22021 8132 22077 8134
rect 22101 8132 22157 8134
rect 22181 8132 22237 8134
rect 22558 9596 22560 9616
rect 22560 9596 22612 9616
rect 22612 9596 22614 9616
rect 22558 9560 22614 9596
rect 21941 7098 21997 7100
rect 22021 7098 22077 7100
rect 22101 7098 22157 7100
rect 22181 7098 22237 7100
rect 21941 7046 21987 7098
rect 21987 7046 21997 7098
rect 22021 7046 22051 7098
rect 22051 7046 22063 7098
rect 22063 7046 22077 7098
rect 22101 7046 22115 7098
rect 22115 7046 22127 7098
rect 22127 7046 22157 7098
rect 22181 7046 22191 7098
rect 22191 7046 22237 7098
rect 21941 7044 21997 7046
rect 22021 7044 22077 7046
rect 22101 7044 22157 7046
rect 22181 7044 22237 7046
rect 21941 6010 21997 6012
rect 22021 6010 22077 6012
rect 22101 6010 22157 6012
rect 22181 6010 22237 6012
rect 21941 5958 21987 6010
rect 21987 5958 21997 6010
rect 22021 5958 22051 6010
rect 22051 5958 22063 6010
rect 22063 5958 22077 6010
rect 22101 5958 22115 6010
rect 22115 5958 22127 6010
rect 22127 5958 22157 6010
rect 22181 5958 22191 6010
rect 22191 5958 22237 6010
rect 21941 5956 21997 5958
rect 22021 5956 22077 5958
rect 22101 5956 22157 5958
rect 22181 5956 22237 5958
rect 21941 4922 21997 4924
rect 22021 4922 22077 4924
rect 22101 4922 22157 4924
rect 22181 4922 22237 4924
rect 21941 4870 21987 4922
rect 21987 4870 21997 4922
rect 22021 4870 22051 4922
rect 22051 4870 22063 4922
rect 22063 4870 22077 4922
rect 22101 4870 22115 4922
rect 22115 4870 22127 4922
rect 22127 4870 22157 4922
rect 22181 4870 22191 4922
rect 22191 4870 22237 4922
rect 21941 4868 21997 4870
rect 22021 4868 22077 4870
rect 22101 4868 22157 4870
rect 22181 4868 22237 4870
rect 26138 14170 26194 14172
rect 26218 14170 26274 14172
rect 26298 14170 26354 14172
rect 26378 14170 26434 14172
rect 26138 14118 26184 14170
rect 26184 14118 26194 14170
rect 26218 14118 26248 14170
rect 26248 14118 26260 14170
rect 26260 14118 26274 14170
rect 26298 14118 26312 14170
rect 26312 14118 26324 14170
rect 26324 14118 26354 14170
rect 26378 14118 26388 14170
rect 26388 14118 26434 14170
rect 26138 14116 26194 14118
rect 26218 14116 26274 14118
rect 26298 14116 26354 14118
rect 26378 14116 26434 14118
rect 26138 13082 26194 13084
rect 26218 13082 26274 13084
rect 26298 13082 26354 13084
rect 26378 13082 26434 13084
rect 26138 13030 26184 13082
rect 26184 13030 26194 13082
rect 26218 13030 26248 13082
rect 26248 13030 26260 13082
rect 26260 13030 26274 13082
rect 26298 13030 26312 13082
rect 26312 13030 26324 13082
rect 26324 13030 26354 13082
rect 26378 13030 26388 13082
rect 26388 13030 26434 13082
rect 26138 13028 26194 13030
rect 26218 13028 26274 13030
rect 26298 13028 26354 13030
rect 26378 13028 26434 13030
rect 26138 11994 26194 11996
rect 26218 11994 26274 11996
rect 26298 11994 26354 11996
rect 26378 11994 26434 11996
rect 26138 11942 26184 11994
rect 26184 11942 26194 11994
rect 26218 11942 26248 11994
rect 26248 11942 26260 11994
rect 26260 11942 26274 11994
rect 26298 11942 26312 11994
rect 26312 11942 26324 11994
rect 26324 11942 26354 11994
rect 26378 11942 26388 11994
rect 26388 11942 26434 11994
rect 26138 11940 26194 11942
rect 26218 11940 26274 11942
rect 26298 11940 26354 11942
rect 26378 11940 26434 11942
rect 26138 10906 26194 10908
rect 26218 10906 26274 10908
rect 26298 10906 26354 10908
rect 26378 10906 26434 10908
rect 26138 10854 26184 10906
rect 26184 10854 26194 10906
rect 26218 10854 26248 10906
rect 26248 10854 26260 10906
rect 26260 10854 26274 10906
rect 26298 10854 26312 10906
rect 26312 10854 26324 10906
rect 26324 10854 26354 10906
rect 26378 10854 26388 10906
rect 26388 10854 26434 10906
rect 26138 10852 26194 10854
rect 26218 10852 26274 10854
rect 26298 10852 26354 10854
rect 26378 10852 26434 10854
rect 26138 9818 26194 9820
rect 26218 9818 26274 9820
rect 26298 9818 26354 9820
rect 26378 9818 26434 9820
rect 26138 9766 26184 9818
rect 26184 9766 26194 9818
rect 26218 9766 26248 9818
rect 26248 9766 26260 9818
rect 26260 9766 26274 9818
rect 26298 9766 26312 9818
rect 26312 9766 26324 9818
rect 26324 9766 26354 9818
rect 26378 9766 26388 9818
rect 26388 9766 26434 9818
rect 26138 9764 26194 9766
rect 26218 9764 26274 9766
rect 26298 9764 26354 9766
rect 26378 9764 26434 9766
rect 26138 8730 26194 8732
rect 26218 8730 26274 8732
rect 26298 8730 26354 8732
rect 26378 8730 26434 8732
rect 26138 8678 26184 8730
rect 26184 8678 26194 8730
rect 26218 8678 26248 8730
rect 26248 8678 26260 8730
rect 26260 8678 26274 8730
rect 26298 8678 26312 8730
rect 26312 8678 26324 8730
rect 26324 8678 26354 8730
rect 26378 8678 26388 8730
rect 26388 8678 26434 8730
rect 26138 8676 26194 8678
rect 26218 8676 26274 8678
rect 26298 8676 26354 8678
rect 26378 8676 26434 8678
rect 26138 7642 26194 7644
rect 26218 7642 26274 7644
rect 26298 7642 26354 7644
rect 26378 7642 26434 7644
rect 26138 7590 26184 7642
rect 26184 7590 26194 7642
rect 26218 7590 26248 7642
rect 26248 7590 26260 7642
rect 26260 7590 26274 7642
rect 26298 7590 26312 7642
rect 26312 7590 26324 7642
rect 26324 7590 26354 7642
rect 26378 7590 26388 7642
rect 26388 7590 26434 7642
rect 26138 7588 26194 7590
rect 26218 7588 26274 7590
rect 26298 7588 26354 7590
rect 26378 7588 26434 7590
rect 26138 6554 26194 6556
rect 26218 6554 26274 6556
rect 26298 6554 26354 6556
rect 26378 6554 26434 6556
rect 26138 6502 26184 6554
rect 26184 6502 26194 6554
rect 26218 6502 26248 6554
rect 26248 6502 26260 6554
rect 26260 6502 26274 6554
rect 26298 6502 26312 6554
rect 26312 6502 26324 6554
rect 26324 6502 26354 6554
rect 26378 6502 26388 6554
rect 26388 6502 26434 6554
rect 26138 6500 26194 6502
rect 26218 6500 26274 6502
rect 26298 6500 26354 6502
rect 26378 6500 26434 6502
rect 26138 5466 26194 5468
rect 26218 5466 26274 5468
rect 26298 5466 26354 5468
rect 26378 5466 26434 5468
rect 26138 5414 26184 5466
rect 26184 5414 26194 5466
rect 26218 5414 26248 5466
rect 26248 5414 26260 5466
rect 26260 5414 26274 5466
rect 26298 5414 26312 5466
rect 26312 5414 26324 5466
rect 26324 5414 26354 5466
rect 26378 5414 26388 5466
rect 26388 5414 26434 5466
rect 26138 5412 26194 5414
rect 26218 5412 26274 5414
rect 26298 5412 26354 5414
rect 26378 5412 26434 5414
rect 26138 4378 26194 4380
rect 26218 4378 26274 4380
rect 26298 4378 26354 4380
rect 26378 4378 26434 4380
rect 26138 4326 26184 4378
rect 26184 4326 26194 4378
rect 26218 4326 26248 4378
rect 26248 4326 26260 4378
rect 26260 4326 26274 4378
rect 26298 4326 26312 4378
rect 26312 4326 26324 4378
rect 26324 4326 26354 4378
rect 26378 4326 26388 4378
rect 26388 4326 26434 4378
rect 26138 4324 26194 4326
rect 26218 4324 26274 4326
rect 26298 4324 26354 4326
rect 26378 4324 26434 4326
rect 30335 22330 30391 22332
rect 30415 22330 30471 22332
rect 30495 22330 30551 22332
rect 30575 22330 30631 22332
rect 30335 22278 30381 22330
rect 30381 22278 30391 22330
rect 30415 22278 30445 22330
rect 30445 22278 30457 22330
rect 30457 22278 30471 22330
rect 30495 22278 30509 22330
rect 30509 22278 30521 22330
rect 30521 22278 30551 22330
rect 30575 22278 30585 22330
rect 30585 22278 30631 22330
rect 30335 22276 30391 22278
rect 30415 22276 30471 22278
rect 30495 22276 30551 22278
rect 30575 22276 30631 22278
rect 30335 21242 30391 21244
rect 30415 21242 30471 21244
rect 30495 21242 30551 21244
rect 30575 21242 30631 21244
rect 30335 21190 30381 21242
rect 30381 21190 30391 21242
rect 30415 21190 30445 21242
rect 30445 21190 30457 21242
rect 30457 21190 30471 21242
rect 30495 21190 30509 21242
rect 30509 21190 30521 21242
rect 30521 21190 30551 21242
rect 30575 21190 30585 21242
rect 30585 21190 30631 21242
rect 30335 21188 30391 21190
rect 30415 21188 30471 21190
rect 30495 21188 30551 21190
rect 30575 21188 30631 21190
rect 30335 20154 30391 20156
rect 30415 20154 30471 20156
rect 30495 20154 30551 20156
rect 30575 20154 30631 20156
rect 30335 20102 30381 20154
rect 30381 20102 30391 20154
rect 30415 20102 30445 20154
rect 30445 20102 30457 20154
rect 30457 20102 30471 20154
rect 30495 20102 30509 20154
rect 30509 20102 30521 20154
rect 30521 20102 30551 20154
rect 30575 20102 30585 20154
rect 30585 20102 30631 20154
rect 30335 20100 30391 20102
rect 30415 20100 30471 20102
rect 30495 20100 30551 20102
rect 30575 20100 30631 20102
rect 30335 19066 30391 19068
rect 30415 19066 30471 19068
rect 30495 19066 30551 19068
rect 30575 19066 30631 19068
rect 30335 19014 30381 19066
rect 30381 19014 30391 19066
rect 30415 19014 30445 19066
rect 30445 19014 30457 19066
rect 30457 19014 30471 19066
rect 30495 19014 30509 19066
rect 30509 19014 30521 19066
rect 30521 19014 30551 19066
rect 30575 19014 30585 19066
rect 30585 19014 30631 19066
rect 30335 19012 30391 19014
rect 30415 19012 30471 19014
rect 30495 19012 30551 19014
rect 30575 19012 30631 19014
rect 30335 17978 30391 17980
rect 30415 17978 30471 17980
rect 30495 17978 30551 17980
rect 30575 17978 30631 17980
rect 30335 17926 30381 17978
rect 30381 17926 30391 17978
rect 30415 17926 30445 17978
rect 30445 17926 30457 17978
rect 30457 17926 30471 17978
rect 30495 17926 30509 17978
rect 30509 17926 30521 17978
rect 30521 17926 30551 17978
rect 30575 17926 30585 17978
rect 30585 17926 30631 17978
rect 30335 17924 30391 17926
rect 30415 17924 30471 17926
rect 30495 17924 30551 17926
rect 30575 17924 30631 17926
rect 30335 16890 30391 16892
rect 30415 16890 30471 16892
rect 30495 16890 30551 16892
rect 30575 16890 30631 16892
rect 30335 16838 30381 16890
rect 30381 16838 30391 16890
rect 30415 16838 30445 16890
rect 30445 16838 30457 16890
rect 30457 16838 30471 16890
rect 30495 16838 30509 16890
rect 30509 16838 30521 16890
rect 30521 16838 30551 16890
rect 30575 16838 30585 16890
rect 30585 16838 30631 16890
rect 30335 16836 30391 16838
rect 30415 16836 30471 16838
rect 30495 16836 30551 16838
rect 30575 16836 30631 16838
rect 30335 15802 30391 15804
rect 30415 15802 30471 15804
rect 30495 15802 30551 15804
rect 30575 15802 30631 15804
rect 30335 15750 30381 15802
rect 30381 15750 30391 15802
rect 30415 15750 30445 15802
rect 30445 15750 30457 15802
rect 30457 15750 30471 15802
rect 30495 15750 30509 15802
rect 30509 15750 30521 15802
rect 30521 15750 30551 15802
rect 30575 15750 30585 15802
rect 30585 15750 30631 15802
rect 30335 15748 30391 15750
rect 30415 15748 30471 15750
rect 30495 15748 30551 15750
rect 30575 15748 30631 15750
rect 34532 33754 34588 33756
rect 34612 33754 34668 33756
rect 34692 33754 34748 33756
rect 34772 33754 34828 33756
rect 34532 33702 34578 33754
rect 34578 33702 34588 33754
rect 34612 33702 34642 33754
rect 34642 33702 34654 33754
rect 34654 33702 34668 33754
rect 34692 33702 34706 33754
rect 34706 33702 34718 33754
rect 34718 33702 34748 33754
rect 34772 33702 34782 33754
rect 34782 33702 34828 33754
rect 34532 33700 34588 33702
rect 34612 33700 34668 33702
rect 34692 33700 34748 33702
rect 34772 33700 34828 33702
rect 34532 32666 34588 32668
rect 34612 32666 34668 32668
rect 34692 32666 34748 32668
rect 34772 32666 34828 32668
rect 34532 32614 34578 32666
rect 34578 32614 34588 32666
rect 34612 32614 34642 32666
rect 34642 32614 34654 32666
rect 34654 32614 34668 32666
rect 34692 32614 34706 32666
rect 34706 32614 34718 32666
rect 34718 32614 34748 32666
rect 34772 32614 34782 32666
rect 34782 32614 34828 32666
rect 34532 32612 34588 32614
rect 34612 32612 34668 32614
rect 34692 32612 34748 32614
rect 34772 32612 34828 32614
rect 34532 31578 34588 31580
rect 34612 31578 34668 31580
rect 34692 31578 34748 31580
rect 34772 31578 34828 31580
rect 34532 31526 34578 31578
rect 34578 31526 34588 31578
rect 34612 31526 34642 31578
rect 34642 31526 34654 31578
rect 34654 31526 34668 31578
rect 34692 31526 34706 31578
rect 34706 31526 34718 31578
rect 34718 31526 34748 31578
rect 34772 31526 34782 31578
rect 34782 31526 34828 31578
rect 34532 31524 34588 31526
rect 34612 31524 34668 31526
rect 34692 31524 34748 31526
rect 34772 31524 34828 31526
rect 34532 30490 34588 30492
rect 34612 30490 34668 30492
rect 34692 30490 34748 30492
rect 34772 30490 34828 30492
rect 34532 30438 34578 30490
rect 34578 30438 34588 30490
rect 34612 30438 34642 30490
rect 34642 30438 34654 30490
rect 34654 30438 34668 30490
rect 34692 30438 34706 30490
rect 34706 30438 34718 30490
rect 34718 30438 34748 30490
rect 34772 30438 34782 30490
rect 34782 30438 34828 30490
rect 34532 30436 34588 30438
rect 34612 30436 34668 30438
rect 34692 30436 34748 30438
rect 34772 30436 34828 30438
rect 34532 29402 34588 29404
rect 34612 29402 34668 29404
rect 34692 29402 34748 29404
rect 34772 29402 34828 29404
rect 34532 29350 34578 29402
rect 34578 29350 34588 29402
rect 34612 29350 34642 29402
rect 34642 29350 34654 29402
rect 34654 29350 34668 29402
rect 34692 29350 34706 29402
rect 34706 29350 34718 29402
rect 34718 29350 34748 29402
rect 34772 29350 34782 29402
rect 34782 29350 34828 29402
rect 34532 29348 34588 29350
rect 34612 29348 34668 29350
rect 34692 29348 34748 29350
rect 34772 29348 34828 29350
rect 34532 28314 34588 28316
rect 34612 28314 34668 28316
rect 34692 28314 34748 28316
rect 34772 28314 34828 28316
rect 34532 28262 34578 28314
rect 34578 28262 34588 28314
rect 34612 28262 34642 28314
rect 34642 28262 34654 28314
rect 34654 28262 34668 28314
rect 34692 28262 34706 28314
rect 34706 28262 34718 28314
rect 34718 28262 34748 28314
rect 34772 28262 34782 28314
rect 34782 28262 34828 28314
rect 34532 28260 34588 28262
rect 34612 28260 34668 28262
rect 34692 28260 34748 28262
rect 34772 28260 34828 28262
rect 34794 27956 34796 27976
rect 34796 27956 34848 27976
rect 34848 27956 34850 27976
rect 34794 27920 34850 27956
rect 32586 26424 32642 26480
rect 34532 27226 34588 27228
rect 34612 27226 34668 27228
rect 34692 27226 34748 27228
rect 34772 27226 34828 27228
rect 34532 27174 34578 27226
rect 34578 27174 34588 27226
rect 34612 27174 34642 27226
rect 34642 27174 34654 27226
rect 34654 27174 34668 27226
rect 34692 27174 34706 27226
rect 34706 27174 34718 27226
rect 34718 27174 34748 27226
rect 34772 27174 34782 27226
rect 34782 27174 34828 27226
rect 34532 27172 34588 27174
rect 34612 27172 34668 27174
rect 34692 27172 34748 27174
rect 34772 27172 34828 27174
rect 34532 26138 34588 26140
rect 34612 26138 34668 26140
rect 34692 26138 34748 26140
rect 34772 26138 34828 26140
rect 34532 26086 34578 26138
rect 34578 26086 34588 26138
rect 34612 26086 34642 26138
rect 34642 26086 34654 26138
rect 34654 26086 34668 26138
rect 34692 26086 34706 26138
rect 34706 26086 34718 26138
rect 34718 26086 34748 26138
rect 34772 26086 34782 26138
rect 34782 26086 34828 26138
rect 34532 26084 34588 26086
rect 34612 26084 34668 26086
rect 34692 26084 34748 26086
rect 34772 26084 34828 26086
rect 30335 14714 30391 14716
rect 30415 14714 30471 14716
rect 30495 14714 30551 14716
rect 30575 14714 30631 14716
rect 30335 14662 30381 14714
rect 30381 14662 30391 14714
rect 30415 14662 30445 14714
rect 30445 14662 30457 14714
rect 30457 14662 30471 14714
rect 30495 14662 30509 14714
rect 30509 14662 30521 14714
rect 30521 14662 30551 14714
rect 30575 14662 30585 14714
rect 30585 14662 30631 14714
rect 30335 14660 30391 14662
rect 30415 14660 30471 14662
rect 30495 14660 30551 14662
rect 30575 14660 30631 14662
rect 30335 13626 30391 13628
rect 30415 13626 30471 13628
rect 30495 13626 30551 13628
rect 30575 13626 30631 13628
rect 30335 13574 30381 13626
rect 30381 13574 30391 13626
rect 30415 13574 30445 13626
rect 30445 13574 30457 13626
rect 30457 13574 30471 13626
rect 30495 13574 30509 13626
rect 30509 13574 30521 13626
rect 30521 13574 30551 13626
rect 30575 13574 30585 13626
rect 30585 13574 30631 13626
rect 30335 13572 30391 13574
rect 30415 13572 30471 13574
rect 30495 13572 30551 13574
rect 30575 13572 30631 13574
rect 30335 12538 30391 12540
rect 30415 12538 30471 12540
rect 30495 12538 30551 12540
rect 30575 12538 30631 12540
rect 30335 12486 30381 12538
rect 30381 12486 30391 12538
rect 30415 12486 30445 12538
rect 30445 12486 30457 12538
rect 30457 12486 30471 12538
rect 30495 12486 30509 12538
rect 30509 12486 30521 12538
rect 30521 12486 30551 12538
rect 30575 12486 30585 12538
rect 30585 12486 30631 12538
rect 30335 12484 30391 12486
rect 30415 12484 30471 12486
rect 30495 12484 30551 12486
rect 30575 12484 30631 12486
rect 30335 11450 30391 11452
rect 30415 11450 30471 11452
rect 30495 11450 30551 11452
rect 30575 11450 30631 11452
rect 30335 11398 30381 11450
rect 30381 11398 30391 11450
rect 30415 11398 30445 11450
rect 30445 11398 30457 11450
rect 30457 11398 30471 11450
rect 30495 11398 30509 11450
rect 30509 11398 30521 11450
rect 30521 11398 30551 11450
rect 30575 11398 30585 11450
rect 30585 11398 30631 11450
rect 30335 11396 30391 11398
rect 30415 11396 30471 11398
rect 30495 11396 30551 11398
rect 30575 11396 30631 11398
rect 30335 10362 30391 10364
rect 30415 10362 30471 10364
rect 30495 10362 30551 10364
rect 30575 10362 30631 10364
rect 30335 10310 30381 10362
rect 30381 10310 30391 10362
rect 30415 10310 30445 10362
rect 30445 10310 30457 10362
rect 30457 10310 30471 10362
rect 30495 10310 30509 10362
rect 30509 10310 30521 10362
rect 30521 10310 30551 10362
rect 30575 10310 30585 10362
rect 30585 10310 30631 10362
rect 30335 10308 30391 10310
rect 30415 10308 30471 10310
rect 30495 10308 30551 10310
rect 30575 10308 30631 10310
rect 30335 9274 30391 9276
rect 30415 9274 30471 9276
rect 30495 9274 30551 9276
rect 30575 9274 30631 9276
rect 30335 9222 30381 9274
rect 30381 9222 30391 9274
rect 30415 9222 30445 9274
rect 30445 9222 30457 9274
rect 30457 9222 30471 9274
rect 30495 9222 30509 9274
rect 30509 9222 30521 9274
rect 30521 9222 30551 9274
rect 30575 9222 30585 9274
rect 30585 9222 30631 9274
rect 30335 9220 30391 9222
rect 30415 9220 30471 9222
rect 30495 9220 30551 9222
rect 30575 9220 30631 9222
rect 30335 8186 30391 8188
rect 30415 8186 30471 8188
rect 30495 8186 30551 8188
rect 30575 8186 30631 8188
rect 30335 8134 30381 8186
rect 30381 8134 30391 8186
rect 30415 8134 30445 8186
rect 30445 8134 30457 8186
rect 30457 8134 30471 8186
rect 30495 8134 30509 8186
rect 30509 8134 30521 8186
rect 30521 8134 30551 8186
rect 30575 8134 30585 8186
rect 30585 8134 30631 8186
rect 30335 8132 30391 8134
rect 30415 8132 30471 8134
rect 30495 8132 30551 8134
rect 30575 8132 30631 8134
rect 30335 7098 30391 7100
rect 30415 7098 30471 7100
rect 30495 7098 30551 7100
rect 30575 7098 30631 7100
rect 30335 7046 30381 7098
rect 30381 7046 30391 7098
rect 30415 7046 30445 7098
rect 30445 7046 30457 7098
rect 30457 7046 30471 7098
rect 30495 7046 30509 7098
rect 30509 7046 30521 7098
rect 30521 7046 30551 7098
rect 30575 7046 30585 7098
rect 30585 7046 30631 7098
rect 30335 7044 30391 7046
rect 30415 7044 30471 7046
rect 30495 7044 30551 7046
rect 30575 7044 30631 7046
rect 30335 6010 30391 6012
rect 30415 6010 30471 6012
rect 30495 6010 30551 6012
rect 30575 6010 30631 6012
rect 30335 5958 30381 6010
rect 30381 5958 30391 6010
rect 30415 5958 30445 6010
rect 30445 5958 30457 6010
rect 30457 5958 30471 6010
rect 30495 5958 30509 6010
rect 30509 5958 30521 6010
rect 30521 5958 30551 6010
rect 30575 5958 30585 6010
rect 30585 5958 30631 6010
rect 30335 5956 30391 5958
rect 30415 5956 30471 5958
rect 30495 5956 30551 5958
rect 30575 5956 30631 5958
rect 34532 25050 34588 25052
rect 34612 25050 34668 25052
rect 34692 25050 34748 25052
rect 34772 25050 34828 25052
rect 34532 24998 34578 25050
rect 34578 24998 34588 25050
rect 34612 24998 34642 25050
rect 34642 24998 34654 25050
rect 34654 24998 34668 25050
rect 34692 24998 34706 25050
rect 34706 24998 34718 25050
rect 34718 24998 34748 25050
rect 34772 24998 34782 25050
rect 34782 24998 34828 25050
rect 34532 24996 34588 24998
rect 34612 24996 34668 24998
rect 34692 24996 34748 24998
rect 34772 24996 34828 24998
rect 34532 23962 34588 23964
rect 34612 23962 34668 23964
rect 34692 23962 34748 23964
rect 34772 23962 34828 23964
rect 34532 23910 34578 23962
rect 34578 23910 34588 23962
rect 34612 23910 34642 23962
rect 34642 23910 34654 23962
rect 34654 23910 34668 23962
rect 34692 23910 34706 23962
rect 34706 23910 34718 23962
rect 34718 23910 34748 23962
rect 34772 23910 34782 23962
rect 34782 23910 34828 23962
rect 34532 23908 34588 23910
rect 34612 23908 34668 23910
rect 34692 23908 34748 23910
rect 34772 23908 34828 23910
rect 34532 22874 34588 22876
rect 34612 22874 34668 22876
rect 34692 22874 34748 22876
rect 34772 22874 34828 22876
rect 34532 22822 34578 22874
rect 34578 22822 34588 22874
rect 34612 22822 34642 22874
rect 34642 22822 34654 22874
rect 34654 22822 34668 22874
rect 34692 22822 34706 22874
rect 34706 22822 34718 22874
rect 34718 22822 34748 22874
rect 34772 22822 34782 22874
rect 34782 22822 34828 22874
rect 34532 22820 34588 22822
rect 34612 22820 34668 22822
rect 34692 22820 34748 22822
rect 34772 22820 34828 22822
rect 34532 21786 34588 21788
rect 34612 21786 34668 21788
rect 34692 21786 34748 21788
rect 34772 21786 34828 21788
rect 34532 21734 34578 21786
rect 34578 21734 34588 21786
rect 34612 21734 34642 21786
rect 34642 21734 34654 21786
rect 34654 21734 34668 21786
rect 34692 21734 34706 21786
rect 34706 21734 34718 21786
rect 34718 21734 34748 21786
rect 34772 21734 34782 21786
rect 34782 21734 34828 21786
rect 34532 21732 34588 21734
rect 34612 21732 34668 21734
rect 34692 21732 34748 21734
rect 34772 21732 34828 21734
rect 34794 21120 34850 21176
rect 34532 20698 34588 20700
rect 34612 20698 34668 20700
rect 34692 20698 34748 20700
rect 34772 20698 34828 20700
rect 34532 20646 34578 20698
rect 34578 20646 34588 20698
rect 34612 20646 34642 20698
rect 34642 20646 34654 20698
rect 34654 20646 34668 20698
rect 34692 20646 34706 20698
rect 34706 20646 34718 20698
rect 34718 20646 34748 20698
rect 34772 20646 34782 20698
rect 34782 20646 34828 20698
rect 34532 20644 34588 20646
rect 34612 20644 34668 20646
rect 34692 20644 34748 20646
rect 34772 20644 34828 20646
rect 34532 19610 34588 19612
rect 34612 19610 34668 19612
rect 34692 19610 34748 19612
rect 34772 19610 34828 19612
rect 34532 19558 34578 19610
rect 34578 19558 34588 19610
rect 34612 19558 34642 19610
rect 34642 19558 34654 19610
rect 34654 19558 34668 19610
rect 34692 19558 34706 19610
rect 34706 19558 34718 19610
rect 34718 19558 34748 19610
rect 34772 19558 34782 19610
rect 34782 19558 34828 19610
rect 34532 19556 34588 19558
rect 34612 19556 34668 19558
rect 34692 19556 34748 19558
rect 34772 19556 34828 19558
rect 34532 18522 34588 18524
rect 34612 18522 34668 18524
rect 34692 18522 34748 18524
rect 34772 18522 34828 18524
rect 34532 18470 34578 18522
rect 34578 18470 34588 18522
rect 34612 18470 34642 18522
rect 34642 18470 34654 18522
rect 34654 18470 34668 18522
rect 34692 18470 34706 18522
rect 34706 18470 34718 18522
rect 34718 18470 34748 18522
rect 34772 18470 34782 18522
rect 34782 18470 34828 18522
rect 34532 18468 34588 18470
rect 34612 18468 34668 18470
rect 34692 18468 34748 18470
rect 34772 18468 34828 18470
rect 34532 17434 34588 17436
rect 34612 17434 34668 17436
rect 34692 17434 34748 17436
rect 34772 17434 34828 17436
rect 34532 17382 34578 17434
rect 34578 17382 34588 17434
rect 34612 17382 34642 17434
rect 34642 17382 34654 17434
rect 34654 17382 34668 17434
rect 34692 17382 34706 17434
rect 34706 17382 34718 17434
rect 34718 17382 34748 17434
rect 34772 17382 34782 17434
rect 34782 17382 34828 17434
rect 34532 17380 34588 17382
rect 34612 17380 34668 17382
rect 34692 17380 34748 17382
rect 34772 17380 34828 17382
rect 34532 16346 34588 16348
rect 34612 16346 34668 16348
rect 34692 16346 34748 16348
rect 34772 16346 34828 16348
rect 34532 16294 34578 16346
rect 34578 16294 34588 16346
rect 34612 16294 34642 16346
rect 34642 16294 34654 16346
rect 34654 16294 34668 16346
rect 34692 16294 34706 16346
rect 34706 16294 34718 16346
rect 34718 16294 34748 16346
rect 34772 16294 34782 16346
rect 34782 16294 34828 16346
rect 34532 16292 34588 16294
rect 34612 16292 34668 16294
rect 34692 16292 34748 16294
rect 34772 16292 34828 16294
rect 34532 15258 34588 15260
rect 34612 15258 34668 15260
rect 34692 15258 34748 15260
rect 34772 15258 34828 15260
rect 34532 15206 34578 15258
rect 34578 15206 34588 15258
rect 34612 15206 34642 15258
rect 34642 15206 34654 15258
rect 34654 15206 34668 15258
rect 34692 15206 34706 15258
rect 34706 15206 34718 15258
rect 34718 15206 34748 15258
rect 34772 15206 34782 15258
rect 34782 15206 34828 15258
rect 34532 15204 34588 15206
rect 34612 15204 34668 15206
rect 34692 15204 34748 15206
rect 34772 15204 34828 15206
rect 34702 14320 34758 14376
rect 34532 14170 34588 14172
rect 34612 14170 34668 14172
rect 34692 14170 34748 14172
rect 34772 14170 34828 14172
rect 34532 14118 34578 14170
rect 34578 14118 34588 14170
rect 34612 14118 34642 14170
rect 34642 14118 34654 14170
rect 34654 14118 34668 14170
rect 34692 14118 34706 14170
rect 34706 14118 34718 14170
rect 34718 14118 34748 14170
rect 34772 14118 34782 14170
rect 34782 14118 34828 14170
rect 34532 14116 34588 14118
rect 34612 14116 34668 14118
rect 34692 14116 34748 14118
rect 34772 14116 34828 14118
rect 34532 13082 34588 13084
rect 34612 13082 34668 13084
rect 34692 13082 34748 13084
rect 34772 13082 34828 13084
rect 34532 13030 34578 13082
rect 34578 13030 34588 13082
rect 34612 13030 34642 13082
rect 34642 13030 34654 13082
rect 34654 13030 34668 13082
rect 34692 13030 34706 13082
rect 34706 13030 34718 13082
rect 34718 13030 34748 13082
rect 34772 13030 34782 13082
rect 34782 13030 34828 13082
rect 34532 13028 34588 13030
rect 34612 13028 34668 13030
rect 34692 13028 34748 13030
rect 34772 13028 34828 13030
rect 34532 11994 34588 11996
rect 34612 11994 34668 11996
rect 34692 11994 34748 11996
rect 34772 11994 34828 11996
rect 34532 11942 34578 11994
rect 34578 11942 34588 11994
rect 34612 11942 34642 11994
rect 34642 11942 34654 11994
rect 34654 11942 34668 11994
rect 34692 11942 34706 11994
rect 34706 11942 34718 11994
rect 34718 11942 34748 11994
rect 34772 11942 34782 11994
rect 34782 11942 34828 11994
rect 34532 11940 34588 11942
rect 34612 11940 34668 11942
rect 34692 11940 34748 11942
rect 34772 11940 34828 11942
rect 34532 10906 34588 10908
rect 34612 10906 34668 10908
rect 34692 10906 34748 10908
rect 34772 10906 34828 10908
rect 34532 10854 34578 10906
rect 34578 10854 34588 10906
rect 34612 10854 34642 10906
rect 34642 10854 34654 10906
rect 34654 10854 34668 10906
rect 34692 10854 34706 10906
rect 34706 10854 34718 10906
rect 34718 10854 34748 10906
rect 34772 10854 34782 10906
rect 34782 10854 34828 10906
rect 34532 10852 34588 10854
rect 34612 10852 34668 10854
rect 34692 10852 34748 10854
rect 34772 10852 34828 10854
rect 34532 9818 34588 9820
rect 34612 9818 34668 9820
rect 34692 9818 34748 9820
rect 34772 9818 34828 9820
rect 34532 9766 34578 9818
rect 34578 9766 34588 9818
rect 34612 9766 34642 9818
rect 34642 9766 34654 9818
rect 34654 9766 34668 9818
rect 34692 9766 34706 9818
rect 34706 9766 34718 9818
rect 34718 9766 34748 9818
rect 34772 9766 34782 9818
rect 34782 9766 34828 9818
rect 34532 9764 34588 9766
rect 34612 9764 34668 9766
rect 34692 9764 34748 9766
rect 34772 9764 34828 9766
rect 34532 8730 34588 8732
rect 34612 8730 34668 8732
rect 34692 8730 34748 8732
rect 34772 8730 34828 8732
rect 34532 8678 34578 8730
rect 34578 8678 34588 8730
rect 34612 8678 34642 8730
rect 34642 8678 34654 8730
rect 34654 8678 34668 8730
rect 34692 8678 34706 8730
rect 34706 8678 34718 8730
rect 34718 8678 34748 8730
rect 34772 8678 34782 8730
rect 34782 8678 34828 8730
rect 34532 8676 34588 8678
rect 34612 8676 34668 8678
rect 34692 8676 34748 8678
rect 34772 8676 34828 8678
rect 34794 8200 34850 8256
rect 30335 4922 30391 4924
rect 30415 4922 30471 4924
rect 30495 4922 30551 4924
rect 30575 4922 30631 4924
rect 30335 4870 30381 4922
rect 30381 4870 30391 4922
rect 30415 4870 30445 4922
rect 30445 4870 30457 4922
rect 30457 4870 30471 4922
rect 30495 4870 30509 4922
rect 30509 4870 30521 4922
rect 30521 4870 30551 4922
rect 30575 4870 30585 4922
rect 30585 4870 30631 4922
rect 30335 4868 30391 4870
rect 30415 4868 30471 4870
rect 30495 4868 30551 4870
rect 30575 4868 30631 4870
rect 34532 7642 34588 7644
rect 34612 7642 34668 7644
rect 34692 7642 34748 7644
rect 34772 7642 34828 7644
rect 34532 7590 34578 7642
rect 34578 7590 34588 7642
rect 34612 7590 34642 7642
rect 34642 7590 34654 7642
rect 34654 7590 34668 7642
rect 34692 7590 34706 7642
rect 34706 7590 34718 7642
rect 34718 7590 34748 7642
rect 34772 7590 34782 7642
rect 34782 7590 34828 7642
rect 34532 7588 34588 7590
rect 34612 7588 34668 7590
rect 34692 7588 34748 7590
rect 34772 7588 34828 7590
rect 34532 6554 34588 6556
rect 34612 6554 34668 6556
rect 34692 6554 34748 6556
rect 34772 6554 34828 6556
rect 34532 6502 34578 6554
rect 34578 6502 34588 6554
rect 34612 6502 34642 6554
rect 34642 6502 34654 6554
rect 34654 6502 34668 6554
rect 34692 6502 34706 6554
rect 34706 6502 34718 6554
rect 34718 6502 34748 6554
rect 34772 6502 34782 6554
rect 34782 6502 34828 6554
rect 34532 6500 34588 6502
rect 34612 6500 34668 6502
rect 34692 6500 34748 6502
rect 34772 6500 34828 6502
rect 34532 5466 34588 5468
rect 34612 5466 34668 5468
rect 34692 5466 34748 5468
rect 34772 5466 34828 5468
rect 34532 5414 34578 5466
rect 34578 5414 34588 5466
rect 34612 5414 34642 5466
rect 34642 5414 34654 5466
rect 34654 5414 34668 5466
rect 34692 5414 34706 5466
rect 34706 5414 34718 5466
rect 34718 5414 34748 5466
rect 34772 5414 34782 5466
rect 34782 5414 34828 5466
rect 34532 5412 34588 5414
rect 34612 5412 34668 5414
rect 34692 5412 34748 5414
rect 34772 5412 34828 5414
rect 34532 4378 34588 4380
rect 34612 4378 34668 4380
rect 34692 4378 34748 4380
rect 34772 4378 34828 4380
rect 34532 4326 34578 4378
rect 34578 4326 34588 4378
rect 34612 4326 34642 4378
rect 34642 4326 34654 4378
rect 34654 4326 34668 4378
rect 34692 4326 34706 4378
rect 34706 4326 34718 4378
rect 34718 4326 34748 4378
rect 34772 4326 34782 4378
rect 34782 4326 34828 4378
rect 34532 4324 34588 4326
rect 34612 4324 34668 4326
rect 34692 4324 34748 4326
rect 34772 4324 34828 4326
rect 21941 3834 21997 3836
rect 22021 3834 22077 3836
rect 22101 3834 22157 3836
rect 22181 3834 22237 3836
rect 21941 3782 21987 3834
rect 21987 3782 21997 3834
rect 22021 3782 22051 3834
rect 22051 3782 22063 3834
rect 22063 3782 22077 3834
rect 22101 3782 22115 3834
rect 22115 3782 22127 3834
rect 22127 3782 22157 3834
rect 22181 3782 22191 3834
rect 22191 3782 22237 3834
rect 21941 3780 21997 3782
rect 22021 3780 22077 3782
rect 22101 3780 22157 3782
rect 22181 3780 22237 3782
rect 30335 3834 30391 3836
rect 30415 3834 30471 3836
rect 30495 3834 30551 3836
rect 30575 3834 30631 3836
rect 30335 3782 30381 3834
rect 30381 3782 30391 3834
rect 30415 3782 30445 3834
rect 30445 3782 30457 3834
rect 30457 3782 30471 3834
rect 30495 3782 30509 3834
rect 30509 3782 30521 3834
rect 30521 3782 30551 3834
rect 30575 3782 30585 3834
rect 30585 3782 30631 3834
rect 30335 3780 30391 3782
rect 30415 3780 30471 3782
rect 30495 3780 30551 3782
rect 30575 3780 30631 3782
rect 17744 3290 17800 3292
rect 17824 3290 17880 3292
rect 17904 3290 17960 3292
rect 17984 3290 18040 3292
rect 17744 3238 17790 3290
rect 17790 3238 17800 3290
rect 17824 3238 17854 3290
rect 17854 3238 17866 3290
rect 17866 3238 17880 3290
rect 17904 3238 17918 3290
rect 17918 3238 17930 3290
rect 17930 3238 17960 3290
rect 17984 3238 17994 3290
rect 17994 3238 18040 3290
rect 17744 3236 17800 3238
rect 17824 3236 17880 3238
rect 17904 3236 17960 3238
rect 17984 3236 18040 3238
rect 21941 2746 21997 2748
rect 22021 2746 22077 2748
rect 22101 2746 22157 2748
rect 22181 2746 22237 2748
rect 21941 2694 21987 2746
rect 21987 2694 21997 2746
rect 22021 2694 22051 2746
rect 22051 2694 22063 2746
rect 22063 2694 22077 2746
rect 22101 2694 22115 2746
rect 22115 2694 22127 2746
rect 22127 2694 22157 2746
rect 22181 2694 22191 2746
rect 22191 2694 22237 2746
rect 21941 2692 21997 2694
rect 22021 2692 22077 2694
rect 22101 2692 22157 2694
rect 22181 2692 22237 2694
rect 26138 3290 26194 3292
rect 26218 3290 26274 3292
rect 26298 3290 26354 3292
rect 26378 3290 26434 3292
rect 26138 3238 26184 3290
rect 26184 3238 26194 3290
rect 26218 3238 26248 3290
rect 26248 3238 26260 3290
rect 26260 3238 26274 3290
rect 26298 3238 26312 3290
rect 26312 3238 26324 3290
rect 26324 3238 26354 3290
rect 26378 3238 26388 3290
rect 26388 3238 26434 3290
rect 26138 3236 26194 3238
rect 26218 3236 26274 3238
rect 26298 3236 26354 3238
rect 26378 3236 26434 3238
rect 30335 2746 30391 2748
rect 30415 2746 30471 2748
rect 30495 2746 30551 2748
rect 30575 2746 30631 2748
rect 30335 2694 30381 2746
rect 30381 2694 30391 2746
rect 30415 2694 30445 2746
rect 30445 2694 30457 2746
rect 30457 2694 30471 2746
rect 30495 2694 30509 2746
rect 30509 2694 30521 2746
rect 30521 2694 30551 2746
rect 30575 2694 30585 2746
rect 30585 2694 30631 2746
rect 30335 2692 30391 2694
rect 30415 2692 30471 2694
rect 30495 2692 30551 2694
rect 30575 2692 30631 2694
rect 34532 3290 34588 3292
rect 34612 3290 34668 3292
rect 34692 3290 34748 3292
rect 34772 3290 34828 3292
rect 34532 3238 34578 3290
rect 34578 3238 34588 3290
rect 34612 3238 34642 3290
rect 34642 3238 34654 3290
rect 34654 3238 34668 3290
rect 34692 3238 34706 3290
rect 34706 3238 34718 3290
rect 34718 3238 34748 3290
rect 34772 3238 34782 3290
rect 34782 3238 34828 3290
rect 34532 3236 34588 3238
rect 34612 3236 34668 3238
rect 34692 3236 34748 3238
rect 34772 3236 34828 3238
rect 9350 2202 9406 2204
rect 9430 2202 9486 2204
rect 9510 2202 9566 2204
rect 9590 2202 9646 2204
rect 9350 2150 9396 2202
rect 9396 2150 9406 2202
rect 9430 2150 9460 2202
rect 9460 2150 9472 2202
rect 9472 2150 9486 2202
rect 9510 2150 9524 2202
rect 9524 2150 9536 2202
rect 9536 2150 9566 2202
rect 9590 2150 9600 2202
rect 9600 2150 9646 2202
rect 9350 2148 9406 2150
rect 9430 2148 9486 2150
rect 9510 2148 9566 2150
rect 9590 2148 9646 2150
rect 17744 2202 17800 2204
rect 17824 2202 17880 2204
rect 17904 2202 17960 2204
rect 17984 2202 18040 2204
rect 17744 2150 17790 2202
rect 17790 2150 17800 2202
rect 17824 2150 17854 2202
rect 17854 2150 17866 2202
rect 17866 2150 17880 2202
rect 17904 2150 17918 2202
rect 17918 2150 17930 2202
rect 17930 2150 17960 2202
rect 17984 2150 17994 2202
rect 17994 2150 18040 2202
rect 17744 2148 17800 2150
rect 17824 2148 17880 2150
rect 17904 2148 17960 2150
rect 17984 2148 18040 2150
rect 26138 2202 26194 2204
rect 26218 2202 26274 2204
rect 26298 2202 26354 2204
rect 26378 2202 26434 2204
rect 26138 2150 26184 2202
rect 26184 2150 26194 2202
rect 26218 2150 26248 2202
rect 26248 2150 26260 2202
rect 26260 2150 26274 2202
rect 26298 2150 26312 2202
rect 26312 2150 26324 2202
rect 26324 2150 26354 2202
rect 26378 2150 26388 2202
rect 26388 2150 26434 2202
rect 26138 2148 26194 2150
rect 26218 2148 26274 2150
rect 26298 2148 26354 2150
rect 26378 2148 26434 2150
rect 34532 2202 34588 2204
rect 34612 2202 34668 2204
rect 34692 2202 34748 2204
rect 34772 2202 34828 2204
rect 34532 2150 34578 2202
rect 34578 2150 34588 2202
rect 34612 2150 34642 2202
rect 34642 2150 34654 2202
rect 34654 2150 34668 2202
rect 34692 2150 34706 2202
rect 34706 2150 34718 2202
rect 34718 2150 34748 2202
rect 34772 2150 34782 2202
rect 34782 2150 34828 2202
rect 34532 2148 34588 2150
rect 34612 2148 34668 2150
rect 34692 2148 34748 2150
rect 34772 2148 34828 2150
rect 34518 1400 34574 1456
<< metal3 >>
rect 5143 35392 5459 35393
rect 5143 35328 5149 35392
rect 5213 35328 5229 35392
rect 5293 35328 5309 35392
rect 5373 35328 5389 35392
rect 5453 35328 5459 35392
rect 5143 35327 5459 35328
rect 13537 35392 13853 35393
rect 13537 35328 13543 35392
rect 13607 35328 13623 35392
rect 13687 35328 13703 35392
rect 13767 35328 13783 35392
rect 13847 35328 13853 35392
rect 13537 35327 13853 35328
rect 21931 35392 22247 35393
rect 21931 35328 21937 35392
rect 22001 35328 22017 35392
rect 22081 35328 22097 35392
rect 22161 35328 22177 35392
rect 22241 35328 22247 35392
rect 21931 35327 22247 35328
rect 30325 35392 30641 35393
rect 30325 35328 30331 35392
rect 30395 35328 30411 35392
rect 30475 35328 30491 35392
rect 30555 35328 30571 35392
rect 30635 35328 30641 35392
rect 30325 35327 30641 35328
rect 9340 34848 9656 34849
rect 9340 34784 9346 34848
rect 9410 34784 9426 34848
rect 9490 34784 9506 34848
rect 9570 34784 9586 34848
rect 9650 34784 9656 34848
rect 9340 34783 9656 34784
rect 17734 34848 18050 34849
rect 17734 34784 17740 34848
rect 17804 34784 17820 34848
rect 17884 34784 17900 34848
rect 17964 34784 17980 34848
rect 18044 34784 18050 34848
rect 17734 34783 18050 34784
rect 26128 34848 26444 34849
rect 26128 34784 26134 34848
rect 26198 34784 26214 34848
rect 26278 34784 26294 34848
rect 26358 34784 26374 34848
rect 26438 34784 26444 34848
rect 26128 34783 26444 34784
rect 34522 34848 34838 34849
rect 34522 34784 34528 34848
rect 34592 34784 34608 34848
rect 34672 34784 34688 34848
rect 34752 34784 34768 34848
rect 34832 34784 34838 34848
rect 34522 34783 34838 34784
rect 35073 34778 35873 34808
rect 35022 34688 35873 34778
rect 31017 34642 31083 34645
rect 35022 34642 35082 34688
rect 31017 34640 35082 34642
rect 31017 34584 31022 34640
rect 31078 34584 35082 34640
rect 31017 34582 35082 34584
rect 31017 34579 31083 34582
rect 5143 34304 5459 34305
rect 5143 34240 5149 34304
rect 5213 34240 5229 34304
rect 5293 34240 5309 34304
rect 5373 34240 5389 34304
rect 5453 34240 5459 34304
rect 5143 34239 5459 34240
rect 13537 34304 13853 34305
rect 13537 34240 13543 34304
rect 13607 34240 13623 34304
rect 13687 34240 13703 34304
rect 13767 34240 13783 34304
rect 13847 34240 13853 34304
rect 13537 34239 13853 34240
rect 21931 34304 22247 34305
rect 21931 34240 21937 34304
rect 22001 34240 22017 34304
rect 22081 34240 22097 34304
rect 22161 34240 22177 34304
rect 22241 34240 22247 34304
rect 21931 34239 22247 34240
rect 30325 34304 30641 34305
rect 30325 34240 30331 34304
rect 30395 34240 30411 34304
rect 30475 34240 30491 34304
rect 30555 34240 30571 34304
rect 30635 34240 30641 34304
rect 30325 34239 30641 34240
rect 9340 33760 9656 33761
rect 9340 33696 9346 33760
rect 9410 33696 9426 33760
rect 9490 33696 9506 33760
rect 9570 33696 9586 33760
rect 9650 33696 9656 33760
rect 9340 33695 9656 33696
rect 17734 33760 18050 33761
rect 17734 33696 17740 33760
rect 17804 33696 17820 33760
rect 17884 33696 17900 33760
rect 17964 33696 17980 33760
rect 18044 33696 18050 33760
rect 17734 33695 18050 33696
rect 26128 33760 26444 33761
rect 26128 33696 26134 33760
rect 26198 33696 26214 33760
rect 26278 33696 26294 33760
rect 26358 33696 26374 33760
rect 26438 33696 26444 33760
rect 26128 33695 26444 33696
rect 34522 33760 34838 33761
rect 34522 33696 34528 33760
rect 34592 33696 34608 33760
rect 34672 33696 34688 33760
rect 34752 33696 34768 33760
rect 34832 33696 34838 33760
rect 34522 33695 34838 33696
rect 5143 33216 5459 33217
rect 5143 33152 5149 33216
rect 5213 33152 5229 33216
rect 5293 33152 5309 33216
rect 5373 33152 5389 33216
rect 5453 33152 5459 33216
rect 5143 33151 5459 33152
rect 13537 33216 13853 33217
rect 13537 33152 13543 33216
rect 13607 33152 13623 33216
rect 13687 33152 13703 33216
rect 13767 33152 13783 33216
rect 13847 33152 13853 33216
rect 13537 33151 13853 33152
rect 21931 33216 22247 33217
rect 21931 33152 21937 33216
rect 22001 33152 22017 33216
rect 22081 33152 22097 33216
rect 22161 33152 22177 33216
rect 22241 33152 22247 33216
rect 21931 33151 22247 33152
rect 30325 33216 30641 33217
rect 30325 33152 30331 33216
rect 30395 33152 30411 33216
rect 30475 33152 30491 33216
rect 30555 33152 30571 33216
rect 30635 33152 30641 33216
rect 30325 33151 30641 33152
rect 0 32738 800 32768
rect 933 32738 999 32741
rect 0 32736 999 32738
rect 0 32680 938 32736
rect 994 32680 999 32736
rect 0 32678 999 32680
rect 0 32648 800 32678
rect 933 32675 999 32678
rect 9340 32672 9656 32673
rect 9340 32608 9346 32672
rect 9410 32608 9426 32672
rect 9490 32608 9506 32672
rect 9570 32608 9586 32672
rect 9650 32608 9656 32672
rect 9340 32607 9656 32608
rect 17734 32672 18050 32673
rect 17734 32608 17740 32672
rect 17804 32608 17820 32672
rect 17884 32608 17900 32672
rect 17964 32608 17980 32672
rect 18044 32608 18050 32672
rect 17734 32607 18050 32608
rect 26128 32672 26444 32673
rect 26128 32608 26134 32672
rect 26198 32608 26214 32672
rect 26278 32608 26294 32672
rect 26358 32608 26374 32672
rect 26438 32608 26444 32672
rect 26128 32607 26444 32608
rect 34522 32672 34838 32673
rect 34522 32608 34528 32672
rect 34592 32608 34608 32672
rect 34672 32608 34688 32672
rect 34752 32608 34768 32672
rect 34832 32608 34838 32672
rect 34522 32607 34838 32608
rect 5143 32128 5459 32129
rect 5143 32064 5149 32128
rect 5213 32064 5229 32128
rect 5293 32064 5309 32128
rect 5373 32064 5389 32128
rect 5453 32064 5459 32128
rect 5143 32063 5459 32064
rect 13537 32128 13853 32129
rect 13537 32064 13543 32128
rect 13607 32064 13623 32128
rect 13687 32064 13703 32128
rect 13767 32064 13783 32128
rect 13847 32064 13853 32128
rect 13537 32063 13853 32064
rect 21931 32128 22247 32129
rect 21931 32064 21937 32128
rect 22001 32064 22017 32128
rect 22081 32064 22097 32128
rect 22161 32064 22177 32128
rect 22241 32064 22247 32128
rect 21931 32063 22247 32064
rect 30325 32128 30641 32129
rect 30325 32064 30331 32128
rect 30395 32064 30411 32128
rect 30475 32064 30491 32128
rect 30555 32064 30571 32128
rect 30635 32064 30641 32128
rect 30325 32063 30641 32064
rect 9340 31584 9656 31585
rect 9340 31520 9346 31584
rect 9410 31520 9426 31584
rect 9490 31520 9506 31584
rect 9570 31520 9586 31584
rect 9650 31520 9656 31584
rect 9340 31519 9656 31520
rect 17734 31584 18050 31585
rect 17734 31520 17740 31584
rect 17804 31520 17820 31584
rect 17884 31520 17900 31584
rect 17964 31520 17980 31584
rect 18044 31520 18050 31584
rect 17734 31519 18050 31520
rect 26128 31584 26444 31585
rect 26128 31520 26134 31584
rect 26198 31520 26214 31584
rect 26278 31520 26294 31584
rect 26358 31520 26374 31584
rect 26438 31520 26444 31584
rect 26128 31519 26444 31520
rect 34522 31584 34838 31585
rect 34522 31520 34528 31584
rect 34592 31520 34608 31584
rect 34672 31520 34688 31584
rect 34752 31520 34768 31584
rect 34832 31520 34838 31584
rect 34522 31519 34838 31520
rect 5143 31040 5459 31041
rect 5143 30976 5149 31040
rect 5213 30976 5229 31040
rect 5293 30976 5309 31040
rect 5373 30976 5389 31040
rect 5453 30976 5459 31040
rect 5143 30975 5459 30976
rect 13537 31040 13853 31041
rect 13537 30976 13543 31040
rect 13607 30976 13623 31040
rect 13687 30976 13703 31040
rect 13767 30976 13783 31040
rect 13847 30976 13853 31040
rect 13537 30975 13853 30976
rect 21931 31040 22247 31041
rect 21931 30976 21937 31040
rect 22001 30976 22017 31040
rect 22081 30976 22097 31040
rect 22161 30976 22177 31040
rect 22241 30976 22247 31040
rect 21931 30975 22247 30976
rect 30325 31040 30641 31041
rect 30325 30976 30331 31040
rect 30395 30976 30411 31040
rect 30475 30976 30491 31040
rect 30555 30976 30571 31040
rect 30635 30976 30641 31040
rect 30325 30975 30641 30976
rect 9340 30496 9656 30497
rect 9340 30432 9346 30496
rect 9410 30432 9426 30496
rect 9490 30432 9506 30496
rect 9570 30432 9586 30496
rect 9650 30432 9656 30496
rect 9340 30431 9656 30432
rect 17734 30496 18050 30497
rect 17734 30432 17740 30496
rect 17804 30432 17820 30496
rect 17884 30432 17900 30496
rect 17964 30432 17980 30496
rect 18044 30432 18050 30496
rect 17734 30431 18050 30432
rect 26128 30496 26444 30497
rect 26128 30432 26134 30496
rect 26198 30432 26214 30496
rect 26278 30432 26294 30496
rect 26358 30432 26374 30496
rect 26438 30432 26444 30496
rect 26128 30431 26444 30432
rect 34522 30496 34838 30497
rect 34522 30432 34528 30496
rect 34592 30432 34608 30496
rect 34672 30432 34688 30496
rect 34752 30432 34768 30496
rect 34832 30432 34838 30496
rect 34522 30431 34838 30432
rect 5143 29952 5459 29953
rect 5143 29888 5149 29952
rect 5213 29888 5229 29952
rect 5293 29888 5309 29952
rect 5373 29888 5389 29952
rect 5453 29888 5459 29952
rect 5143 29887 5459 29888
rect 13537 29952 13853 29953
rect 13537 29888 13543 29952
rect 13607 29888 13623 29952
rect 13687 29888 13703 29952
rect 13767 29888 13783 29952
rect 13847 29888 13853 29952
rect 13537 29887 13853 29888
rect 21931 29952 22247 29953
rect 21931 29888 21937 29952
rect 22001 29888 22017 29952
rect 22081 29888 22097 29952
rect 22161 29888 22177 29952
rect 22241 29888 22247 29952
rect 21931 29887 22247 29888
rect 30325 29952 30641 29953
rect 30325 29888 30331 29952
rect 30395 29888 30411 29952
rect 30475 29888 30491 29952
rect 30555 29888 30571 29952
rect 30635 29888 30641 29952
rect 30325 29887 30641 29888
rect 9121 29610 9187 29613
rect 10225 29610 10291 29613
rect 9121 29608 10291 29610
rect 9121 29552 9126 29608
rect 9182 29552 10230 29608
rect 10286 29552 10291 29608
rect 9121 29550 10291 29552
rect 9121 29547 9187 29550
rect 10225 29547 10291 29550
rect 9340 29408 9656 29409
rect 9340 29344 9346 29408
rect 9410 29344 9426 29408
rect 9490 29344 9506 29408
rect 9570 29344 9586 29408
rect 9650 29344 9656 29408
rect 9340 29343 9656 29344
rect 17734 29408 18050 29409
rect 17734 29344 17740 29408
rect 17804 29344 17820 29408
rect 17884 29344 17900 29408
rect 17964 29344 17980 29408
rect 18044 29344 18050 29408
rect 17734 29343 18050 29344
rect 26128 29408 26444 29409
rect 26128 29344 26134 29408
rect 26198 29344 26214 29408
rect 26278 29344 26294 29408
rect 26358 29344 26374 29408
rect 26438 29344 26444 29408
rect 26128 29343 26444 29344
rect 34522 29408 34838 29409
rect 34522 29344 34528 29408
rect 34592 29344 34608 29408
rect 34672 29344 34688 29408
rect 34752 29344 34768 29408
rect 34832 29344 34838 29408
rect 34522 29343 34838 29344
rect 5143 28864 5459 28865
rect 5143 28800 5149 28864
rect 5213 28800 5229 28864
rect 5293 28800 5309 28864
rect 5373 28800 5389 28864
rect 5453 28800 5459 28864
rect 5143 28799 5459 28800
rect 13537 28864 13853 28865
rect 13537 28800 13543 28864
rect 13607 28800 13623 28864
rect 13687 28800 13703 28864
rect 13767 28800 13783 28864
rect 13847 28800 13853 28864
rect 13537 28799 13853 28800
rect 21931 28864 22247 28865
rect 21931 28800 21937 28864
rect 22001 28800 22017 28864
rect 22081 28800 22097 28864
rect 22161 28800 22177 28864
rect 22241 28800 22247 28864
rect 21931 28799 22247 28800
rect 30325 28864 30641 28865
rect 30325 28800 30331 28864
rect 30395 28800 30411 28864
rect 30475 28800 30491 28864
rect 30555 28800 30571 28864
rect 30635 28800 30641 28864
rect 30325 28799 30641 28800
rect 9340 28320 9656 28321
rect 9340 28256 9346 28320
rect 9410 28256 9426 28320
rect 9490 28256 9506 28320
rect 9570 28256 9586 28320
rect 9650 28256 9656 28320
rect 9340 28255 9656 28256
rect 17734 28320 18050 28321
rect 17734 28256 17740 28320
rect 17804 28256 17820 28320
rect 17884 28256 17900 28320
rect 17964 28256 17980 28320
rect 18044 28256 18050 28320
rect 17734 28255 18050 28256
rect 26128 28320 26444 28321
rect 26128 28256 26134 28320
rect 26198 28256 26214 28320
rect 26278 28256 26294 28320
rect 26358 28256 26374 28320
rect 26438 28256 26444 28320
rect 26128 28255 26444 28256
rect 34522 28320 34838 28321
rect 34522 28256 34528 28320
rect 34592 28256 34608 28320
rect 34672 28256 34688 28320
rect 34752 28256 34768 28320
rect 34832 28256 34838 28320
rect 34522 28255 34838 28256
rect 34789 27978 34855 27981
rect 35073 27978 35873 28008
rect 34789 27976 35873 27978
rect 34789 27920 34794 27976
rect 34850 27920 35873 27976
rect 34789 27918 35873 27920
rect 34789 27915 34855 27918
rect 35073 27888 35873 27918
rect 5143 27776 5459 27777
rect 5143 27712 5149 27776
rect 5213 27712 5229 27776
rect 5293 27712 5309 27776
rect 5373 27712 5389 27776
rect 5453 27712 5459 27776
rect 5143 27711 5459 27712
rect 13537 27776 13853 27777
rect 13537 27712 13543 27776
rect 13607 27712 13623 27776
rect 13687 27712 13703 27776
rect 13767 27712 13783 27776
rect 13847 27712 13853 27776
rect 13537 27711 13853 27712
rect 21931 27776 22247 27777
rect 21931 27712 21937 27776
rect 22001 27712 22017 27776
rect 22081 27712 22097 27776
rect 22161 27712 22177 27776
rect 22241 27712 22247 27776
rect 21931 27711 22247 27712
rect 30325 27776 30641 27777
rect 30325 27712 30331 27776
rect 30395 27712 30411 27776
rect 30475 27712 30491 27776
rect 30555 27712 30571 27776
rect 30635 27712 30641 27776
rect 30325 27711 30641 27712
rect 9340 27232 9656 27233
rect 9340 27168 9346 27232
rect 9410 27168 9426 27232
rect 9490 27168 9506 27232
rect 9570 27168 9586 27232
rect 9650 27168 9656 27232
rect 9340 27167 9656 27168
rect 17734 27232 18050 27233
rect 17734 27168 17740 27232
rect 17804 27168 17820 27232
rect 17884 27168 17900 27232
rect 17964 27168 17980 27232
rect 18044 27168 18050 27232
rect 17734 27167 18050 27168
rect 26128 27232 26444 27233
rect 26128 27168 26134 27232
rect 26198 27168 26214 27232
rect 26278 27168 26294 27232
rect 26358 27168 26374 27232
rect 26438 27168 26444 27232
rect 26128 27167 26444 27168
rect 34522 27232 34838 27233
rect 34522 27168 34528 27232
rect 34592 27168 34608 27232
rect 34672 27168 34688 27232
rect 34752 27168 34768 27232
rect 34832 27168 34838 27232
rect 34522 27167 34838 27168
rect 5143 26688 5459 26689
rect 5143 26624 5149 26688
rect 5213 26624 5229 26688
rect 5293 26624 5309 26688
rect 5373 26624 5389 26688
rect 5453 26624 5459 26688
rect 5143 26623 5459 26624
rect 13537 26688 13853 26689
rect 13537 26624 13543 26688
rect 13607 26624 13623 26688
rect 13687 26624 13703 26688
rect 13767 26624 13783 26688
rect 13847 26624 13853 26688
rect 13537 26623 13853 26624
rect 21931 26688 22247 26689
rect 21931 26624 21937 26688
rect 22001 26624 22017 26688
rect 22081 26624 22097 26688
rect 22161 26624 22177 26688
rect 22241 26624 22247 26688
rect 21931 26623 22247 26624
rect 30325 26688 30641 26689
rect 30325 26624 30331 26688
rect 30395 26624 30411 26688
rect 30475 26624 30491 26688
rect 30555 26624 30571 26688
rect 30635 26624 30641 26688
rect 30325 26623 30641 26624
rect 25037 26482 25103 26485
rect 32581 26482 32647 26485
rect 25037 26480 32647 26482
rect 25037 26424 25042 26480
rect 25098 26424 32586 26480
rect 32642 26424 32647 26480
rect 25037 26422 32647 26424
rect 25037 26419 25103 26422
rect 32581 26419 32647 26422
rect 1393 26210 1459 26213
rect 798 26208 1459 26210
rect 798 26152 1398 26208
rect 1454 26152 1459 26208
rect 798 26150 1459 26152
rect 798 25968 858 26150
rect 1393 26147 1459 26150
rect 9340 26144 9656 26145
rect 9340 26080 9346 26144
rect 9410 26080 9426 26144
rect 9490 26080 9506 26144
rect 9570 26080 9586 26144
rect 9650 26080 9656 26144
rect 9340 26079 9656 26080
rect 17734 26144 18050 26145
rect 17734 26080 17740 26144
rect 17804 26080 17820 26144
rect 17884 26080 17900 26144
rect 17964 26080 17980 26144
rect 18044 26080 18050 26144
rect 17734 26079 18050 26080
rect 26128 26144 26444 26145
rect 26128 26080 26134 26144
rect 26198 26080 26214 26144
rect 26278 26080 26294 26144
rect 26358 26080 26374 26144
rect 26438 26080 26444 26144
rect 26128 26079 26444 26080
rect 34522 26144 34838 26145
rect 34522 26080 34528 26144
rect 34592 26080 34608 26144
rect 34672 26080 34688 26144
rect 34752 26080 34768 26144
rect 34832 26080 34838 26144
rect 34522 26079 34838 26080
rect 0 25878 858 25968
rect 0 25848 800 25878
rect 5143 25600 5459 25601
rect 5143 25536 5149 25600
rect 5213 25536 5229 25600
rect 5293 25536 5309 25600
rect 5373 25536 5389 25600
rect 5453 25536 5459 25600
rect 5143 25535 5459 25536
rect 13537 25600 13853 25601
rect 13537 25536 13543 25600
rect 13607 25536 13623 25600
rect 13687 25536 13703 25600
rect 13767 25536 13783 25600
rect 13847 25536 13853 25600
rect 13537 25535 13853 25536
rect 21931 25600 22247 25601
rect 21931 25536 21937 25600
rect 22001 25536 22017 25600
rect 22081 25536 22097 25600
rect 22161 25536 22177 25600
rect 22241 25536 22247 25600
rect 21931 25535 22247 25536
rect 30325 25600 30641 25601
rect 30325 25536 30331 25600
rect 30395 25536 30411 25600
rect 30475 25536 30491 25600
rect 30555 25536 30571 25600
rect 30635 25536 30641 25600
rect 30325 25535 30641 25536
rect 9340 25056 9656 25057
rect 9340 24992 9346 25056
rect 9410 24992 9426 25056
rect 9490 24992 9506 25056
rect 9570 24992 9586 25056
rect 9650 24992 9656 25056
rect 9340 24991 9656 24992
rect 17734 25056 18050 25057
rect 17734 24992 17740 25056
rect 17804 24992 17820 25056
rect 17884 24992 17900 25056
rect 17964 24992 17980 25056
rect 18044 24992 18050 25056
rect 17734 24991 18050 24992
rect 26128 25056 26444 25057
rect 26128 24992 26134 25056
rect 26198 24992 26214 25056
rect 26278 24992 26294 25056
rect 26358 24992 26374 25056
rect 26438 24992 26444 25056
rect 26128 24991 26444 24992
rect 34522 25056 34838 25057
rect 34522 24992 34528 25056
rect 34592 24992 34608 25056
rect 34672 24992 34688 25056
rect 34752 24992 34768 25056
rect 34832 24992 34838 25056
rect 34522 24991 34838 24992
rect 5143 24512 5459 24513
rect 5143 24448 5149 24512
rect 5213 24448 5229 24512
rect 5293 24448 5309 24512
rect 5373 24448 5389 24512
rect 5453 24448 5459 24512
rect 5143 24447 5459 24448
rect 13537 24512 13853 24513
rect 13537 24448 13543 24512
rect 13607 24448 13623 24512
rect 13687 24448 13703 24512
rect 13767 24448 13783 24512
rect 13847 24448 13853 24512
rect 13537 24447 13853 24448
rect 21931 24512 22247 24513
rect 21931 24448 21937 24512
rect 22001 24448 22017 24512
rect 22081 24448 22097 24512
rect 22161 24448 22177 24512
rect 22241 24448 22247 24512
rect 21931 24447 22247 24448
rect 30325 24512 30641 24513
rect 30325 24448 30331 24512
rect 30395 24448 30411 24512
rect 30475 24448 30491 24512
rect 30555 24448 30571 24512
rect 30635 24448 30641 24512
rect 30325 24447 30641 24448
rect 9340 23968 9656 23969
rect 9340 23904 9346 23968
rect 9410 23904 9426 23968
rect 9490 23904 9506 23968
rect 9570 23904 9586 23968
rect 9650 23904 9656 23968
rect 9340 23903 9656 23904
rect 17734 23968 18050 23969
rect 17734 23904 17740 23968
rect 17804 23904 17820 23968
rect 17884 23904 17900 23968
rect 17964 23904 17980 23968
rect 18044 23904 18050 23968
rect 17734 23903 18050 23904
rect 26128 23968 26444 23969
rect 26128 23904 26134 23968
rect 26198 23904 26214 23968
rect 26278 23904 26294 23968
rect 26358 23904 26374 23968
rect 26438 23904 26444 23968
rect 26128 23903 26444 23904
rect 34522 23968 34838 23969
rect 34522 23904 34528 23968
rect 34592 23904 34608 23968
rect 34672 23904 34688 23968
rect 34752 23904 34768 23968
rect 34832 23904 34838 23968
rect 34522 23903 34838 23904
rect 5143 23424 5459 23425
rect 5143 23360 5149 23424
rect 5213 23360 5229 23424
rect 5293 23360 5309 23424
rect 5373 23360 5389 23424
rect 5453 23360 5459 23424
rect 5143 23359 5459 23360
rect 13537 23424 13853 23425
rect 13537 23360 13543 23424
rect 13607 23360 13623 23424
rect 13687 23360 13703 23424
rect 13767 23360 13783 23424
rect 13847 23360 13853 23424
rect 13537 23359 13853 23360
rect 21931 23424 22247 23425
rect 21931 23360 21937 23424
rect 22001 23360 22017 23424
rect 22081 23360 22097 23424
rect 22161 23360 22177 23424
rect 22241 23360 22247 23424
rect 21931 23359 22247 23360
rect 30325 23424 30641 23425
rect 30325 23360 30331 23424
rect 30395 23360 30411 23424
rect 30475 23360 30491 23424
rect 30555 23360 30571 23424
rect 30635 23360 30641 23424
rect 30325 23359 30641 23360
rect 9340 22880 9656 22881
rect 9340 22816 9346 22880
rect 9410 22816 9426 22880
rect 9490 22816 9506 22880
rect 9570 22816 9586 22880
rect 9650 22816 9656 22880
rect 9340 22815 9656 22816
rect 17734 22880 18050 22881
rect 17734 22816 17740 22880
rect 17804 22816 17820 22880
rect 17884 22816 17900 22880
rect 17964 22816 17980 22880
rect 18044 22816 18050 22880
rect 17734 22815 18050 22816
rect 26128 22880 26444 22881
rect 26128 22816 26134 22880
rect 26198 22816 26214 22880
rect 26278 22816 26294 22880
rect 26358 22816 26374 22880
rect 26438 22816 26444 22880
rect 26128 22815 26444 22816
rect 34522 22880 34838 22881
rect 34522 22816 34528 22880
rect 34592 22816 34608 22880
rect 34672 22816 34688 22880
rect 34752 22816 34768 22880
rect 34832 22816 34838 22880
rect 34522 22815 34838 22816
rect 5143 22336 5459 22337
rect 5143 22272 5149 22336
rect 5213 22272 5229 22336
rect 5293 22272 5309 22336
rect 5373 22272 5389 22336
rect 5453 22272 5459 22336
rect 5143 22271 5459 22272
rect 13537 22336 13853 22337
rect 13537 22272 13543 22336
rect 13607 22272 13623 22336
rect 13687 22272 13703 22336
rect 13767 22272 13783 22336
rect 13847 22272 13853 22336
rect 13537 22271 13853 22272
rect 21931 22336 22247 22337
rect 21931 22272 21937 22336
rect 22001 22272 22017 22336
rect 22081 22272 22097 22336
rect 22161 22272 22177 22336
rect 22241 22272 22247 22336
rect 21931 22271 22247 22272
rect 30325 22336 30641 22337
rect 30325 22272 30331 22336
rect 30395 22272 30411 22336
rect 30475 22272 30491 22336
rect 30555 22272 30571 22336
rect 30635 22272 30641 22336
rect 30325 22271 30641 22272
rect 9340 21792 9656 21793
rect 9340 21728 9346 21792
rect 9410 21728 9426 21792
rect 9490 21728 9506 21792
rect 9570 21728 9586 21792
rect 9650 21728 9656 21792
rect 9340 21727 9656 21728
rect 17734 21792 18050 21793
rect 17734 21728 17740 21792
rect 17804 21728 17820 21792
rect 17884 21728 17900 21792
rect 17964 21728 17980 21792
rect 18044 21728 18050 21792
rect 17734 21727 18050 21728
rect 26128 21792 26444 21793
rect 26128 21728 26134 21792
rect 26198 21728 26214 21792
rect 26278 21728 26294 21792
rect 26358 21728 26374 21792
rect 26438 21728 26444 21792
rect 26128 21727 26444 21728
rect 34522 21792 34838 21793
rect 34522 21728 34528 21792
rect 34592 21728 34608 21792
rect 34672 21728 34688 21792
rect 34752 21728 34768 21792
rect 34832 21728 34838 21792
rect 34522 21727 34838 21728
rect 5143 21248 5459 21249
rect 5143 21184 5149 21248
rect 5213 21184 5229 21248
rect 5293 21184 5309 21248
rect 5373 21184 5389 21248
rect 5453 21184 5459 21248
rect 5143 21183 5459 21184
rect 13537 21248 13853 21249
rect 13537 21184 13543 21248
rect 13607 21184 13623 21248
rect 13687 21184 13703 21248
rect 13767 21184 13783 21248
rect 13847 21184 13853 21248
rect 13537 21183 13853 21184
rect 21931 21248 22247 21249
rect 21931 21184 21937 21248
rect 22001 21184 22017 21248
rect 22081 21184 22097 21248
rect 22161 21184 22177 21248
rect 22241 21184 22247 21248
rect 21931 21183 22247 21184
rect 30325 21248 30641 21249
rect 30325 21184 30331 21248
rect 30395 21184 30411 21248
rect 30475 21184 30491 21248
rect 30555 21184 30571 21248
rect 30635 21184 30641 21248
rect 30325 21183 30641 21184
rect 34789 21178 34855 21181
rect 35073 21178 35873 21208
rect 34789 21176 35873 21178
rect 34789 21120 34794 21176
rect 34850 21120 35873 21176
rect 34789 21118 35873 21120
rect 34789 21115 34855 21118
rect 35073 21088 35873 21118
rect 9340 20704 9656 20705
rect 9340 20640 9346 20704
rect 9410 20640 9426 20704
rect 9490 20640 9506 20704
rect 9570 20640 9586 20704
rect 9650 20640 9656 20704
rect 9340 20639 9656 20640
rect 17734 20704 18050 20705
rect 17734 20640 17740 20704
rect 17804 20640 17820 20704
rect 17884 20640 17900 20704
rect 17964 20640 17980 20704
rect 18044 20640 18050 20704
rect 17734 20639 18050 20640
rect 26128 20704 26444 20705
rect 26128 20640 26134 20704
rect 26198 20640 26214 20704
rect 26278 20640 26294 20704
rect 26358 20640 26374 20704
rect 26438 20640 26444 20704
rect 26128 20639 26444 20640
rect 34522 20704 34838 20705
rect 34522 20640 34528 20704
rect 34592 20640 34608 20704
rect 34672 20640 34688 20704
rect 34752 20640 34768 20704
rect 34832 20640 34838 20704
rect 34522 20639 34838 20640
rect 21541 20498 21607 20501
rect 24393 20498 24459 20501
rect 21541 20496 24459 20498
rect 21541 20440 21546 20496
rect 21602 20440 24398 20496
rect 24454 20440 24459 20496
rect 21541 20438 24459 20440
rect 21541 20435 21607 20438
rect 24393 20435 24459 20438
rect 5717 20362 5783 20365
rect 12249 20362 12315 20365
rect 5717 20360 12315 20362
rect 5717 20304 5722 20360
rect 5778 20304 12254 20360
rect 12310 20304 12315 20360
rect 5717 20302 12315 20304
rect 5717 20299 5783 20302
rect 12249 20299 12315 20302
rect 5143 20160 5459 20161
rect 5143 20096 5149 20160
rect 5213 20096 5229 20160
rect 5293 20096 5309 20160
rect 5373 20096 5389 20160
rect 5453 20096 5459 20160
rect 5143 20095 5459 20096
rect 13537 20160 13853 20161
rect 13537 20096 13543 20160
rect 13607 20096 13623 20160
rect 13687 20096 13703 20160
rect 13767 20096 13783 20160
rect 13847 20096 13853 20160
rect 13537 20095 13853 20096
rect 21931 20160 22247 20161
rect 21931 20096 21937 20160
rect 22001 20096 22017 20160
rect 22081 20096 22097 20160
rect 22161 20096 22177 20160
rect 22241 20096 22247 20160
rect 21931 20095 22247 20096
rect 30325 20160 30641 20161
rect 30325 20096 30331 20160
rect 30395 20096 30411 20160
rect 30475 20096 30491 20160
rect 30555 20096 30571 20160
rect 30635 20096 30641 20160
rect 30325 20095 30641 20096
rect 0 19818 800 19848
rect 933 19818 999 19821
rect 0 19816 999 19818
rect 0 19760 938 19816
rect 994 19760 999 19816
rect 0 19758 999 19760
rect 0 19728 800 19758
rect 933 19755 999 19758
rect 5993 19818 6059 19821
rect 11973 19818 12039 19821
rect 5993 19816 12039 19818
rect 5993 19760 5998 19816
rect 6054 19760 11978 19816
rect 12034 19760 12039 19816
rect 5993 19758 12039 19760
rect 5993 19755 6059 19758
rect 11973 19755 12039 19758
rect 9340 19616 9656 19617
rect 9340 19552 9346 19616
rect 9410 19552 9426 19616
rect 9490 19552 9506 19616
rect 9570 19552 9586 19616
rect 9650 19552 9656 19616
rect 9340 19551 9656 19552
rect 17734 19616 18050 19617
rect 17734 19552 17740 19616
rect 17804 19552 17820 19616
rect 17884 19552 17900 19616
rect 17964 19552 17980 19616
rect 18044 19552 18050 19616
rect 17734 19551 18050 19552
rect 26128 19616 26444 19617
rect 26128 19552 26134 19616
rect 26198 19552 26214 19616
rect 26278 19552 26294 19616
rect 26358 19552 26374 19616
rect 26438 19552 26444 19616
rect 26128 19551 26444 19552
rect 34522 19616 34838 19617
rect 34522 19552 34528 19616
rect 34592 19552 34608 19616
rect 34672 19552 34688 19616
rect 34752 19552 34768 19616
rect 34832 19552 34838 19616
rect 34522 19551 34838 19552
rect 3141 19410 3207 19413
rect 8477 19410 8543 19413
rect 3141 19408 8543 19410
rect 3141 19352 3146 19408
rect 3202 19352 8482 19408
rect 8538 19352 8543 19408
rect 3141 19350 8543 19352
rect 3141 19347 3207 19350
rect 8477 19347 8543 19350
rect 11697 19410 11763 19413
rect 12893 19410 12959 19413
rect 11697 19408 12959 19410
rect 11697 19352 11702 19408
rect 11758 19352 12898 19408
rect 12954 19352 12959 19408
rect 11697 19350 12959 19352
rect 11697 19347 11763 19350
rect 12893 19347 12959 19350
rect 5143 19072 5459 19073
rect 5143 19008 5149 19072
rect 5213 19008 5229 19072
rect 5293 19008 5309 19072
rect 5373 19008 5389 19072
rect 5453 19008 5459 19072
rect 5143 19007 5459 19008
rect 13537 19072 13853 19073
rect 13537 19008 13543 19072
rect 13607 19008 13623 19072
rect 13687 19008 13703 19072
rect 13767 19008 13783 19072
rect 13847 19008 13853 19072
rect 13537 19007 13853 19008
rect 21931 19072 22247 19073
rect 21931 19008 21937 19072
rect 22001 19008 22017 19072
rect 22081 19008 22097 19072
rect 22161 19008 22177 19072
rect 22241 19008 22247 19072
rect 21931 19007 22247 19008
rect 30325 19072 30641 19073
rect 30325 19008 30331 19072
rect 30395 19008 30411 19072
rect 30475 19008 30491 19072
rect 30555 19008 30571 19072
rect 30635 19008 30641 19072
rect 30325 19007 30641 19008
rect 4613 18866 4679 18869
rect 8753 18866 8819 18869
rect 4613 18864 8819 18866
rect 4613 18808 4618 18864
rect 4674 18808 8758 18864
rect 8814 18808 8819 18864
rect 4613 18806 8819 18808
rect 4613 18803 4679 18806
rect 8753 18803 8819 18806
rect 9673 18730 9739 18733
rect 12065 18730 12131 18733
rect 9673 18728 12131 18730
rect 9673 18672 9678 18728
rect 9734 18672 12070 18728
rect 12126 18672 12131 18728
rect 9673 18670 12131 18672
rect 9673 18667 9739 18670
rect 12065 18667 12131 18670
rect 9340 18528 9656 18529
rect 9340 18464 9346 18528
rect 9410 18464 9426 18528
rect 9490 18464 9506 18528
rect 9570 18464 9586 18528
rect 9650 18464 9656 18528
rect 9340 18463 9656 18464
rect 17734 18528 18050 18529
rect 17734 18464 17740 18528
rect 17804 18464 17820 18528
rect 17884 18464 17900 18528
rect 17964 18464 17980 18528
rect 18044 18464 18050 18528
rect 17734 18463 18050 18464
rect 26128 18528 26444 18529
rect 26128 18464 26134 18528
rect 26198 18464 26214 18528
rect 26278 18464 26294 18528
rect 26358 18464 26374 18528
rect 26438 18464 26444 18528
rect 26128 18463 26444 18464
rect 34522 18528 34838 18529
rect 34522 18464 34528 18528
rect 34592 18464 34608 18528
rect 34672 18464 34688 18528
rect 34752 18464 34768 18528
rect 34832 18464 34838 18528
rect 34522 18463 34838 18464
rect 5143 17984 5459 17985
rect 5143 17920 5149 17984
rect 5213 17920 5229 17984
rect 5293 17920 5309 17984
rect 5373 17920 5389 17984
rect 5453 17920 5459 17984
rect 5143 17919 5459 17920
rect 13537 17984 13853 17985
rect 13537 17920 13543 17984
rect 13607 17920 13623 17984
rect 13687 17920 13703 17984
rect 13767 17920 13783 17984
rect 13847 17920 13853 17984
rect 13537 17919 13853 17920
rect 21931 17984 22247 17985
rect 21931 17920 21937 17984
rect 22001 17920 22017 17984
rect 22081 17920 22097 17984
rect 22161 17920 22177 17984
rect 22241 17920 22247 17984
rect 21931 17919 22247 17920
rect 30325 17984 30641 17985
rect 30325 17920 30331 17984
rect 30395 17920 30411 17984
rect 30475 17920 30491 17984
rect 30555 17920 30571 17984
rect 30635 17920 30641 17984
rect 30325 17919 30641 17920
rect 7097 17778 7163 17781
rect 8937 17778 9003 17781
rect 7097 17776 9003 17778
rect 7097 17720 7102 17776
rect 7158 17720 8942 17776
rect 8998 17720 9003 17776
rect 7097 17718 9003 17720
rect 7097 17715 7163 17718
rect 8937 17715 9003 17718
rect 9070 17716 9076 17780
rect 9140 17778 9146 17780
rect 9305 17778 9371 17781
rect 9140 17776 9371 17778
rect 9140 17720 9310 17776
rect 9366 17720 9371 17776
rect 9140 17718 9371 17720
rect 9140 17716 9146 17718
rect 9305 17715 9371 17718
rect 9340 17440 9656 17441
rect 9340 17376 9346 17440
rect 9410 17376 9426 17440
rect 9490 17376 9506 17440
rect 9570 17376 9586 17440
rect 9650 17376 9656 17440
rect 9340 17375 9656 17376
rect 17734 17440 18050 17441
rect 17734 17376 17740 17440
rect 17804 17376 17820 17440
rect 17884 17376 17900 17440
rect 17964 17376 17980 17440
rect 18044 17376 18050 17440
rect 17734 17375 18050 17376
rect 26128 17440 26444 17441
rect 26128 17376 26134 17440
rect 26198 17376 26214 17440
rect 26278 17376 26294 17440
rect 26358 17376 26374 17440
rect 26438 17376 26444 17440
rect 26128 17375 26444 17376
rect 34522 17440 34838 17441
rect 34522 17376 34528 17440
rect 34592 17376 34608 17440
rect 34672 17376 34688 17440
rect 34752 17376 34768 17440
rect 34832 17376 34838 17440
rect 34522 17375 34838 17376
rect 3601 17234 3667 17237
rect 7373 17234 7439 17237
rect 3601 17232 7439 17234
rect 3601 17176 3606 17232
rect 3662 17176 7378 17232
rect 7434 17176 7439 17232
rect 3601 17174 7439 17176
rect 3601 17171 3667 17174
rect 7373 17171 7439 17174
rect 5143 16896 5459 16897
rect 5143 16832 5149 16896
rect 5213 16832 5229 16896
rect 5293 16832 5309 16896
rect 5373 16832 5389 16896
rect 5453 16832 5459 16896
rect 5143 16831 5459 16832
rect 13537 16896 13853 16897
rect 13537 16832 13543 16896
rect 13607 16832 13623 16896
rect 13687 16832 13703 16896
rect 13767 16832 13783 16896
rect 13847 16832 13853 16896
rect 13537 16831 13853 16832
rect 21931 16896 22247 16897
rect 21931 16832 21937 16896
rect 22001 16832 22017 16896
rect 22081 16832 22097 16896
rect 22161 16832 22177 16896
rect 22241 16832 22247 16896
rect 21931 16831 22247 16832
rect 30325 16896 30641 16897
rect 30325 16832 30331 16896
rect 30395 16832 30411 16896
rect 30475 16832 30491 16896
rect 30555 16832 30571 16896
rect 30635 16832 30641 16896
rect 30325 16831 30641 16832
rect 7925 16826 7991 16829
rect 9305 16826 9371 16829
rect 7925 16824 9371 16826
rect 7925 16768 7930 16824
rect 7986 16768 9310 16824
rect 9366 16768 9371 16824
rect 7925 16766 9371 16768
rect 7925 16763 7991 16766
rect 9305 16763 9371 16766
rect 4429 16690 4495 16693
rect 7741 16690 7807 16693
rect 8845 16690 8911 16693
rect 4429 16688 8911 16690
rect 4429 16632 4434 16688
rect 4490 16632 7746 16688
rect 7802 16632 8850 16688
rect 8906 16632 8911 16688
rect 4429 16630 8911 16632
rect 4429 16627 4495 16630
rect 7741 16627 7807 16630
rect 8845 16627 8911 16630
rect 6821 16554 6887 16557
rect 9397 16554 9463 16557
rect 6821 16552 9463 16554
rect 6821 16496 6826 16552
rect 6882 16496 9402 16552
rect 9458 16496 9463 16552
rect 6821 16494 9463 16496
rect 6821 16491 6887 16494
rect 9397 16491 9463 16494
rect 8293 16420 8359 16421
rect 8293 16416 8340 16420
rect 8404 16418 8410 16420
rect 8293 16360 8298 16416
rect 8293 16356 8340 16360
rect 8404 16358 8450 16418
rect 8404 16356 8410 16358
rect 8518 16356 8524 16420
rect 8588 16418 8594 16420
rect 8753 16418 8819 16421
rect 8588 16416 8819 16418
rect 8588 16360 8758 16416
rect 8814 16360 8819 16416
rect 8588 16358 8819 16360
rect 8588 16356 8594 16358
rect 8293 16355 8359 16356
rect 8753 16355 8819 16358
rect 9340 16352 9656 16353
rect 9340 16288 9346 16352
rect 9410 16288 9426 16352
rect 9490 16288 9506 16352
rect 9570 16288 9586 16352
rect 9650 16288 9656 16352
rect 9340 16287 9656 16288
rect 17734 16352 18050 16353
rect 17734 16288 17740 16352
rect 17804 16288 17820 16352
rect 17884 16288 17900 16352
rect 17964 16288 17980 16352
rect 18044 16288 18050 16352
rect 17734 16287 18050 16288
rect 26128 16352 26444 16353
rect 26128 16288 26134 16352
rect 26198 16288 26214 16352
rect 26278 16288 26294 16352
rect 26358 16288 26374 16352
rect 26438 16288 26444 16352
rect 26128 16287 26444 16288
rect 34522 16352 34838 16353
rect 34522 16288 34528 16352
rect 34592 16288 34608 16352
rect 34672 16288 34688 16352
rect 34752 16288 34768 16352
rect 34832 16288 34838 16352
rect 34522 16287 34838 16288
rect 8109 16282 8175 16285
rect 8753 16282 8819 16285
rect 8109 16280 8819 16282
rect 8109 16224 8114 16280
rect 8170 16224 8758 16280
rect 8814 16224 8819 16280
rect 8109 16222 8819 16224
rect 8109 16219 8175 16222
rect 8753 16219 8819 16222
rect 8569 16146 8635 16149
rect 11789 16146 11855 16149
rect 8569 16144 11855 16146
rect 8569 16088 8574 16144
rect 8630 16088 11794 16144
rect 11850 16088 11855 16144
rect 8569 16086 11855 16088
rect 8569 16083 8635 16086
rect 11789 16083 11855 16086
rect 9070 15948 9076 16012
rect 9140 16010 9146 16012
rect 9213 16010 9279 16013
rect 9140 16008 9279 16010
rect 9140 15952 9218 16008
rect 9274 15952 9279 16008
rect 9140 15950 9279 15952
rect 9140 15948 9146 15950
rect 9213 15947 9279 15950
rect 5143 15808 5459 15809
rect 5143 15744 5149 15808
rect 5213 15744 5229 15808
rect 5293 15744 5309 15808
rect 5373 15744 5389 15808
rect 5453 15744 5459 15808
rect 5143 15743 5459 15744
rect 13537 15808 13853 15809
rect 13537 15744 13543 15808
rect 13607 15744 13623 15808
rect 13687 15744 13703 15808
rect 13767 15744 13783 15808
rect 13847 15744 13853 15808
rect 13537 15743 13853 15744
rect 21931 15808 22247 15809
rect 21931 15744 21937 15808
rect 22001 15744 22017 15808
rect 22081 15744 22097 15808
rect 22161 15744 22177 15808
rect 22241 15744 22247 15808
rect 21931 15743 22247 15744
rect 30325 15808 30641 15809
rect 30325 15744 30331 15808
rect 30395 15744 30411 15808
rect 30475 15744 30491 15808
rect 30555 15744 30571 15808
rect 30635 15744 30641 15808
rect 30325 15743 30641 15744
rect 9673 15602 9739 15605
rect 11513 15602 11579 15605
rect 9673 15600 11579 15602
rect 9673 15544 9678 15600
rect 9734 15544 11518 15600
rect 11574 15544 11579 15600
rect 9673 15542 11579 15544
rect 9673 15539 9739 15542
rect 11513 15539 11579 15542
rect 6913 15466 6979 15469
rect 14825 15466 14891 15469
rect 6913 15464 14891 15466
rect 6913 15408 6918 15464
rect 6974 15408 14830 15464
rect 14886 15408 14891 15464
rect 6913 15406 14891 15408
rect 6913 15403 6979 15406
rect 14825 15403 14891 15406
rect 19977 15466 20043 15469
rect 22645 15466 22711 15469
rect 23289 15466 23355 15469
rect 19977 15464 23355 15466
rect 19977 15408 19982 15464
rect 20038 15408 22650 15464
rect 22706 15408 23294 15464
rect 23350 15408 23355 15464
rect 19977 15406 23355 15408
rect 19977 15403 20043 15406
rect 22645 15403 22711 15406
rect 23289 15403 23355 15406
rect 9765 15330 9831 15333
rect 12157 15330 12223 15333
rect 9765 15328 12223 15330
rect 9765 15272 9770 15328
rect 9826 15272 12162 15328
rect 12218 15272 12223 15328
rect 9765 15270 12223 15272
rect 9765 15267 9831 15270
rect 12157 15267 12223 15270
rect 9340 15264 9656 15265
rect 9340 15200 9346 15264
rect 9410 15200 9426 15264
rect 9490 15200 9506 15264
rect 9570 15200 9586 15264
rect 9650 15200 9656 15264
rect 9340 15199 9656 15200
rect 17734 15264 18050 15265
rect 17734 15200 17740 15264
rect 17804 15200 17820 15264
rect 17884 15200 17900 15264
rect 17964 15200 17980 15264
rect 18044 15200 18050 15264
rect 17734 15199 18050 15200
rect 26128 15264 26444 15265
rect 26128 15200 26134 15264
rect 26198 15200 26214 15264
rect 26278 15200 26294 15264
rect 26358 15200 26374 15264
rect 26438 15200 26444 15264
rect 26128 15199 26444 15200
rect 34522 15264 34838 15265
rect 34522 15200 34528 15264
rect 34592 15200 34608 15264
rect 34672 15200 34688 15264
rect 34752 15200 34768 15264
rect 34832 15200 34838 15264
rect 34522 15199 34838 15200
rect 5809 15194 5875 15197
rect 7925 15194 7991 15197
rect 5809 15192 7991 15194
rect 5809 15136 5814 15192
rect 5870 15136 7930 15192
rect 7986 15136 7991 15192
rect 5809 15134 7991 15136
rect 5809 15131 5875 15134
rect 7925 15131 7991 15134
rect 11881 15058 11947 15061
rect 13445 15058 13511 15061
rect 11881 15056 13511 15058
rect 11881 15000 11886 15056
rect 11942 15000 13450 15056
rect 13506 15000 13511 15056
rect 11881 14998 13511 15000
rect 11881 14995 11947 14998
rect 13445 14995 13511 14998
rect 7005 14922 7071 14925
rect 12801 14922 12867 14925
rect 7005 14920 12867 14922
rect 7005 14864 7010 14920
rect 7066 14864 12806 14920
rect 12862 14864 12867 14920
rect 7005 14862 12867 14864
rect 7005 14859 7071 14862
rect 12801 14859 12867 14862
rect 8569 14788 8635 14789
rect 8518 14724 8524 14788
rect 8588 14786 8635 14788
rect 8588 14784 8680 14786
rect 8630 14728 8680 14784
rect 8588 14726 8680 14728
rect 8588 14724 8635 14726
rect 8569 14723 8635 14724
rect 5143 14720 5459 14721
rect 5143 14656 5149 14720
rect 5213 14656 5229 14720
rect 5293 14656 5309 14720
rect 5373 14656 5389 14720
rect 5453 14656 5459 14720
rect 5143 14655 5459 14656
rect 13537 14720 13853 14721
rect 13537 14656 13543 14720
rect 13607 14656 13623 14720
rect 13687 14656 13703 14720
rect 13767 14656 13783 14720
rect 13847 14656 13853 14720
rect 13537 14655 13853 14656
rect 21931 14720 22247 14721
rect 21931 14656 21937 14720
rect 22001 14656 22017 14720
rect 22081 14656 22097 14720
rect 22161 14656 22177 14720
rect 22241 14656 22247 14720
rect 21931 14655 22247 14656
rect 30325 14720 30641 14721
rect 30325 14656 30331 14720
rect 30395 14656 30411 14720
rect 30475 14656 30491 14720
rect 30555 14656 30571 14720
rect 30635 14656 30641 14720
rect 30325 14655 30641 14656
rect 34697 14378 34763 14381
rect 35073 14378 35873 14408
rect 34697 14376 35873 14378
rect 34697 14320 34702 14376
rect 34758 14320 35873 14376
rect 34697 14318 35873 14320
rect 34697 14315 34763 14318
rect 35073 14288 35873 14318
rect 9340 14176 9656 14177
rect 9340 14112 9346 14176
rect 9410 14112 9426 14176
rect 9490 14112 9506 14176
rect 9570 14112 9586 14176
rect 9650 14112 9656 14176
rect 9340 14111 9656 14112
rect 17734 14176 18050 14177
rect 17734 14112 17740 14176
rect 17804 14112 17820 14176
rect 17884 14112 17900 14176
rect 17964 14112 17980 14176
rect 18044 14112 18050 14176
rect 17734 14111 18050 14112
rect 26128 14176 26444 14177
rect 26128 14112 26134 14176
rect 26198 14112 26214 14176
rect 26278 14112 26294 14176
rect 26358 14112 26374 14176
rect 26438 14112 26444 14176
rect 26128 14111 26444 14112
rect 34522 14176 34838 14177
rect 34522 14112 34528 14176
rect 34592 14112 34608 14176
rect 34672 14112 34688 14176
rect 34752 14112 34768 14176
rect 34832 14112 34838 14176
rect 34522 14111 34838 14112
rect 4245 13970 4311 13973
rect 4613 13970 4679 13973
rect 4245 13968 4679 13970
rect 4245 13912 4250 13968
rect 4306 13912 4618 13968
rect 4674 13912 4679 13968
rect 4245 13910 4679 13912
rect 4245 13907 4311 13910
rect 4613 13907 4679 13910
rect 11237 13970 11303 13973
rect 13353 13970 13419 13973
rect 11237 13968 13419 13970
rect 11237 13912 11242 13968
rect 11298 13912 13358 13968
rect 13414 13912 13419 13968
rect 11237 13910 13419 13912
rect 11237 13907 11303 13910
rect 13353 13907 13419 13910
rect 5143 13632 5459 13633
rect 5143 13568 5149 13632
rect 5213 13568 5229 13632
rect 5293 13568 5309 13632
rect 5373 13568 5389 13632
rect 5453 13568 5459 13632
rect 5143 13567 5459 13568
rect 13537 13632 13853 13633
rect 13537 13568 13543 13632
rect 13607 13568 13623 13632
rect 13687 13568 13703 13632
rect 13767 13568 13783 13632
rect 13847 13568 13853 13632
rect 13537 13567 13853 13568
rect 21931 13632 22247 13633
rect 21931 13568 21937 13632
rect 22001 13568 22017 13632
rect 22081 13568 22097 13632
rect 22161 13568 22177 13632
rect 22241 13568 22247 13632
rect 21931 13567 22247 13568
rect 30325 13632 30641 13633
rect 30325 13568 30331 13632
rect 30395 13568 30411 13632
rect 30475 13568 30491 13632
rect 30555 13568 30571 13632
rect 30635 13568 30641 13632
rect 30325 13567 30641 13568
rect 8293 13428 8359 13429
rect 8293 13424 8340 13428
rect 8404 13426 8410 13428
rect 11237 13426 11303 13429
rect 8404 13424 11303 13426
rect 8293 13368 8298 13424
rect 8404 13368 11242 13424
rect 11298 13368 11303 13424
rect 8293 13364 8340 13368
rect 8404 13366 11303 13368
rect 8404 13364 8410 13366
rect 8293 13363 8359 13364
rect 11237 13363 11303 13366
rect 9340 13088 9656 13089
rect 0 13018 800 13048
rect 9340 13024 9346 13088
rect 9410 13024 9426 13088
rect 9490 13024 9506 13088
rect 9570 13024 9586 13088
rect 9650 13024 9656 13088
rect 9340 13023 9656 13024
rect 17734 13088 18050 13089
rect 17734 13024 17740 13088
rect 17804 13024 17820 13088
rect 17884 13024 17900 13088
rect 17964 13024 17980 13088
rect 18044 13024 18050 13088
rect 17734 13023 18050 13024
rect 26128 13088 26444 13089
rect 26128 13024 26134 13088
rect 26198 13024 26214 13088
rect 26278 13024 26294 13088
rect 26358 13024 26374 13088
rect 26438 13024 26444 13088
rect 26128 13023 26444 13024
rect 34522 13088 34838 13089
rect 34522 13024 34528 13088
rect 34592 13024 34608 13088
rect 34672 13024 34688 13088
rect 34752 13024 34768 13088
rect 34832 13024 34838 13088
rect 34522 13023 34838 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 5143 12544 5459 12545
rect 5143 12480 5149 12544
rect 5213 12480 5229 12544
rect 5293 12480 5309 12544
rect 5373 12480 5389 12544
rect 5453 12480 5459 12544
rect 5143 12479 5459 12480
rect 13537 12544 13853 12545
rect 13537 12480 13543 12544
rect 13607 12480 13623 12544
rect 13687 12480 13703 12544
rect 13767 12480 13783 12544
rect 13847 12480 13853 12544
rect 13537 12479 13853 12480
rect 21931 12544 22247 12545
rect 21931 12480 21937 12544
rect 22001 12480 22017 12544
rect 22081 12480 22097 12544
rect 22161 12480 22177 12544
rect 22241 12480 22247 12544
rect 21931 12479 22247 12480
rect 30325 12544 30641 12545
rect 30325 12480 30331 12544
rect 30395 12480 30411 12544
rect 30475 12480 30491 12544
rect 30555 12480 30571 12544
rect 30635 12480 30641 12544
rect 30325 12479 30641 12480
rect 7465 12474 7531 12477
rect 9305 12474 9371 12477
rect 7465 12472 9371 12474
rect 7465 12416 7470 12472
rect 7526 12416 9310 12472
rect 9366 12416 9371 12472
rect 7465 12414 9371 12416
rect 7465 12411 7531 12414
rect 9305 12411 9371 12414
rect 5441 12202 5507 12205
rect 12709 12202 12775 12205
rect 5441 12200 12775 12202
rect 5441 12144 5446 12200
rect 5502 12144 12714 12200
rect 12770 12144 12775 12200
rect 5441 12142 12775 12144
rect 5441 12139 5507 12142
rect 12709 12139 12775 12142
rect 9340 12000 9656 12001
rect 9340 11936 9346 12000
rect 9410 11936 9426 12000
rect 9490 11936 9506 12000
rect 9570 11936 9586 12000
rect 9650 11936 9656 12000
rect 9340 11935 9656 11936
rect 17734 12000 18050 12001
rect 17734 11936 17740 12000
rect 17804 11936 17820 12000
rect 17884 11936 17900 12000
rect 17964 11936 17980 12000
rect 18044 11936 18050 12000
rect 17734 11935 18050 11936
rect 26128 12000 26444 12001
rect 26128 11936 26134 12000
rect 26198 11936 26214 12000
rect 26278 11936 26294 12000
rect 26358 11936 26374 12000
rect 26438 11936 26444 12000
rect 26128 11935 26444 11936
rect 34522 12000 34838 12001
rect 34522 11936 34528 12000
rect 34592 11936 34608 12000
rect 34672 11936 34688 12000
rect 34752 11936 34768 12000
rect 34832 11936 34838 12000
rect 34522 11935 34838 11936
rect 10317 11930 10383 11933
rect 10182 11928 10383 11930
rect 10182 11872 10322 11928
rect 10378 11872 10383 11928
rect 10182 11870 10383 11872
rect 5073 11794 5139 11797
rect 10182 11794 10242 11870
rect 10317 11867 10383 11870
rect 11881 11930 11947 11933
rect 13169 11930 13235 11933
rect 13721 11930 13787 11933
rect 11881 11928 13787 11930
rect 11881 11872 11886 11928
rect 11942 11872 13174 11928
rect 13230 11872 13726 11928
rect 13782 11872 13787 11928
rect 11881 11870 13787 11872
rect 11881 11867 11947 11870
rect 13169 11867 13235 11870
rect 13721 11867 13787 11870
rect 5073 11792 10242 11794
rect 5073 11736 5078 11792
rect 5134 11736 10242 11792
rect 5073 11734 10242 11736
rect 10409 11794 10475 11797
rect 11881 11794 11947 11797
rect 10409 11792 11947 11794
rect 10409 11736 10414 11792
rect 10470 11736 11886 11792
rect 11942 11736 11947 11792
rect 10409 11734 11947 11736
rect 5073 11731 5139 11734
rect 10409 11731 10475 11734
rect 11881 11731 11947 11734
rect 8385 11658 8451 11661
rect 9397 11658 9463 11661
rect 8385 11656 9463 11658
rect 8385 11600 8390 11656
rect 8446 11600 9402 11656
rect 9458 11600 9463 11656
rect 8385 11598 9463 11600
rect 8385 11595 8451 11598
rect 9397 11595 9463 11598
rect 8385 11522 8451 11525
rect 9765 11522 9831 11525
rect 8385 11520 9831 11522
rect 8385 11464 8390 11520
rect 8446 11464 9770 11520
rect 9826 11464 9831 11520
rect 8385 11462 9831 11464
rect 8385 11459 8451 11462
rect 9765 11459 9831 11462
rect 5143 11456 5459 11457
rect 5143 11392 5149 11456
rect 5213 11392 5229 11456
rect 5293 11392 5309 11456
rect 5373 11392 5389 11456
rect 5453 11392 5459 11456
rect 5143 11391 5459 11392
rect 13537 11456 13853 11457
rect 13537 11392 13543 11456
rect 13607 11392 13623 11456
rect 13687 11392 13703 11456
rect 13767 11392 13783 11456
rect 13847 11392 13853 11456
rect 13537 11391 13853 11392
rect 21931 11456 22247 11457
rect 21931 11392 21937 11456
rect 22001 11392 22017 11456
rect 22081 11392 22097 11456
rect 22161 11392 22177 11456
rect 22241 11392 22247 11456
rect 21931 11391 22247 11392
rect 30325 11456 30641 11457
rect 30325 11392 30331 11456
rect 30395 11392 30411 11456
rect 30475 11392 30491 11456
rect 30555 11392 30571 11456
rect 30635 11392 30641 11456
rect 30325 11391 30641 11392
rect 9121 11386 9187 11389
rect 10041 11386 10107 11389
rect 9121 11384 10107 11386
rect 9121 11328 9126 11384
rect 9182 11328 10046 11384
rect 10102 11328 10107 11384
rect 9121 11326 10107 11328
rect 9121 11323 9187 11326
rect 10041 11323 10107 11326
rect 6821 11114 6887 11117
rect 12525 11114 12591 11117
rect 6821 11112 12591 11114
rect 6821 11056 6826 11112
rect 6882 11056 12530 11112
rect 12586 11056 12591 11112
rect 6821 11054 12591 11056
rect 6821 11051 6887 11054
rect 12525 11051 12591 11054
rect 6269 10978 6335 10981
rect 8569 10978 8635 10981
rect 6269 10976 8635 10978
rect 6269 10920 6274 10976
rect 6330 10920 8574 10976
rect 8630 10920 8635 10976
rect 6269 10918 8635 10920
rect 6269 10915 6335 10918
rect 8569 10915 8635 10918
rect 9340 10912 9656 10913
rect 9340 10848 9346 10912
rect 9410 10848 9426 10912
rect 9490 10848 9506 10912
rect 9570 10848 9586 10912
rect 9650 10848 9656 10912
rect 9340 10847 9656 10848
rect 17734 10912 18050 10913
rect 17734 10848 17740 10912
rect 17804 10848 17820 10912
rect 17884 10848 17900 10912
rect 17964 10848 17980 10912
rect 18044 10848 18050 10912
rect 17734 10847 18050 10848
rect 26128 10912 26444 10913
rect 26128 10848 26134 10912
rect 26198 10848 26214 10912
rect 26278 10848 26294 10912
rect 26358 10848 26374 10912
rect 26438 10848 26444 10912
rect 26128 10847 26444 10848
rect 34522 10912 34838 10913
rect 34522 10848 34528 10912
rect 34592 10848 34608 10912
rect 34672 10848 34688 10912
rect 34752 10848 34768 10912
rect 34832 10848 34838 10912
rect 34522 10847 34838 10848
rect 5143 10368 5459 10369
rect 5143 10304 5149 10368
rect 5213 10304 5229 10368
rect 5293 10304 5309 10368
rect 5373 10304 5389 10368
rect 5453 10304 5459 10368
rect 5143 10303 5459 10304
rect 13537 10368 13853 10369
rect 13537 10304 13543 10368
rect 13607 10304 13623 10368
rect 13687 10304 13703 10368
rect 13767 10304 13783 10368
rect 13847 10304 13853 10368
rect 13537 10303 13853 10304
rect 21931 10368 22247 10369
rect 21931 10304 21937 10368
rect 22001 10304 22017 10368
rect 22081 10304 22097 10368
rect 22161 10304 22177 10368
rect 22241 10304 22247 10368
rect 21931 10303 22247 10304
rect 30325 10368 30641 10369
rect 30325 10304 30331 10368
rect 30395 10304 30411 10368
rect 30475 10304 30491 10368
rect 30555 10304 30571 10368
rect 30635 10304 30641 10368
rect 30325 10303 30641 10304
rect 9340 9824 9656 9825
rect 9340 9760 9346 9824
rect 9410 9760 9426 9824
rect 9490 9760 9506 9824
rect 9570 9760 9586 9824
rect 9650 9760 9656 9824
rect 9340 9759 9656 9760
rect 17734 9824 18050 9825
rect 17734 9760 17740 9824
rect 17804 9760 17820 9824
rect 17884 9760 17900 9824
rect 17964 9760 17980 9824
rect 18044 9760 18050 9824
rect 17734 9759 18050 9760
rect 26128 9824 26444 9825
rect 26128 9760 26134 9824
rect 26198 9760 26214 9824
rect 26278 9760 26294 9824
rect 26358 9760 26374 9824
rect 26438 9760 26444 9824
rect 26128 9759 26444 9760
rect 34522 9824 34838 9825
rect 34522 9760 34528 9824
rect 34592 9760 34608 9824
rect 34672 9760 34688 9824
rect 34752 9760 34768 9824
rect 34832 9760 34838 9824
rect 34522 9759 34838 9760
rect 10869 9754 10935 9757
rect 12433 9754 12499 9757
rect 13537 9754 13603 9757
rect 10869 9752 13603 9754
rect 10869 9696 10874 9752
rect 10930 9696 12438 9752
rect 12494 9696 13542 9752
rect 13598 9696 13603 9752
rect 10869 9694 13603 9696
rect 10869 9691 10935 9694
rect 12433 9691 12499 9694
rect 13537 9691 13603 9694
rect 12157 9618 12223 9621
rect 13721 9618 13787 9621
rect 12157 9616 13787 9618
rect 12157 9560 12162 9616
rect 12218 9560 13726 9616
rect 13782 9560 13787 9616
rect 12157 9558 13787 9560
rect 12157 9555 12223 9558
rect 13721 9555 13787 9558
rect 20161 9618 20227 9621
rect 22553 9618 22619 9621
rect 20161 9616 22619 9618
rect 20161 9560 20166 9616
rect 20222 9560 22558 9616
rect 22614 9560 22619 9616
rect 20161 9558 22619 9560
rect 20161 9555 20227 9558
rect 22553 9555 22619 9558
rect 15193 9482 15259 9485
rect 15837 9482 15903 9485
rect 15193 9480 15903 9482
rect 15193 9424 15198 9480
rect 15254 9424 15842 9480
rect 15898 9424 15903 9480
rect 15193 9422 15903 9424
rect 15193 9419 15259 9422
rect 15837 9419 15903 9422
rect 5143 9280 5459 9281
rect 5143 9216 5149 9280
rect 5213 9216 5229 9280
rect 5293 9216 5309 9280
rect 5373 9216 5389 9280
rect 5453 9216 5459 9280
rect 5143 9215 5459 9216
rect 13537 9280 13853 9281
rect 13537 9216 13543 9280
rect 13607 9216 13623 9280
rect 13687 9216 13703 9280
rect 13767 9216 13783 9280
rect 13847 9216 13853 9280
rect 13537 9215 13853 9216
rect 21931 9280 22247 9281
rect 21931 9216 21937 9280
rect 22001 9216 22017 9280
rect 22081 9216 22097 9280
rect 22161 9216 22177 9280
rect 22241 9216 22247 9280
rect 21931 9215 22247 9216
rect 30325 9280 30641 9281
rect 30325 9216 30331 9280
rect 30395 9216 30411 9280
rect 30475 9216 30491 9280
rect 30555 9216 30571 9280
rect 30635 9216 30641 9280
rect 30325 9215 30641 9216
rect 9340 8736 9656 8737
rect 9340 8672 9346 8736
rect 9410 8672 9426 8736
rect 9490 8672 9506 8736
rect 9570 8672 9586 8736
rect 9650 8672 9656 8736
rect 9340 8671 9656 8672
rect 17734 8736 18050 8737
rect 17734 8672 17740 8736
rect 17804 8672 17820 8736
rect 17884 8672 17900 8736
rect 17964 8672 17980 8736
rect 18044 8672 18050 8736
rect 17734 8671 18050 8672
rect 26128 8736 26444 8737
rect 26128 8672 26134 8736
rect 26198 8672 26214 8736
rect 26278 8672 26294 8736
rect 26358 8672 26374 8736
rect 26438 8672 26444 8736
rect 26128 8671 26444 8672
rect 34522 8736 34838 8737
rect 34522 8672 34528 8736
rect 34592 8672 34608 8736
rect 34672 8672 34688 8736
rect 34752 8672 34768 8736
rect 34832 8672 34838 8736
rect 34522 8671 34838 8672
rect 34789 8258 34855 8261
rect 35073 8258 35873 8288
rect 34789 8256 35873 8258
rect 34789 8200 34794 8256
rect 34850 8200 35873 8256
rect 34789 8198 35873 8200
rect 34789 8195 34855 8198
rect 5143 8192 5459 8193
rect 5143 8128 5149 8192
rect 5213 8128 5229 8192
rect 5293 8128 5309 8192
rect 5373 8128 5389 8192
rect 5453 8128 5459 8192
rect 5143 8127 5459 8128
rect 13537 8192 13853 8193
rect 13537 8128 13543 8192
rect 13607 8128 13623 8192
rect 13687 8128 13703 8192
rect 13767 8128 13783 8192
rect 13847 8128 13853 8192
rect 13537 8127 13853 8128
rect 21931 8192 22247 8193
rect 21931 8128 21937 8192
rect 22001 8128 22017 8192
rect 22081 8128 22097 8192
rect 22161 8128 22177 8192
rect 22241 8128 22247 8192
rect 21931 8127 22247 8128
rect 30325 8192 30641 8193
rect 30325 8128 30331 8192
rect 30395 8128 30411 8192
rect 30475 8128 30491 8192
rect 30555 8128 30571 8192
rect 30635 8128 30641 8192
rect 35073 8168 35873 8198
rect 30325 8127 30641 8128
rect 9340 7648 9656 7649
rect 9340 7584 9346 7648
rect 9410 7584 9426 7648
rect 9490 7584 9506 7648
rect 9570 7584 9586 7648
rect 9650 7584 9656 7648
rect 9340 7583 9656 7584
rect 17734 7648 18050 7649
rect 17734 7584 17740 7648
rect 17804 7584 17820 7648
rect 17884 7584 17900 7648
rect 17964 7584 17980 7648
rect 18044 7584 18050 7648
rect 17734 7583 18050 7584
rect 26128 7648 26444 7649
rect 26128 7584 26134 7648
rect 26198 7584 26214 7648
rect 26278 7584 26294 7648
rect 26358 7584 26374 7648
rect 26438 7584 26444 7648
rect 26128 7583 26444 7584
rect 34522 7648 34838 7649
rect 34522 7584 34528 7648
rect 34592 7584 34608 7648
rect 34672 7584 34688 7648
rect 34752 7584 34768 7648
rect 34832 7584 34838 7648
rect 34522 7583 34838 7584
rect 5143 7104 5459 7105
rect 5143 7040 5149 7104
rect 5213 7040 5229 7104
rect 5293 7040 5309 7104
rect 5373 7040 5389 7104
rect 5453 7040 5459 7104
rect 5143 7039 5459 7040
rect 13537 7104 13853 7105
rect 13537 7040 13543 7104
rect 13607 7040 13623 7104
rect 13687 7040 13703 7104
rect 13767 7040 13783 7104
rect 13847 7040 13853 7104
rect 13537 7039 13853 7040
rect 21931 7104 22247 7105
rect 21931 7040 21937 7104
rect 22001 7040 22017 7104
rect 22081 7040 22097 7104
rect 22161 7040 22177 7104
rect 22241 7040 22247 7104
rect 21931 7039 22247 7040
rect 30325 7104 30641 7105
rect 30325 7040 30331 7104
rect 30395 7040 30411 7104
rect 30475 7040 30491 7104
rect 30555 7040 30571 7104
rect 30635 7040 30641 7104
rect 30325 7039 30641 7040
rect 9340 6560 9656 6561
rect 9340 6496 9346 6560
rect 9410 6496 9426 6560
rect 9490 6496 9506 6560
rect 9570 6496 9586 6560
rect 9650 6496 9656 6560
rect 9340 6495 9656 6496
rect 17734 6560 18050 6561
rect 17734 6496 17740 6560
rect 17804 6496 17820 6560
rect 17884 6496 17900 6560
rect 17964 6496 17980 6560
rect 18044 6496 18050 6560
rect 17734 6495 18050 6496
rect 26128 6560 26444 6561
rect 26128 6496 26134 6560
rect 26198 6496 26214 6560
rect 26278 6496 26294 6560
rect 26358 6496 26374 6560
rect 26438 6496 26444 6560
rect 26128 6495 26444 6496
rect 34522 6560 34838 6561
rect 34522 6496 34528 6560
rect 34592 6496 34608 6560
rect 34672 6496 34688 6560
rect 34752 6496 34768 6560
rect 34832 6496 34838 6560
rect 34522 6495 34838 6496
rect 0 6218 800 6248
rect 933 6218 999 6221
rect 0 6216 999 6218
rect 0 6160 938 6216
rect 994 6160 999 6216
rect 0 6158 999 6160
rect 0 6128 800 6158
rect 933 6155 999 6158
rect 5143 6016 5459 6017
rect 5143 5952 5149 6016
rect 5213 5952 5229 6016
rect 5293 5952 5309 6016
rect 5373 5952 5389 6016
rect 5453 5952 5459 6016
rect 5143 5951 5459 5952
rect 13537 6016 13853 6017
rect 13537 5952 13543 6016
rect 13607 5952 13623 6016
rect 13687 5952 13703 6016
rect 13767 5952 13783 6016
rect 13847 5952 13853 6016
rect 13537 5951 13853 5952
rect 21931 6016 22247 6017
rect 21931 5952 21937 6016
rect 22001 5952 22017 6016
rect 22081 5952 22097 6016
rect 22161 5952 22177 6016
rect 22241 5952 22247 6016
rect 21931 5951 22247 5952
rect 30325 6016 30641 6017
rect 30325 5952 30331 6016
rect 30395 5952 30411 6016
rect 30475 5952 30491 6016
rect 30555 5952 30571 6016
rect 30635 5952 30641 6016
rect 30325 5951 30641 5952
rect 9340 5472 9656 5473
rect 9340 5408 9346 5472
rect 9410 5408 9426 5472
rect 9490 5408 9506 5472
rect 9570 5408 9586 5472
rect 9650 5408 9656 5472
rect 9340 5407 9656 5408
rect 17734 5472 18050 5473
rect 17734 5408 17740 5472
rect 17804 5408 17820 5472
rect 17884 5408 17900 5472
rect 17964 5408 17980 5472
rect 18044 5408 18050 5472
rect 17734 5407 18050 5408
rect 26128 5472 26444 5473
rect 26128 5408 26134 5472
rect 26198 5408 26214 5472
rect 26278 5408 26294 5472
rect 26358 5408 26374 5472
rect 26438 5408 26444 5472
rect 26128 5407 26444 5408
rect 34522 5472 34838 5473
rect 34522 5408 34528 5472
rect 34592 5408 34608 5472
rect 34672 5408 34688 5472
rect 34752 5408 34768 5472
rect 34832 5408 34838 5472
rect 34522 5407 34838 5408
rect 5143 4928 5459 4929
rect 5143 4864 5149 4928
rect 5213 4864 5229 4928
rect 5293 4864 5309 4928
rect 5373 4864 5389 4928
rect 5453 4864 5459 4928
rect 5143 4863 5459 4864
rect 13537 4928 13853 4929
rect 13537 4864 13543 4928
rect 13607 4864 13623 4928
rect 13687 4864 13703 4928
rect 13767 4864 13783 4928
rect 13847 4864 13853 4928
rect 13537 4863 13853 4864
rect 21931 4928 22247 4929
rect 21931 4864 21937 4928
rect 22001 4864 22017 4928
rect 22081 4864 22097 4928
rect 22161 4864 22177 4928
rect 22241 4864 22247 4928
rect 21931 4863 22247 4864
rect 30325 4928 30641 4929
rect 30325 4864 30331 4928
rect 30395 4864 30411 4928
rect 30475 4864 30491 4928
rect 30555 4864 30571 4928
rect 30635 4864 30641 4928
rect 30325 4863 30641 4864
rect 9340 4384 9656 4385
rect 9340 4320 9346 4384
rect 9410 4320 9426 4384
rect 9490 4320 9506 4384
rect 9570 4320 9586 4384
rect 9650 4320 9656 4384
rect 9340 4319 9656 4320
rect 17734 4384 18050 4385
rect 17734 4320 17740 4384
rect 17804 4320 17820 4384
rect 17884 4320 17900 4384
rect 17964 4320 17980 4384
rect 18044 4320 18050 4384
rect 17734 4319 18050 4320
rect 26128 4384 26444 4385
rect 26128 4320 26134 4384
rect 26198 4320 26214 4384
rect 26278 4320 26294 4384
rect 26358 4320 26374 4384
rect 26438 4320 26444 4384
rect 26128 4319 26444 4320
rect 34522 4384 34838 4385
rect 34522 4320 34528 4384
rect 34592 4320 34608 4384
rect 34672 4320 34688 4384
rect 34752 4320 34768 4384
rect 34832 4320 34838 4384
rect 34522 4319 34838 4320
rect 5143 3840 5459 3841
rect 5143 3776 5149 3840
rect 5213 3776 5229 3840
rect 5293 3776 5309 3840
rect 5373 3776 5389 3840
rect 5453 3776 5459 3840
rect 5143 3775 5459 3776
rect 13537 3840 13853 3841
rect 13537 3776 13543 3840
rect 13607 3776 13623 3840
rect 13687 3776 13703 3840
rect 13767 3776 13783 3840
rect 13847 3776 13853 3840
rect 13537 3775 13853 3776
rect 21931 3840 22247 3841
rect 21931 3776 21937 3840
rect 22001 3776 22017 3840
rect 22081 3776 22097 3840
rect 22161 3776 22177 3840
rect 22241 3776 22247 3840
rect 21931 3775 22247 3776
rect 30325 3840 30641 3841
rect 30325 3776 30331 3840
rect 30395 3776 30411 3840
rect 30475 3776 30491 3840
rect 30555 3776 30571 3840
rect 30635 3776 30641 3840
rect 30325 3775 30641 3776
rect 9340 3296 9656 3297
rect 9340 3232 9346 3296
rect 9410 3232 9426 3296
rect 9490 3232 9506 3296
rect 9570 3232 9586 3296
rect 9650 3232 9656 3296
rect 9340 3231 9656 3232
rect 17734 3296 18050 3297
rect 17734 3232 17740 3296
rect 17804 3232 17820 3296
rect 17884 3232 17900 3296
rect 17964 3232 17980 3296
rect 18044 3232 18050 3296
rect 17734 3231 18050 3232
rect 26128 3296 26444 3297
rect 26128 3232 26134 3296
rect 26198 3232 26214 3296
rect 26278 3232 26294 3296
rect 26358 3232 26374 3296
rect 26438 3232 26444 3296
rect 26128 3231 26444 3232
rect 34522 3296 34838 3297
rect 34522 3232 34528 3296
rect 34592 3232 34608 3296
rect 34672 3232 34688 3296
rect 34752 3232 34768 3296
rect 34832 3232 34838 3296
rect 34522 3231 34838 3232
rect 5143 2752 5459 2753
rect 5143 2688 5149 2752
rect 5213 2688 5229 2752
rect 5293 2688 5309 2752
rect 5373 2688 5389 2752
rect 5453 2688 5459 2752
rect 5143 2687 5459 2688
rect 13537 2752 13853 2753
rect 13537 2688 13543 2752
rect 13607 2688 13623 2752
rect 13687 2688 13703 2752
rect 13767 2688 13783 2752
rect 13847 2688 13853 2752
rect 13537 2687 13853 2688
rect 21931 2752 22247 2753
rect 21931 2688 21937 2752
rect 22001 2688 22017 2752
rect 22081 2688 22097 2752
rect 22161 2688 22177 2752
rect 22241 2688 22247 2752
rect 21931 2687 22247 2688
rect 30325 2752 30641 2753
rect 30325 2688 30331 2752
rect 30395 2688 30411 2752
rect 30475 2688 30491 2752
rect 30555 2688 30571 2752
rect 30635 2688 30641 2752
rect 30325 2687 30641 2688
rect 9340 2208 9656 2209
rect 9340 2144 9346 2208
rect 9410 2144 9426 2208
rect 9490 2144 9506 2208
rect 9570 2144 9586 2208
rect 9650 2144 9656 2208
rect 9340 2143 9656 2144
rect 17734 2208 18050 2209
rect 17734 2144 17740 2208
rect 17804 2144 17820 2208
rect 17884 2144 17900 2208
rect 17964 2144 17980 2208
rect 18044 2144 18050 2208
rect 17734 2143 18050 2144
rect 26128 2208 26444 2209
rect 26128 2144 26134 2208
rect 26198 2144 26214 2208
rect 26278 2144 26294 2208
rect 26358 2144 26374 2208
rect 26438 2144 26444 2208
rect 26128 2143 26444 2144
rect 34522 2208 34838 2209
rect 34522 2144 34528 2208
rect 34592 2144 34608 2208
rect 34672 2144 34688 2208
rect 34752 2144 34768 2208
rect 34832 2144 34838 2208
rect 34522 2143 34838 2144
rect 34513 1458 34579 1461
rect 35073 1458 35873 1488
rect 34513 1456 35873 1458
rect 34513 1400 34518 1456
rect 34574 1400 35873 1456
rect 34513 1398 35873 1400
rect 34513 1395 34579 1398
rect 35073 1368 35873 1398
<< via3 >>
rect 5149 35388 5213 35392
rect 5149 35332 5153 35388
rect 5153 35332 5209 35388
rect 5209 35332 5213 35388
rect 5149 35328 5213 35332
rect 5229 35388 5293 35392
rect 5229 35332 5233 35388
rect 5233 35332 5289 35388
rect 5289 35332 5293 35388
rect 5229 35328 5293 35332
rect 5309 35388 5373 35392
rect 5309 35332 5313 35388
rect 5313 35332 5369 35388
rect 5369 35332 5373 35388
rect 5309 35328 5373 35332
rect 5389 35388 5453 35392
rect 5389 35332 5393 35388
rect 5393 35332 5449 35388
rect 5449 35332 5453 35388
rect 5389 35328 5453 35332
rect 13543 35388 13607 35392
rect 13543 35332 13547 35388
rect 13547 35332 13603 35388
rect 13603 35332 13607 35388
rect 13543 35328 13607 35332
rect 13623 35388 13687 35392
rect 13623 35332 13627 35388
rect 13627 35332 13683 35388
rect 13683 35332 13687 35388
rect 13623 35328 13687 35332
rect 13703 35388 13767 35392
rect 13703 35332 13707 35388
rect 13707 35332 13763 35388
rect 13763 35332 13767 35388
rect 13703 35328 13767 35332
rect 13783 35388 13847 35392
rect 13783 35332 13787 35388
rect 13787 35332 13843 35388
rect 13843 35332 13847 35388
rect 13783 35328 13847 35332
rect 21937 35388 22001 35392
rect 21937 35332 21941 35388
rect 21941 35332 21997 35388
rect 21997 35332 22001 35388
rect 21937 35328 22001 35332
rect 22017 35388 22081 35392
rect 22017 35332 22021 35388
rect 22021 35332 22077 35388
rect 22077 35332 22081 35388
rect 22017 35328 22081 35332
rect 22097 35388 22161 35392
rect 22097 35332 22101 35388
rect 22101 35332 22157 35388
rect 22157 35332 22161 35388
rect 22097 35328 22161 35332
rect 22177 35388 22241 35392
rect 22177 35332 22181 35388
rect 22181 35332 22237 35388
rect 22237 35332 22241 35388
rect 22177 35328 22241 35332
rect 30331 35388 30395 35392
rect 30331 35332 30335 35388
rect 30335 35332 30391 35388
rect 30391 35332 30395 35388
rect 30331 35328 30395 35332
rect 30411 35388 30475 35392
rect 30411 35332 30415 35388
rect 30415 35332 30471 35388
rect 30471 35332 30475 35388
rect 30411 35328 30475 35332
rect 30491 35388 30555 35392
rect 30491 35332 30495 35388
rect 30495 35332 30551 35388
rect 30551 35332 30555 35388
rect 30491 35328 30555 35332
rect 30571 35388 30635 35392
rect 30571 35332 30575 35388
rect 30575 35332 30631 35388
rect 30631 35332 30635 35388
rect 30571 35328 30635 35332
rect 9346 34844 9410 34848
rect 9346 34788 9350 34844
rect 9350 34788 9406 34844
rect 9406 34788 9410 34844
rect 9346 34784 9410 34788
rect 9426 34844 9490 34848
rect 9426 34788 9430 34844
rect 9430 34788 9486 34844
rect 9486 34788 9490 34844
rect 9426 34784 9490 34788
rect 9506 34844 9570 34848
rect 9506 34788 9510 34844
rect 9510 34788 9566 34844
rect 9566 34788 9570 34844
rect 9506 34784 9570 34788
rect 9586 34844 9650 34848
rect 9586 34788 9590 34844
rect 9590 34788 9646 34844
rect 9646 34788 9650 34844
rect 9586 34784 9650 34788
rect 17740 34844 17804 34848
rect 17740 34788 17744 34844
rect 17744 34788 17800 34844
rect 17800 34788 17804 34844
rect 17740 34784 17804 34788
rect 17820 34844 17884 34848
rect 17820 34788 17824 34844
rect 17824 34788 17880 34844
rect 17880 34788 17884 34844
rect 17820 34784 17884 34788
rect 17900 34844 17964 34848
rect 17900 34788 17904 34844
rect 17904 34788 17960 34844
rect 17960 34788 17964 34844
rect 17900 34784 17964 34788
rect 17980 34844 18044 34848
rect 17980 34788 17984 34844
rect 17984 34788 18040 34844
rect 18040 34788 18044 34844
rect 17980 34784 18044 34788
rect 26134 34844 26198 34848
rect 26134 34788 26138 34844
rect 26138 34788 26194 34844
rect 26194 34788 26198 34844
rect 26134 34784 26198 34788
rect 26214 34844 26278 34848
rect 26214 34788 26218 34844
rect 26218 34788 26274 34844
rect 26274 34788 26278 34844
rect 26214 34784 26278 34788
rect 26294 34844 26358 34848
rect 26294 34788 26298 34844
rect 26298 34788 26354 34844
rect 26354 34788 26358 34844
rect 26294 34784 26358 34788
rect 26374 34844 26438 34848
rect 26374 34788 26378 34844
rect 26378 34788 26434 34844
rect 26434 34788 26438 34844
rect 26374 34784 26438 34788
rect 34528 34844 34592 34848
rect 34528 34788 34532 34844
rect 34532 34788 34588 34844
rect 34588 34788 34592 34844
rect 34528 34784 34592 34788
rect 34608 34844 34672 34848
rect 34608 34788 34612 34844
rect 34612 34788 34668 34844
rect 34668 34788 34672 34844
rect 34608 34784 34672 34788
rect 34688 34844 34752 34848
rect 34688 34788 34692 34844
rect 34692 34788 34748 34844
rect 34748 34788 34752 34844
rect 34688 34784 34752 34788
rect 34768 34844 34832 34848
rect 34768 34788 34772 34844
rect 34772 34788 34828 34844
rect 34828 34788 34832 34844
rect 34768 34784 34832 34788
rect 5149 34300 5213 34304
rect 5149 34244 5153 34300
rect 5153 34244 5209 34300
rect 5209 34244 5213 34300
rect 5149 34240 5213 34244
rect 5229 34300 5293 34304
rect 5229 34244 5233 34300
rect 5233 34244 5289 34300
rect 5289 34244 5293 34300
rect 5229 34240 5293 34244
rect 5309 34300 5373 34304
rect 5309 34244 5313 34300
rect 5313 34244 5369 34300
rect 5369 34244 5373 34300
rect 5309 34240 5373 34244
rect 5389 34300 5453 34304
rect 5389 34244 5393 34300
rect 5393 34244 5449 34300
rect 5449 34244 5453 34300
rect 5389 34240 5453 34244
rect 13543 34300 13607 34304
rect 13543 34244 13547 34300
rect 13547 34244 13603 34300
rect 13603 34244 13607 34300
rect 13543 34240 13607 34244
rect 13623 34300 13687 34304
rect 13623 34244 13627 34300
rect 13627 34244 13683 34300
rect 13683 34244 13687 34300
rect 13623 34240 13687 34244
rect 13703 34300 13767 34304
rect 13703 34244 13707 34300
rect 13707 34244 13763 34300
rect 13763 34244 13767 34300
rect 13703 34240 13767 34244
rect 13783 34300 13847 34304
rect 13783 34244 13787 34300
rect 13787 34244 13843 34300
rect 13843 34244 13847 34300
rect 13783 34240 13847 34244
rect 21937 34300 22001 34304
rect 21937 34244 21941 34300
rect 21941 34244 21997 34300
rect 21997 34244 22001 34300
rect 21937 34240 22001 34244
rect 22017 34300 22081 34304
rect 22017 34244 22021 34300
rect 22021 34244 22077 34300
rect 22077 34244 22081 34300
rect 22017 34240 22081 34244
rect 22097 34300 22161 34304
rect 22097 34244 22101 34300
rect 22101 34244 22157 34300
rect 22157 34244 22161 34300
rect 22097 34240 22161 34244
rect 22177 34300 22241 34304
rect 22177 34244 22181 34300
rect 22181 34244 22237 34300
rect 22237 34244 22241 34300
rect 22177 34240 22241 34244
rect 30331 34300 30395 34304
rect 30331 34244 30335 34300
rect 30335 34244 30391 34300
rect 30391 34244 30395 34300
rect 30331 34240 30395 34244
rect 30411 34300 30475 34304
rect 30411 34244 30415 34300
rect 30415 34244 30471 34300
rect 30471 34244 30475 34300
rect 30411 34240 30475 34244
rect 30491 34300 30555 34304
rect 30491 34244 30495 34300
rect 30495 34244 30551 34300
rect 30551 34244 30555 34300
rect 30491 34240 30555 34244
rect 30571 34300 30635 34304
rect 30571 34244 30575 34300
rect 30575 34244 30631 34300
rect 30631 34244 30635 34300
rect 30571 34240 30635 34244
rect 9346 33756 9410 33760
rect 9346 33700 9350 33756
rect 9350 33700 9406 33756
rect 9406 33700 9410 33756
rect 9346 33696 9410 33700
rect 9426 33756 9490 33760
rect 9426 33700 9430 33756
rect 9430 33700 9486 33756
rect 9486 33700 9490 33756
rect 9426 33696 9490 33700
rect 9506 33756 9570 33760
rect 9506 33700 9510 33756
rect 9510 33700 9566 33756
rect 9566 33700 9570 33756
rect 9506 33696 9570 33700
rect 9586 33756 9650 33760
rect 9586 33700 9590 33756
rect 9590 33700 9646 33756
rect 9646 33700 9650 33756
rect 9586 33696 9650 33700
rect 17740 33756 17804 33760
rect 17740 33700 17744 33756
rect 17744 33700 17800 33756
rect 17800 33700 17804 33756
rect 17740 33696 17804 33700
rect 17820 33756 17884 33760
rect 17820 33700 17824 33756
rect 17824 33700 17880 33756
rect 17880 33700 17884 33756
rect 17820 33696 17884 33700
rect 17900 33756 17964 33760
rect 17900 33700 17904 33756
rect 17904 33700 17960 33756
rect 17960 33700 17964 33756
rect 17900 33696 17964 33700
rect 17980 33756 18044 33760
rect 17980 33700 17984 33756
rect 17984 33700 18040 33756
rect 18040 33700 18044 33756
rect 17980 33696 18044 33700
rect 26134 33756 26198 33760
rect 26134 33700 26138 33756
rect 26138 33700 26194 33756
rect 26194 33700 26198 33756
rect 26134 33696 26198 33700
rect 26214 33756 26278 33760
rect 26214 33700 26218 33756
rect 26218 33700 26274 33756
rect 26274 33700 26278 33756
rect 26214 33696 26278 33700
rect 26294 33756 26358 33760
rect 26294 33700 26298 33756
rect 26298 33700 26354 33756
rect 26354 33700 26358 33756
rect 26294 33696 26358 33700
rect 26374 33756 26438 33760
rect 26374 33700 26378 33756
rect 26378 33700 26434 33756
rect 26434 33700 26438 33756
rect 26374 33696 26438 33700
rect 34528 33756 34592 33760
rect 34528 33700 34532 33756
rect 34532 33700 34588 33756
rect 34588 33700 34592 33756
rect 34528 33696 34592 33700
rect 34608 33756 34672 33760
rect 34608 33700 34612 33756
rect 34612 33700 34668 33756
rect 34668 33700 34672 33756
rect 34608 33696 34672 33700
rect 34688 33756 34752 33760
rect 34688 33700 34692 33756
rect 34692 33700 34748 33756
rect 34748 33700 34752 33756
rect 34688 33696 34752 33700
rect 34768 33756 34832 33760
rect 34768 33700 34772 33756
rect 34772 33700 34828 33756
rect 34828 33700 34832 33756
rect 34768 33696 34832 33700
rect 5149 33212 5213 33216
rect 5149 33156 5153 33212
rect 5153 33156 5209 33212
rect 5209 33156 5213 33212
rect 5149 33152 5213 33156
rect 5229 33212 5293 33216
rect 5229 33156 5233 33212
rect 5233 33156 5289 33212
rect 5289 33156 5293 33212
rect 5229 33152 5293 33156
rect 5309 33212 5373 33216
rect 5309 33156 5313 33212
rect 5313 33156 5369 33212
rect 5369 33156 5373 33212
rect 5309 33152 5373 33156
rect 5389 33212 5453 33216
rect 5389 33156 5393 33212
rect 5393 33156 5449 33212
rect 5449 33156 5453 33212
rect 5389 33152 5453 33156
rect 13543 33212 13607 33216
rect 13543 33156 13547 33212
rect 13547 33156 13603 33212
rect 13603 33156 13607 33212
rect 13543 33152 13607 33156
rect 13623 33212 13687 33216
rect 13623 33156 13627 33212
rect 13627 33156 13683 33212
rect 13683 33156 13687 33212
rect 13623 33152 13687 33156
rect 13703 33212 13767 33216
rect 13703 33156 13707 33212
rect 13707 33156 13763 33212
rect 13763 33156 13767 33212
rect 13703 33152 13767 33156
rect 13783 33212 13847 33216
rect 13783 33156 13787 33212
rect 13787 33156 13843 33212
rect 13843 33156 13847 33212
rect 13783 33152 13847 33156
rect 21937 33212 22001 33216
rect 21937 33156 21941 33212
rect 21941 33156 21997 33212
rect 21997 33156 22001 33212
rect 21937 33152 22001 33156
rect 22017 33212 22081 33216
rect 22017 33156 22021 33212
rect 22021 33156 22077 33212
rect 22077 33156 22081 33212
rect 22017 33152 22081 33156
rect 22097 33212 22161 33216
rect 22097 33156 22101 33212
rect 22101 33156 22157 33212
rect 22157 33156 22161 33212
rect 22097 33152 22161 33156
rect 22177 33212 22241 33216
rect 22177 33156 22181 33212
rect 22181 33156 22237 33212
rect 22237 33156 22241 33212
rect 22177 33152 22241 33156
rect 30331 33212 30395 33216
rect 30331 33156 30335 33212
rect 30335 33156 30391 33212
rect 30391 33156 30395 33212
rect 30331 33152 30395 33156
rect 30411 33212 30475 33216
rect 30411 33156 30415 33212
rect 30415 33156 30471 33212
rect 30471 33156 30475 33212
rect 30411 33152 30475 33156
rect 30491 33212 30555 33216
rect 30491 33156 30495 33212
rect 30495 33156 30551 33212
rect 30551 33156 30555 33212
rect 30491 33152 30555 33156
rect 30571 33212 30635 33216
rect 30571 33156 30575 33212
rect 30575 33156 30631 33212
rect 30631 33156 30635 33212
rect 30571 33152 30635 33156
rect 9346 32668 9410 32672
rect 9346 32612 9350 32668
rect 9350 32612 9406 32668
rect 9406 32612 9410 32668
rect 9346 32608 9410 32612
rect 9426 32668 9490 32672
rect 9426 32612 9430 32668
rect 9430 32612 9486 32668
rect 9486 32612 9490 32668
rect 9426 32608 9490 32612
rect 9506 32668 9570 32672
rect 9506 32612 9510 32668
rect 9510 32612 9566 32668
rect 9566 32612 9570 32668
rect 9506 32608 9570 32612
rect 9586 32668 9650 32672
rect 9586 32612 9590 32668
rect 9590 32612 9646 32668
rect 9646 32612 9650 32668
rect 9586 32608 9650 32612
rect 17740 32668 17804 32672
rect 17740 32612 17744 32668
rect 17744 32612 17800 32668
rect 17800 32612 17804 32668
rect 17740 32608 17804 32612
rect 17820 32668 17884 32672
rect 17820 32612 17824 32668
rect 17824 32612 17880 32668
rect 17880 32612 17884 32668
rect 17820 32608 17884 32612
rect 17900 32668 17964 32672
rect 17900 32612 17904 32668
rect 17904 32612 17960 32668
rect 17960 32612 17964 32668
rect 17900 32608 17964 32612
rect 17980 32668 18044 32672
rect 17980 32612 17984 32668
rect 17984 32612 18040 32668
rect 18040 32612 18044 32668
rect 17980 32608 18044 32612
rect 26134 32668 26198 32672
rect 26134 32612 26138 32668
rect 26138 32612 26194 32668
rect 26194 32612 26198 32668
rect 26134 32608 26198 32612
rect 26214 32668 26278 32672
rect 26214 32612 26218 32668
rect 26218 32612 26274 32668
rect 26274 32612 26278 32668
rect 26214 32608 26278 32612
rect 26294 32668 26358 32672
rect 26294 32612 26298 32668
rect 26298 32612 26354 32668
rect 26354 32612 26358 32668
rect 26294 32608 26358 32612
rect 26374 32668 26438 32672
rect 26374 32612 26378 32668
rect 26378 32612 26434 32668
rect 26434 32612 26438 32668
rect 26374 32608 26438 32612
rect 34528 32668 34592 32672
rect 34528 32612 34532 32668
rect 34532 32612 34588 32668
rect 34588 32612 34592 32668
rect 34528 32608 34592 32612
rect 34608 32668 34672 32672
rect 34608 32612 34612 32668
rect 34612 32612 34668 32668
rect 34668 32612 34672 32668
rect 34608 32608 34672 32612
rect 34688 32668 34752 32672
rect 34688 32612 34692 32668
rect 34692 32612 34748 32668
rect 34748 32612 34752 32668
rect 34688 32608 34752 32612
rect 34768 32668 34832 32672
rect 34768 32612 34772 32668
rect 34772 32612 34828 32668
rect 34828 32612 34832 32668
rect 34768 32608 34832 32612
rect 5149 32124 5213 32128
rect 5149 32068 5153 32124
rect 5153 32068 5209 32124
rect 5209 32068 5213 32124
rect 5149 32064 5213 32068
rect 5229 32124 5293 32128
rect 5229 32068 5233 32124
rect 5233 32068 5289 32124
rect 5289 32068 5293 32124
rect 5229 32064 5293 32068
rect 5309 32124 5373 32128
rect 5309 32068 5313 32124
rect 5313 32068 5369 32124
rect 5369 32068 5373 32124
rect 5309 32064 5373 32068
rect 5389 32124 5453 32128
rect 5389 32068 5393 32124
rect 5393 32068 5449 32124
rect 5449 32068 5453 32124
rect 5389 32064 5453 32068
rect 13543 32124 13607 32128
rect 13543 32068 13547 32124
rect 13547 32068 13603 32124
rect 13603 32068 13607 32124
rect 13543 32064 13607 32068
rect 13623 32124 13687 32128
rect 13623 32068 13627 32124
rect 13627 32068 13683 32124
rect 13683 32068 13687 32124
rect 13623 32064 13687 32068
rect 13703 32124 13767 32128
rect 13703 32068 13707 32124
rect 13707 32068 13763 32124
rect 13763 32068 13767 32124
rect 13703 32064 13767 32068
rect 13783 32124 13847 32128
rect 13783 32068 13787 32124
rect 13787 32068 13843 32124
rect 13843 32068 13847 32124
rect 13783 32064 13847 32068
rect 21937 32124 22001 32128
rect 21937 32068 21941 32124
rect 21941 32068 21997 32124
rect 21997 32068 22001 32124
rect 21937 32064 22001 32068
rect 22017 32124 22081 32128
rect 22017 32068 22021 32124
rect 22021 32068 22077 32124
rect 22077 32068 22081 32124
rect 22017 32064 22081 32068
rect 22097 32124 22161 32128
rect 22097 32068 22101 32124
rect 22101 32068 22157 32124
rect 22157 32068 22161 32124
rect 22097 32064 22161 32068
rect 22177 32124 22241 32128
rect 22177 32068 22181 32124
rect 22181 32068 22237 32124
rect 22237 32068 22241 32124
rect 22177 32064 22241 32068
rect 30331 32124 30395 32128
rect 30331 32068 30335 32124
rect 30335 32068 30391 32124
rect 30391 32068 30395 32124
rect 30331 32064 30395 32068
rect 30411 32124 30475 32128
rect 30411 32068 30415 32124
rect 30415 32068 30471 32124
rect 30471 32068 30475 32124
rect 30411 32064 30475 32068
rect 30491 32124 30555 32128
rect 30491 32068 30495 32124
rect 30495 32068 30551 32124
rect 30551 32068 30555 32124
rect 30491 32064 30555 32068
rect 30571 32124 30635 32128
rect 30571 32068 30575 32124
rect 30575 32068 30631 32124
rect 30631 32068 30635 32124
rect 30571 32064 30635 32068
rect 9346 31580 9410 31584
rect 9346 31524 9350 31580
rect 9350 31524 9406 31580
rect 9406 31524 9410 31580
rect 9346 31520 9410 31524
rect 9426 31580 9490 31584
rect 9426 31524 9430 31580
rect 9430 31524 9486 31580
rect 9486 31524 9490 31580
rect 9426 31520 9490 31524
rect 9506 31580 9570 31584
rect 9506 31524 9510 31580
rect 9510 31524 9566 31580
rect 9566 31524 9570 31580
rect 9506 31520 9570 31524
rect 9586 31580 9650 31584
rect 9586 31524 9590 31580
rect 9590 31524 9646 31580
rect 9646 31524 9650 31580
rect 9586 31520 9650 31524
rect 17740 31580 17804 31584
rect 17740 31524 17744 31580
rect 17744 31524 17800 31580
rect 17800 31524 17804 31580
rect 17740 31520 17804 31524
rect 17820 31580 17884 31584
rect 17820 31524 17824 31580
rect 17824 31524 17880 31580
rect 17880 31524 17884 31580
rect 17820 31520 17884 31524
rect 17900 31580 17964 31584
rect 17900 31524 17904 31580
rect 17904 31524 17960 31580
rect 17960 31524 17964 31580
rect 17900 31520 17964 31524
rect 17980 31580 18044 31584
rect 17980 31524 17984 31580
rect 17984 31524 18040 31580
rect 18040 31524 18044 31580
rect 17980 31520 18044 31524
rect 26134 31580 26198 31584
rect 26134 31524 26138 31580
rect 26138 31524 26194 31580
rect 26194 31524 26198 31580
rect 26134 31520 26198 31524
rect 26214 31580 26278 31584
rect 26214 31524 26218 31580
rect 26218 31524 26274 31580
rect 26274 31524 26278 31580
rect 26214 31520 26278 31524
rect 26294 31580 26358 31584
rect 26294 31524 26298 31580
rect 26298 31524 26354 31580
rect 26354 31524 26358 31580
rect 26294 31520 26358 31524
rect 26374 31580 26438 31584
rect 26374 31524 26378 31580
rect 26378 31524 26434 31580
rect 26434 31524 26438 31580
rect 26374 31520 26438 31524
rect 34528 31580 34592 31584
rect 34528 31524 34532 31580
rect 34532 31524 34588 31580
rect 34588 31524 34592 31580
rect 34528 31520 34592 31524
rect 34608 31580 34672 31584
rect 34608 31524 34612 31580
rect 34612 31524 34668 31580
rect 34668 31524 34672 31580
rect 34608 31520 34672 31524
rect 34688 31580 34752 31584
rect 34688 31524 34692 31580
rect 34692 31524 34748 31580
rect 34748 31524 34752 31580
rect 34688 31520 34752 31524
rect 34768 31580 34832 31584
rect 34768 31524 34772 31580
rect 34772 31524 34828 31580
rect 34828 31524 34832 31580
rect 34768 31520 34832 31524
rect 5149 31036 5213 31040
rect 5149 30980 5153 31036
rect 5153 30980 5209 31036
rect 5209 30980 5213 31036
rect 5149 30976 5213 30980
rect 5229 31036 5293 31040
rect 5229 30980 5233 31036
rect 5233 30980 5289 31036
rect 5289 30980 5293 31036
rect 5229 30976 5293 30980
rect 5309 31036 5373 31040
rect 5309 30980 5313 31036
rect 5313 30980 5369 31036
rect 5369 30980 5373 31036
rect 5309 30976 5373 30980
rect 5389 31036 5453 31040
rect 5389 30980 5393 31036
rect 5393 30980 5449 31036
rect 5449 30980 5453 31036
rect 5389 30976 5453 30980
rect 13543 31036 13607 31040
rect 13543 30980 13547 31036
rect 13547 30980 13603 31036
rect 13603 30980 13607 31036
rect 13543 30976 13607 30980
rect 13623 31036 13687 31040
rect 13623 30980 13627 31036
rect 13627 30980 13683 31036
rect 13683 30980 13687 31036
rect 13623 30976 13687 30980
rect 13703 31036 13767 31040
rect 13703 30980 13707 31036
rect 13707 30980 13763 31036
rect 13763 30980 13767 31036
rect 13703 30976 13767 30980
rect 13783 31036 13847 31040
rect 13783 30980 13787 31036
rect 13787 30980 13843 31036
rect 13843 30980 13847 31036
rect 13783 30976 13847 30980
rect 21937 31036 22001 31040
rect 21937 30980 21941 31036
rect 21941 30980 21997 31036
rect 21997 30980 22001 31036
rect 21937 30976 22001 30980
rect 22017 31036 22081 31040
rect 22017 30980 22021 31036
rect 22021 30980 22077 31036
rect 22077 30980 22081 31036
rect 22017 30976 22081 30980
rect 22097 31036 22161 31040
rect 22097 30980 22101 31036
rect 22101 30980 22157 31036
rect 22157 30980 22161 31036
rect 22097 30976 22161 30980
rect 22177 31036 22241 31040
rect 22177 30980 22181 31036
rect 22181 30980 22237 31036
rect 22237 30980 22241 31036
rect 22177 30976 22241 30980
rect 30331 31036 30395 31040
rect 30331 30980 30335 31036
rect 30335 30980 30391 31036
rect 30391 30980 30395 31036
rect 30331 30976 30395 30980
rect 30411 31036 30475 31040
rect 30411 30980 30415 31036
rect 30415 30980 30471 31036
rect 30471 30980 30475 31036
rect 30411 30976 30475 30980
rect 30491 31036 30555 31040
rect 30491 30980 30495 31036
rect 30495 30980 30551 31036
rect 30551 30980 30555 31036
rect 30491 30976 30555 30980
rect 30571 31036 30635 31040
rect 30571 30980 30575 31036
rect 30575 30980 30631 31036
rect 30631 30980 30635 31036
rect 30571 30976 30635 30980
rect 9346 30492 9410 30496
rect 9346 30436 9350 30492
rect 9350 30436 9406 30492
rect 9406 30436 9410 30492
rect 9346 30432 9410 30436
rect 9426 30492 9490 30496
rect 9426 30436 9430 30492
rect 9430 30436 9486 30492
rect 9486 30436 9490 30492
rect 9426 30432 9490 30436
rect 9506 30492 9570 30496
rect 9506 30436 9510 30492
rect 9510 30436 9566 30492
rect 9566 30436 9570 30492
rect 9506 30432 9570 30436
rect 9586 30492 9650 30496
rect 9586 30436 9590 30492
rect 9590 30436 9646 30492
rect 9646 30436 9650 30492
rect 9586 30432 9650 30436
rect 17740 30492 17804 30496
rect 17740 30436 17744 30492
rect 17744 30436 17800 30492
rect 17800 30436 17804 30492
rect 17740 30432 17804 30436
rect 17820 30492 17884 30496
rect 17820 30436 17824 30492
rect 17824 30436 17880 30492
rect 17880 30436 17884 30492
rect 17820 30432 17884 30436
rect 17900 30492 17964 30496
rect 17900 30436 17904 30492
rect 17904 30436 17960 30492
rect 17960 30436 17964 30492
rect 17900 30432 17964 30436
rect 17980 30492 18044 30496
rect 17980 30436 17984 30492
rect 17984 30436 18040 30492
rect 18040 30436 18044 30492
rect 17980 30432 18044 30436
rect 26134 30492 26198 30496
rect 26134 30436 26138 30492
rect 26138 30436 26194 30492
rect 26194 30436 26198 30492
rect 26134 30432 26198 30436
rect 26214 30492 26278 30496
rect 26214 30436 26218 30492
rect 26218 30436 26274 30492
rect 26274 30436 26278 30492
rect 26214 30432 26278 30436
rect 26294 30492 26358 30496
rect 26294 30436 26298 30492
rect 26298 30436 26354 30492
rect 26354 30436 26358 30492
rect 26294 30432 26358 30436
rect 26374 30492 26438 30496
rect 26374 30436 26378 30492
rect 26378 30436 26434 30492
rect 26434 30436 26438 30492
rect 26374 30432 26438 30436
rect 34528 30492 34592 30496
rect 34528 30436 34532 30492
rect 34532 30436 34588 30492
rect 34588 30436 34592 30492
rect 34528 30432 34592 30436
rect 34608 30492 34672 30496
rect 34608 30436 34612 30492
rect 34612 30436 34668 30492
rect 34668 30436 34672 30492
rect 34608 30432 34672 30436
rect 34688 30492 34752 30496
rect 34688 30436 34692 30492
rect 34692 30436 34748 30492
rect 34748 30436 34752 30492
rect 34688 30432 34752 30436
rect 34768 30492 34832 30496
rect 34768 30436 34772 30492
rect 34772 30436 34828 30492
rect 34828 30436 34832 30492
rect 34768 30432 34832 30436
rect 5149 29948 5213 29952
rect 5149 29892 5153 29948
rect 5153 29892 5209 29948
rect 5209 29892 5213 29948
rect 5149 29888 5213 29892
rect 5229 29948 5293 29952
rect 5229 29892 5233 29948
rect 5233 29892 5289 29948
rect 5289 29892 5293 29948
rect 5229 29888 5293 29892
rect 5309 29948 5373 29952
rect 5309 29892 5313 29948
rect 5313 29892 5369 29948
rect 5369 29892 5373 29948
rect 5309 29888 5373 29892
rect 5389 29948 5453 29952
rect 5389 29892 5393 29948
rect 5393 29892 5449 29948
rect 5449 29892 5453 29948
rect 5389 29888 5453 29892
rect 13543 29948 13607 29952
rect 13543 29892 13547 29948
rect 13547 29892 13603 29948
rect 13603 29892 13607 29948
rect 13543 29888 13607 29892
rect 13623 29948 13687 29952
rect 13623 29892 13627 29948
rect 13627 29892 13683 29948
rect 13683 29892 13687 29948
rect 13623 29888 13687 29892
rect 13703 29948 13767 29952
rect 13703 29892 13707 29948
rect 13707 29892 13763 29948
rect 13763 29892 13767 29948
rect 13703 29888 13767 29892
rect 13783 29948 13847 29952
rect 13783 29892 13787 29948
rect 13787 29892 13843 29948
rect 13843 29892 13847 29948
rect 13783 29888 13847 29892
rect 21937 29948 22001 29952
rect 21937 29892 21941 29948
rect 21941 29892 21997 29948
rect 21997 29892 22001 29948
rect 21937 29888 22001 29892
rect 22017 29948 22081 29952
rect 22017 29892 22021 29948
rect 22021 29892 22077 29948
rect 22077 29892 22081 29948
rect 22017 29888 22081 29892
rect 22097 29948 22161 29952
rect 22097 29892 22101 29948
rect 22101 29892 22157 29948
rect 22157 29892 22161 29948
rect 22097 29888 22161 29892
rect 22177 29948 22241 29952
rect 22177 29892 22181 29948
rect 22181 29892 22237 29948
rect 22237 29892 22241 29948
rect 22177 29888 22241 29892
rect 30331 29948 30395 29952
rect 30331 29892 30335 29948
rect 30335 29892 30391 29948
rect 30391 29892 30395 29948
rect 30331 29888 30395 29892
rect 30411 29948 30475 29952
rect 30411 29892 30415 29948
rect 30415 29892 30471 29948
rect 30471 29892 30475 29948
rect 30411 29888 30475 29892
rect 30491 29948 30555 29952
rect 30491 29892 30495 29948
rect 30495 29892 30551 29948
rect 30551 29892 30555 29948
rect 30491 29888 30555 29892
rect 30571 29948 30635 29952
rect 30571 29892 30575 29948
rect 30575 29892 30631 29948
rect 30631 29892 30635 29948
rect 30571 29888 30635 29892
rect 9346 29404 9410 29408
rect 9346 29348 9350 29404
rect 9350 29348 9406 29404
rect 9406 29348 9410 29404
rect 9346 29344 9410 29348
rect 9426 29404 9490 29408
rect 9426 29348 9430 29404
rect 9430 29348 9486 29404
rect 9486 29348 9490 29404
rect 9426 29344 9490 29348
rect 9506 29404 9570 29408
rect 9506 29348 9510 29404
rect 9510 29348 9566 29404
rect 9566 29348 9570 29404
rect 9506 29344 9570 29348
rect 9586 29404 9650 29408
rect 9586 29348 9590 29404
rect 9590 29348 9646 29404
rect 9646 29348 9650 29404
rect 9586 29344 9650 29348
rect 17740 29404 17804 29408
rect 17740 29348 17744 29404
rect 17744 29348 17800 29404
rect 17800 29348 17804 29404
rect 17740 29344 17804 29348
rect 17820 29404 17884 29408
rect 17820 29348 17824 29404
rect 17824 29348 17880 29404
rect 17880 29348 17884 29404
rect 17820 29344 17884 29348
rect 17900 29404 17964 29408
rect 17900 29348 17904 29404
rect 17904 29348 17960 29404
rect 17960 29348 17964 29404
rect 17900 29344 17964 29348
rect 17980 29404 18044 29408
rect 17980 29348 17984 29404
rect 17984 29348 18040 29404
rect 18040 29348 18044 29404
rect 17980 29344 18044 29348
rect 26134 29404 26198 29408
rect 26134 29348 26138 29404
rect 26138 29348 26194 29404
rect 26194 29348 26198 29404
rect 26134 29344 26198 29348
rect 26214 29404 26278 29408
rect 26214 29348 26218 29404
rect 26218 29348 26274 29404
rect 26274 29348 26278 29404
rect 26214 29344 26278 29348
rect 26294 29404 26358 29408
rect 26294 29348 26298 29404
rect 26298 29348 26354 29404
rect 26354 29348 26358 29404
rect 26294 29344 26358 29348
rect 26374 29404 26438 29408
rect 26374 29348 26378 29404
rect 26378 29348 26434 29404
rect 26434 29348 26438 29404
rect 26374 29344 26438 29348
rect 34528 29404 34592 29408
rect 34528 29348 34532 29404
rect 34532 29348 34588 29404
rect 34588 29348 34592 29404
rect 34528 29344 34592 29348
rect 34608 29404 34672 29408
rect 34608 29348 34612 29404
rect 34612 29348 34668 29404
rect 34668 29348 34672 29404
rect 34608 29344 34672 29348
rect 34688 29404 34752 29408
rect 34688 29348 34692 29404
rect 34692 29348 34748 29404
rect 34748 29348 34752 29404
rect 34688 29344 34752 29348
rect 34768 29404 34832 29408
rect 34768 29348 34772 29404
rect 34772 29348 34828 29404
rect 34828 29348 34832 29404
rect 34768 29344 34832 29348
rect 5149 28860 5213 28864
rect 5149 28804 5153 28860
rect 5153 28804 5209 28860
rect 5209 28804 5213 28860
rect 5149 28800 5213 28804
rect 5229 28860 5293 28864
rect 5229 28804 5233 28860
rect 5233 28804 5289 28860
rect 5289 28804 5293 28860
rect 5229 28800 5293 28804
rect 5309 28860 5373 28864
rect 5309 28804 5313 28860
rect 5313 28804 5369 28860
rect 5369 28804 5373 28860
rect 5309 28800 5373 28804
rect 5389 28860 5453 28864
rect 5389 28804 5393 28860
rect 5393 28804 5449 28860
rect 5449 28804 5453 28860
rect 5389 28800 5453 28804
rect 13543 28860 13607 28864
rect 13543 28804 13547 28860
rect 13547 28804 13603 28860
rect 13603 28804 13607 28860
rect 13543 28800 13607 28804
rect 13623 28860 13687 28864
rect 13623 28804 13627 28860
rect 13627 28804 13683 28860
rect 13683 28804 13687 28860
rect 13623 28800 13687 28804
rect 13703 28860 13767 28864
rect 13703 28804 13707 28860
rect 13707 28804 13763 28860
rect 13763 28804 13767 28860
rect 13703 28800 13767 28804
rect 13783 28860 13847 28864
rect 13783 28804 13787 28860
rect 13787 28804 13843 28860
rect 13843 28804 13847 28860
rect 13783 28800 13847 28804
rect 21937 28860 22001 28864
rect 21937 28804 21941 28860
rect 21941 28804 21997 28860
rect 21997 28804 22001 28860
rect 21937 28800 22001 28804
rect 22017 28860 22081 28864
rect 22017 28804 22021 28860
rect 22021 28804 22077 28860
rect 22077 28804 22081 28860
rect 22017 28800 22081 28804
rect 22097 28860 22161 28864
rect 22097 28804 22101 28860
rect 22101 28804 22157 28860
rect 22157 28804 22161 28860
rect 22097 28800 22161 28804
rect 22177 28860 22241 28864
rect 22177 28804 22181 28860
rect 22181 28804 22237 28860
rect 22237 28804 22241 28860
rect 22177 28800 22241 28804
rect 30331 28860 30395 28864
rect 30331 28804 30335 28860
rect 30335 28804 30391 28860
rect 30391 28804 30395 28860
rect 30331 28800 30395 28804
rect 30411 28860 30475 28864
rect 30411 28804 30415 28860
rect 30415 28804 30471 28860
rect 30471 28804 30475 28860
rect 30411 28800 30475 28804
rect 30491 28860 30555 28864
rect 30491 28804 30495 28860
rect 30495 28804 30551 28860
rect 30551 28804 30555 28860
rect 30491 28800 30555 28804
rect 30571 28860 30635 28864
rect 30571 28804 30575 28860
rect 30575 28804 30631 28860
rect 30631 28804 30635 28860
rect 30571 28800 30635 28804
rect 9346 28316 9410 28320
rect 9346 28260 9350 28316
rect 9350 28260 9406 28316
rect 9406 28260 9410 28316
rect 9346 28256 9410 28260
rect 9426 28316 9490 28320
rect 9426 28260 9430 28316
rect 9430 28260 9486 28316
rect 9486 28260 9490 28316
rect 9426 28256 9490 28260
rect 9506 28316 9570 28320
rect 9506 28260 9510 28316
rect 9510 28260 9566 28316
rect 9566 28260 9570 28316
rect 9506 28256 9570 28260
rect 9586 28316 9650 28320
rect 9586 28260 9590 28316
rect 9590 28260 9646 28316
rect 9646 28260 9650 28316
rect 9586 28256 9650 28260
rect 17740 28316 17804 28320
rect 17740 28260 17744 28316
rect 17744 28260 17800 28316
rect 17800 28260 17804 28316
rect 17740 28256 17804 28260
rect 17820 28316 17884 28320
rect 17820 28260 17824 28316
rect 17824 28260 17880 28316
rect 17880 28260 17884 28316
rect 17820 28256 17884 28260
rect 17900 28316 17964 28320
rect 17900 28260 17904 28316
rect 17904 28260 17960 28316
rect 17960 28260 17964 28316
rect 17900 28256 17964 28260
rect 17980 28316 18044 28320
rect 17980 28260 17984 28316
rect 17984 28260 18040 28316
rect 18040 28260 18044 28316
rect 17980 28256 18044 28260
rect 26134 28316 26198 28320
rect 26134 28260 26138 28316
rect 26138 28260 26194 28316
rect 26194 28260 26198 28316
rect 26134 28256 26198 28260
rect 26214 28316 26278 28320
rect 26214 28260 26218 28316
rect 26218 28260 26274 28316
rect 26274 28260 26278 28316
rect 26214 28256 26278 28260
rect 26294 28316 26358 28320
rect 26294 28260 26298 28316
rect 26298 28260 26354 28316
rect 26354 28260 26358 28316
rect 26294 28256 26358 28260
rect 26374 28316 26438 28320
rect 26374 28260 26378 28316
rect 26378 28260 26434 28316
rect 26434 28260 26438 28316
rect 26374 28256 26438 28260
rect 34528 28316 34592 28320
rect 34528 28260 34532 28316
rect 34532 28260 34588 28316
rect 34588 28260 34592 28316
rect 34528 28256 34592 28260
rect 34608 28316 34672 28320
rect 34608 28260 34612 28316
rect 34612 28260 34668 28316
rect 34668 28260 34672 28316
rect 34608 28256 34672 28260
rect 34688 28316 34752 28320
rect 34688 28260 34692 28316
rect 34692 28260 34748 28316
rect 34748 28260 34752 28316
rect 34688 28256 34752 28260
rect 34768 28316 34832 28320
rect 34768 28260 34772 28316
rect 34772 28260 34828 28316
rect 34828 28260 34832 28316
rect 34768 28256 34832 28260
rect 5149 27772 5213 27776
rect 5149 27716 5153 27772
rect 5153 27716 5209 27772
rect 5209 27716 5213 27772
rect 5149 27712 5213 27716
rect 5229 27772 5293 27776
rect 5229 27716 5233 27772
rect 5233 27716 5289 27772
rect 5289 27716 5293 27772
rect 5229 27712 5293 27716
rect 5309 27772 5373 27776
rect 5309 27716 5313 27772
rect 5313 27716 5369 27772
rect 5369 27716 5373 27772
rect 5309 27712 5373 27716
rect 5389 27772 5453 27776
rect 5389 27716 5393 27772
rect 5393 27716 5449 27772
rect 5449 27716 5453 27772
rect 5389 27712 5453 27716
rect 13543 27772 13607 27776
rect 13543 27716 13547 27772
rect 13547 27716 13603 27772
rect 13603 27716 13607 27772
rect 13543 27712 13607 27716
rect 13623 27772 13687 27776
rect 13623 27716 13627 27772
rect 13627 27716 13683 27772
rect 13683 27716 13687 27772
rect 13623 27712 13687 27716
rect 13703 27772 13767 27776
rect 13703 27716 13707 27772
rect 13707 27716 13763 27772
rect 13763 27716 13767 27772
rect 13703 27712 13767 27716
rect 13783 27772 13847 27776
rect 13783 27716 13787 27772
rect 13787 27716 13843 27772
rect 13843 27716 13847 27772
rect 13783 27712 13847 27716
rect 21937 27772 22001 27776
rect 21937 27716 21941 27772
rect 21941 27716 21997 27772
rect 21997 27716 22001 27772
rect 21937 27712 22001 27716
rect 22017 27772 22081 27776
rect 22017 27716 22021 27772
rect 22021 27716 22077 27772
rect 22077 27716 22081 27772
rect 22017 27712 22081 27716
rect 22097 27772 22161 27776
rect 22097 27716 22101 27772
rect 22101 27716 22157 27772
rect 22157 27716 22161 27772
rect 22097 27712 22161 27716
rect 22177 27772 22241 27776
rect 22177 27716 22181 27772
rect 22181 27716 22237 27772
rect 22237 27716 22241 27772
rect 22177 27712 22241 27716
rect 30331 27772 30395 27776
rect 30331 27716 30335 27772
rect 30335 27716 30391 27772
rect 30391 27716 30395 27772
rect 30331 27712 30395 27716
rect 30411 27772 30475 27776
rect 30411 27716 30415 27772
rect 30415 27716 30471 27772
rect 30471 27716 30475 27772
rect 30411 27712 30475 27716
rect 30491 27772 30555 27776
rect 30491 27716 30495 27772
rect 30495 27716 30551 27772
rect 30551 27716 30555 27772
rect 30491 27712 30555 27716
rect 30571 27772 30635 27776
rect 30571 27716 30575 27772
rect 30575 27716 30631 27772
rect 30631 27716 30635 27772
rect 30571 27712 30635 27716
rect 9346 27228 9410 27232
rect 9346 27172 9350 27228
rect 9350 27172 9406 27228
rect 9406 27172 9410 27228
rect 9346 27168 9410 27172
rect 9426 27228 9490 27232
rect 9426 27172 9430 27228
rect 9430 27172 9486 27228
rect 9486 27172 9490 27228
rect 9426 27168 9490 27172
rect 9506 27228 9570 27232
rect 9506 27172 9510 27228
rect 9510 27172 9566 27228
rect 9566 27172 9570 27228
rect 9506 27168 9570 27172
rect 9586 27228 9650 27232
rect 9586 27172 9590 27228
rect 9590 27172 9646 27228
rect 9646 27172 9650 27228
rect 9586 27168 9650 27172
rect 17740 27228 17804 27232
rect 17740 27172 17744 27228
rect 17744 27172 17800 27228
rect 17800 27172 17804 27228
rect 17740 27168 17804 27172
rect 17820 27228 17884 27232
rect 17820 27172 17824 27228
rect 17824 27172 17880 27228
rect 17880 27172 17884 27228
rect 17820 27168 17884 27172
rect 17900 27228 17964 27232
rect 17900 27172 17904 27228
rect 17904 27172 17960 27228
rect 17960 27172 17964 27228
rect 17900 27168 17964 27172
rect 17980 27228 18044 27232
rect 17980 27172 17984 27228
rect 17984 27172 18040 27228
rect 18040 27172 18044 27228
rect 17980 27168 18044 27172
rect 26134 27228 26198 27232
rect 26134 27172 26138 27228
rect 26138 27172 26194 27228
rect 26194 27172 26198 27228
rect 26134 27168 26198 27172
rect 26214 27228 26278 27232
rect 26214 27172 26218 27228
rect 26218 27172 26274 27228
rect 26274 27172 26278 27228
rect 26214 27168 26278 27172
rect 26294 27228 26358 27232
rect 26294 27172 26298 27228
rect 26298 27172 26354 27228
rect 26354 27172 26358 27228
rect 26294 27168 26358 27172
rect 26374 27228 26438 27232
rect 26374 27172 26378 27228
rect 26378 27172 26434 27228
rect 26434 27172 26438 27228
rect 26374 27168 26438 27172
rect 34528 27228 34592 27232
rect 34528 27172 34532 27228
rect 34532 27172 34588 27228
rect 34588 27172 34592 27228
rect 34528 27168 34592 27172
rect 34608 27228 34672 27232
rect 34608 27172 34612 27228
rect 34612 27172 34668 27228
rect 34668 27172 34672 27228
rect 34608 27168 34672 27172
rect 34688 27228 34752 27232
rect 34688 27172 34692 27228
rect 34692 27172 34748 27228
rect 34748 27172 34752 27228
rect 34688 27168 34752 27172
rect 34768 27228 34832 27232
rect 34768 27172 34772 27228
rect 34772 27172 34828 27228
rect 34828 27172 34832 27228
rect 34768 27168 34832 27172
rect 5149 26684 5213 26688
rect 5149 26628 5153 26684
rect 5153 26628 5209 26684
rect 5209 26628 5213 26684
rect 5149 26624 5213 26628
rect 5229 26684 5293 26688
rect 5229 26628 5233 26684
rect 5233 26628 5289 26684
rect 5289 26628 5293 26684
rect 5229 26624 5293 26628
rect 5309 26684 5373 26688
rect 5309 26628 5313 26684
rect 5313 26628 5369 26684
rect 5369 26628 5373 26684
rect 5309 26624 5373 26628
rect 5389 26684 5453 26688
rect 5389 26628 5393 26684
rect 5393 26628 5449 26684
rect 5449 26628 5453 26684
rect 5389 26624 5453 26628
rect 13543 26684 13607 26688
rect 13543 26628 13547 26684
rect 13547 26628 13603 26684
rect 13603 26628 13607 26684
rect 13543 26624 13607 26628
rect 13623 26684 13687 26688
rect 13623 26628 13627 26684
rect 13627 26628 13683 26684
rect 13683 26628 13687 26684
rect 13623 26624 13687 26628
rect 13703 26684 13767 26688
rect 13703 26628 13707 26684
rect 13707 26628 13763 26684
rect 13763 26628 13767 26684
rect 13703 26624 13767 26628
rect 13783 26684 13847 26688
rect 13783 26628 13787 26684
rect 13787 26628 13843 26684
rect 13843 26628 13847 26684
rect 13783 26624 13847 26628
rect 21937 26684 22001 26688
rect 21937 26628 21941 26684
rect 21941 26628 21997 26684
rect 21997 26628 22001 26684
rect 21937 26624 22001 26628
rect 22017 26684 22081 26688
rect 22017 26628 22021 26684
rect 22021 26628 22077 26684
rect 22077 26628 22081 26684
rect 22017 26624 22081 26628
rect 22097 26684 22161 26688
rect 22097 26628 22101 26684
rect 22101 26628 22157 26684
rect 22157 26628 22161 26684
rect 22097 26624 22161 26628
rect 22177 26684 22241 26688
rect 22177 26628 22181 26684
rect 22181 26628 22237 26684
rect 22237 26628 22241 26684
rect 22177 26624 22241 26628
rect 30331 26684 30395 26688
rect 30331 26628 30335 26684
rect 30335 26628 30391 26684
rect 30391 26628 30395 26684
rect 30331 26624 30395 26628
rect 30411 26684 30475 26688
rect 30411 26628 30415 26684
rect 30415 26628 30471 26684
rect 30471 26628 30475 26684
rect 30411 26624 30475 26628
rect 30491 26684 30555 26688
rect 30491 26628 30495 26684
rect 30495 26628 30551 26684
rect 30551 26628 30555 26684
rect 30491 26624 30555 26628
rect 30571 26684 30635 26688
rect 30571 26628 30575 26684
rect 30575 26628 30631 26684
rect 30631 26628 30635 26684
rect 30571 26624 30635 26628
rect 9346 26140 9410 26144
rect 9346 26084 9350 26140
rect 9350 26084 9406 26140
rect 9406 26084 9410 26140
rect 9346 26080 9410 26084
rect 9426 26140 9490 26144
rect 9426 26084 9430 26140
rect 9430 26084 9486 26140
rect 9486 26084 9490 26140
rect 9426 26080 9490 26084
rect 9506 26140 9570 26144
rect 9506 26084 9510 26140
rect 9510 26084 9566 26140
rect 9566 26084 9570 26140
rect 9506 26080 9570 26084
rect 9586 26140 9650 26144
rect 9586 26084 9590 26140
rect 9590 26084 9646 26140
rect 9646 26084 9650 26140
rect 9586 26080 9650 26084
rect 17740 26140 17804 26144
rect 17740 26084 17744 26140
rect 17744 26084 17800 26140
rect 17800 26084 17804 26140
rect 17740 26080 17804 26084
rect 17820 26140 17884 26144
rect 17820 26084 17824 26140
rect 17824 26084 17880 26140
rect 17880 26084 17884 26140
rect 17820 26080 17884 26084
rect 17900 26140 17964 26144
rect 17900 26084 17904 26140
rect 17904 26084 17960 26140
rect 17960 26084 17964 26140
rect 17900 26080 17964 26084
rect 17980 26140 18044 26144
rect 17980 26084 17984 26140
rect 17984 26084 18040 26140
rect 18040 26084 18044 26140
rect 17980 26080 18044 26084
rect 26134 26140 26198 26144
rect 26134 26084 26138 26140
rect 26138 26084 26194 26140
rect 26194 26084 26198 26140
rect 26134 26080 26198 26084
rect 26214 26140 26278 26144
rect 26214 26084 26218 26140
rect 26218 26084 26274 26140
rect 26274 26084 26278 26140
rect 26214 26080 26278 26084
rect 26294 26140 26358 26144
rect 26294 26084 26298 26140
rect 26298 26084 26354 26140
rect 26354 26084 26358 26140
rect 26294 26080 26358 26084
rect 26374 26140 26438 26144
rect 26374 26084 26378 26140
rect 26378 26084 26434 26140
rect 26434 26084 26438 26140
rect 26374 26080 26438 26084
rect 34528 26140 34592 26144
rect 34528 26084 34532 26140
rect 34532 26084 34588 26140
rect 34588 26084 34592 26140
rect 34528 26080 34592 26084
rect 34608 26140 34672 26144
rect 34608 26084 34612 26140
rect 34612 26084 34668 26140
rect 34668 26084 34672 26140
rect 34608 26080 34672 26084
rect 34688 26140 34752 26144
rect 34688 26084 34692 26140
rect 34692 26084 34748 26140
rect 34748 26084 34752 26140
rect 34688 26080 34752 26084
rect 34768 26140 34832 26144
rect 34768 26084 34772 26140
rect 34772 26084 34828 26140
rect 34828 26084 34832 26140
rect 34768 26080 34832 26084
rect 5149 25596 5213 25600
rect 5149 25540 5153 25596
rect 5153 25540 5209 25596
rect 5209 25540 5213 25596
rect 5149 25536 5213 25540
rect 5229 25596 5293 25600
rect 5229 25540 5233 25596
rect 5233 25540 5289 25596
rect 5289 25540 5293 25596
rect 5229 25536 5293 25540
rect 5309 25596 5373 25600
rect 5309 25540 5313 25596
rect 5313 25540 5369 25596
rect 5369 25540 5373 25596
rect 5309 25536 5373 25540
rect 5389 25596 5453 25600
rect 5389 25540 5393 25596
rect 5393 25540 5449 25596
rect 5449 25540 5453 25596
rect 5389 25536 5453 25540
rect 13543 25596 13607 25600
rect 13543 25540 13547 25596
rect 13547 25540 13603 25596
rect 13603 25540 13607 25596
rect 13543 25536 13607 25540
rect 13623 25596 13687 25600
rect 13623 25540 13627 25596
rect 13627 25540 13683 25596
rect 13683 25540 13687 25596
rect 13623 25536 13687 25540
rect 13703 25596 13767 25600
rect 13703 25540 13707 25596
rect 13707 25540 13763 25596
rect 13763 25540 13767 25596
rect 13703 25536 13767 25540
rect 13783 25596 13847 25600
rect 13783 25540 13787 25596
rect 13787 25540 13843 25596
rect 13843 25540 13847 25596
rect 13783 25536 13847 25540
rect 21937 25596 22001 25600
rect 21937 25540 21941 25596
rect 21941 25540 21997 25596
rect 21997 25540 22001 25596
rect 21937 25536 22001 25540
rect 22017 25596 22081 25600
rect 22017 25540 22021 25596
rect 22021 25540 22077 25596
rect 22077 25540 22081 25596
rect 22017 25536 22081 25540
rect 22097 25596 22161 25600
rect 22097 25540 22101 25596
rect 22101 25540 22157 25596
rect 22157 25540 22161 25596
rect 22097 25536 22161 25540
rect 22177 25596 22241 25600
rect 22177 25540 22181 25596
rect 22181 25540 22237 25596
rect 22237 25540 22241 25596
rect 22177 25536 22241 25540
rect 30331 25596 30395 25600
rect 30331 25540 30335 25596
rect 30335 25540 30391 25596
rect 30391 25540 30395 25596
rect 30331 25536 30395 25540
rect 30411 25596 30475 25600
rect 30411 25540 30415 25596
rect 30415 25540 30471 25596
rect 30471 25540 30475 25596
rect 30411 25536 30475 25540
rect 30491 25596 30555 25600
rect 30491 25540 30495 25596
rect 30495 25540 30551 25596
rect 30551 25540 30555 25596
rect 30491 25536 30555 25540
rect 30571 25596 30635 25600
rect 30571 25540 30575 25596
rect 30575 25540 30631 25596
rect 30631 25540 30635 25596
rect 30571 25536 30635 25540
rect 9346 25052 9410 25056
rect 9346 24996 9350 25052
rect 9350 24996 9406 25052
rect 9406 24996 9410 25052
rect 9346 24992 9410 24996
rect 9426 25052 9490 25056
rect 9426 24996 9430 25052
rect 9430 24996 9486 25052
rect 9486 24996 9490 25052
rect 9426 24992 9490 24996
rect 9506 25052 9570 25056
rect 9506 24996 9510 25052
rect 9510 24996 9566 25052
rect 9566 24996 9570 25052
rect 9506 24992 9570 24996
rect 9586 25052 9650 25056
rect 9586 24996 9590 25052
rect 9590 24996 9646 25052
rect 9646 24996 9650 25052
rect 9586 24992 9650 24996
rect 17740 25052 17804 25056
rect 17740 24996 17744 25052
rect 17744 24996 17800 25052
rect 17800 24996 17804 25052
rect 17740 24992 17804 24996
rect 17820 25052 17884 25056
rect 17820 24996 17824 25052
rect 17824 24996 17880 25052
rect 17880 24996 17884 25052
rect 17820 24992 17884 24996
rect 17900 25052 17964 25056
rect 17900 24996 17904 25052
rect 17904 24996 17960 25052
rect 17960 24996 17964 25052
rect 17900 24992 17964 24996
rect 17980 25052 18044 25056
rect 17980 24996 17984 25052
rect 17984 24996 18040 25052
rect 18040 24996 18044 25052
rect 17980 24992 18044 24996
rect 26134 25052 26198 25056
rect 26134 24996 26138 25052
rect 26138 24996 26194 25052
rect 26194 24996 26198 25052
rect 26134 24992 26198 24996
rect 26214 25052 26278 25056
rect 26214 24996 26218 25052
rect 26218 24996 26274 25052
rect 26274 24996 26278 25052
rect 26214 24992 26278 24996
rect 26294 25052 26358 25056
rect 26294 24996 26298 25052
rect 26298 24996 26354 25052
rect 26354 24996 26358 25052
rect 26294 24992 26358 24996
rect 26374 25052 26438 25056
rect 26374 24996 26378 25052
rect 26378 24996 26434 25052
rect 26434 24996 26438 25052
rect 26374 24992 26438 24996
rect 34528 25052 34592 25056
rect 34528 24996 34532 25052
rect 34532 24996 34588 25052
rect 34588 24996 34592 25052
rect 34528 24992 34592 24996
rect 34608 25052 34672 25056
rect 34608 24996 34612 25052
rect 34612 24996 34668 25052
rect 34668 24996 34672 25052
rect 34608 24992 34672 24996
rect 34688 25052 34752 25056
rect 34688 24996 34692 25052
rect 34692 24996 34748 25052
rect 34748 24996 34752 25052
rect 34688 24992 34752 24996
rect 34768 25052 34832 25056
rect 34768 24996 34772 25052
rect 34772 24996 34828 25052
rect 34828 24996 34832 25052
rect 34768 24992 34832 24996
rect 5149 24508 5213 24512
rect 5149 24452 5153 24508
rect 5153 24452 5209 24508
rect 5209 24452 5213 24508
rect 5149 24448 5213 24452
rect 5229 24508 5293 24512
rect 5229 24452 5233 24508
rect 5233 24452 5289 24508
rect 5289 24452 5293 24508
rect 5229 24448 5293 24452
rect 5309 24508 5373 24512
rect 5309 24452 5313 24508
rect 5313 24452 5369 24508
rect 5369 24452 5373 24508
rect 5309 24448 5373 24452
rect 5389 24508 5453 24512
rect 5389 24452 5393 24508
rect 5393 24452 5449 24508
rect 5449 24452 5453 24508
rect 5389 24448 5453 24452
rect 13543 24508 13607 24512
rect 13543 24452 13547 24508
rect 13547 24452 13603 24508
rect 13603 24452 13607 24508
rect 13543 24448 13607 24452
rect 13623 24508 13687 24512
rect 13623 24452 13627 24508
rect 13627 24452 13683 24508
rect 13683 24452 13687 24508
rect 13623 24448 13687 24452
rect 13703 24508 13767 24512
rect 13703 24452 13707 24508
rect 13707 24452 13763 24508
rect 13763 24452 13767 24508
rect 13703 24448 13767 24452
rect 13783 24508 13847 24512
rect 13783 24452 13787 24508
rect 13787 24452 13843 24508
rect 13843 24452 13847 24508
rect 13783 24448 13847 24452
rect 21937 24508 22001 24512
rect 21937 24452 21941 24508
rect 21941 24452 21997 24508
rect 21997 24452 22001 24508
rect 21937 24448 22001 24452
rect 22017 24508 22081 24512
rect 22017 24452 22021 24508
rect 22021 24452 22077 24508
rect 22077 24452 22081 24508
rect 22017 24448 22081 24452
rect 22097 24508 22161 24512
rect 22097 24452 22101 24508
rect 22101 24452 22157 24508
rect 22157 24452 22161 24508
rect 22097 24448 22161 24452
rect 22177 24508 22241 24512
rect 22177 24452 22181 24508
rect 22181 24452 22237 24508
rect 22237 24452 22241 24508
rect 22177 24448 22241 24452
rect 30331 24508 30395 24512
rect 30331 24452 30335 24508
rect 30335 24452 30391 24508
rect 30391 24452 30395 24508
rect 30331 24448 30395 24452
rect 30411 24508 30475 24512
rect 30411 24452 30415 24508
rect 30415 24452 30471 24508
rect 30471 24452 30475 24508
rect 30411 24448 30475 24452
rect 30491 24508 30555 24512
rect 30491 24452 30495 24508
rect 30495 24452 30551 24508
rect 30551 24452 30555 24508
rect 30491 24448 30555 24452
rect 30571 24508 30635 24512
rect 30571 24452 30575 24508
rect 30575 24452 30631 24508
rect 30631 24452 30635 24508
rect 30571 24448 30635 24452
rect 9346 23964 9410 23968
rect 9346 23908 9350 23964
rect 9350 23908 9406 23964
rect 9406 23908 9410 23964
rect 9346 23904 9410 23908
rect 9426 23964 9490 23968
rect 9426 23908 9430 23964
rect 9430 23908 9486 23964
rect 9486 23908 9490 23964
rect 9426 23904 9490 23908
rect 9506 23964 9570 23968
rect 9506 23908 9510 23964
rect 9510 23908 9566 23964
rect 9566 23908 9570 23964
rect 9506 23904 9570 23908
rect 9586 23964 9650 23968
rect 9586 23908 9590 23964
rect 9590 23908 9646 23964
rect 9646 23908 9650 23964
rect 9586 23904 9650 23908
rect 17740 23964 17804 23968
rect 17740 23908 17744 23964
rect 17744 23908 17800 23964
rect 17800 23908 17804 23964
rect 17740 23904 17804 23908
rect 17820 23964 17884 23968
rect 17820 23908 17824 23964
rect 17824 23908 17880 23964
rect 17880 23908 17884 23964
rect 17820 23904 17884 23908
rect 17900 23964 17964 23968
rect 17900 23908 17904 23964
rect 17904 23908 17960 23964
rect 17960 23908 17964 23964
rect 17900 23904 17964 23908
rect 17980 23964 18044 23968
rect 17980 23908 17984 23964
rect 17984 23908 18040 23964
rect 18040 23908 18044 23964
rect 17980 23904 18044 23908
rect 26134 23964 26198 23968
rect 26134 23908 26138 23964
rect 26138 23908 26194 23964
rect 26194 23908 26198 23964
rect 26134 23904 26198 23908
rect 26214 23964 26278 23968
rect 26214 23908 26218 23964
rect 26218 23908 26274 23964
rect 26274 23908 26278 23964
rect 26214 23904 26278 23908
rect 26294 23964 26358 23968
rect 26294 23908 26298 23964
rect 26298 23908 26354 23964
rect 26354 23908 26358 23964
rect 26294 23904 26358 23908
rect 26374 23964 26438 23968
rect 26374 23908 26378 23964
rect 26378 23908 26434 23964
rect 26434 23908 26438 23964
rect 26374 23904 26438 23908
rect 34528 23964 34592 23968
rect 34528 23908 34532 23964
rect 34532 23908 34588 23964
rect 34588 23908 34592 23964
rect 34528 23904 34592 23908
rect 34608 23964 34672 23968
rect 34608 23908 34612 23964
rect 34612 23908 34668 23964
rect 34668 23908 34672 23964
rect 34608 23904 34672 23908
rect 34688 23964 34752 23968
rect 34688 23908 34692 23964
rect 34692 23908 34748 23964
rect 34748 23908 34752 23964
rect 34688 23904 34752 23908
rect 34768 23964 34832 23968
rect 34768 23908 34772 23964
rect 34772 23908 34828 23964
rect 34828 23908 34832 23964
rect 34768 23904 34832 23908
rect 5149 23420 5213 23424
rect 5149 23364 5153 23420
rect 5153 23364 5209 23420
rect 5209 23364 5213 23420
rect 5149 23360 5213 23364
rect 5229 23420 5293 23424
rect 5229 23364 5233 23420
rect 5233 23364 5289 23420
rect 5289 23364 5293 23420
rect 5229 23360 5293 23364
rect 5309 23420 5373 23424
rect 5309 23364 5313 23420
rect 5313 23364 5369 23420
rect 5369 23364 5373 23420
rect 5309 23360 5373 23364
rect 5389 23420 5453 23424
rect 5389 23364 5393 23420
rect 5393 23364 5449 23420
rect 5449 23364 5453 23420
rect 5389 23360 5453 23364
rect 13543 23420 13607 23424
rect 13543 23364 13547 23420
rect 13547 23364 13603 23420
rect 13603 23364 13607 23420
rect 13543 23360 13607 23364
rect 13623 23420 13687 23424
rect 13623 23364 13627 23420
rect 13627 23364 13683 23420
rect 13683 23364 13687 23420
rect 13623 23360 13687 23364
rect 13703 23420 13767 23424
rect 13703 23364 13707 23420
rect 13707 23364 13763 23420
rect 13763 23364 13767 23420
rect 13703 23360 13767 23364
rect 13783 23420 13847 23424
rect 13783 23364 13787 23420
rect 13787 23364 13843 23420
rect 13843 23364 13847 23420
rect 13783 23360 13847 23364
rect 21937 23420 22001 23424
rect 21937 23364 21941 23420
rect 21941 23364 21997 23420
rect 21997 23364 22001 23420
rect 21937 23360 22001 23364
rect 22017 23420 22081 23424
rect 22017 23364 22021 23420
rect 22021 23364 22077 23420
rect 22077 23364 22081 23420
rect 22017 23360 22081 23364
rect 22097 23420 22161 23424
rect 22097 23364 22101 23420
rect 22101 23364 22157 23420
rect 22157 23364 22161 23420
rect 22097 23360 22161 23364
rect 22177 23420 22241 23424
rect 22177 23364 22181 23420
rect 22181 23364 22237 23420
rect 22237 23364 22241 23420
rect 22177 23360 22241 23364
rect 30331 23420 30395 23424
rect 30331 23364 30335 23420
rect 30335 23364 30391 23420
rect 30391 23364 30395 23420
rect 30331 23360 30395 23364
rect 30411 23420 30475 23424
rect 30411 23364 30415 23420
rect 30415 23364 30471 23420
rect 30471 23364 30475 23420
rect 30411 23360 30475 23364
rect 30491 23420 30555 23424
rect 30491 23364 30495 23420
rect 30495 23364 30551 23420
rect 30551 23364 30555 23420
rect 30491 23360 30555 23364
rect 30571 23420 30635 23424
rect 30571 23364 30575 23420
rect 30575 23364 30631 23420
rect 30631 23364 30635 23420
rect 30571 23360 30635 23364
rect 9346 22876 9410 22880
rect 9346 22820 9350 22876
rect 9350 22820 9406 22876
rect 9406 22820 9410 22876
rect 9346 22816 9410 22820
rect 9426 22876 9490 22880
rect 9426 22820 9430 22876
rect 9430 22820 9486 22876
rect 9486 22820 9490 22876
rect 9426 22816 9490 22820
rect 9506 22876 9570 22880
rect 9506 22820 9510 22876
rect 9510 22820 9566 22876
rect 9566 22820 9570 22876
rect 9506 22816 9570 22820
rect 9586 22876 9650 22880
rect 9586 22820 9590 22876
rect 9590 22820 9646 22876
rect 9646 22820 9650 22876
rect 9586 22816 9650 22820
rect 17740 22876 17804 22880
rect 17740 22820 17744 22876
rect 17744 22820 17800 22876
rect 17800 22820 17804 22876
rect 17740 22816 17804 22820
rect 17820 22876 17884 22880
rect 17820 22820 17824 22876
rect 17824 22820 17880 22876
rect 17880 22820 17884 22876
rect 17820 22816 17884 22820
rect 17900 22876 17964 22880
rect 17900 22820 17904 22876
rect 17904 22820 17960 22876
rect 17960 22820 17964 22876
rect 17900 22816 17964 22820
rect 17980 22876 18044 22880
rect 17980 22820 17984 22876
rect 17984 22820 18040 22876
rect 18040 22820 18044 22876
rect 17980 22816 18044 22820
rect 26134 22876 26198 22880
rect 26134 22820 26138 22876
rect 26138 22820 26194 22876
rect 26194 22820 26198 22876
rect 26134 22816 26198 22820
rect 26214 22876 26278 22880
rect 26214 22820 26218 22876
rect 26218 22820 26274 22876
rect 26274 22820 26278 22876
rect 26214 22816 26278 22820
rect 26294 22876 26358 22880
rect 26294 22820 26298 22876
rect 26298 22820 26354 22876
rect 26354 22820 26358 22876
rect 26294 22816 26358 22820
rect 26374 22876 26438 22880
rect 26374 22820 26378 22876
rect 26378 22820 26434 22876
rect 26434 22820 26438 22876
rect 26374 22816 26438 22820
rect 34528 22876 34592 22880
rect 34528 22820 34532 22876
rect 34532 22820 34588 22876
rect 34588 22820 34592 22876
rect 34528 22816 34592 22820
rect 34608 22876 34672 22880
rect 34608 22820 34612 22876
rect 34612 22820 34668 22876
rect 34668 22820 34672 22876
rect 34608 22816 34672 22820
rect 34688 22876 34752 22880
rect 34688 22820 34692 22876
rect 34692 22820 34748 22876
rect 34748 22820 34752 22876
rect 34688 22816 34752 22820
rect 34768 22876 34832 22880
rect 34768 22820 34772 22876
rect 34772 22820 34828 22876
rect 34828 22820 34832 22876
rect 34768 22816 34832 22820
rect 5149 22332 5213 22336
rect 5149 22276 5153 22332
rect 5153 22276 5209 22332
rect 5209 22276 5213 22332
rect 5149 22272 5213 22276
rect 5229 22332 5293 22336
rect 5229 22276 5233 22332
rect 5233 22276 5289 22332
rect 5289 22276 5293 22332
rect 5229 22272 5293 22276
rect 5309 22332 5373 22336
rect 5309 22276 5313 22332
rect 5313 22276 5369 22332
rect 5369 22276 5373 22332
rect 5309 22272 5373 22276
rect 5389 22332 5453 22336
rect 5389 22276 5393 22332
rect 5393 22276 5449 22332
rect 5449 22276 5453 22332
rect 5389 22272 5453 22276
rect 13543 22332 13607 22336
rect 13543 22276 13547 22332
rect 13547 22276 13603 22332
rect 13603 22276 13607 22332
rect 13543 22272 13607 22276
rect 13623 22332 13687 22336
rect 13623 22276 13627 22332
rect 13627 22276 13683 22332
rect 13683 22276 13687 22332
rect 13623 22272 13687 22276
rect 13703 22332 13767 22336
rect 13703 22276 13707 22332
rect 13707 22276 13763 22332
rect 13763 22276 13767 22332
rect 13703 22272 13767 22276
rect 13783 22332 13847 22336
rect 13783 22276 13787 22332
rect 13787 22276 13843 22332
rect 13843 22276 13847 22332
rect 13783 22272 13847 22276
rect 21937 22332 22001 22336
rect 21937 22276 21941 22332
rect 21941 22276 21997 22332
rect 21997 22276 22001 22332
rect 21937 22272 22001 22276
rect 22017 22332 22081 22336
rect 22017 22276 22021 22332
rect 22021 22276 22077 22332
rect 22077 22276 22081 22332
rect 22017 22272 22081 22276
rect 22097 22332 22161 22336
rect 22097 22276 22101 22332
rect 22101 22276 22157 22332
rect 22157 22276 22161 22332
rect 22097 22272 22161 22276
rect 22177 22332 22241 22336
rect 22177 22276 22181 22332
rect 22181 22276 22237 22332
rect 22237 22276 22241 22332
rect 22177 22272 22241 22276
rect 30331 22332 30395 22336
rect 30331 22276 30335 22332
rect 30335 22276 30391 22332
rect 30391 22276 30395 22332
rect 30331 22272 30395 22276
rect 30411 22332 30475 22336
rect 30411 22276 30415 22332
rect 30415 22276 30471 22332
rect 30471 22276 30475 22332
rect 30411 22272 30475 22276
rect 30491 22332 30555 22336
rect 30491 22276 30495 22332
rect 30495 22276 30551 22332
rect 30551 22276 30555 22332
rect 30491 22272 30555 22276
rect 30571 22332 30635 22336
rect 30571 22276 30575 22332
rect 30575 22276 30631 22332
rect 30631 22276 30635 22332
rect 30571 22272 30635 22276
rect 9346 21788 9410 21792
rect 9346 21732 9350 21788
rect 9350 21732 9406 21788
rect 9406 21732 9410 21788
rect 9346 21728 9410 21732
rect 9426 21788 9490 21792
rect 9426 21732 9430 21788
rect 9430 21732 9486 21788
rect 9486 21732 9490 21788
rect 9426 21728 9490 21732
rect 9506 21788 9570 21792
rect 9506 21732 9510 21788
rect 9510 21732 9566 21788
rect 9566 21732 9570 21788
rect 9506 21728 9570 21732
rect 9586 21788 9650 21792
rect 9586 21732 9590 21788
rect 9590 21732 9646 21788
rect 9646 21732 9650 21788
rect 9586 21728 9650 21732
rect 17740 21788 17804 21792
rect 17740 21732 17744 21788
rect 17744 21732 17800 21788
rect 17800 21732 17804 21788
rect 17740 21728 17804 21732
rect 17820 21788 17884 21792
rect 17820 21732 17824 21788
rect 17824 21732 17880 21788
rect 17880 21732 17884 21788
rect 17820 21728 17884 21732
rect 17900 21788 17964 21792
rect 17900 21732 17904 21788
rect 17904 21732 17960 21788
rect 17960 21732 17964 21788
rect 17900 21728 17964 21732
rect 17980 21788 18044 21792
rect 17980 21732 17984 21788
rect 17984 21732 18040 21788
rect 18040 21732 18044 21788
rect 17980 21728 18044 21732
rect 26134 21788 26198 21792
rect 26134 21732 26138 21788
rect 26138 21732 26194 21788
rect 26194 21732 26198 21788
rect 26134 21728 26198 21732
rect 26214 21788 26278 21792
rect 26214 21732 26218 21788
rect 26218 21732 26274 21788
rect 26274 21732 26278 21788
rect 26214 21728 26278 21732
rect 26294 21788 26358 21792
rect 26294 21732 26298 21788
rect 26298 21732 26354 21788
rect 26354 21732 26358 21788
rect 26294 21728 26358 21732
rect 26374 21788 26438 21792
rect 26374 21732 26378 21788
rect 26378 21732 26434 21788
rect 26434 21732 26438 21788
rect 26374 21728 26438 21732
rect 34528 21788 34592 21792
rect 34528 21732 34532 21788
rect 34532 21732 34588 21788
rect 34588 21732 34592 21788
rect 34528 21728 34592 21732
rect 34608 21788 34672 21792
rect 34608 21732 34612 21788
rect 34612 21732 34668 21788
rect 34668 21732 34672 21788
rect 34608 21728 34672 21732
rect 34688 21788 34752 21792
rect 34688 21732 34692 21788
rect 34692 21732 34748 21788
rect 34748 21732 34752 21788
rect 34688 21728 34752 21732
rect 34768 21788 34832 21792
rect 34768 21732 34772 21788
rect 34772 21732 34828 21788
rect 34828 21732 34832 21788
rect 34768 21728 34832 21732
rect 5149 21244 5213 21248
rect 5149 21188 5153 21244
rect 5153 21188 5209 21244
rect 5209 21188 5213 21244
rect 5149 21184 5213 21188
rect 5229 21244 5293 21248
rect 5229 21188 5233 21244
rect 5233 21188 5289 21244
rect 5289 21188 5293 21244
rect 5229 21184 5293 21188
rect 5309 21244 5373 21248
rect 5309 21188 5313 21244
rect 5313 21188 5369 21244
rect 5369 21188 5373 21244
rect 5309 21184 5373 21188
rect 5389 21244 5453 21248
rect 5389 21188 5393 21244
rect 5393 21188 5449 21244
rect 5449 21188 5453 21244
rect 5389 21184 5453 21188
rect 13543 21244 13607 21248
rect 13543 21188 13547 21244
rect 13547 21188 13603 21244
rect 13603 21188 13607 21244
rect 13543 21184 13607 21188
rect 13623 21244 13687 21248
rect 13623 21188 13627 21244
rect 13627 21188 13683 21244
rect 13683 21188 13687 21244
rect 13623 21184 13687 21188
rect 13703 21244 13767 21248
rect 13703 21188 13707 21244
rect 13707 21188 13763 21244
rect 13763 21188 13767 21244
rect 13703 21184 13767 21188
rect 13783 21244 13847 21248
rect 13783 21188 13787 21244
rect 13787 21188 13843 21244
rect 13843 21188 13847 21244
rect 13783 21184 13847 21188
rect 21937 21244 22001 21248
rect 21937 21188 21941 21244
rect 21941 21188 21997 21244
rect 21997 21188 22001 21244
rect 21937 21184 22001 21188
rect 22017 21244 22081 21248
rect 22017 21188 22021 21244
rect 22021 21188 22077 21244
rect 22077 21188 22081 21244
rect 22017 21184 22081 21188
rect 22097 21244 22161 21248
rect 22097 21188 22101 21244
rect 22101 21188 22157 21244
rect 22157 21188 22161 21244
rect 22097 21184 22161 21188
rect 22177 21244 22241 21248
rect 22177 21188 22181 21244
rect 22181 21188 22237 21244
rect 22237 21188 22241 21244
rect 22177 21184 22241 21188
rect 30331 21244 30395 21248
rect 30331 21188 30335 21244
rect 30335 21188 30391 21244
rect 30391 21188 30395 21244
rect 30331 21184 30395 21188
rect 30411 21244 30475 21248
rect 30411 21188 30415 21244
rect 30415 21188 30471 21244
rect 30471 21188 30475 21244
rect 30411 21184 30475 21188
rect 30491 21244 30555 21248
rect 30491 21188 30495 21244
rect 30495 21188 30551 21244
rect 30551 21188 30555 21244
rect 30491 21184 30555 21188
rect 30571 21244 30635 21248
rect 30571 21188 30575 21244
rect 30575 21188 30631 21244
rect 30631 21188 30635 21244
rect 30571 21184 30635 21188
rect 9346 20700 9410 20704
rect 9346 20644 9350 20700
rect 9350 20644 9406 20700
rect 9406 20644 9410 20700
rect 9346 20640 9410 20644
rect 9426 20700 9490 20704
rect 9426 20644 9430 20700
rect 9430 20644 9486 20700
rect 9486 20644 9490 20700
rect 9426 20640 9490 20644
rect 9506 20700 9570 20704
rect 9506 20644 9510 20700
rect 9510 20644 9566 20700
rect 9566 20644 9570 20700
rect 9506 20640 9570 20644
rect 9586 20700 9650 20704
rect 9586 20644 9590 20700
rect 9590 20644 9646 20700
rect 9646 20644 9650 20700
rect 9586 20640 9650 20644
rect 17740 20700 17804 20704
rect 17740 20644 17744 20700
rect 17744 20644 17800 20700
rect 17800 20644 17804 20700
rect 17740 20640 17804 20644
rect 17820 20700 17884 20704
rect 17820 20644 17824 20700
rect 17824 20644 17880 20700
rect 17880 20644 17884 20700
rect 17820 20640 17884 20644
rect 17900 20700 17964 20704
rect 17900 20644 17904 20700
rect 17904 20644 17960 20700
rect 17960 20644 17964 20700
rect 17900 20640 17964 20644
rect 17980 20700 18044 20704
rect 17980 20644 17984 20700
rect 17984 20644 18040 20700
rect 18040 20644 18044 20700
rect 17980 20640 18044 20644
rect 26134 20700 26198 20704
rect 26134 20644 26138 20700
rect 26138 20644 26194 20700
rect 26194 20644 26198 20700
rect 26134 20640 26198 20644
rect 26214 20700 26278 20704
rect 26214 20644 26218 20700
rect 26218 20644 26274 20700
rect 26274 20644 26278 20700
rect 26214 20640 26278 20644
rect 26294 20700 26358 20704
rect 26294 20644 26298 20700
rect 26298 20644 26354 20700
rect 26354 20644 26358 20700
rect 26294 20640 26358 20644
rect 26374 20700 26438 20704
rect 26374 20644 26378 20700
rect 26378 20644 26434 20700
rect 26434 20644 26438 20700
rect 26374 20640 26438 20644
rect 34528 20700 34592 20704
rect 34528 20644 34532 20700
rect 34532 20644 34588 20700
rect 34588 20644 34592 20700
rect 34528 20640 34592 20644
rect 34608 20700 34672 20704
rect 34608 20644 34612 20700
rect 34612 20644 34668 20700
rect 34668 20644 34672 20700
rect 34608 20640 34672 20644
rect 34688 20700 34752 20704
rect 34688 20644 34692 20700
rect 34692 20644 34748 20700
rect 34748 20644 34752 20700
rect 34688 20640 34752 20644
rect 34768 20700 34832 20704
rect 34768 20644 34772 20700
rect 34772 20644 34828 20700
rect 34828 20644 34832 20700
rect 34768 20640 34832 20644
rect 5149 20156 5213 20160
rect 5149 20100 5153 20156
rect 5153 20100 5209 20156
rect 5209 20100 5213 20156
rect 5149 20096 5213 20100
rect 5229 20156 5293 20160
rect 5229 20100 5233 20156
rect 5233 20100 5289 20156
rect 5289 20100 5293 20156
rect 5229 20096 5293 20100
rect 5309 20156 5373 20160
rect 5309 20100 5313 20156
rect 5313 20100 5369 20156
rect 5369 20100 5373 20156
rect 5309 20096 5373 20100
rect 5389 20156 5453 20160
rect 5389 20100 5393 20156
rect 5393 20100 5449 20156
rect 5449 20100 5453 20156
rect 5389 20096 5453 20100
rect 13543 20156 13607 20160
rect 13543 20100 13547 20156
rect 13547 20100 13603 20156
rect 13603 20100 13607 20156
rect 13543 20096 13607 20100
rect 13623 20156 13687 20160
rect 13623 20100 13627 20156
rect 13627 20100 13683 20156
rect 13683 20100 13687 20156
rect 13623 20096 13687 20100
rect 13703 20156 13767 20160
rect 13703 20100 13707 20156
rect 13707 20100 13763 20156
rect 13763 20100 13767 20156
rect 13703 20096 13767 20100
rect 13783 20156 13847 20160
rect 13783 20100 13787 20156
rect 13787 20100 13843 20156
rect 13843 20100 13847 20156
rect 13783 20096 13847 20100
rect 21937 20156 22001 20160
rect 21937 20100 21941 20156
rect 21941 20100 21997 20156
rect 21997 20100 22001 20156
rect 21937 20096 22001 20100
rect 22017 20156 22081 20160
rect 22017 20100 22021 20156
rect 22021 20100 22077 20156
rect 22077 20100 22081 20156
rect 22017 20096 22081 20100
rect 22097 20156 22161 20160
rect 22097 20100 22101 20156
rect 22101 20100 22157 20156
rect 22157 20100 22161 20156
rect 22097 20096 22161 20100
rect 22177 20156 22241 20160
rect 22177 20100 22181 20156
rect 22181 20100 22237 20156
rect 22237 20100 22241 20156
rect 22177 20096 22241 20100
rect 30331 20156 30395 20160
rect 30331 20100 30335 20156
rect 30335 20100 30391 20156
rect 30391 20100 30395 20156
rect 30331 20096 30395 20100
rect 30411 20156 30475 20160
rect 30411 20100 30415 20156
rect 30415 20100 30471 20156
rect 30471 20100 30475 20156
rect 30411 20096 30475 20100
rect 30491 20156 30555 20160
rect 30491 20100 30495 20156
rect 30495 20100 30551 20156
rect 30551 20100 30555 20156
rect 30491 20096 30555 20100
rect 30571 20156 30635 20160
rect 30571 20100 30575 20156
rect 30575 20100 30631 20156
rect 30631 20100 30635 20156
rect 30571 20096 30635 20100
rect 9346 19612 9410 19616
rect 9346 19556 9350 19612
rect 9350 19556 9406 19612
rect 9406 19556 9410 19612
rect 9346 19552 9410 19556
rect 9426 19612 9490 19616
rect 9426 19556 9430 19612
rect 9430 19556 9486 19612
rect 9486 19556 9490 19612
rect 9426 19552 9490 19556
rect 9506 19612 9570 19616
rect 9506 19556 9510 19612
rect 9510 19556 9566 19612
rect 9566 19556 9570 19612
rect 9506 19552 9570 19556
rect 9586 19612 9650 19616
rect 9586 19556 9590 19612
rect 9590 19556 9646 19612
rect 9646 19556 9650 19612
rect 9586 19552 9650 19556
rect 17740 19612 17804 19616
rect 17740 19556 17744 19612
rect 17744 19556 17800 19612
rect 17800 19556 17804 19612
rect 17740 19552 17804 19556
rect 17820 19612 17884 19616
rect 17820 19556 17824 19612
rect 17824 19556 17880 19612
rect 17880 19556 17884 19612
rect 17820 19552 17884 19556
rect 17900 19612 17964 19616
rect 17900 19556 17904 19612
rect 17904 19556 17960 19612
rect 17960 19556 17964 19612
rect 17900 19552 17964 19556
rect 17980 19612 18044 19616
rect 17980 19556 17984 19612
rect 17984 19556 18040 19612
rect 18040 19556 18044 19612
rect 17980 19552 18044 19556
rect 26134 19612 26198 19616
rect 26134 19556 26138 19612
rect 26138 19556 26194 19612
rect 26194 19556 26198 19612
rect 26134 19552 26198 19556
rect 26214 19612 26278 19616
rect 26214 19556 26218 19612
rect 26218 19556 26274 19612
rect 26274 19556 26278 19612
rect 26214 19552 26278 19556
rect 26294 19612 26358 19616
rect 26294 19556 26298 19612
rect 26298 19556 26354 19612
rect 26354 19556 26358 19612
rect 26294 19552 26358 19556
rect 26374 19612 26438 19616
rect 26374 19556 26378 19612
rect 26378 19556 26434 19612
rect 26434 19556 26438 19612
rect 26374 19552 26438 19556
rect 34528 19612 34592 19616
rect 34528 19556 34532 19612
rect 34532 19556 34588 19612
rect 34588 19556 34592 19612
rect 34528 19552 34592 19556
rect 34608 19612 34672 19616
rect 34608 19556 34612 19612
rect 34612 19556 34668 19612
rect 34668 19556 34672 19612
rect 34608 19552 34672 19556
rect 34688 19612 34752 19616
rect 34688 19556 34692 19612
rect 34692 19556 34748 19612
rect 34748 19556 34752 19612
rect 34688 19552 34752 19556
rect 34768 19612 34832 19616
rect 34768 19556 34772 19612
rect 34772 19556 34828 19612
rect 34828 19556 34832 19612
rect 34768 19552 34832 19556
rect 5149 19068 5213 19072
rect 5149 19012 5153 19068
rect 5153 19012 5209 19068
rect 5209 19012 5213 19068
rect 5149 19008 5213 19012
rect 5229 19068 5293 19072
rect 5229 19012 5233 19068
rect 5233 19012 5289 19068
rect 5289 19012 5293 19068
rect 5229 19008 5293 19012
rect 5309 19068 5373 19072
rect 5309 19012 5313 19068
rect 5313 19012 5369 19068
rect 5369 19012 5373 19068
rect 5309 19008 5373 19012
rect 5389 19068 5453 19072
rect 5389 19012 5393 19068
rect 5393 19012 5449 19068
rect 5449 19012 5453 19068
rect 5389 19008 5453 19012
rect 13543 19068 13607 19072
rect 13543 19012 13547 19068
rect 13547 19012 13603 19068
rect 13603 19012 13607 19068
rect 13543 19008 13607 19012
rect 13623 19068 13687 19072
rect 13623 19012 13627 19068
rect 13627 19012 13683 19068
rect 13683 19012 13687 19068
rect 13623 19008 13687 19012
rect 13703 19068 13767 19072
rect 13703 19012 13707 19068
rect 13707 19012 13763 19068
rect 13763 19012 13767 19068
rect 13703 19008 13767 19012
rect 13783 19068 13847 19072
rect 13783 19012 13787 19068
rect 13787 19012 13843 19068
rect 13843 19012 13847 19068
rect 13783 19008 13847 19012
rect 21937 19068 22001 19072
rect 21937 19012 21941 19068
rect 21941 19012 21997 19068
rect 21997 19012 22001 19068
rect 21937 19008 22001 19012
rect 22017 19068 22081 19072
rect 22017 19012 22021 19068
rect 22021 19012 22077 19068
rect 22077 19012 22081 19068
rect 22017 19008 22081 19012
rect 22097 19068 22161 19072
rect 22097 19012 22101 19068
rect 22101 19012 22157 19068
rect 22157 19012 22161 19068
rect 22097 19008 22161 19012
rect 22177 19068 22241 19072
rect 22177 19012 22181 19068
rect 22181 19012 22237 19068
rect 22237 19012 22241 19068
rect 22177 19008 22241 19012
rect 30331 19068 30395 19072
rect 30331 19012 30335 19068
rect 30335 19012 30391 19068
rect 30391 19012 30395 19068
rect 30331 19008 30395 19012
rect 30411 19068 30475 19072
rect 30411 19012 30415 19068
rect 30415 19012 30471 19068
rect 30471 19012 30475 19068
rect 30411 19008 30475 19012
rect 30491 19068 30555 19072
rect 30491 19012 30495 19068
rect 30495 19012 30551 19068
rect 30551 19012 30555 19068
rect 30491 19008 30555 19012
rect 30571 19068 30635 19072
rect 30571 19012 30575 19068
rect 30575 19012 30631 19068
rect 30631 19012 30635 19068
rect 30571 19008 30635 19012
rect 9346 18524 9410 18528
rect 9346 18468 9350 18524
rect 9350 18468 9406 18524
rect 9406 18468 9410 18524
rect 9346 18464 9410 18468
rect 9426 18524 9490 18528
rect 9426 18468 9430 18524
rect 9430 18468 9486 18524
rect 9486 18468 9490 18524
rect 9426 18464 9490 18468
rect 9506 18524 9570 18528
rect 9506 18468 9510 18524
rect 9510 18468 9566 18524
rect 9566 18468 9570 18524
rect 9506 18464 9570 18468
rect 9586 18524 9650 18528
rect 9586 18468 9590 18524
rect 9590 18468 9646 18524
rect 9646 18468 9650 18524
rect 9586 18464 9650 18468
rect 17740 18524 17804 18528
rect 17740 18468 17744 18524
rect 17744 18468 17800 18524
rect 17800 18468 17804 18524
rect 17740 18464 17804 18468
rect 17820 18524 17884 18528
rect 17820 18468 17824 18524
rect 17824 18468 17880 18524
rect 17880 18468 17884 18524
rect 17820 18464 17884 18468
rect 17900 18524 17964 18528
rect 17900 18468 17904 18524
rect 17904 18468 17960 18524
rect 17960 18468 17964 18524
rect 17900 18464 17964 18468
rect 17980 18524 18044 18528
rect 17980 18468 17984 18524
rect 17984 18468 18040 18524
rect 18040 18468 18044 18524
rect 17980 18464 18044 18468
rect 26134 18524 26198 18528
rect 26134 18468 26138 18524
rect 26138 18468 26194 18524
rect 26194 18468 26198 18524
rect 26134 18464 26198 18468
rect 26214 18524 26278 18528
rect 26214 18468 26218 18524
rect 26218 18468 26274 18524
rect 26274 18468 26278 18524
rect 26214 18464 26278 18468
rect 26294 18524 26358 18528
rect 26294 18468 26298 18524
rect 26298 18468 26354 18524
rect 26354 18468 26358 18524
rect 26294 18464 26358 18468
rect 26374 18524 26438 18528
rect 26374 18468 26378 18524
rect 26378 18468 26434 18524
rect 26434 18468 26438 18524
rect 26374 18464 26438 18468
rect 34528 18524 34592 18528
rect 34528 18468 34532 18524
rect 34532 18468 34588 18524
rect 34588 18468 34592 18524
rect 34528 18464 34592 18468
rect 34608 18524 34672 18528
rect 34608 18468 34612 18524
rect 34612 18468 34668 18524
rect 34668 18468 34672 18524
rect 34608 18464 34672 18468
rect 34688 18524 34752 18528
rect 34688 18468 34692 18524
rect 34692 18468 34748 18524
rect 34748 18468 34752 18524
rect 34688 18464 34752 18468
rect 34768 18524 34832 18528
rect 34768 18468 34772 18524
rect 34772 18468 34828 18524
rect 34828 18468 34832 18524
rect 34768 18464 34832 18468
rect 5149 17980 5213 17984
rect 5149 17924 5153 17980
rect 5153 17924 5209 17980
rect 5209 17924 5213 17980
rect 5149 17920 5213 17924
rect 5229 17980 5293 17984
rect 5229 17924 5233 17980
rect 5233 17924 5289 17980
rect 5289 17924 5293 17980
rect 5229 17920 5293 17924
rect 5309 17980 5373 17984
rect 5309 17924 5313 17980
rect 5313 17924 5369 17980
rect 5369 17924 5373 17980
rect 5309 17920 5373 17924
rect 5389 17980 5453 17984
rect 5389 17924 5393 17980
rect 5393 17924 5449 17980
rect 5449 17924 5453 17980
rect 5389 17920 5453 17924
rect 13543 17980 13607 17984
rect 13543 17924 13547 17980
rect 13547 17924 13603 17980
rect 13603 17924 13607 17980
rect 13543 17920 13607 17924
rect 13623 17980 13687 17984
rect 13623 17924 13627 17980
rect 13627 17924 13683 17980
rect 13683 17924 13687 17980
rect 13623 17920 13687 17924
rect 13703 17980 13767 17984
rect 13703 17924 13707 17980
rect 13707 17924 13763 17980
rect 13763 17924 13767 17980
rect 13703 17920 13767 17924
rect 13783 17980 13847 17984
rect 13783 17924 13787 17980
rect 13787 17924 13843 17980
rect 13843 17924 13847 17980
rect 13783 17920 13847 17924
rect 21937 17980 22001 17984
rect 21937 17924 21941 17980
rect 21941 17924 21997 17980
rect 21997 17924 22001 17980
rect 21937 17920 22001 17924
rect 22017 17980 22081 17984
rect 22017 17924 22021 17980
rect 22021 17924 22077 17980
rect 22077 17924 22081 17980
rect 22017 17920 22081 17924
rect 22097 17980 22161 17984
rect 22097 17924 22101 17980
rect 22101 17924 22157 17980
rect 22157 17924 22161 17980
rect 22097 17920 22161 17924
rect 22177 17980 22241 17984
rect 22177 17924 22181 17980
rect 22181 17924 22237 17980
rect 22237 17924 22241 17980
rect 22177 17920 22241 17924
rect 30331 17980 30395 17984
rect 30331 17924 30335 17980
rect 30335 17924 30391 17980
rect 30391 17924 30395 17980
rect 30331 17920 30395 17924
rect 30411 17980 30475 17984
rect 30411 17924 30415 17980
rect 30415 17924 30471 17980
rect 30471 17924 30475 17980
rect 30411 17920 30475 17924
rect 30491 17980 30555 17984
rect 30491 17924 30495 17980
rect 30495 17924 30551 17980
rect 30551 17924 30555 17980
rect 30491 17920 30555 17924
rect 30571 17980 30635 17984
rect 30571 17924 30575 17980
rect 30575 17924 30631 17980
rect 30631 17924 30635 17980
rect 30571 17920 30635 17924
rect 9076 17716 9140 17780
rect 9346 17436 9410 17440
rect 9346 17380 9350 17436
rect 9350 17380 9406 17436
rect 9406 17380 9410 17436
rect 9346 17376 9410 17380
rect 9426 17436 9490 17440
rect 9426 17380 9430 17436
rect 9430 17380 9486 17436
rect 9486 17380 9490 17436
rect 9426 17376 9490 17380
rect 9506 17436 9570 17440
rect 9506 17380 9510 17436
rect 9510 17380 9566 17436
rect 9566 17380 9570 17436
rect 9506 17376 9570 17380
rect 9586 17436 9650 17440
rect 9586 17380 9590 17436
rect 9590 17380 9646 17436
rect 9646 17380 9650 17436
rect 9586 17376 9650 17380
rect 17740 17436 17804 17440
rect 17740 17380 17744 17436
rect 17744 17380 17800 17436
rect 17800 17380 17804 17436
rect 17740 17376 17804 17380
rect 17820 17436 17884 17440
rect 17820 17380 17824 17436
rect 17824 17380 17880 17436
rect 17880 17380 17884 17436
rect 17820 17376 17884 17380
rect 17900 17436 17964 17440
rect 17900 17380 17904 17436
rect 17904 17380 17960 17436
rect 17960 17380 17964 17436
rect 17900 17376 17964 17380
rect 17980 17436 18044 17440
rect 17980 17380 17984 17436
rect 17984 17380 18040 17436
rect 18040 17380 18044 17436
rect 17980 17376 18044 17380
rect 26134 17436 26198 17440
rect 26134 17380 26138 17436
rect 26138 17380 26194 17436
rect 26194 17380 26198 17436
rect 26134 17376 26198 17380
rect 26214 17436 26278 17440
rect 26214 17380 26218 17436
rect 26218 17380 26274 17436
rect 26274 17380 26278 17436
rect 26214 17376 26278 17380
rect 26294 17436 26358 17440
rect 26294 17380 26298 17436
rect 26298 17380 26354 17436
rect 26354 17380 26358 17436
rect 26294 17376 26358 17380
rect 26374 17436 26438 17440
rect 26374 17380 26378 17436
rect 26378 17380 26434 17436
rect 26434 17380 26438 17436
rect 26374 17376 26438 17380
rect 34528 17436 34592 17440
rect 34528 17380 34532 17436
rect 34532 17380 34588 17436
rect 34588 17380 34592 17436
rect 34528 17376 34592 17380
rect 34608 17436 34672 17440
rect 34608 17380 34612 17436
rect 34612 17380 34668 17436
rect 34668 17380 34672 17436
rect 34608 17376 34672 17380
rect 34688 17436 34752 17440
rect 34688 17380 34692 17436
rect 34692 17380 34748 17436
rect 34748 17380 34752 17436
rect 34688 17376 34752 17380
rect 34768 17436 34832 17440
rect 34768 17380 34772 17436
rect 34772 17380 34828 17436
rect 34828 17380 34832 17436
rect 34768 17376 34832 17380
rect 5149 16892 5213 16896
rect 5149 16836 5153 16892
rect 5153 16836 5209 16892
rect 5209 16836 5213 16892
rect 5149 16832 5213 16836
rect 5229 16892 5293 16896
rect 5229 16836 5233 16892
rect 5233 16836 5289 16892
rect 5289 16836 5293 16892
rect 5229 16832 5293 16836
rect 5309 16892 5373 16896
rect 5309 16836 5313 16892
rect 5313 16836 5369 16892
rect 5369 16836 5373 16892
rect 5309 16832 5373 16836
rect 5389 16892 5453 16896
rect 5389 16836 5393 16892
rect 5393 16836 5449 16892
rect 5449 16836 5453 16892
rect 5389 16832 5453 16836
rect 13543 16892 13607 16896
rect 13543 16836 13547 16892
rect 13547 16836 13603 16892
rect 13603 16836 13607 16892
rect 13543 16832 13607 16836
rect 13623 16892 13687 16896
rect 13623 16836 13627 16892
rect 13627 16836 13683 16892
rect 13683 16836 13687 16892
rect 13623 16832 13687 16836
rect 13703 16892 13767 16896
rect 13703 16836 13707 16892
rect 13707 16836 13763 16892
rect 13763 16836 13767 16892
rect 13703 16832 13767 16836
rect 13783 16892 13847 16896
rect 13783 16836 13787 16892
rect 13787 16836 13843 16892
rect 13843 16836 13847 16892
rect 13783 16832 13847 16836
rect 21937 16892 22001 16896
rect 21937 16836 21941 16892
rect 21941 16836 21997 16892
rect 21997 16836 22001 16892
rect 21937 16832 22001 16836
rect 22017 16892 22081 16896
rect 22017 16836 22021 16892
rect 22021 16836 22077 16892
rect 22077 16836 22081 16892
rect 22017 16832 22081 16836
rect 22097 16892 22161 16896
rect 22097 16836 22101 16892
rect 22101 16836 22157 16892
rect 22157 16836 22161 16892
rect 22097 16832 22161 16836
rect 22177 16892 22241 16896
rect 22177 16836 22181 16892
rect 22181 16836 22237 16892
rect 22237 16836 22241 16892
rect 22177 16832 22241 16836
rect 30331 16892 30395 16896
rect 30331 16836 30335 16892
rect 30335 16836 30391 16892
rect 30391 16836 30395 16892
rect 30331 16832 30395 16836
rect 30411 16892 30475 16896
rect 30411 16836 30415 16892
rect 30415 16836 30471 16892
rect 30471 16836 30475 16892
rect 30411 16832 30475 16836
rect 30491 16892 30555 16896
rect 30491 16836 30495 16892
rect 30495 16836 30551 16892
rect 30551 16836 30555 16892
rect 30491 16832 30555 16836
rect 30571 16892 30635 16896
rect 30571 16836 30575 16892
rect 30575 16836 30631 16892
rect 30631 16836 30635 16892
rect 30571 16832 30635 16836
rect 8340 16416 8404 16420
rect 8340 16360 8354 16416
rect 8354 16360 8404 16416
rect 8340 16356 8404 16360
rect 8524 16356 8588 16420
rect 9346 16348 9410 16352
rect 9346 16292 9350 16348
rect 9350 16292 9406 16348
rect 9406 16292 9410 16348
rect 9346 16288 9410 16292
rect 9426 16348 9490 16352
rect 9426 16292 9430 16348
rect 9430 16292 9486 16348
rect 9486 16292 9490 16348
rect 9426 16288 9490 16292
rect 9506 16348 9570 16352
rect 9506 16292 9510 16348
rect 9510 16292 9566 16348
rect 9566 16292 9570 16348
rect 9506 16288 9570 16292
rect 9586 16348 9650 16352
rect 9586 16292 9590 16348
rect 9590 16292 9646 16348
rect 9646 16292 9650 16348
rect 9586 16288 9650 16292
rect 17740 16348 17804 16352
rect 17740 16292 17744 16348
rect 17744 16292 17800 16348
rect 17800 16292 17804 16348
rect 17740 16288 17804 16292
rect 17820 16348 17884 16352
rect 17820 16292 17824 16348
rect 17824 16292 17880 16348
rect 17880 16292 17884 16348
rect 17820 16288 17884 16292
rect 17900 16348 17964 16352
rect 17900 16292 17904 16348
rect 17904 16292 17960 16348
rect 17960 16292 17964 16348
rect 17900 16288 17964 16292
rect 17980 16348 18044 16352
rect 17980 16292 17984 16348
rect 17984 16292 18040 16348
rect 18040 16292 18044 16348
rect 17980 16288 18044 16292
rect 26134 16348 26198 16352
rect 26134 16292 26138 16348
rect 26138 16292 26194 16348
rect 26194 16292 26198 16348
rect 26134 16288 26198 16292
rect 26214 16348 26278 16352
rect 26214 16292 26218 16348
rect 26218 16292 26274 16348
rect 26274 16292 26278 16348
rect 26214 16288 26278 16292
rect 26294 16348 26358 16352
rect 26294 16292 26298 16348
rect 26298 16292 26354 16348
rect 26354 16292 26358 16348
rect 26294 16288 26358 16292
rect 26374 16348 26438 16352
rect 26374 16292 26378 16348
rect 26378 16292 26434 16348
rect 26434 16292 26438 16348
rect 26374 16288 26438 16292
rect 34528 16348 34592 16352
rect 34528 16292 34532 16348
rect 34532 16292 34588 16348
rect 34588 16292 34592 16348
rect 34528 16288 34592 16292
rect 34608 16348 34672 16352
rect 34608 16292 34612 16348
rect 34612 16292 34668 16348
rect 34668 16292 34672 16348
rect 34608 16288 34672 16292
rect 34688 16348 34752 16352
rect 34688 16292 34692 16348
rect 34692 16292 34748 16348
rect 34748 16292 34752 16348
rect 34688 16288 34752 16292
rect 34768 16348 34832 16352
rect 34768 16292 34772 16348
rect 34772 16292 34828 16348
rect 34828 16292 34832 16348
rect 34768 16288 34832 16292
rect 9076 15948 9140 16012
rect 5149 15804 5213 15808
rect 5149 15748 5153 15804
rect 5153 15748 5209 15804
rect 5209 15748 5213 15804
rect 5149 15744 5213 15748
rect 5229 15804 5293 15808
rect 5229 15748 5233 15804
rect 5233 15748 5289 15804
rect 5289 15748 5293 15804
rect 5229 15744 5293 15748
rect 5309 15804 5373 15808
rect 5309 15748 5313 15804
rect 5313 15748 5369 15804
rect 5369 15748 5373 15804
rect 5309 15744 5373 15748
rect 5389 15804 5453 15808
rect 5389 15748 5393 15804
rect 5393 15748 5449 15804
rect 5449 15748 5453 15804
rect 5389 15744 5453 15748
rect 13543 15804 13607 15808
rect 13543 15748 13547 15804
rect 13547 15748 13603 15804
rect 13603 15748 13607 15804
rect 13543 15744 13607 15748
rect 13623 15804 13687 15808
rect 13623 15748 13627 15804
rect 13627 15748 13683 15804
rect 13683 15748 13687 15804
rect 13623 15744 13687 15748
rect 13703 15804 13767 15808
rect 13703 15748 13707 15804
rect 13707 15748 13763 15804
rect 13763 15748 13767 15804
rect 13703 15744 13767 15748
rect 13783 15804 13847 15808
rect 13783 15748 13787 15804
rect 13787 15748 13843 15804
rect 13843 15748 13847 15804
rect 13783 15744 13847 15748
rect 21937 15804 22001 15808
rect 21937 15748 21941 15804
rect 21941 15748 21997 15804
rect 21997 15748 22001 15804
rect 21937 15744 22001 15748
rect 22017 15804 22081 15808
rect 22017 15748 22021 15804
rect 22021 15748 22077 15804
rect 22077 15748 22081 15804
rect 22017 15744 22081 15748
rect 22097 15804 22161 15808
rect 22097 15748 22101 15804
rect 22101 15748 22157 15804
rect 22157 15748 22161 15804
rect 22097 15744 22161 15748
rect 22177 15804 22241 15808
rect 22177 15748 22181 15804
rect 22181 15748 22237 15804
rect 22237 15748 22241 15804
rect 22177 15744 22241 15748
rect 30331 15804 30395 15808
rect 30331 15748 30335 15804
rect 30335 15748 30391 15804
rect 30391 15748 30395 15804
rect 30331 15744 30395 15748
rect 30411 15804 30475 15808
rect 30411 15748 30415 15804
rect 30415 15748 30471 15804
rect 30471 15748 30475 15804
rect 30411 15744 30475 15748
rect 30491 15804 30555 15808
rect 30491 15748 30495 15804
rect 30495 15748 30551 15804
rect 30551 15748 30555 15804
rect 30491 15744 30555 15748
rect 30571 15804 30635 15808
rect 30571 15748 30575 15804
rect 30575 15748 30631 15804
rect 30631 15748 30635 15804
rect 30571 15744 30635 15748
rect 9346 15260 9410 15264
rect 9346 15204 9350 15260
rect 9350 15204 9406 15260
rect 9406 15204 9410 15260
rect 9346 15200 9410 15204
rect 9426 15260 9490 15264
rect 9426 15204 9430 15260
rect 9430 15204 9486 15260
rect 9486 15204 9490 15260
rect 9426 15200 9490 15204
rect 9506 15260 9570 15264
rect 9506 15204 9510 15260
rect 9510 15204 9566 15260
rect 9566 15204 9570 15260
rect 9506 15200 9570 15204
rect 9586 15260 9650 15264
rect 9586 15204 9590 15260
rect 9590 15204 9646 15260
rect 9646 15204 9650 15260
rect 9586 15200 9650 15204
rect 17740 15260 17804 15264
rect 17740 15204 17744 15260
rect 17744 15204 17800 15260
rect 17800 15204 17804 15260
rect 17740 15200 17804 15204
rect 17820 15260 17884 15264
rect 17820 15204 17824 15260
rect 17824 15204 17880 15260
rect 17880 15204 17884 15260
rect 17820 15200 17884 15204
rect 17900 15260 17964 15264
rect 17900 15204 17904 15260
rect 17904 15204 17960 15260
rect 17960 15204 17964 15260
rect 17900 15200 17964 15204
rect 17980 15260 18044 15264
rect 17980 15204 17984 15260
rect 17984 15204 18040 15260
rect 18040 15204 18044 15260
rect 17980 15200 18044 15204
rect 26134 15260 26198 15264
rect 26134 15204 26138 15260
rect 26138 15204 26194 15260
rect 26194 15204 26198 15260
rect 26134 15200 26198 15204
rect 26214 15260 26278 15264
rect 26214 15204 26218 15260
rect 26218 15204 26274 15260
rect 26274 15204 26278 15260
rect 26214 15200 26278 15204
rect 26294 15260 26358 15264
rect 26294 15204 26298 15260
rect 26298 15204 26354 15260
rect 26354 15204 26358 15260
rect 26294 15200 26358 15204
rect 26374 15260 26438 15264
rect 26374 15204 26378 15260
rect 26378 15204 26434 15260
rect 26434 15204 26438 15260
rect 26374 15200 26438 15204
rect 34528 15260 34592 15264
rect 34528 15204 34532 15260
rect 34532 15204 34588 15260
rect 34588 15204 34592 15260
rect 34528 15200 34592 15204
rect 34608 15260 34672 15264
rect 34608 15204 34612 15260
rect 34612 15204 34668 15260
rect 34668 15204 34672 15260
rect 34608 15200 34672 15204
rect 34688 15260 34752 15264
rect 34688 15204 34692 15260
rect 34692 15204 34748 15260
rect 34748 15204 34752 15260
rect 34688 15200 34752 15204
rect 34768 15260 34832 15264
rect 34768 15204 34772 15260
rect 34772 15204 34828 15260
rect 34828 15204 34832 15260
rect 34768 15200 34832 15204
rect 8524 14784 8588 14788
rect 8524 14728 8574 14784
rect 8574 14728 8588 14784
rect 8524 14724 8588 14728
rect 5149 14716 5213 14720
rect 5149 14660 5153 14716
rect 5153 14660 5209 14716
rect 5209 14660 5213 14716
rect 5149 14656 5213 14660
rect 5229 14716 5293 14720
rect 5229 14660 5233 14716
rect 5233 14660 5289 14716
rect 5289 14660 5293 14716
rect 5229 14656 5293 14660
rect 5309 14716 5373 14720
rect 5309 14660 5313 14716
rect 5313 14660 5369 14716
rect 5369 14660 5373 14716
rect 5309 14656 5373 14660
rect 5389 14716 5453 14720
rect 5389 14660 5393 14716
rect 5393 14660 5449 14716
rect 5449 14660 5453 14716
rect 5389 14656 5453 14660
rect 13543 14716 13607 14720
rect 13543 14660 13547 14716
rect 13547 14660 13603 14716
rect 13603 14660 13607 14716
rect 13543 14656 13607 14660
rect 13623 14716 13687 14720
rect 13623 14660 13627 14716
rect 13627 14660 13683 14716
rect 13683 14660 13687 14716
rect 13623 14656 13687 14660
rect 13703 14716 13767 14720
rect 13703 14660 13707 14716
rect 13707 14660 13763 14716
rect 13763 14660 13767 14716
rect 13703 14656 13767 14660
rect 13783 14716 13847 14720
rect 13783 14660 13787 14716
rect 13787 14660 13843 14716
rect 13843 14660 13847 14716
rect 13783 14656 13847 14660
rect 21937 14716 22001 14720
rect 21937 14660 21941 14716
rect 21941 14660 21997 14716
rect 21997 14660 22001 14716
rect 21937 14656 22001 14660
rect 22017 14716 22081 14720
rect 22017 14660 22021 14716
rect 22021 14660 22077 14716
rect 22077 14660 22081 14716
rect 22017 14656 22081 14660
rect 22097 14716 22161 14720
rect 22097 14660 22101 14716
rect 22101 14660 22157 14716
rect 22157 14660 22161 14716
rect 22097 14656 22161 14660
rect 22177 14716 22241 14720
rect 22177 14660 22181 14716
rect 22181 14660 22237 14716
rect 22237 14660 22241 14716
rect 22177 14656 22241 14660
rect 30331 14716 30395 14720
rect 30331 14660 30335 14716
rect 30335 14660 30391 14716
rect 30391 14660 30395 14716
rect 30331 14656 30395 14660
rect 30411 14716 30475 14720
rect 30411 14660 30415 14716
rect 30415 14660 30471 14716
rect 30471 14660 30475 14716
rect 30411 14656 30475 14660
rect 30491 14716 30555 14720
rect 30491 14660 30495 14716
rect 30495 14660 30551 14716
rect 30551 14660 30555 14716
rect 30491 14656 30555 14660
rect 30571 14716 30635 14720
rect 30571 14660 30575 14716
rect 30575 14660 30631 14716
rect 30631 14660 30635 14716
rect 30571 14656 30635 14660
rect 9346 14172 9410 14176
rect 9346 14116 9350 14172
rect 9350 14116 9406 14172
rect 9406 14116 9410 14172
rect 9346 14112 9410 14116
rect 9426 14172 9490 14176
rect 9426 14116 9430 14172
rect 9430 14116 9486 14172
rect 9486 14116 9490 14172
rect 9426 14112 9490 14116
rect 9506 14172 9570 14176
rect 9506 14116 9510 14172
rect 9510 14116 9566 14172
rect 9566 14116 9570 14172
rect 9506 14112 9570 14116
rect 9586 14172 9650 14176
rect 9586 14116 9590 14172
rect 9590 14116 9646 14172
rect 9646 14116 9650 14172
rect 9586 14112 9650 14116
rect 17740 14172 17804 14176
rect 17740 14116 17744 14172
rect 17744 14116 17800 14172
rect 17800 14116 17804 14172
rect 17740 14112 17804 14116
rect 17820 14172 17884 14176
rect 17820 14116 17824 14172
rect 17824 14116 17880 14172
rect 17880 14116 17884 14172
rect 17820 14112 17884 14116
rect 17900 14172 17964 14176
rect 17900 14116 17904 14172
rect 17904 14116 17960 14172
rect 17960 14116 17964 14172
rect 17900 14112 17964 14116
rect 17980 14172 18044 14176
rect 17980 14116 17984 14172
rect 17984 14116 18040 14172
rect 18040 14116 18044 14172
rect 17980 14112 18044 14116
rect 26134 14172 26198 14176
rect 26134 14116 26138 14172
rect 26138 14116 26194 14172
rect 26194 14116 26198 14172
rect 26134 14112 26198 14116
rect 26214 14172 26278 14176
rect 26214 14116 26218 14172
rect 26218 14116 26274 14172
rect 26274 14116 26278 14172
rect 26214 14112 26278 14116
rect 26294 14172 26358 14176
rect 26294 14116 26298 14172
rect 26298 14116 26354 14172
rect 26354 14116 26358 14172
rect 26294 14112 26358 14116
rect 26374 14172 26438 14176
rect 26374 14116 26378 14172
rect 26378 14116 26434 14172
rect 26434 14116 26438 14172
rect 26374 14112 26438 14116
rect 34528 14172 34592 14176
rect 34528 14116 34532 14172
rect 34532 14116 34588 14172
rect 34588 14116 34592 14172
rect 34528 14112 34592 14116
rect 34608 14172 34672 14176
rect 34608 14116 34612 14172
rect 34612 14116 34668 14172
rect 34668 14116 34672 14172
rect 34608 14112 34672 14116
rect 34688 14172 34752 14176
rect 34688 14116 34692 14172
rect 34692 14116 34748 14172
rect 34748 14116 34752 14172
rect 34688 14112 34752 14116
rect 34768 14172 34832 14176
rect 34768 14116 34772 14172
rect 34772 14116 34828 14172
rect 34828 14116 34832 14172
rect 34768 14112 34832 14116
rect 5149 13628 5213 13632
rect 5149 13572 5153 13628
rect 5153 13572 5209 13628
rect 5209 13572 5213 13628
rect 5149 13568 5213 13572
rect 5229 13628 5293 13632
rect 5229 13572 5233 13628
rect 5233 13572 5289 13628
rect 5289 13572 5293 13628
rect 5229 13568 5293 13572
rect 5309 13628 5373 13632
rect 5309 13572 5313 13628
rect 5313 13572 5369 13628
rect 5369 13572 5373 13628
rect 5309 13568 5373 13572
rect 5389 13628 5453 13632
rect 5389 13572 5393 13628
rect 5393 13572 5449 13628
rect 5449 13572 5453 13628
rect 5389 13568 5453 13572
rect 13543 13628 13607 13632
rect 13543 13572 13547 13628
rect 13547 13572 13603 13628
rect 13603 13572 13607 13628
rect 13543 13568 13607 13572
rect 13623 13628 13687 13632
rect 13623 13572 13627 13628
rect 13627 13572 13683 13628
rect 13683 13572 13687 13628
rect 13623 13568 13687 13572
rect 13703 13628 13767 13632
rect 13703 13572 13707 13628
rect 13707 13572 13763 13628
rect 13763 13572 13767 13628
rect 13703 13568 13767 13572
rect 13783 13628 13847 13632
rect 13783 13572 13787 13628
rect 13787 13572 13843 13628
rect 13843 13572 13847 13628
rect 13783 13568 13847 13572
rect 21937 13628 22001 13632
rect 21937 13572 21941 13628
rect 21941 13572 21997 13628
rect 21997 13572 22001 13628
rect 21937 13568 22001 13572
rect 22017 13628 22081 13632
rect 22017 13572 22021 13628
rect 22021 13572 22077 13628
rect 22077 13572 22081 13628
rect 22017 13568 22081 13572
rect 22097 13628 22161 13632
rect 22097 13572 22101 13628
rect 22101 13572 22157 13628
rect 22157 13572 22161 13628
rect 22097 13568 22161 13572
rect 22177 13628 22241 13632
rect 22177 13572 22181 13628
rect 22181 13572 22237 13628
rect 22237 13572 22241 13628
rect 22177 13568 22241 13572
rect 30331 13628 30395 13632
rect 30331 13572 30335 13628
rect 30335 13572 30391 13628
rect 30391 13572 30395 13628
rect 30331 13568 30395 13572
rect 30411 13628 30475 13632
rect 30411 13572 30415 13628
rect 30415 13572 30471 13628
rect 30471 13572 30475 13628
rect 30411 13568 30475 13572
rect 30491 13628 30555 13632
rect 30491 13572 30495 13628
rect 30495 13572 30551 13628
rect 30551 13572 30555 13628
rect 30491 13568 30555 13572
rect 30571 13628 30635 13632
rect 30571 13572 30575 13628
rect 30575 13572 30631 13628
rect 30631 13572 30635 13628
rect 30571 13568 30635 13572
rect 8340 13424 8404 13428
rect 8340 13368 8354 13424
rect 8354 13368 8404 13424
rect 8340 13364 8404 13368
rect 9346 13084 9410 13088
rect 9346 13028 9350 13084
rect 9350 13028 9406 13084
rect 9406 13028 9410 13084
rect 9346 13024 9410 13028
rect 9426 13084 9490 13088
rect 9426 13028 9430 13084
rect 9430 13028 9486 13084
rect 9486 13028 9490 13084
rect 9426 13024 9490 13028
rect 9506 13084 9570 13088
rect 9506 13028 9510 13084
rect 9510 13028 9566 13084
rect 9566 13028 9570 13084
rect 9506 13024 9570 13028
rect 9586 13084 9650 13088
rect 9586 13028 9590 13084
rect 9590 13028 9646 13084
rect 9646 13028 9650 13084
rect 9586 13024 9650 13028
rect 17740 13084 17804 13088
rect 17740 13028 17744 13084
rect 17744 13028 17800 13084
rect 17800 13028 17804 13084
rect 17740 13024 17804 13028
rect 17820 13084 17884 13088
rect 17820 13028 17824 13084
rect 17824 13028 17880 13084
rect 17880 13028 17884 13084
rect 17820 13024 17884 13028
rect 17900 13084 17964 13088
rect 17900 13028 17904 13084
rect 17904 13028 17960 13084
rect 17960 13028 17964 13084
rect 17900 13024 17964 13028
rect 17980 13084 18044 13088
rect 17980 13028 17984 13084
rect 17984 13028 18040 13084
rect 18040 13028 18044 13084
rect 17980 13024 18044 13028
rect 26134 13084 26198 13088
rect 26134 13028 26138 13084
rect 26138 13028 26194 13084
rect 26194 13028 26198 13084
rect 26134 13024 26198 13028
rect 26214 13084 26278 13088
rect 26214 13028 26218 13084
rect 26218 13028 26274 13084
rect 26274 13028 26278 13084
rect 26214 13024 26278 13028
rect 26294 13084 26358 13088
rect 26294 13028 26298 13084
rect 26298 13028 26354 13084
rect 26354 13028 26358 13084
rect 26294 13024 26358 13028
rect 26374 13084 26438 13088
rect 26374 13028 26378 13084
rect 26378 13028 26434 13084
rect 26434 13028 26438 13084
rect 26374 13024 26438 13028
rect 34528 13084 34592 13088
rect 34528 13028 34532 13084
rect 34532 13028 34588 13084
rect 34588 13028 34592 13084
rect 34528 13024 34592 13028
rect 34608 13084 34672 13088
rect 34608 13028 34612 13084
rect 34612 13028 34668 13084
rect 34668 13028 34672 13084
rect 34608 13024 34672 13028
rect 34688 13084 34752 13088
rect 34688 13028 34692 13084
rect 34692 13028 34748 13084
rect 34748 13028 34752 13084
rect 34688 13024 34752 13028
rect 34768 13084 34832 13088
rect 34768 13028 34772 13084
rect 34772 13028 34828 13084
rect 34828 13028 34832 13084
rect 34768 13024 34832 13028
rect 5149 12540 5213 12544
rect 5149 12484 5153 12540
rect 5153 12484 5209 12540
rect 5209 12484 5213 12540
rect 5149 12480 5213 12484
rect 5229 12540 5293 12544
rect 5229 12484 5233 12540
rect 5233 12484 5289 12540
rect 5289 12484 5293 12540
rect 5229 12480 5293 12484
rect 5309 12540 5373 12544
rect 5309 12484 5313 12540
rect 5313 12484 5369 12540
rect 5369 12484 5373 12540
rect 5309 12480 5373 12484
rect 5389 12540 5453 12544
rect 5389 12484 5393 12540
rect 5393 12484 5449 12540
rect 5449 12484 5453 12540
rect 5389 12480 5453 12484
rect 13543 12540 13607 12544
rect 13543 12484 13547 12540
rect 13547 12484 13603 12540
rect 13603 12484 13607 12540
rect 13543 12480 13607 12484
rect 13623 12540 13687 12544
rect 13623 12484 13627 12540
rect 13627 12484 13683 12540
rect 13683 12484 13687 12540
rect 13623 12480 13687 12484
rect 13703 12540 13767 12544
rect 13703 12484 13707 12540
rect 13707 12484 13763 12540
rect 13763 12484 13767 12540
rect 13703 12480 13767 12484
rect 13783 12540 13847 12544
rect 13783 12484 13787 12540
rect 13787 12484 13843 12540
rect 13843 12484 13847 12540
rect 13783 12480 13847 12484
rect 21937 12540 22001 12544
rect 21937 12484 21941 12540
rect 21941 12484 21997 12540
rect 21997 12484 22001 12540
rect 21937 12480 22001 12484
rect 22017 12540 22081 12544
rect 22017 12484 22021 12540
rect 22021 12484 22077 12540
rect 22077 12484 22081 12540
rect 22017 12480 22081 12484
rect 22097 12540 22161 12544
rect 22097 12484 22101 12540
rect 22101 12484 22157 12540
rect 22157 12484 22161 12540
rect 22097 12480 22161 12484
rect 22177 12540 22241 12544
rect 22177 12484 22181 12540
rect 22181 12484 22237 12540
rect 22237 12484 22241 12540
rect 22177 12480 22241 12484
rect 30331 12540 30395 12544
rect 30331 12484 30335 12540
rect 30335 12484 30391 12540
rect 30391 12484 30395 12540
rect 30331 12480 30395 12484
rect 30411 12540 30475 12544
rect 30411 12484 30415 12540
rect 30415 12484 30471 12540
rect 30471 12484 30475 12540
rect 30411 12480 30475 12484
rect 30491 12540 30555 12544
rect 30491 12484 30495 12540
rect 30495 12484 30551 12540
rect 30551 12484 30555 12540
rect 30491 12480 30555 12484
rect 30571 12540 30635 12544
rect 30571 12484 30575 12540
rect 30575 12484 30631 12540
rect 30631 12484 30635 12540
rect 30571 12480 30635 12484
rect 9346 11996 9410 12000
rect 9346 11940 9350 11996
rect 9350 11940 9406 11996
rect 9406 11940 9410 11996
rect 9346 11936 9410 11940
rect 9426 11996 9490 12000
rect 9426 11940 9430 11996
rect 9430 11940 9486 11996
rect 9486 11940 9490 11996
rect 9426 11936 9490 11940
rect 9506 11996 9570 12000
rect 9506 11940 9510 11996
rect 9510 11940 9566 11996
rect 9566 11940 9570 11996
rect 9506 11936 9570 11940
rect 9586 11996 9650 12000
rect 9586 11940 9590 11996
rect 9590 11940 9646 11996
rect 9646 11940 9650 11996
rect 9586 11936 9650 11940
rect 17740 11996 17804 12000
rect 17740 11940 17744 11996
rect 17744 11940 17800 11996
rect 17800 11940 17804 11996
rect 17740 11936 17804 11940
rect 17820 11996 17884 12000
rect 17820 11940 17824 11996
rect 17824 11940 17880 11996
rect 17880 11940 17884 11996
rect 17820 11936 17884 11940
rect 17900 11996 17964 12000
rect 17900 11940 17904 11996
rect 17904 11940 17960 11996
rect 17960 11940 17964 11996
rect 17900 11936 17964 11940
rect 17980 11996 18044 12000
rect 17980 11940 17984 11996
rect 17984 11940 18040 11996
rect 18040 11940 18044 11996
rect 17980 11936 18044 11940
rect 26134 11996 26198 12000
rect 26134 11940 26138 11996
rect 26138 11940 26194 11996
rect 26194 11940 26198 11996
rect 26134 11936 26198 11940
rect 26214 11996 26278 12000
rect 26214 11940 26218 11996
rect 26218 11940 26274 11996
rect 26274 11940 26278 11996
rect 26214 11936 26278 11940
rect 26294 11996 26358 12000
rect 26294 11940 26298 11996
rect 26298 11940 26354 11996
rect 26354 11940 26358 11996
rect 26294 11936 26358 11940
rect 26374 11996 26438 12000
rect 26374 11940 26378 11996
rect 26378 11940 26434 11996
rect 26434 11940 26438 11996
rect 26374 11936 26438 11940
rect 34528 11996 34592 12000
rect 34528 11940 34532 11996
rect 34532 11940 34588 11996
rect 34588 11940 34592 11996
rect 34528 11936 34592 11940
rect 34608 11996 34672 12000
rect 34608 11940 34612 11996
rect 34612 11940 34668 11996
rect 34668 11940 34672 11996
rect 34608 11936 34672 11940
rect 34688 11996 34752 12000
rect 34688 11940 34692 11996
rect 34692 11940 34748 11996
rect 34748 11940 34752 11996
rect 34688 11936 34752 11940
rect 34768 11996 34832 12000
rect 34768 11940 34772 11996
rect 34772 11940 34828 11996
rect 34828 11940 34832 11996
rect 34768 11936 34832 11940
rect 5149 11452 5213 11456
rect 5149 11396 5153 11452
rect 5153 11396 5209 11452
rect 5209 11396 5213 11452
rect 5149 11392 5213 11396
rect 5229 11452 5293 11456
rect 5229 11396 5233 11452
rect 5233 11396 5289 11452
rect 5289 11396 5293 11452
rect 5229 11392 5293 11396
rect 5309 11452 5373 11456
rect 5309 11396 5313 11452
rect 5313 11396 5369 11452
rect 5369 11396 5373 11452
rect 5309 11392 5373 11396
rect 5389 11452 5453 11456
rect 5389 11396 5393 11452
rect 5393 11396 5449 11452
rect 5449 11396 5453 11452
rect 5389 11392 5453 11396
rect 13543 11452 13607 11456
rect 13543 11396 13547 11452
rect 13547 11396 13603 11452
rect 13603 11396 13607 11452
rect 13543 11392 13607 11396
rect 13623 11452 13687 11456
rect 13623 11396 13627 11452
rect 13627 11396 13683 11452
rect 13683 11396 13687 11452
rect 13623 11392 13687 11396
rect 13703 11452 13767 11456
rect 13703 11396 13707 11452
rect 13707 11396 13763 11452
rect 13763 11396 13767 11452
rect 13703 11392 13767 11396
rect 13783 11452 13847 11456
rect 13783 11396 13787 11452
rect 13787 11396 13843 11452
rect 13843 11396 13847 11452
rect 13783 11392 13847 11396
rect 21937 11452 22001 11456
rect 21937 11396 21941 11452
rect 21941 11396 21997 11452
rect 21997 11396 22001 11452
rect 21937 11392 22001 11396
rect 22017 11452 22081 11456
rect 22017 11396 22021 11452
rect 22021 11396 22077 11452
rect 22077 11396 22081 11452
rect 22017 11392 22081 11396
rect 22097 11452 22161 11456
rect 22097 11396 22101 11452
rect 22101 11396 22157 11452
rect 22157 11396 22161 11452
rect 22097 11392 22161 11396
rect 22177 11452 22241 11456
rect 22177 11396 22181 11452
rect 22181 11396 22237 11452
rect 22237 11396 22241 11452
rect 22177 11392 22241 11396
rect 30331 11452 30395 11456
rect 30331 11396 30335 11452
rect 30335 11396 30391 11452
rect 30391 11396 30395 11452
rect 30331 11392 30395 11396
rect 30411 11452 30475 11456
rect 30411 11396 30415 11452
rect 30415 11396 30471 11452
rect 30471 11396 30475 11452
rect 30411 11392 30475 11396
rect 30491 11452 30555 11456
rect 30491 11396 30495 11452
rect 30495 11396 30551 11452
rect 30551 11396 30555 11452
rect 30491 11392 30555 11396
rect 30571 11452 30635 11456
rect 30571 11396 30575 11452
rect 30575 11396 30631 11452
rect 30631 11396 30635 11452
rect 30571 11392 30635 11396
rect 9346 10908 9410 10912
rect 9346 10852 9350 10908
rect 9350 10852 9406 10908
rect 9406 10852 9410 10908
rect 9346 10848 9410 10852
rect 9426 10908 9490 10912
rect 9426 10852 9430 10908
rect 9430 10852 9486 10908
rect 9486 10852 9490 10908
rect 9426 10848 9490 10852
rect 9506 10908 9570 10912
rect 9506 10852 9510 10908
rect 9510 10852 9566 10908
rect 9566 10852 9570 10908
rect 9506 10848 9570 10852
rect 9586 10908 9650 10912
rect 9586 10852 9590 10908
rect 9590 10852 9646 10908
rect 9646 10852 9650 10908
rect 9586 10848 9650 10852
rect 17740 10908 17804 10912
rect 17740 10852 17744 10908
rect 17744 10852 17800 10908
rect 17800 10852 17804 10908
rect 17740 10848 17804 10852
rect 17820 10908 17884 10912
rect 17820 10852 17824 10908
rect 17824 10852 17880 10908
rect 17880 10852 17884 10908
rect 17820 10848 17884 10852
rect 17900 10908 17964 10912
rect 17900 10852 17904 10908
rect 17904 10852 17960 10908
rect 17960 10852 17964 10908
rect 17900 10848 17964 10852
rect 17980 10908 18044 10912
rect 17980 10852 17984 10908
rect 17984 10852 18040 10908
rect 18040 10852 18044 10908
rect 17980 10848 18044 10852
rect 26134 10908 26198 10912
rect 26134 10852 26138 10908
rect 26138 10852 26194 10908
rect 26194 10852 26198 10908
rect 26134 10848 26198 10852
rect 26214 10908 26278 10912
rect 26214 10852 26218 10908
rect 26218 10852 26274 10908
rect 26274 10852 26278 10908
rect 26214 10848 26278 10852
rect 26294 10908 26358 10912
rect 26294 10852 26298 10908
rect 26298 10852 26354 10908
rect 26354 10852 26358 10908
rect 26294 10848 26358 10852
rect 26374 10908 26438 10912
rect 26374 10852 26378 10908
rect 26378 10852 26434 10908
rect 26434 10852 26438 10908
rect 26374 10848 26438 10852
rect 34528 10908 34592 10912
rect 34528 10852 34532 10908
rect 34532 10852 34588 10908
rect 34588 10852 34592 10908
rect 34528 10848 34592 10852
rect 34608 10908 34672 10912
rect 34608 10852 34612 10908
rect 34612 10852 34668 10908
rect 34668 10852 34672 10908
rect 34608 10848 34672 10852
rect 34688 10908 34752 10912
rect 34688 10852 34692 10908
rect 34692 10852 34748 10908
rect 34748 10852 34752 10908
rect 34688 10848 34752 10852
rect 34768 10908 34832 10912
rect 34768 10852 34772 10908
rect 34772 10852 34828 10908
rect 34828 10852 34832 10908
rect 34768 10848 34832 10852
rect 5149 10364 5213 10368
rect 5149 10308 5153 10364
rect 5153 10308 5209 10364
rect 5209 10308 5213 10364
rect 5149 10304 5213 10308
rect 5229 10364 5293 10368
rect 5229 10308 5233 10364
rect 5233 10308 5289 10364
rect 5289 10308 5293 10364
rect 5229 10304 5293 10308
rect 5309 10364 5373 10368
rect 5309 10308 5313 10364
rect 5313 10308 5369 10364
rect 5369 10308 5373 10364
rect 5309 10304 5373 10308
rect 5389 10364 5453 10368
rect 5389 10308 5393 10364
rect 5393 10308 5449 10364
rect 5449 10308 5453 10364
rect 5389 10304 5453 10308
rect 13543 10364 13607 10368
rect 13543 10308 13547 10364
rect 13547 10308 13603 10364
rect 13603 10308 13607 10364
rect 13543 10304 13607 10308
rect 13623 10364 13687 10368
rect 13623 10308 13627 10364
rect 13627 10308 13683 10364
rect 13683 10308 13687 10364
rect 13623 10304 13687 10308
rect 13703 10364 13767 10368
rect 13703 10308 13707 10364
rect 13707 10308 13763 10364
rect 13763 10308 13767 10364
rect 13703 10304 13767 10308
rect 13783 10364 13847 10368
rect 13783 10308 13787 10364
rect 13787 10308 13843 10364
rect 13843 10308 13847 10364
rect 13783 10304 13847 10308
rect 21937 10364 22001 10368
rect 21937 10308 21941 10364
rect 21941 10308 21997 10364
rect 21997 10308 22001 10364
rect 21937 10304 22001 10308
rect 22017 10364 22081 10368
rect 22017 10308 22021 10364
rect 22021 10308 22077 10364
rect 22077 10308 22081 10364
rect 22017 10304 22081 10308
rect 22097 10364 22161 10368
rect 22097 10308 22101 10364
rect 22101 10308 22157 10364
rect 22157 10308 22161 10364
rect 22097 10304 22161 10308
rect 22177 10364 22241 10368
rect 22177 10308 22181 10364
rect 22181 10308 22237 10364
rect 22237 10308 22241 10364
rect 22177 10304 22241 10308
rect 30331 10364 30395 10368
rect 30331 10308 30335 10364
rect 30335 10308 30391 10364
rect 30391 10308 30395 10364
rect 30331 10304 30395 10308
rect 30411 10364 30475 10368
rect 30411 10308 30415 10364
rect 30415 10308 30471 10364
rect 30471 10308 30475 10364
rect 30411 10304 30475 10308
rect 30491 10364 30555 10368
rect 30491 10308 30495 10364
rect 30495 10308 30551 10364
rect 30551 10308 30555 10364
rect 30491 10304 30555 10308
rect 30571 10364 30635 10368
rect 30571 10308 30575 10364
rect 30575 10308 30631 10364
rect 30631 10308 30635 10364
rect 30571 10304 30635 10308
rect 9346 9820 9410 9824
rect 9346 9764 9350 9820
rect 9350 9764 9406 9820
rect 9406 9764 9410 9820
rect 9346 9760 9410 9764
rect 9426 9820 9490 9824
rect 9426 9764 9430 9820
rect 9430 9764 9486 9820
rect 9486 9764 9490 9820
rect 9426 9760 9490 9764
rect 9506 9820 9570 9824
rect 9506 9764 9510 9820
rect 9510 9764 9566 9820
rect 9566 9764 9570 9820
rect 9506 9760 9570 9764
rect 9586 9820 9650 9824
rect 9586 9764 9590 9820
rect 9590 9764 9646 9820
rect 9646 9764 9650 9820
rect 9586 9760 9650 9764
rect 17740 9820 17804 9824
rect 17740 9764 17744 9820
rect 17744 9764 17800 9820
rect 17800 9764 17804 9820
rect 17740 9760 17804 9764
rect 17820 9820 17884 9824
rect 17820 9764 17824 9820
rect 17824 9764 17880 9820
rect 17880 9764 17884 9820
rect 17820 9760 17884 9764
rect 17900 9820 17964 9824
rect 17900 9764 17904 9820
rect 17904 9764 17960 9820
rect 17960 9764 17964 9820
rect 17900 9760 17964 9764
rect 17980 9820 18044 9824
rect 17980 9764 17984 9820
rect 17984 9764 18040 9820
rect 18040 9764 18044 9820
rect 17980 9760 18044 9764
rect 26134 9820 26198 9824
rect 26134 9764 26138 9820
rect 26138 9764 26194 9820
rect 26194 9764 26198 9820
rect 26134 9760 26198 9764
rect 26214 9820 26278 9824
rect 26214 9764 26218 9820
rect 26218 9764 26274 9820
rect 26274 9764 26278 9820
rect 26214 9760 26278 9764
rect 26294 9820 26358 9824
rect 26294 9764 26298 9820
rect 26298 9764 26354 9820
rect 26354 9764 26358 9820
rect 26294 9760 26358 9764
rect 26374 9820 26438 9824
rect 26374 9764 26378 9820
rect 26378 9764 26434 9820
rect 26434 9764 26438 9820
rect 26374 9760 26438 9764
rect 34528 9820 34592 9824
rect 34528 9764 34532 9820
rect 34532 9764 34588 9820
rect 34588 9764 34592 9820
rect 34528 9760 34592 9764
rect 34608 9820 34672 9824
rect 34608 9764 34612 9820
rect 34612 9764 34668 9820
rect 34668 9764 34672 9820
rect 34608 9760 34672 9764
rect 34688 9820 34752 9824
rect 34688 9764 34692 9820
rect 34692 9764 34748 9820
rect 34748 9764 34752 9820
rect 34688 9760 34752 9764
rect 34768 9820 34832 9824
rect 34768 9764 34772 9820
rect 34772 9764 34828 9820
rect 34828 9764 34832 9820
rect 34768 9760 34832 9764
rect 5149 9276 5213 9280
rect 5149 9220 5153 9276
rect 5153 9220 5209 9276
rect 5209 9220 5213 9276
rect 5149 9216 5213 9220
rect 5229 9276 5293 9280
rect 5229 9220 5233 9276
rect 5233 9220 5289 9276
rect 5289 9220 5293 9276
rect 5229 9216 5293 9220
rect 5309 9276 5373 9280
rect 5309 9220 5313 9276
rect 5313 9220 5369 9276
rect 5369 9220 5373 9276
rect 5309 9216 5373 9220
rect 5389 9276 5453 9280
rect 5389 9220 5393 9276
rect 5393 9220 5449 9276
rect 5449 9220 5453 9276
rect 5389 9216 5453 9220
rect 13543 9276 13607 9280
rect 13543 9220 13547 9276
rect 13547 9220 13603 9276
rect 13603 9220 13607 9276
rect 13543 9216 13607 9220
rect 13623 9276 13687 9280
rect 13623 9220 13627 9276
rect 13627 9220 13683 9276
rect 13683 9220 13687 9276
rect 13623 9216 13687 9220
rect 13703 9276 13767 9280
rect 13703 9220 13707 9276
rect 13707 9220 13763 9276
rect 13763 9220 13767 9276
rect 13703 9216 13767 9220
rect 13783 9276 13847 9280
rect 13783 9220 13787 9276
rect 13787 9220 13843 9276
rect 13843 9220 13847 9276
rect 13783 9216 13847 9220
rect 21937 9276 22001 9280
rect 21937 9220 21941 9276
rect 21941 9220 21997 9276
rect 21997 9220 22001 9276
rect 21937 9216 22001 9220
rect 22017 9276 22081 9280
rect 22017 9220 22021 9276
rect 22021 9220 22077 9276
rect 22077 9220 22081 9276
rect 22017 9216 22081 9220
rect 22097 9276 22161 9280
rect 22097 9220 22101 9276
rect 22101 9220 22157 9276
rect 22157 9220 22161 9276
rect 22097 9216 22161 9220
rect 22177 9276 22241 9280
rect 22177 9220 22181 9276
rect 22181 9220 22237 9276
rect 22237 9220 22241 9276
rect 22177 9216 22241 9220
rect 30331 9276 30395 9280
rect 30331 9220 30335 9276
rect 30335 9220 30391 9276
rect 30391 9220 30395 9276
rect 30331 9216 30395 9220
rect 30411 9276 30475 9280
rect 30411 9220 30415 9276
rect 30415 9220 30471 9276
rect 30471 9220 30475 9276
rect 30411 9216 30475 9220
rect 30491 9276 30555 9280
rect 30491 9220 30495 9276
rect 30495 9220 30551 9276
rect 30551 9220 30555 9276
rect 30491 9216 30555 9220
rect 30571 9276 30635 9280
rect 30571 9220 30575 9276
rect 30575 9220 30631 9276
rect 30631 9220 30635 9276
rect 30571 9216 30635 9220
rect 9346 8732 9410 8736
rect 9346 8676 9350 8732
rect 9350 8676 9406 8732
rect 9406 8676 9410 8732
rect 9346 8672 9410 8676
rect 9426 8732 9490 8736
rect 9426 8676 9430 8732
rect 9430 8676 9486 8732
rect 9486 8676 9490 8732
rect 9426 8672 9490 8676
rect 9506 8732 9570 8736
rect 9506 8676 9510 8732
rect 9510 8676 9566 8732
rect 9566 8676 9570 8732
rect 9506 8672 9570 8676
rect 9586 8732 9650 8736
rect 9586 8676 9590 8732
rect 9590 8676 9646 8732
rect 9646 8676 9650 8732
rect 9586 8672 9650 8676
rect 17740 8732 17804 8736
rect 17740 8676 17744 8732
rect 17744 8676 17800 8732
rect 17800 8676 17804 8732
rect 17740 8672 17804 8676
rect 17820 8732 17884 8736
rect 17820 8676 17824 8732
rect 17824 8676 17880 8732
rect 17880 8676 17884 8732
rect 17820 8672 17884 8676
rect 17900 8732 17964 8736
rect 17900 8676 17904 8732
rect 17904 8676 17960 8732
rect 17960 8676 17964 8732
rect 17900 8672 17964 8676
rect 17980 8732 18044 8736
rect 17980 8676 17984 8732
rect 17984 8676 18040 8732
rect 18040 8676 18044 8732
rect 17980 8672 18044 8676
rect 26134 8732 26198 8736
rect 26134 8676 26138 8732
rect 26138 8676 26194 8732
rect 26194 8676 26198 8732
rect 26134 8672 26198 8676
rect 26214 8732 26278 8736
rect 26214 8676 26218 8732
rect 26218 8676 26274 8732
rect 26274 8676 26278 8732
rect 26214 8672 26278 8676
rect 26294 8732 26358 8736
rect 26294 8676 26298 8732
rect 26298 8676 26354 8732
rect 26354 8676 26358 8732
rect 26294 8672 26358 8676
rect 26374 8732 26438 8736
rect 26374 8676 26378 8732
rect 26378 8676 26434 8732
rect 26434 8676 26438 8732
rect 26374 8672 26438 8676
rect 34528 8732 34592 8736
rect 34528 8676 34532 8732
rect 34532 8676 34588 8732
rect 34588 8676 34592 8732
rect 34528 8672 34592 8676
rect 34608 8732 34672 8736
rect 34608 8676 34612 8732
rect 34612 8676 34668 8732
rect 34668 8676 34672 8732
rect 34608 8672 34672 8676
rect 34688 8732 34752 8736
rect 34688 8676 34692 8732
rect 34692 8676 34748 8732
rect 34748 8676 34752 8732
rect 34688 8672 34752 8676
rect 34768 8732 34832 8736
rect 34768 8676 34772 8732
rect 34772 8676 34828 8732
rect 34828 8676 34832 8732
rect 34768 8672 34832 8676
rect 5149 8188 5213 8192
rect 5149 8132 5153 8188
rect 5153 8132 5209 8188
rect 5209 8132 5213 8188
rect 5149 8128 5213 8132
rect 5229 8188 5293 8192
rect 5229 8132 5233 8188
rect 5233 8132 5289 8188
rect 5289 8132 5293 8188
rect 5229 8128 5293 8132
rect 5309 8188 5373 8192
rect 5309 8132 5313 8188
rect 5313 8132 5369 8188
rect 5369 8132 5373 8188
rect 5309 8128 5373 8132
rect 5389 8188 5453 8192
rect 5389 8132 5393 8188
rect 5393 8132 5449 8188
rect 5449 8132 5453 8188
rect 5389 8128 5453 8132
rect 13543 8188 13607 8192
rect 13543 8132 13547 8188
rect 13547 8132 13603 8188
rect 13603 8132 13607 8188
rect 13543 8128 13607 8132
rect 13623 8188 13687 8192
rect 13623 8132 13627 8188
rect 13627 8132 13683 8188
rect 13683 8132 13687 8188
rect 13623 8128 13687 8132
rect 13703 8188 13767 8192
rect 13703 8132 13707 8188
rect 13707 8132 13763 8188
rect 13763 8132 13767 8188
rect 13703 8128 13767 8132
rect 13783 8188 13847 8192
rect 13783 8132 13787 8188
rect 13787 8132 13843 8188
rect 13843 8132 13847 8188
rect 13783 8128 13847 8132
rect 21937 8188 22001 8192
rect 21937 8132 21941 8188
rect 21941 8132 21997 8188
rect 21997 8132 22001 8188
rect 21937 8128 22001 8132
rect 22017 8188 22081 8192
rect 22017 8132 22021 8188
rect 22021 8132 22077 8188
rect 22077 8132 22081 8188
rect 22017 8128 22081 8132
rect 22097 8188 22161 8192
rect 22097 8132 22101 8188
rect 22101 8132 22157 8188
rect 22157 8132 22161 8188
rect 22097 8128 22161 8132
rect 22177 8188 22241 8192
rect 22177 8132 22181 8188
rect 22181 8132 22237 8188
rect 22237 8132 22241 8188
rect 22177 8128 22241 8132
rect 30331 8188 30395 8192
rect 30331 8132 30335 8188
rect 30335 8132 30391 8188
rect 30391 8132 30395 8188
rect 30331 8128 30395 8132
rect 30411 8188 30475 8192
rect 30411 8132 30415 8188
rect 30415 8132 30471 8188
rect 30471 8132 30475 8188
rect 30411 8128 30475 8132
rect 30491 8188 30555 8192
rect 30491 8132 30495 8188
rect 30495 8132 30551 8188
rect 30551 8132 30555 8188
rect 30491 8128 30555 8132
rect 30571 8188 30635 8192
rect 30571 8132 30575 8188
rect 30575 8132 30631 8188
rect 30631 8132 30635 8188
rect 30571 8128 30635 8132
rect 9346 7644 9410 7648
rect 9346 7588 9350 7644
rect 9350 7588 9406 7644
rect 9406 7588 9410 7644
rect 9346 7584 9410 7588
rect 9426 7644 9490 7648
rect 9426 7588 9430 7644
rect 9430 7588 9486 7644
rect 9486 7588 9490 7644
rect 9426 7584 9490 7588
rect 9506 7644 9570 7648
rect 9506 7588 9510 7644
rect 9510 7588 9566 7644
rect 9566 7588 9570 7644
rect 9506 7584 9570 7588
rect 9586 7644 9650 7648
rect 9586 7588 9590 7644
rect 9590 7588 9646 7644
rect 9646 7588 9650 7644
rect 9586 7584 9650 7588
rect 17740 7644 17804 7648
rect 17740 7588 17744 7644
rect 17744 7588 17800 7644
rect 17800 7588 17804 7644
rect 17740 7584 17804 7588
rect 17820 7644 17884 7648
rect 17820 7588 17824 7644
rect 17824 7588 17880 7644
rect 17880 7588 17884 7644
rect 17820 7584 17884 7588
rect 17900 7644 17964 7648
rect 17900 7588 17904 7644
rect 17904 7588 17960 7644
rect 17960 7588 17964 7644
rect 17900 7584 17964 7588
rect 17980 7644 18044 7648
rect 17980 7588 17984 7644
rect 17984 7588 18040 7644
rect 18040 7588 18044 7644
rect 17980 7584 18044 7588
rect 26134 7644 26198 7648
rect 26134 7588 26138 7644
rect 26138 7588 26194 7644
rect 26194 7588 26198 7644
rect 26134 7584 26198 7588
rect 26214 7644 26278 7648
rect 26214 7588 26218 7644
rect 26218 7588 26274 7644
rect 26274 7588 26278 7644
rect 26214 7584 26278 7588
rect 26294 7644 26358 7648
rect 26294 7588 26298 7644
rect 26298 7588 26354 7644
rect 26354 7588 26358 7644
rect 26294 7584 26358 7588
rect 26374 7644 26438 7648
rect 26374 7588 26378 7644
rect 26378 7588 26434 7644
rect 26434 7588 26438 7644
rect 26374 7584 26438 7588
rect 34528 7644 34592 7648
rect 34528 7588 34532 7644
rect 34532 7588 34588 7644
rect 34588 7588 34592 7644
rect 34528 7584 34592 7588
rect 34608 7644 34672 7648
rect 34608 7588 34612 7644
rect 34612 7588 34668 7644
rect 34668 7588 34672 7644
rect 34608 7584 34672 7588
rect 34688 7644 34752 7648
rect 34688 7588 34692 7644
rect 34692 7588 34748 7644
rect 34748 7588 34752 7644
rect 34688 7584 34752 7588
rect 34768 7644 34832 7648
rect 34768 7588 34772 7644
rect 34772 7588 34828 7644
rect 34828 7588 34832 7644
rect 34768 7584 34832 7588
rect 5149 7100 5213 7104
rect 5149 7044 5153 7100
rect 5153 7044 5209 7100
rect 5209 7044 5213 7100
rect 5149 7040 5213 7044
rect 5229 7100 5293 7104
rect 5229 7044 5233 7100
rect 5233 7044 5289 7100
rect 5289 7044 5293 7100
rect 5229 7040 5293 7044
rect 5309 7100 5373 7104
rect 5309 7044 5313 7100
rect 5313 7044 5369 7100
rect 5369 7044 5373 7100
rect 5309 7040 5373 7044
rect 5389 7100 5453 7104
rect 5389 7044 5393 7100
rect 5393 7044 5449 7100
rect 5449 7044 5453 7100
rect 5389 7040 5453 7044
rect 13543 7100 13607 7104
rect 13543 7044 13547 7100
rect 13547 7044 13603 7100
rect 13603 7044 13607 7100
rect 13543 7040 13607 7044
rect 13623 7100 13687 7104
rect 13623 7044 13627 7100
rect 13627 7044 13683 7100
rect 13683 7044 13687 7100
rect 13623 7040 13687 7044
rect 13703 7100 13767 7104
rect 13703 7044 13707 7100
rect 13707 7044 13763 7100
rect 13763 7044 13767 7100
rect 13703 7040 13767 7044
rect 13783 7100 13847 7104
rect 13783 7044 13787 7100
rect 13787 7044 13843 7100
rect 13843 7044 13847 7100
rect 13783 7040 13847 7044
rect 21937 7100 22001 7104
rect 21937 7044 21941 7100
rect 21941 7044 21997 7100
rect 21997 7044 22001 7100
rect 21937 7040 22001 7044
rect 22017 7100 22081 7104
rect 22017 7044 22021 7100
rect 22021 7044 22077 7100
rect 22077 7044 22081 7100
rect 22017 7040 22081 7044
rect 22097 7100 22161 7104
rect 22097 7044 22101 7100
rect 22101 7044 22157 7100
rect 22157 7044 22161 7100
rect 22097 7040 22161 7044
rect 22177 7100 22241 7104
rect 22177 7044 22181 7100
rect 22181 7044 22237 7100
rect 22237 7044 22241 7100
rect 22177 7040 22241 7044
rect 30331 7100 30395 7104
rect 30331 7044 30335 7100
rect 30335 7044 30391 7100
rect 30391 7044 30395 7100
rect 30331 7040 30395 7044
rect 30411 7100 30475 7104
rect 30411 7044 30415 7100
rect 30415 7044 30471 7100
rect 30471 7044 30475 7100
rect 30411 7040 30475 7044
rect 30491 7100 30555 7104
rect 30491 7044 30495 7100
rect 30495 7044 30551 7100
rect 30551 7044 30555 7100
rect 30491 7040 30555 7044
rect 30571 7100 30635 7104
rect 30571 7044 30575 7100
rect 30575 7044 30631 7100
rect 30631 7044 30635 7100
rect 30571 7040 30635 7044
rect 9346 6556 9410 6560
rect 9346 6500 9350 6556
rect 9350 6500 9406 6556
rect 9406 6500 9410 6556
rect 9346 6496 9410 6500
rect 9426 6556 9490 6560
rect 9426 6500 9430 6556
rect 9430 6500 9486 6556
rect 9486 6500 9490 6556
rect 9426 6496 9490 6500
rect 9506 6556 9570 6560
rect 9506 6500 9510 6556
rect 9510 6500 9566 6556
rect 9566 6500 9570 6556
rect 9506 6496 9570 6500
rect 9586 6556 9650 6560
rect 9586 6500 9590 6556
rect 9590 6500 9646 6556
rect 9646 6500 9650 6556
rect 9586 6496 9650 6500
rect 17740 6556 17804 6560
rect 17740 6500 17744 6556
rect 17744 6500 17800 6556
rect 17800 6500 17804 6556
rect 17740 6496 17804 6500
rect 17820 6556 17884 6560
rect 17820 6500 17824 6556
rect 17824 6500 17880 6556
rect 17880 6500 17884 6556
rect 17820 6496 17884 6500
rect 17900 6556 17964 6560
rect 17900 6500 17904 6556
rect 17904 6500 17960 6556
rect 17960 6500 17964 6556
rect 17900 6496 17964 6500
rect 17980 6556 18044 6560
rect 17980 6500 17984 6556
rect 17984 6500 18040 6556
rect 18040 6500 18044 6556
rect 17980 6496 18044 6500
rect 26134 6556 26198 6560
rect 26134 6500 26138 6556
rect 26138 6500 26194 6556
rect 26194 6500 26198 6556
rect 26134 6496 26198 6500
rect 26214 6556 26278 6560
rect 26214 6500 26218 6556
rect 26218 6500 26274 6556
rect 26274 6500 26278 6556
rect 26214 6496 26278 6500
rect 26294 6556 26358 6560
rect 26294 6500 26298 6556
rect 26298 6500 26354 6556
rect 26354 6500 26358 6556
rect 26294 6496 26358 6500
rect 26374 6556 26438 6560
rect 26374 6500 26378 6556
rect 26378 6500 26434 6556
rect 26434 6500 26438 6556
rect 26374 6496 26438 6500
rect 34528 6556 34592 6560
rect 34528 6500 34532 6556
rect 34532 6500 34588 6556
rect 34588 6500 34592 6556
rect 34528 6496 34592 6500
rect 34608 6556 34672 6560
rect 34608 6500 34612 6556
rect 34612 6500 34668 6556
rect 34668 6500 34672 6556
rect 34608 6496 34672 6500
rect 34688 6556 34752 6560
rect 34688 6500 34692 6556
rect 34692 6500 34748 6556
rect 34748 6500 34752 6556
rect 34688 6496 34752 6500
rect 34768 6556 34832 6560
rect 34768 6500 34772 6556
rect 34772 6500 34828 6556
rect 34828 6500 34832 6556
rect 34768 6496 34832 6500
rect 5149 6012 5213 6016
rect 5149 5956 5153 6012
rect 5153 5956 5209 6012
rect 5209 5956 5213 6012
rect 5149 5952 5213 5956
rect 5229 6012 5293 6016
rect 5229 5956 5233 6012
rect 5233 5956 5289 6012
rect 5289 5956 5293 6012
rect 5229 5952 5293 5956
rect 5309 6012 5373 6016
rect 5309 5956 5313 6012
rect 5313 5956 5369 6012
rect 5369 5956 5373 6012
rect 5309 5952 5373 5956
rect 5389 6012 5453 6016
rect 5389 5956 5393 6012
rect 5393 5956 5449 6012
rect 5449 5956 5453 6012
rect 5389 5952 5453 5956
rect 13543 6012 13607 6016
rect 13543 5956 13547 6012
rect 13547 5956 13603 6012
rect 13603 5956 13607 6012
rect 13543 5952 13607 5956
rect 13623 6012 13687 6016
rect 13623 5956 13627 6012
rect 13627 5956 13683 6012
rect 13683 5956 13687 6012
rect 13623 5952 13687 5956
rect 13703 6012 13767 6016
rect 13703 5956 13707 6012
rect 13707 5956 13763 6012
rect 13763 5956 13767 6012
rect 13703 5952 13767 5956
rect 13783 6012 13847 6016
rect 13783 5956 13787 6012
rect 13787 5956 13843 6012
rect 13843 5956 13847 6012
rect 13783 5952 13847 5956
rect 21937 6012 22001 6016
rect 21937 5956 21941 6012
rect 21941 5956 21997 6012
rect 21997 5956 22001 6012
rect 21937 5952 22001 5956
rect 22017 6012 22081 6016
rect 22017 5956 22021 6012
rect 22021 5956 22077 6012
rect 22077 5956 22081 6012
rect 22017 5952 22081 5956
rect 22097 6012 22161 6016
rect 22097 5956 22101 6012
rect 22101 5956 22157 6012
rect 22157 5956 22161 6012
rect 22097 5952 22161 5956
rect 22177 6012 22241 6016
rect 22177 5956 22181 6012
rect 22181 5956 22237 6012
rect 22237 5956 22241 6012
rect 22177 5952 22241 5956
rect 30331 6012 30395 6016
rect 30331 5956 30335 6012
rect 30335 5956 30391 6012
rect 30391 5956 30395 6012
rect 30331 5952 30395 5956
rect 30411 6012 30475 6016
rect 30411 5956 30415 6012
rect 30415 5956 30471 6012
rect 30471 5956 30475 6012
rect 30411 5952 30475 5956
rect 30491 6012 30555 6016
rect 30491 5956 30495 6012
rect 30495 5956 30551 6012
rect 30551 5956 30555 6012
rect 30491 5952 30555 5956
rect 30571 6012 30635 6016
rect 30571 5956 30575 6012
rect 30575 5956 30631 6012
rect 30631 5956 30635 6012
rect 30571 5952 30635 5956
rect 9346 5468 9410 5472
rect 9346 5412 9350 5468
rect 9350 5412 9406 5468
rect 9406 5412 9410 5468
rect 9346 5408 9410 5412
rect 9426 5468 9490 5472
rect 9426 5412 9430 5468
rect 9430 5412 9486 5468
rect 9486 5412 9490 5468
rect 9426 5408 9490 5412
rect 9506 5468 9570 5472
rect 9506 5412 9510 5468
rect 9510 5412 9566 5468
rect 9566 5412 9570 5468
rect 9506 5408 9570 5412
rect 9586 5468 9650 5472
rect 9586 5412 9590 5468
rect 9590 5412 9646 5468
rect 9646 5412 9650 5468
rect 9586 5408 9650 5412
rect 17740 5468 17804 5472
rect 17740 5412 17744 5468
rect 17744 5412 17800 5468
rect 17800 5412 17804 5468
rect 17740 5408 17804 5412
rect 17820 5468 17884 5472
rect 17820 5412 17824 5468
rect 17824 5412 17880 5468
rect 17880 5412 17884 5468
rect 17820 5408 17884 5412
rect 17900 5468 17964 5472
rect 17900 5412 17904 5468
rect 17904 5412 17960 5468
rect 17960 5412 17964 5468
rect 17900 5408 17964 5412
rect 17980 5468 18044 5472
rect 17980 5412 17984 5468
rect 17984 5412 18040 5468
rect 18040 5412 18044 5468
rect 17980 5408 18044 5412
rect 26134 5468 26198 5472
rect 26134 5412 26138 5468
rect 26138 5412 26194 5468
rect 26194 5412 26198 5468
rect 26134 5408 26198 5412
rect 26214 5468 26278 5472
rect 26214 5412 26218 5468
rect 26218 5412 26274 5468
rect 26274 5412 26278 5468
rect 26214 5408 26278 5412
rect 26294 5468 26358 5472
rect 26294 5412 26298 5468
rect 26298 5412 26354 5468
rect 26354 5412 26358 5468
rect 26294 5408 26358 5412
rect 26374 5468 26438 5472
rect 26374 5412 26378 5468
rect 26378 5412 26434 5468
rect 26434 5412 26438 5468
rect 26374 5408 26438 5412
rect 34528 5468 34592 5472
rect 34528 5412 34532 5468
rect 34532 5412 34588 5468
rect 34588 5412 34592 5468
rect 34528 5408 34592 5412
rect 34608 5468 34672 5472
rect 34608 5412 34612 5468
rect 34612 5412 34668 5468
rect 34668 5412 34672 5468
rect 34608 5408 34672 5412
rect 34688 5468 34752 5472
rect 34688 5412 34692 5468
rect 34692 5412 34748 5468
rect 34748 5412 34752 5468
rect 34688 5408 34752 5412
rect 34768 5468 34832 5472
rect 34768 5412 34772 5468
rect 34772 5412 34828 5468
rect 34828 5412 34832 5468
rect 34768 5408 34832 5412
rect 5149 4924 5213 4928
rect 5149 4868 5153 4924
rect 5153 4868 5209 4924
rect 5209 4868 5213 4924
rect 5149 4864 5213 4868
rect 5229 4924 5293 4928
rect 5229 4868 5233 4924
rect 5233 4868 5289 4924
rect 5289 4868 5293 4924
rect 5229 4864 5293 4868
rect 5309 4924 5373 4928
rect 5309 4868 5313 4924
rect 5313 4868 5369 4924
rect 5369 4868 5373 4924
rect 5309 4864 5373 4868
rect 5389 4924 5453 4928
rect 5389 4868 5393 4924
rect 5393 4868 5449 4924
rect 5449 4868 5453 4924
rect 5389 4864 5453 4868
rect 13543 4924 13607 4928
rect 13543 4868 13547 4924
rect 13547 4868 13603 4924
rect 13603 4868 13607 4924
rect 13543 4864 13607 4868
rect 13623 4924 13687 4928
rect 13623 4868 13627 4924
rect 13627 4868 13683 4924
rect 13683 4868 13687 4924
rect 13623 4864 13687 4868
rect 13703 4924 13767 4928
rect 13703 4868 13707 4924
rect 13707 4868 13763 4924
rect 13763 4868 13767 4924
rect 13703 4864 13767 4868
rect 13783 4924 13847 4928
rect 13783 4868 13787 4924
rect 13787 4868 13843 4924
rect 13843 4868 13847 4924
rect 13783 4864 13847 4868
rect 21937 4924 22001 4928
rect 21937 4868 21941 4924
rect 21941 4868 21997 4924
rect 21997 4868 22001 4924
rect 21937 4864 22001 4868
rect 22017 4924 22081 4928
rect 22017 4868 22021 4924
rect 22021 4868 22077 4924
rect 22077 4868 22081 4924
rect 22017 4864 22081 4868
rect 22097 4924 22161 4928
rect 22097 4868 22101 4924
rect 22101 4868 22157 4924
rect 22157 4868 22161 4924
rect 22097 4864 22161 4868
rect 22177 4924 22241 4928
rect 22177 4868 22181 4924
rect 22181 4868 22237 4924
rect 22237 4868 22241 4924
rect 22177 4864 22241 4868
rect 30331 4924 30395 4928
rect 30331 4868 30335 4924
rect 30335 4868 30391 4924
rect 30391 4868 30395 4924
rect 30331 4864 30395 4868
rect 30411 4924 30475 4928
rect 30411 4868 30415 4924
rect 30415 4868 30471 4924
rect 30471 4868 30475 4924
rect 30411 4864 30475 4868
rect 30491 4924 30555 4928
rect 30491 4868 30495 4924
rect 30495 4868 30551 4924
rect 30551 4868 30555 4924
rect 30491 4864 30555 4868
rect 30571 4924 30635 4928
rect 30571 4868 30575 4924
rect 30575 4868 30631 4924
rect 30631 4868 30635 4924
rect 30571 4864 30635 4868
rect 9346 4380 9410 4384
rect 9346 4324 9350 4380
rect 9350 4324 9406 4380
rect 9406 4324 9410 4380
rect 9346 4320 9410 4324
rect 9426 4380 9490 4384
rect 9426 4324 9430 4380
rect 9430 4324 9486 4380
rect 9486 4324 9490 4380
rect 9426 4320 9490 4324
rect 9506 4380 9570 4384
rect 9506 4324 9510 4380
rect 9510 4324 9566 4380
rect 9566 4324 9570 4380
rect 9506 4320 9570 4324
rect 9586 4380 9650 4384
rect 9586 4324 9590 4380
rect 9590 4324 9646 4380
rect 9646 4324 9650 4380
rect 9586 4320 9650 4324
rect 17740 4380 17804 4384
rect 17740 4324 17744 4380
rect 17744 4324 17800 4380
rect 17800 4324 17804 4380
rect 17740 4320 17804 4324
rect 17820 4380 17884 4384
rect 17820 4324 17824 4380
rect 17824 4324 17880 4380
rect 17880 4324 17884 4380
rect 17820 4320 17884 4324
rect 17900 4380 17964 4384
rect 17900 4324 17904 4380
rect 17904 4324 17960 4380
rect 17960 4324 17964 4380
rect 17900 4320 17964 4324
rect 17980 4380 18044 4384
rect 17980 4324 17984 4380
rect 17984 4324 18040 4380
rect 18040 4324 18044 4380
rect 17980 4320 18044 4324
rect 26134 4380 26198 4384
rect 26134 4324 26138 4380
rect 26138 4324 26194 4380
rect 26194 4324 26198 4380
rect 26134 4320 26198 4324
rect 26214 4380 26278 4384
rect 26214 4324 26218 4380
rect 26218 4324 26274 4380
rect 26274 4324 26278 4380
rect 26214 4320 26278 4324
rect 26294 4380 26358 4384
rect 26294 4324 26298 4380
rect 26298 4324 26354 4380
rect 26354 4324 26358 4380
rect 26294 4320 26358 4324
rect 26374 4380 26438 4384
rect 26374 4324 26378 4380
rect 26378 4324 26434 4380
rect 26434 4324 26438 4380
rect 26374 4320 26438 4324
rect 34528 4380 34592 4384
rect 34528 4324 34532 4380
rect 34532 4324 34588 4380
rect 34588 4324 34592 4380
rect 34528 4320 34592 4324
rect 34608 4380 34672 4384
rect 34608 4324 34612 4380
rect 34612 4324 34668 4380
rect 34668 4324 34672 4380
rect 34608 4320 34672 4324
rect 34688 4380 34752 4384
rect 34688 4324 34692 4380
rect 34692 4324 34748 4380
rect 34748 4324 34752 4380
rect 34688 4320 34752 4324
rect 34768 4380 34832 4384
rect 34768 4324 34772 4380
rect 34772 4324 34828 4380
rect 34828 4324 34832 4380
rect 34768 4320 34832 4324
rect 5149 3836 5213 3840
rect 5149 3780 5153 3836
rect 5153 3780 5209 3836
rect 5209 3780 5213 3836
rect 5149 3776 5213 3780
rect 5229 3836 5293 3840
rect 5229 3780 5233 3836
rect 5233 3780 5289 3836
rect 5289 3780 5293 3836
rect 5229 3776 5293 3780
rect 5309 3836 5373 3840
rect 5309 3780 5313 3836
rect 5313 3780 5369 3836
rect 5369 3780 5373 3836
rect 5309 3776 5373 3780
rect 5389 3836 5453 3840
rect 5389 3780 5393 3836
rect 5393 3780 5449 3836
rect 5449 3780 5453 3836
rect 5389 3776 5453 3780
rect 13543 3836 13607 3840
rect 13543 3780 13547 3836
rect 13547 3780 13603 3836
rect 13603 3780 13607 3836
rect 13543 3776 13607 3780
rect 13623 3836 13687 3840
rect 13623 3780 13627 3836
rect 13627 3780 13683 3836
rect 13683 3780 13687 3836
rect 13623 3776 13687 3780
rect 13703 3836 13767 3840
rect 13703 3780 13707 3836
rect 13707 3780 13763 3836
rect 13763 3780 13767 3836
rect 13703 3776 13767 3780
rect 13783 3836 13847 3840
rect 13783 3780 13787 3836
rect 13787 3780 13843 3836
rect 13843 3780 13847 3836
rect 13783 3776 13847 3780
rect 21937 3836 22001 3840
rect 21937 3780 21941 3836
rect 21941 3780 21997 3836
rect 21997 3780 22001 3836
rect 21937 3776 22001 3780
rect 22017 3836 22081 3840
rect 22017 3780 22021 3836
rect 22021 3780 22077 3836
rect 22077 3780 22081 3836
rect 22017 3776 22081 3780
rect 22097 3836 22161 3840
rect 22097 3780 22101 3836
rect 22101 3780 22157 3836
rect 22157 3780 22161 3836
rect 22097 3776 22161 3780
rect 22177 3836 22241 3840
rect 22177 3780 22181 3836
rect 22181 3780 22237 3836
rect 22237 3780 22241 3836
rect 22177 3776 22241 3780
rect 30331 3836 30395 3840
rect 30331 3780 30335 3836
rect 30335 3780 30391 3836
rect 30391 3780 30395 3836
rect 30331 3776 30395 3780
rect 30411 3836 30475 3840
rect 30411 3780 30415 3836
rect 30415 3780 30471 3836
rect 30471 3780 30475 3836
rect 30411 3776 30475 3780
rect 30491 3836 30555 3840
rect 30491 3780 30495 3836
rect 30495 3780 30551 3836
rect 30551 3780 30555 3836
rect 30491 3776 30555 3780
rect 30571 3836 30635 3840
rect 30571 3780 30575 3836
rect 30575 3780 30631 3836
rect 30631 3780 30635 3836
rect 30571 3776 30635 3780
rect 9346 3292 9410 3296
rect 9346 3236 9350 3292
rect 9350 3236 9406 3292
rect 9406 3236 9410 3292
rect 9346 3232 9410 3236
rect 9426 3292 9490 3296
rect 9426 3236 9430 3292
rect 9430 3236 9486 3292
rect 9486 3236 9490 3292
rect 9426 3232 9490 3236
rect 9506 3292 9570 3296
rect 9506 3236 9510 3292
rect 9510 3236 9566 3292
rect 9566 3236 9570 3292
rect 9506 3232 9570 3236
rect 9586 3292 9650 3296
rect 9586 3236 9590 3292
rect 9590 3236 9646 3292
rect 9646 3236 9650 3292
rect 9586 3232 9650 3236
rect 17740 3292 17804 3296
rect 17740 3236 17744 3292
rect 17744 3236 17800 3292
rect 17800 3236 17804 3292
rect 17740 3232 17804 3236
rect 17820 3292 17884 3296
rect 17820 3236 17824 3292
rect 17824 3236 17880 3292
rect 17880 3236 17884 3292
rect 17820 3232 17884 3236
rect 17900 3292 17964 3296
rect 17900 3236 17904 3292
rect 17904 3236 17960 3292
rect 17960 3236 17964 3292
rect 17900 3232 17964 3236
rect 17980 3292 18044 3296
rect 17980 3236 17984 3292
rect 17984 3236 18040 3292
rect 18040 3236 18044 3292
rect 17980 3232 18044 3236
rect 26134 3292 26198 3296
rect 26134 3236 26138 3292
rect 26138 3236 26194 3292
rect 26194 3236 26198 3292
rect 26134 3232 26198 3236
rect 26214 3292 26278 3296
rect 26214 3236 26218 3292
rect 26218 3236 26274 3292
rect 26274 3236 26278 3292
rect 26214 3232 26278 3236
rect 26294 3292 26358 3296
rect 26294 3236 26298 3292
rect 26298 3236 26354 3292
rect 26354 3236 26358 3292
rect 26294 3232 26358 3236
rect 26374 3292 26438 3296
rect 26374 3236 26378 3292
rect 26378 3236 26434 3292
rect 26434 3236 26438 3292
rect 26374 3232 26438 3236
rect 34528 3292 34592 3296
rect 34528 3236 34532 3292
rect 34532 3236 34588 3292
rect 34588 3236 34592 3292
rect 34528 3232 34592 3236
rect 34608 3292 34672 3296
rect 34608 3236 34612 3292
rect 34612 3236 34668 3292
rect 34668 3236 34672 3292
rect 34608 3232 34672 3236
rect 34688 3292 34752 3296
rect 34688 3236 34692 3292
rect 34692 3236 34748 3292
rect 34748 3236 34752 3292
rect 34688 3232 34752 3236
rect 34768 3292 34832 3296
rect 34768 3236 34772 3292
rect 34772 3236 34828 3292
rect 34828 3236 34832 3292
rect 34768 3232 34832 3236
rect 5149 2748 5213 2752
rect 5149 2692 5153 2748
rect 5153 2692 5209 2748
rect 5209 2692 5213 2748
rect 5149 2688 5213 2692
rect 5229 2748 5293 2752
rect 5229 2692 5233 2748
rect 5233 2692 5289 2748
rect 5289 2692 5293 2748
rect 5229 2688 5293 2692
rect 5309 2748 5373 2752
rect 5309 2692 5313 2748
rect 5313 2692 5369 2748
rect 5369 2692 5373 2748
rect 5309 2688 5373 2692
rect 5389 2748 5453 2752
rect 5389 2692 5393 2748
rect 5393 2692 5449 2748
rect 5449 2692 5453 2748
rect 5389 2688 5453 2692
rect 13543 2748 13607 2752
rect 13543 2692 13547 2748
rect 13547 2692 13603 2748
rect 13603 2692 13607 2748
rect 13543 2688 13607 2692
rect 13623 2748 13687 2752
rect 13623 2692 13627 2748
rect 13627 2692 13683 2748
rect 13683 2692 13687 2748
rect 13623 2688 13687 2692
rect 13703 2748 13767 2752
rect 13703 2692 13707 2748
rect 13707 2692 13763 2748
rect 13763 2692 13767 2748
rect 13703 2688 13767 2692
rect 13783 2748 13847 2752
rect 13783 2692 13787 2748
rect 13787 2692 13843 2748
rect 13843 2692 13847 2748
rect 13783 2688 13847 2692
rect 21937 2748 22001 2752
rect 21937 2692 21941 2748
rect 21941 2692 21997 2748
rect 21997 2692 22001 2748
rect 21937 2688 22001 2692
rect 22017 2748 22081 2752
rect 22017 2692 22021 2748
rect 22021 2692 22077 2748
rect 22077 2692 22081 2748
rect 22017 2688 22081 2692
rect 22097 2748 22161 2752
rect 22097 2692 22101 2748
rect 22101 2692 22157 2748
rect 22157 2692 22161 2748
rect 22097 2688 22161 2692
rect 22177 2748 22241 2752
rect 22177 2692 22181 2748
rect 22181 2692 22237 2748
rect 22237 2692 22241 2748
rect 22177 2688 22241 2692
rect 30331 2748 30395 2752
rect 30331 2692 30335 2748
rect 30335 2692 30391 2748
rect 30391 2692 30395 2748
rect 30331 2688 30395 2692
rect 30411 2748 30475 2752
rect 30411 2692 30415 2748
rect 30415 2692 30471 2748
rect 30471 2692 30475 2748
rect 30411 2688 30475 2692
rect 30491 2748 30555 2752
rect 30491 2692 30495 2748
rect 30495 2692 30551 2748
rect 30551 2692 30555 2748
rect 30491 2688 30555 2692
rect 30571 2748 30635 2752
rect 30571 2692 30575 2748
rect 30575 2692 30631 2748
rect 30631 2692 30635 2748
rect 30571 2688 30635 2692
rect 9346 2204 9410 2208
rect 9346 2148 9350 2204
rect 9350 2148 9406 2204
rect 9406 2148 9410 2204
rect 9346 2144 9410 2148
rect 9426 2204 9490 2208
rect 9426 2148 9430 2204
rect 9430 2148 9486 2204
rect 9486 2148 9490 2204
rect 9426 2144 9490 2148
rect 9506 2204 9570 2208
rect 9506 2148 9510 2204
rect 9510 2148 9566 2204
rect 9566 2148 9570 2204
rect 9506 2144 9570 2148
rect 9586 2204 9650 2208
rect 9586 2148 9590 2204
rect 9590 2148 9646 2204
rect 9646 2148 9650 2204
rect 9586 2144 9650 2148
rect 17740 2204 17804 2208
rect 17740 2148 17744 2204
rect 17744 2148 17800 2204
rect 17800 2148 17804 2204
rect 17740 2144 17804 2148
rect 17820 2204 17884 2208
rect 17820 2148 17824 2204
rect 17824 2148 17880 2204
rect 17880 2148 17884 2204
rect 17820 2144 17884 2148
rect 17900 2204 17964 2208
rect 17900 2148 17904 2204
rect 17904 2148 17960 2204
rect 17960 2148 17964 2204
rect 17900 2144 17964 2148
rect 17980 2204 18044 2208
rect 17980 2148 17984 2204
rect 17984 2148 18040 2204
rect 18040 2148 18044 2204
rect 17980 2144 18044 2148
rect 26134 2204 26198 2208
rect 26134 2148 26138 2204
rect 26138 2148 26194 2204
rect 26194 2148 26198 2204
rect 26134 2144 26198 2148
rect 26214 2204 26278 2208
rect 26214 2148 26218 2204
rect 26218 2148 26274 2204
rect 26274 2148 26278 2204
rect 26214 2144 26278 2148
rect 26294 2204 26358 2208
rect 26294 2148 26298 2204
rect 26298 2148 26354 2204
rect 26354 2148 26358 2204
rect 26294 2144 26358 2148
rect 26374 2204 26438 2208
rect 26374 2148 26378 2204
rect 26378 2148 26434 2204
rect 26434 2148 26438 2204
rect 26374 2144 26438 2148
rect 34528 2204 34592 2208
rect 34528 2148 34532 2204
rect 34532 2148 34588 2204
rect 34588 2148 34592 2204
rect 34528 2144 34592 2148
rect 34608 2204 34672 2208
rect 34608 2148 34612 2204
rect 34612 2148 34668 2204
rect 34668 2148 34672 2204
rect 34608 2144 34672 2148
rect 34688 2204 34752 2208
rect 34688 2148 34692 2204
rect 34692 2148 34748 2204
rect 34748 2148 34752 2204
rect 34688 2144 34752 2148
rect 34768 2204 34832 2208
rect 34768 2148 34772 2204
rect 34772 2148 34828 2204
rect 34828 2148 34832 2204
rect 34768 2144 34832 2148
<< metal4 >>
rect 5141 35392 5461 35408
rect 5141 35328 5149 35392
rect 5213 35328 5229 35392
rect 5293 35328 5309 35392
rect 5373 35328 5389 35392
rect 5453 35328 5461 35392
rect 5141 34304 5461 35328
rect 5141 34240 5149 34304
rect 5213 34240 5229 34304
rect 5293 34240 5309 34304
rect 5373 34240 5389 34304
rect 5453 34240 5461 34304
rect 5141 33216 5461 34240
rect 5141 33152 5149 33216
rect 5213 33152 5229 33216
rect 5293 33152 5309 33216
rect 5373 33152 5389 33216
rect 5453 33152 5461 33216
rect 5141 32128 5461 33152
rect 5141 32064 5149 32128
rect 5213 32064 5229 32128
rect 5293 32064 5309 32128
rect 5373 32064 5389 32128
rect 5453 32064 5461 32128
rect 5141 31040 5461 32064
rect 5141 30976 5149 31040
rect 5213 30976 5229 31040
rect 5293 30976 5309 31040
rect 5373 30976 5389 31040
rect 5453 30976 5461 31040
rect 5141 29952 5461 30976
rect 5141 29888 5149 29952
rect 5213 29888 5229 29952
rect 5293 29888 5309 29952
rect 5373 29888 5389 29952
rect 5453 29888 5461 29952
rect 5141 28864 5461 29888
rect 5141 28800 5149 28864
rect 5213 28800 5229 28864
rect 5293 28800 5309 28864
rect 5373 28800 5389 28864
rect 5453 28800 5461 28864
rect 5141 27776 5461 28800
rect 5141 27712 5149 27776
rect 5213 27712 5229 27776
rect 5293 27712 5309 27776
rect 5373 27712 5389 27776
rect 5453 27712 5461 27776
rect 5141 26688 5461 27712
rect 5141 26624 5149 26688
rect 5213 26624 5229 26688
rect 5293 26624 5309 26688
rect 5373 26624 5389 26688
rect 5453 26624 5461 26688
rect 5141 25600 5461 26624
rect 5141 25536 5149 25600
rect 5213 25536 5229 25600
rect 5293 25536 5309 25600
rect 5373 25536 5389 25600
rect 5453 25536 5461 25600
rect 5141 24512 5461 25536
rect 5141 24448 5149 24512
rect 5213 24448 5229 24512
rect 5293 24448 5309 24512
rect 5373 24448 5389 24512
rect 5453 24448 5461 24512
rect 5141 23424 5461 24448
rect 5141 23360 5149 23424
rect 5213 23360 5229 23424
rect 5293 23360 5309 23424
rect 5373 23360 5389 23424
rect 5453 23360 5461 23424
rect 5141 22336 5461 23360
rect 5141 22272 5149 22336
rect 5213 22272 5229 22336
rect 5293 22272 5309 22336
rect 5373 22272 5389 22336
rect 5453 22272 5461 22336
rect 5141 21248 5461 22272
rect 5141 21184 5149 21248
rect 5213 21184 5229 21248
rect 5293 21184 5309 21248
rect 5373 21184 5389 21248
rect 5453 21184 5461 21248
rect 5141 20160 5461 21184
rect 5141 20096 5149 20160
rect 5213 20096 5229 20160
rect 5293 20096 5309 20160
rect 5373 20096 5389 20160
rect 5453 20096 5461 20160
rect 5141 19072 5461 20096
rect 5141 19008 5149 19072
rect 5213 19008 5229 19072
rect 5293 19008 5309 19072
rect 5373 19008 5389 19072
rect 5453 19008 5461 19072
rect 5141 17984 5461 19008
rect 5141 17920 5149 17984
rect 5213 17920 5229 17984
rect 5293 17920 5309 17984
rect 5373 17920 5389 17984
rect 5453 17920 5461 17984
rect 5141 16896 5461 17920
rect 9338 34848 9658 35408
rect 9338 34784 9346 34848
rect 9410 34784 9426 34848
rect 9490 34784 9506 34848
rect 9570 34784 9586 34848
rect 9650 34784 9658 34848
rect 9338 33760 9658 34784
rect 9338 33696 9346 33760
rect 9410 33696 9426 33760
rect 9490 33696 9506 33760
rect 9570 33696 9586 33760
rect 9650 33696 9658 33760
rect 9338 32672 9658 33696
rect 9338 32608 9346 32672
rect 9410 32608 9426 32672
rect 9490 32608 9506 32672
rect 9570 32608 9586 32672
rect 9650 32608 9658 32672
rect 9338 31584 9658 32608
rect 9338 31520 9346 31584
rect 9410 31520 9426 31584
rect 9490 31520 9506 31584
rect 9570 31520 9586 31584
rect 9650 31520 9658 31584
rect 9338 30496 9658 31520
rect 9338 30432 9346 30496
rect 9410 30432 9426 30496
rect 9490 30432 9506 30496
rect 9570 30432 9586 30496
rect 9650 30432 9658 30496
rect 9338 29408 9658 30432
rect 9338 29344 9346 29408
rect 9410 29344 9426 29408
rect 9490 29344 9506 29408
rect 9570 29344 9586 29408
rect 9650 29344 9658 29408
rect 9338 28320 9658 29344
rect 9338 28256 9346 28320
rect 9410 28256 9426 28320
rect 9490 28256 9506 28320
rect 9570 28256 9586 28320
rect 9650 28256 9658 28320
rect 9338 27232 9658 28256
rect 9338 27168 9346 27232
rect 9410 27168 9426 27232
rect 9490 27168 9506 27232
rect 9570 27168 9586 27232
rect 9650 27168 9658 27232
rect 9338 26144 9658 27168
rect 9338 26080 9346 26144
rect 9410 26080 9426 26144
rect 9490 26080 9506 26144
rect 9570 26080 9586 26144
rect 9650 26080 9658 26144
rect 9338 25056 9658 26080
rect 9338 24992 9346 25056
rect 9410 24992 9426 25056
rect 9490 24992 9506 25056
rect 9570 24992 9586 25056
rect 9650 24992 9658 25056
rect 9338 23968 9658 24992
rect 9338 23904 9346 23968
rect 9410 23904 9426 23968
rect 9490 23904 9506 23968
rect 9570 23904 9586 23968
rect 9650 23904 9658 23968
rect 9338 22880 9658 23904
rect 9338 22816 9346 22880
rect 9410 22816 9426 22880
rect 9490 22816 9506 22880
rect 9570 22816 9586 22880
rect 9650 22816 9658 22880
rect 9338 21792 9658 22816
rect 9338 21728 9346 21792
rect 9410 21728 9426 21792
rect 9490 21728 9506 21792
rect 9570 21728 9586 21792
rect 9650 21728 9658 21792
rect 9338 20704 9658 21728
rect 9338 20640 9346 20704
rect 9410 20640 9426 20704
rect 9490 20640 9506 20704
rect 9570 20640 9586 20704
rect 9650 20640 9658 20704
rect 9338 19616 9658 20640
rect 9338 19552 9346 19616
rect 9410 19552 9426 19616
rect 9490 19552 9506 19616
rect 9570 19552 9586 19616
rect 9650 19552 9658 19616
rect 9338 18528 9658 19552
rect 9338 18464 9346 18528
rect 9410 18464 9426 18528
rect 9490 18464 9506 18528
rect 9570 18464 9586 18528
rect 9650 18464 9658 18528
rect 9075 17780 9141 17781
rect 9075 17716 9076 17780
rect 9140 17716 9141 17780
rect 9075 17715 9141 17716
rect 5141 16832 5149 16896
rect 5213 16832 5229 16896
rect 5293 16832 5309 16896
rect 5373 16832 5389 16896
rect 5453 16832 5461 16896
rect 5141 15808 5461 16832
rect 8339 16420 8405 16421
rect 8339 16356 8340 16420
rect 8404 16356 8405 16420
rect 8339 16355 8405 16356
rect 8523 16420 8589 16421
rect 8523 16356 8524 16420
rect 8588 16356 8589 16420
rect 8523 16355 8589 16356
rect 5141 15744 5149 15808
rect 5213 15744 5229 15808
rect 5293 15744 5309 15808
rect 5373 15744 5389 15808
rect 5453 15744 5461 15808
rect 5141 14720 5461 15744
rect 5141 14656 5149 14720
rect 5213 14656 5229 14720
rect 5293 14656 5309 14720
rect 5373 14656 5389 14720
rect 5453 14656 5461 14720
rect 5141 13632 5461 14656
rect 5141 13568 5149 13632
rect 5213 13568 5229 13632
rect 5293 13568 5309 13632
rect 5373 13568 5389 13632
rect 5453 13568 5461 13632
rect 5141 12544 5461 13568
rect 8342 13429 8402 16355
rect 8526 14789 8586 16355
rect 9078 16013 9138 17715
rect 9338 17440 9658 18464
rect 9338 17376 9346 17440
rect 9410 17376 9426 17440
rect 9490 17376 9506 17440
rect 9570 17376 9586 17440
rect 9650 17376 9658 17440
rect 9338 16352 9658 17376
rect 9338 16288 9346 16352
rect 9410 16288 9426 16352
rect 9490 16288 9506 16352
rect 9570 16288 9586 16352
rect 9650 16288 9658 16352
rect 9075 16012 9141 16013
rect 9075 15948 9076 16012
rect 9140 15948 9141 16012
rect 9075 15947 9141 15948
rect 9338 15264 9658 16288
rect 9338 15200 9346 15264
rect 9410 15200 9426 15264
rect 9490 15200 9506 15264
rect 9570 15200 9586 15264
rect 9650 15200 9658 15264
rect 8523 14788 8589 14789
rect 8523 14724 8524 14788
rect 8588 14724 8589 14788
rect 8523 14723 8589 14724
rect 9338 14176 9658 15200
rect 9338 14112 9346 14176
rect 9410 14112 9426 14176
rect 9490 14112 9506 14176
rect 9570 14112 9586 14176
rect 9650 14112 9658 14176
rect 8339 13428 8405 13429
rect 8339 13364 8340 13428
rect 8404 13364 8405 13428
rect 8339 13363 8405 13364
rect 5141 12480 5149 12544
rect 5213 12480 5229 12544
rect 5293 12480 5309 12544
rect 5373 12480 5389 12544
rect 5453 12480 5461 12544
rect 5141 11456 5461 12480
rect 5141 11392 5149 11456
rect 5213 11392 5229 11456
rect 5293 11392 5309 11456
rect 5373 11392 5389 11456
rect 5453 11392 5461 11456
rect 5141 10368 5461 11392
rect 5141 10304 5149 10368
rect 5213 10304 5229 10368
rect 5293 10304 5309 10368
rect 5373 10304 5389 10368
rect 5453 10304 5461 10368
rect 5141 9280 5461 10304
rect 5141 9216 5149 9280
rect 5213 9216 5229 9280
rect 5293 9216 5309 9280
rect 5373 9216 5389 9280
rect 5453 9216 5461 9280
rect 5141 8192 5461 9216
rect 5141 8128 5149 8192
rect 5213 8128 5229 8192
rect 5293 8128 5309 8192
rect 5373 8128 5389 8192
rect 5453 8128 5461 8192
rect 5141 7104 5461 8128
rect 5141 7040 5149 7104
rect 5213 7040 5229 7104
rect 5293 7040 5309 7104
rect 5373 7040 5389 7104
rect 5453 7040 5461 7104
rect 5141 6016 5461 7040
rect 5141 5952 5149 6016
rect 5213 5952 5229 6016
rect 5293 5952 5309 6016
rect 5373 5952 5389 6016
rect 5453 5952 5461 6016
rect 5141 4928 5461 5952
rect 5141 4864 5149 4928
rect 5213 4864 5229 4928
rect 5293 4864 5309 4928
rect 5373 4864 5389 4928
rect 5453 4864 5461 4928
rect 5141 3840 5461 4864
rect 5141 3776 5149 3840
rect 5213 3776 5229 3840
rect 5293 3776 5309 3840
rect 5373 3776 5389 3840
rect 5453 3776 5461 3840
rect 5141 2752 5461 3776
rect 5141 2688 5149 2752
rect 5213 2688 5229 2752
rect 5293 2688 5309 2752
rect 5373 2688 5389 2752
rect 5453 2688 5461 2752
rect 5141 2128 5461 2688
rect 9338 13088 9658 14112
rect 9338 13024 9346 13088
rect 9410 13024 9426 13088
rect 9490 13024 9506 13088
rect 9570 13024 9586 13088
rect 9650 13024 9658 13088
rect 9338 12000 9658 13024
rect 9338 11936 9346 12000
rect 9410 11936 9426 12000
rect 9490 11936 9506 12000
rect 9570 11936 9586 12000
rect 9650 11936 9658 12000
rect 9338 10912 9658 11936
rect 9338 10848 9346 10912
rect 9410 10848 9426 10912
rect 9490 10848 9506 10912
rect 9570 10848 9586 10912
rect 9650 10848 9658 10912
rect 9338 9824 9658 10848
rect 9338 9760 9346 9824
rect 9410 9760 9426 9824
rect 9490 9760 9506 9824
rect 9570 9760 9586 9824
rect 9650 9760 9658 9824
rect 9338 8736 9658 9760
rect 9338 8672 9346 8736
rect 9410 8672 9426 8736
rect 9490 8672 9506 8736
rect 9570 8672 9586 8736
rect 9650 8672 9658 8736
rect 9338 7648 9658 8672
rect 9338 7584 9346 7648
rect 9410 7584 9426 7648
rect 9490 7584 9506 7648
rect 9570 7584 9586 7648
rect 9650 7584 9658 7648
rect 9338 6560 9658 7584
rect 9338 6496 9346 6560
rect 9410 6496 9426 6560
rect 9490 6496 9506 6560
rect 9570 6496 9586 6560
rect 9650 6496 9658 6560
rect 9338 5472 9658 6496
rect 9338 5408 9346 5472
rect 9410 5408 9426 5472
rect 9490 5408 9506 5472
rect 9570 5408 9586 5472
rect 9650 5408 9658 5472
rect 9338 4384 9658 5408
rect 9338 4320 9346 4384
rect 9410 4320 9426 4384
rect 9490 4320 9506 4384
rect 9570 4320 9586 4384
rect 9650 4320 9658 4384
rect 9338 3296 9658 4320
rect 9338 3232 9346 3296
rect 9410 3232 9426 3296
rect 9490 3232 9506 3296
rect 9570 3232 9586 3296
rect 9650 3232 9658 3296
rect 9338 2208 9658 3232
rect 9338 2144 9346 2208
rect 9410 2144 9426 2208
rect 9490 2144 9506 2208
rect 9570 2144 9586 2208
rect 9650 2144 9658 2208
rect 9338 2128 9658 2144
rect 13535 35392 13855 35408
rect 13535 35328 13543 35392
rect 13607 35328 13623 35392
rect 13687 35328 13703 35392
rect 13767 35328 13783 35392
rect 13847 35328 13855 35392
rect 13535 34304 13855 35328
rect 13535 34240 13543 34304
rect 13607 34240 13623 34304
rect 13687 34240 13703 34304
rect 13767 34240 13783 34304
rect 13847 34240 13855 34304
rect 13535 33216 13855 34240
rect 13535 33152 13543 33216
rect 13607 33152 13623 33216
rect 13687 33152 13703 33216
rect 13767 33152 13783 33216
rect 13847 33152 13855 33216
rect 13535 32128 13855 33152
rect 13535 32064 13543 32128
rect 13607 32064 13623 32128
rect 13687 32064 13703 32128
rect 13767 32064 13783 32128
rect 13847 32064 13855 32128
rect 13535 31040 13855 32064
rect 13535 30976 13543 31040
rect 13607 30976 13623 31040
rect 13687 30976 13703 31040
rect 13767 30976 13783 31040
rect 13847 30976 13855 31040
rect 13535 29952 13855 30976
rect 13535 29888 13543 29952
rect 13607 29888 13623 29952
rect 13687 29888 13703 29952
rect 13767 29888 13783 29952
rect 13847 29888 13855 29952
rect 13535 28864 13855 29888
rect 13535 28800 13543 28864
rect 13607 28800 13623 28864
rect 13687 28800 13703 28864
rect 13767 28800 13783 28864
rect 13847 28800 13855 28864
rect 13535 27776 13855 28800
rect 13535 27712 13543 27776
rect 13607 27712 13623 27776
rect 13687 27712 13703 27776
rect 13767 27712 13783 27776
rect 13847 27712 13855 27776
rect 13535 26688 13855 27712
rect 13535 26624 13543 26688
rect 13607 26624 13623 26688
rect 13687 26624 13703 26688
rect 13767 26624 13783 26688
rect 13847 26624 13855 26688
rect 13535 25600 13855 26624
rect 13535 25536 13543 25600
rect 13607 25536 13623 25600
rect 13687 25536 13703 25600
rect 13767 25536 13783 25600
rect 13847 25536 13855 25600
rect 13535 24512 13855 25536
rect 13535 24448 13543 24512
rect 13607 24448 13623 24512
rect 13687 24448 13703 24512
rect 13767 24448 13783 24512
rect 13847 24448 13855 24512
rect 13535 23424 13855 24448
rect 13535 23360 13543 23424
rect 13607 23360 13623 23424
rect 13687 23360 13703 23424
rect 13767 23360 13783 23424
rect 13847 23360 13855 23424
rect 13535 22336 13855 23360
rect 13535 22272 13543 22336
rect 13607 22272 13623 22336
rect 13687 22272 13703 22336
rect 13767 22272 13783 22336
rect 13847 22272 13855 22336
rect 13535 21248 13855 22272
rect 13535 21184 13543 21248
rect 13607 21184 13623 21248
rect 13687 21184 13703 21248
rect 13767 21184 13783 21248
rect 13847 21184 13855 21248
rect 13535 20160 13855 21184
rect 13535 20096 13543 20160
rect 13607 20096 13623 20160
rect 13687 20096 13703 20160
rect 13767 20096 13783 20160
rect 13847 20096 13855 20160
rect 13535 19072 13855 20096
rect 13535 19008 13543 19072
rect 13607 19008 13623 19072
rect 13687 19008 13703 19072
rect 13767 19008 13783 19072
rect 13847 19008 13855 19072
rect 13535 17984 13855 19008
rect 13535 17920 13543 17984
rect 13607 17920 13623 17984
rect 13687 17920 13703 17984
rect 13767 17920 13783 17984
rect 13847 17920 13855 17984
rect 13535 16896 13855 17920
rect 13535 16832 13543 16896
rect 13607 16832 13623 16896
rect 13687 16832 13703 16896
rect 13767 16832 13783 16896
rect 13847 16832 13855 16896
rect 13535 15808 13855 16832
rect 13535 15744 13543 15808
rect 13607 15744 13623 15808
rect 13687 15744 13703 15808
rect 13767 15744 13783 15808
rect 13847 15744 13855 15808
rect 13535 14720 13855 15744
rect 13535 14656 13543 14720
rect 13607 14656 13623 14720
rect 13687 14656 13703 14720
rect 13767 14656 13783 14720
rect 13847 14656 13855 14720
rect 13535 13632 13855 14656
rect 13535 13568 13543 13632
rect 13607 13568 13623 13632
rect 13687 13568 13703 13632
rect 13767 13568 13783 13632
rect 13847 13568 13855 13632
rect 13535 12544 13855 13568
rect 13535 12480 13543 12544
rect 13607 12480 13623 12544
rect 13687 12480 13703 12544
rect 13767 12480 13783 12544
rect 13847 12480 13855 12544
rect 13535 11456 13855 12480
rect 13535 11392 13543 11456
rect 13607 11392 13623 11456
rect 13687 11392 13703 11456
rect 13767 11392 13783 11456
rect 13847 11392 13855 11456
rect 13535 10368 13855 11392
rect 13535 10304 13543 10368
rect 13607 10304 13623 10368
rect 13687 10304 13703 10368
rect 13767 10304 13783 10368
rect 13847 10304 13855 10368
rect 13535 9280 13855 10304
rect 13535 9216 13543 9280
rect 13607 9216 13623 9280
rect 13687 9216 13703 9280
rect 13767 9216 13783 9280
rect 13847 9216 13855 9280
rect 13535 8192 13855 9216
rect 13535 8128 13543 8192
rect 13607 8128 13623 8192
rect 13687 8128 13703 8192
rect 13767 8128 13783 8192
rect 13847 8128 13855 8192
rect 13535 7104 13855 8128
rect 13535 7040 13543 7104
rect 13607 7040 13623 7104
rect 13687 7040 13703 7104
rect 13767 7040 13783 7104
rect 13847 7040 13855 7104
rect 13535 6016 13855 7040
rect 13535 5952 13543 6016
rect 13607 5952 13623 6016
rect 13687 5952 13703 6016
rect 13767 5952 13783 6016
rect 13847 5952 13855 6016
rect 13535 4928 13855 5952
rect 13535 4864 13543 4928
rect 13607 4864 13623 4928
rect 13687 4864 13703 4928
rect 13767 4864 13783 4928
rect 13847 4864 13855 4928
rect 13535 3840 13855 4864
rect 13535 3776 13543 3840
rect 13607 3776 13623 3840
rect 13687 3776 13703 3840
rect 13767 3776 13783 3840
rect 13847 3776 13855 3840
rect 13535 2752 13855 3776
rect 13535 2688 13543 2752
rect 13607 2688 13623 2752
rect 13687 2688 13703 2752
rect 13767 2688 13783 2752
rect 13847 2688 13855 2752
rect 13535 2128 13855 2688
rect 17732 34848 18052 35408
rect 17732 34784 17740 34848
rect 17804 34784 17820 34848
rect 17884 34784 17900 34848
rect 17964 34784 17980 34848
rect 18044 34784 18052 34848
rect 17732 33760 18052 34784
rect 17732 33696 17740 33760
rect 17804 33696 17820 33760
rect 17884 33696 17900 33760
rect 17964 33696 17980 33760
rect 18044 33696 18052 33760
rect 17732 32672 18052 33696
rect 17732 32608 17740 32672
rect 17804 32608 17820 32672
rect 17884 32608 17900 32672
rect 17964 32608 17980 32672
rect 18044 32608 18052 32672
rect 17732 31584 18052 32608
rect 17732 31520 17740 31584
rect 17804 31520 17820 31584
rect 17884 31520 17900 31584
rect 17964 31520 17980 31584
rect 18044 31520 18052 31584
rect 17732 30496 18052 31520
rect 17732 30432 17740 30496
rect 17804 30432 17820 30496
rect 17884 30432 17900 30496
rect 17964 30432 17980 30496
rect 18044 30432 18052 30496
rect 17732 29408 18052 30432
rect 17732 29344 17740 29408
rect 17804 29344 17820 29408
rect 17884 29344 17900 29408
rect 17964 29344 17980 29408
rect 18044 29344 18052 29408
rect 17732 28320 18052 29344
rect 17732 28256 17740 28320
rect 17804 28256 17820 28320
rect 17884 28256 17900 28320
rect 17964 28256 17980 28320
rect 18044 28256 18052 28320
rect 17732 27232 18052 28256
rect 17732 27168 17740 27232
rect 17804 27168 17820 27232
rect 17884 27168 17900 27232
rect 17964 27168 17980 27232
rect 18044 27168 18052 27232
rect 17732 26144 18052 27168
rect 17732 26080 17740 26144
rect 17804 26080 17820 26144
rect 17884 26080 17900 26144
rect 17964 26080 17980 26144
rect 18044 26080 18052 26144
rect 17732 25056 18052 26080
rect 17732 24992 17740 25056
rect 17804 24992 17820 25056
rect 17884 24992 17900 25056
rect 17964 24992 17980 25056
rect 18044 24992 18052 25056
rect 17732 23968 18052 24992
rect 17732 23904 17740 23968
rect 17804 23904 17820 23968
rect 17884 23904 17900 23968
rect 17964 23904 17980 23968
rect 18044 23904 18052 23968
rect 17732 22880 18052 23904
rect 17732 22816 17740 22880
rect 17804 22816 17820 22880
rect 17884 22816 17900 22880
rect 17964 22816 17980 22880
rect 18044 22816 18052 22880
rect 17732 21792 18052 22816
rect 17732 21728 17740 21792
rect 17804 21728 17820 21792
rect 17884 21728 17900 21792
rect 17964 21728 17980 21792
rect 18044 21728 18052 21792
rect 17732 20704 18052 21728
rect 17732 20640 17740 20704
rect 17804 20640 17820 20704
rect 17884 20640 17900 20704
rect 17964 20640 17980 20704
rect 18044 20640 18052 20704
rect 17732 19616 18052 20640
rect 17732 19552 17740 19616
rect 17804 19552 17820 19616
rect 17884 19552 17900 19616
rect 17964 19552 17980 19616
rect 18044 19552 18052 19616
rect 17732 18528 18052 19552
rect 17732 18464 17740 18528
rect 17804 18464 17820 18528
rect 17884 18464 17900 18528
rect 17964 18464 17980 18528
rect 18044 18464 18052 18528
rect 17732 17440 18052 18464
rect 17732 17376 17740 17440
rect 17804 17376 17820 17440
rect 17884 17376 17900 17440
rect 17964 17376 17980 17440
rect 18044 17376 18052 17440
rect 17732 16352 18052 17376
rect 17732 16288 17740 16352
rect 17804 16288 17820 16352
rect 17884 16288 17900 16352
rect 17964 16288 17980 16352
rect 18044 16288 18052 16352
rect 17732 15264 18052 16288
rect 17732 15200 17740 15264
rect 17804 15200 17820 15264
rect 17884 15200 17900 15264
rect 17964 15200 17980 15264
rect 18044 15200 18052 15264
rect 17732 14176 18052 15200
rect 17732 14112 17740 14176
rect 17804 14112 17820 14176
rect 17884 14112 17900 14176
rect 17964 14112 17980 14176
rect 18044 14112 18052 14176
rect 17732 13088 18052 14112
rect 17732 13024 17740 13088
rect 17804 13024 17820 13088
rect 17884 13024 17900 13088
rect 17964 13024 17980 13088
rect 18044 13024 18052 13088
rect 17732 12000 18052 13024
rect 17732 11936 17740 12000
rect 17804 11936 17820 12000
rect 17884 11936 17900 12000
rect 17964 11936 17980 12000
rect 18044 11936 18052 12000
rect 17732 10912 18052 11936
rect 17732 10848 17740 10912
rect 17804 10848 17820 10912
rect 17884 10848 17900 10912
rect 17964 10848 17980 10912
rect 18044 10848 18052 10912
rect 17732 9824 18052 10848
rect 17732 9760 17740 9824
rect 17804 9760 17820 9824
rect 17884 9760 17900 9824
rect 17964 9760 17980 9824
rect 18044 9760 18052 9824
rect 17732 8736 18052 9760
rect 17732 8672 17740 8736
rect 17804 8672 17820 8736
rect 17884 8672 17900 8736
rect 17964 8672 17980 8736
rect 18044 8672 18052 8736
rect 17732 7648 18052 8672
rect 17732 7584 17740 7648
rect 17804 7584 17820 7648
rect 17884 7584 17900 7648
rect 17964 7584 17980 7648
rect 18044 7584 18052 7648
rect 17732 6560 18052 7584
rect 17732 6496 17740 6560
rect 17804 6496 17820 6560
rect 17884 6496 17900 6560
rect 17964 6496 17980 6560
rect 18044 6496 18052 6560
rect 17732 5472 18052 6496
rect 17732 5408 17740 5472
rect 17804 5408 17820 5472
rect 17884 5408 17900 5472
rect 17964 5408 17980 5472
rect 18044 5408 18052 5472
rect 17732 4384 18052 5408
rect 17732 4320 17740 4384
rect 17804 4320 17820 4384
rect 17884 4320 17900 4384
rect 17964 4320 17980 4384
rect 18044 4320 18052 4384
rect 17732 3296 18052 4320
rect 17732 3232 17740 3296
rect 17804 3232 17820 3296
rect 17884 3232 17900 3296
rect 17964 3232 17980 3296
rect 18044 3232 18052 3296
rect 17732 2208 18052 3232
rect 17732 2144 17740 2208
rect 17804 2144 17820 2208
rect 17884 2144 17900 2208
rect 17964 2144 17980 2208
rect 18044 2144 18052 2208
rect 17732 2128 18052 2144
rect 21929 35392 22249 35408
rect 21929 35328 21937 35392
rect 22001 35328 22017 35392
rect 22081 35328 22097 35392
rect 22161 35328 22177 35392
rect 22241 35328 22249 35392
rect 21929 34304 22249 35328
rect 21929 34240 21937 34304
rect 22001 34240 22017 34304
rect 22081 34240 22097 34304
rect 22161 34240 22177 34304
rect 22241 34240 22249 34304
rect 21929 33216 22249 34240
rect 21929 33152 21937 33216
rect 22001 33152 22017 33216
rect 22081 33152 22097 33216
rect 22161 33152 22177 33216
rect 22241 33152 22249 33216
rect 21929 32128 22249 33152
rect 21929 32064 21937 32128
rect 22001 32064 22017 32128
rect 22081 32064 22097 32128
rect 22161 32064 22177 32128
rect 22241 32064 22249 32128
rect 21929 31040 22249 32064
rect 21929 30976 21937 31040
rect 22001 30976 22017 31040
rect 22081 30976 22097 31040
rect 22161 30976 22177 31040
rect 22241 30976 22249 31040
rect 21929 29952 22249 30976
rect 21929 29888 21937 29952
rect 22001 29888 22017 29952
rect 22081 29888 22097 29952
rect 22161 29888 22177 29952
rect 22241 29888 22249 29952
rect 21929 28864 22249 29888
rect 21929 28800 21937 28864
rect 22001 28800 22017 28864
rect 22081 28800 22097 28864
rect 22161 28800 22177 28864
rect 22241 28800 22249 28864
rect 21929 27776 22249 28800
rect 21929 27712 21937 27776
rect 22001 27712 22017 27776
rect 22081 27712 22097 27776
rect 22161 27712 22177 27776
rect 22241 27712 22249 27776
rect 21929 26688 22249 27712
rect 21929 26624 21937 26688
rect 22001 26624 22017 26688
rect 22081 26624 22097 26688
rect 22161 26624 22177 26688
rect 22241 26624 22249 26688
rect 21929 25600 22249 26624
rect 21929 25536 21937 25600
rect 22001 25536 22017 25600
rect 22081 25536 22097 25600
rect 22161 25536 22177 25600
rect 22241 25536 22249 25600
rect 21929 24512 22249 25536
rect 21929 24448 21937 24512
rect 22001 24448 22017 24512
rect 22081 24448 22097 24512
rect 22161 24448 22177 24512
rect 22241 24448 22249 24512
rect 21929 23424 22249 24448
rect 21929 23360 21937 23424
rect 22001 23360 22017 23424
rect 22081 23360 22097 23424
rect 22161 23360 22177 23424
rect 22241 23360 22249 23424
rect 21929 22336 22249 23360
rect 21929 22272 21937 22336
rect 22001 22272 22017 22336
rect 22081 22272 22097 22336
rect 22161 22272 22177 22336
rect 22241 22272 22249 22336
rect 21929 21248 22249 22272
rect 21929 21184 21937 21248
rect 22001 21184 22017 21248
rect 22081 21184 22097 21248
rect 22161 21184 22177 21248
rect 22241 21184 22249 21248
rect 21929 20160 22249 21184
rect 21929 20096 21937 20160
rect 22001 20096 22017 20160
rect 22081 20096 22097 20160
rect 22161 20096 22177 20160
rect 22241 20096 22249 20160
rect 21929 19072 22249 20096
rect 21929 19008 21937 19072
rect 22001 19008 22017 19072
rect 22081 19008 22097 19072
rect 22161 19008 22177 19072
rect 22241 19008 22249 19072
rect 21929 17984 22249 19008
rect 21929 17920 21937 17984
rect 22001 17920 22017 17984
rect 22081 17920 22097 17984
rect 22161 17920 22177 17984
rect 22241 17920 22249 17984
rect 21929 16896 22249 17920
rect 21929 16832 21937 16896
rect 22001 16832 22017 16896
rect 22081 16832 22097 16896
rect 22161 16832 22177 16896
rect 22241 16832 22249 16896
rect 21929 15808 22249 16832
rect 21929 15744 21937 15808
rect 22001 15744 22017 15808
rect 22081 15744 22097 15808
rect 22161 15744 22177 15808
rect 22241 15744 22249 15808
rect 21929 14720 22249 15744
rect 21929 14656 21937 14720
rect 22001 14656 22017 14720
rect 22081 14656 22097 14720
rect 22161 14656 22177 14720
rect 22241 14656 22249 14720
rect 21929 13632 22249 14656
rect 21929 13568 21937 13632
rect 22001 13568 22017 13632
rect 22081 13568 22097 13632
rect 22161 13568 22177 13632
rect 22241 13568 22249 13632
rect 21929 12544 22249 13568
rect 21929 12480 21937 12544
rect 22001 12480 22017 12544
rect 22081 12480 22097 12544
rect 22161 12480 22177 12544
rect 22241 12480 22249 12544
rect 21929 11456 22249 12480
rect 21929 11392 21937 11456
rect 22001 11392 22017 11456
rect 22081 11392 22097 11456
rect 22161 11392 22177 11456
rect 22241 11392 22249 11456
rect 21929 10368 22249 11392
rect 21929 10304 21937 10368
rect 22001 10304 22017 10368
rect 22081 10304 22097 10368
rect 22161 10304 22177 10368
rect 22241 10304 22249 10368
rect 21929 9280 22249 10304
rect 21929 9216 21937 9280
rect 22001 9216 22017 9280
rect 22081 9216 22097 9280
rect 22161 9216 22177 9280
rect 22241 9216 22249 9280
rect 21929 8192 22249 9216
rect 21929 8128 21937 8192
rect 22001 8128 22017 8192
rect 22081 8128 22097 8192
rect 22161 8128 22177 8192
rect 22241 8128 22249 8192
rect 21929 7104 22249 8128
rect 21929 7040 21937 7104
rect 22001 7040 22017 7104
rect 22081 7040 22097 7104
rect 22161 7040 22177 7104
rect 22241 7040 22249 7104
rect 21929 6016 22249 7040
rect 21929 5952 21937 6016
rect 22001 5952 22017 6016
rect 22081 5952 22097 6016
rect 22161 5952 22177 6016
rect 22241 5952 22249 6016
rect 21929 4928 22249 5952
rect 21929 4864 21937 4928
rect 22001 4864 22017 4928
rect 22081 4864 22097 4928
rect 22161 4864 22177 4928
rect 22241 4864 22249 4928
rect 21929 3840 22249 4864
rect 21929 3776 21937 3840
rect 22001 3776 22017 3840
rect 22081 3776 22097 3840
rect 22161 3776 22177 3840
rect 22241 3776 22249 3840
rect 21929 2752 22249 3776
rect 21929 2688 21937 2752
rect 22001 2688 22017 2752
rect 22081 2688 22097 2752
rect 22161 2688 22177 2752
rect 22241 2688 22249 2752
rect 21929 2128 22249 2688
rect 26126 34848 26446 35408
rect 26126 34784 26134 34848
rect 26198 34784 26214 34848
rect 26278 34784 26294 34848
rect 26358 34784 26374 34848
rect 26438 34784 26446 34848
rect 26126 33760 26446 34784
rect 26126 33696 26134 33760
rect 26198 33696 26214 33760
rect 26278 33696 26294 33760
rect 26358 33696 26374 33760
rect 26438 33696 26446 33760
rect 26126 32672 26446 33696
rect 26126 32608 26134 32672
rect 26198 32608 26214 32672
rect 26278 32608 26294 32672
rect 26358 32608 26374 32672
rect 26438 32608 26446 32672
rect 26126 31584 26446 32608
rect 26126 31520 26134 31584
rect 26198 31520 26214 31584
rect 26278 31520 26294 31584
rect 26358 31520 26374 31584
rect 26438 31520 26446 31584
rect 26126 30496 26446 31520
rect 26126 30432 26134 30496
rect 26198 30432 26214 30496
rect 26278 30432 26294 30496
rect 26358 30432 26374 30496
rect 26438 30432 26446 30496
rect 26126 29408 26446 30432
rect 26126 29344 26134 29408
rect 26198 29344 26214 29408
rect 26278 29344 26294 29408
rect 26358 29344 26374 29408
rect 26438 29344 26446 29408
rect 26126 28320 26446 29344
rect 26126 28256 26134 28320
rect 26198 28256 26214 28320
rect 26278 28256 26294 28320
rect 26358 28256 26374 28320
rect 26438 28256 26446 28320
rect 26126 27232 26446 28256
rect 26126 27168 26134 27232
rect 26198 27168 26214 27232
rect 26278 27168 26294 27232
rect 26358 27168 26374 27232
rect 26438 27168 26446 27232
rect 26126 26144 26446 27168
rect 26126 26080 26134 26144
rect 26198 26080 26214 26144
rect 26278 26080 26294 26144
rect 26358 26080 26374 26144
rect 26438 26080 26446 26144
rect 26126 25056 26446 26080
rect 26126 24992 26134 25056
rect 26198 24992 26214 25056
rect 26278 24992 26294 25056
rect 26358 24992 26374 25056
rect 26438 24992 26446 25056
rect 26126 23968 26446 24992
rect 26126 23904 26134 23968
rect 26198 23904 26214 23968
rect 26278 23904 26294 23968
rect 26358 23904 26374 23968
rect 26438 23904 26446 23968
rect 26126 22880 26446 23904
rect 26126 22816 26134 22880
rect 26198 22816 26214 22880
rect 26278 22816 26294 22880
rect 26358 22816 26374 22880
rect 26438 22816 26446 22880
rect 26126 21792 26446 22816
rect 26126 21728 26134 21792
rect 26198 21728 26214 21792
rect 26278 21728 26294 21792
rect 26358 21728 26374 21792
rect 26438 21728 26446 21792
rect 26126 20704 26446 21728
rect 26126 20640 26134 20704
rect 26198 20640 26214 20704
rect 26278 20640 26294 20704
rect 26358 20640 26374 20704
rect 26438 20640 26446 20704
rect 26126 19616 26446 20640
rect 26126 19552 26134 19616
rect 26198 19552 26214 19616
rect 26278 19552 26294 19616
rect 26358 19552 26374 19616
rect 26438 19552 26446 19616
rect 26126 18528 26446 19552
rect 26126 18464 26134 18528
rect 26198 18464 26214 18528
rect 26278 18464 26294 18528
rect 26358 18464 26374 18528
rect 26438 18464 26446 18528
rect 26126 17440 26446 18464
rect 26126 17376 26134 17440
rect 26198 17376 26214 17440
rect 26278 17376 26294 17440
rect 26358 17376 26374 17440
rect 26438 17376 26446 17440
rect 26126 16352 26446 17376
rect 26126 16288 26134 16352
rect 26198 16288 26214 16352
rect 26278 16288 26294 16352
rect 26358 16288 26374 16352
rect 26438 16288 26446 16352
rect 26126 15264 26446 16288
rect 26126 15200 26134 15264
rect 26198 15200 26214 15264
rect 26278 15200 26294 15264
rect 26358 15200 26374 15264
rect 26438 15200 26446 15264
rect 26126 14176 26446 15200
rect 26126 14112 26134 14176
rect 26198 14112 26214 14176
rect 26278 14112 26294 14176
rect 26358 14112 26374 14176
rect 26438 14112 26446 14176
rect 26126 13088 26446 14112
rect 26126 13024 26134 13088
rect 26198 13024 26214 13088
rect 26278 13024 26294 13088
rect 26358 13024 26374 13088
rect 26438 13024 26446 13088
rect 26126 12000 26446 13024
rect 26126 11936 26134 12000
rect 26198 11936 26214 12000
rect 26278 11936 26294 12000
rect 26358 11936 26374 12000
rect 26438 11936 26446 12000
rect 26126 10912 26446 11936
rect 26126 10848 26134 10912
rect 26198 10848 26214 10912
rect 26278 10848 26294 10912
rect 26358 10848 26374 10912
rect 26438 10848 26446 10912
rect 26126 9824 26446 10848
rect 26126 9760 26134 9824
rect 26198 9760 26214 9824
rect 26278 9760 26294 9824
rect 26358 9760 26374 9824
rect 26438 9760 26446 9824
rect 26126 8736 26446 9760
rect 26126 8672 26134 8736
rect 26198 8672 26214 8736
rect 26278 8672 26294 8736
rect 26358 8672 26374 8736
rect 26438 8672 26446 8736
rect 26126 7648 26446 8672
rect 26126 7584 26134 7648
rect 26198 7584 26214 7648
rect 26278 7584 26294 7648
rect 26358 7584 26374 7648
rect 26438 7584 26446 7648
rect 26126 6560 26446 7584
rect 26126 6496 26134 6560
rect 26198 6496 26214 6560
rect 26278 6496 26294 6560
rect 26358 6496 26374 6560
rect 26438 6496 26446 6560
rect 26126 5472 26446 6496
rect 26126 5408 26134 5472
rect 26198 5408 26214 5472
rect 26278 5408 26294 5472
rect 26358 5408 26374 5472
rect 26438 5408 26446 5472
rect 26126 4384 26446 5408
rect 26126 4320 26134 4384
rect 26198 4320 26214 4384
rect 26278 4320 26294 4384
rect 26358 4320 26374 4384
rect 26438 4320 26446 4384
rect 26126 3296 26446 4320
rect 26126 3232 26134 3296
rect 26198 3232 26214 3296
rect 26278 3232 26294 3296
rect 26358 3232 26374 3296
rect 26438 3232 26446 3296
rect 26126 2208 26446 3232
rect 26126 2144 26134 2208
rect 26198 2144 26214 2208
rect 26278 2144 26294 2208
rect 26358 2144 26374 2208
rect 26438 2144 26446 2208
rect 26126 2128 26446 2144
rect 30323 35392 30643 35408
rect 30323 35328 30331 35392
rect 30395 35328 30411 35392
rect 30475 35328 30491 35392
rect 30555 35328 30571 35392
rect 30635 35328 30643 35392
rect 30323 34304 30643 35328
rect 30323 34240 30331 34304
rect 30395 34240 30411 34304
rect 30475 34240 30491 34304
rect 30555 34240 30571 34304
rect 30635 34240 30643 34304
rect 30323 33216 30643 34240
rect 30323 33152 30331 33216
rect 30395 33152 30411 33216
rect 30475 33152 30491 33216
rect 30555 33152 30571 33216
rect 30635 33152 30643 33216
rect 30323 32128 30643 33152
rect 30323 32064 30331 32128
rect 30395 32064 30411 32128
rect 30475 32064 30491 32128
rect 30555 32064 30571 32128
rect 30635 32064 30643 32128
rect 30323 31040 30643 32064
rect 30323 30976 30331 31040
rect 30395 30976 30411 31040
rect 30475 30976 30491 31040
rect 30555 30976 30571 31040
rect 30635 30976 30643 31040
rect 30323 29952 30643 30976
rect 30323 29888 30331 29952
rect 30395 29888 30411 29952
rect 30475 29888 30491 29952
rect 30555 29888 30571 29952
rect 30635 29888 30643 29952
rect 30323 28864 30643 29888
rect 30323 28800 30331 28864
rect 30395 28800 30411 28864
rect 30475 28800 30491 28864
rect 30555 28800 30571 28864
rect 30635 28800 30643 28864
rect 30323 27776 30643 28800
rect 30323 27712 30331 27776
rect 30395 27712 30411 27776
rect 30475 27712 30491 27776
rect 30555 27712 30571 27776
rect 30635 27712 30643 27776
rect 30323 26688 30643 27712
rect 30323 26624 30331 26688
rect 30395 26624 30411 26688
rect 30475 26624 30491 26688
rect 30555 26624 30571 26688
rect 30635 26624 30643 26688
rect 30323 25600 30643 26624
rect 30323 25536 30331 25600
rect 30395 25536 30411 25600
rect 30475 25536 30491 25600
rect 30555 25536 30571 25600
rect 30635 25536 30643 25600
rect 30323 24512 30643 25536
rect 30323 24448 30331 24512
rect 30395 24448 30411 24512
rect 30475 24448 30491 24512
rect 30555 24448 30571 24512
rect 30635 24448 30643 24512
rect 30323 23424 30643 24448
rect 30323 23360 30331 23424
rect 30395 23360 30411 23424
rect 30475 23360 30491 23424
rect 30555 23360 30571 23424
rect 30635 23360 30643 23424
rect 30323 22336 30643 23360
rect 30323 22272 30331 22336
rect 30395 22272 30411 22336
rect 30475 22272 30491 22336
rect 30555 22272 30571 22336
rect 30635 22272 30643 22336
rect 30323 21248 30643 22272
rect 30323 21184 30331 21248
rect 30395 21184 30411 21248
rect 30475 21184 30491 21248
rect 30555 21184 30571 21248
rect 30635 21184 30643 21248
rect 30323 20160 30643 21184
rect 30323 20096 30331 20160
rect 30395 20096 30411 20160
rect 30475 20096 30491 20160
rect 30555 20096 30571 20160
rect 30635 20096 30643 20160
rect 30323 19072 30643 20096
rect 30323 19008 30331 19072
rect 30395 19008 30411 19072
rect 30475 19008 30491 19072
rect 30555 19008 30571 19072
rect 30635 19008 30643 19072
rect 30323 17984 30643 19008
rect 30323 17920 30331 17984
rect 30395 17920 30411 17984
rect 30475 17920 30491 17984
rect 30555 17920 30571 17984
rect 30635 17920 30643 17984
rect 30323 16896 30643 17920
rect 30323 16832 30331 16896
rect 30395 16832 30411 16896
rect 30475 16832 30491 16896
rect 30555 16832 30571 16896
rect 30635 16832 30643 16896
rect 30323 15808 30643 16832
rect 30323 15744 30331 15808
rect 30395 15744 30411 15808
rect 30475 15744 30491 15808
rect 30555 15744 30571 15808
rect 30635 15744 30643 15808
rect 30323 14720 30643 15744
rect 30323 14656 30331 14720
rect 30395 14656 30411 14720
rect 30475 14656 30491 14720
rect 30555 14656 30571 14720
rect 30635 14656 30643 14720
rect 30323 13632 30643 14656
rect 30323 13568 30331 13632
rect 30395 13568 30411 13632
rect 30475 13568 30491 13632
rect 30555 13568 30571 13632
rect 30635 13568 30643 13632
rect 30323 12544 30643 13568
rect 30323 12480 30331 12544
rect 30395 12480 30411 12544
rect 30475 12480 30491 12544
rect 30555 12480 30571 12544
rect 30635 12480 30643 12544
rect 30323 11456 30643 12480
rect 30323 11392 30331 11456
rect 30395 11392 30411 11456
rect 30475 11392 30491 11456
rect 30555 11392 30571 11456
rect 30635 11392 30643 11456
rect 30323 10368 30643 11392
rect 30323 10304 30331 10368
rect 30395 10304 30411 10368
rect 30475 10304 30491 10368
rect 30555 10304 30571 10368
rect 30635 10304 30643 10368
rect 30323 9280 30643 10304
rect 30323 9216 30331 9280
rect 30395 9216 30411 9280
rect 30475 9216 30491 9280
rect 30555 9216 30571 9280
rect 30635 9216 30643 9280
rect 30323 8192 30643 9216
rect 30323 8128 30331 8192
rect 30395 8128 30411 8192
rect 30475 8128 30491 8192
rect 30555 8128 30571 8192
rect 30635 8128 30643 8192
rect 30323 7104 30643 8128
rect 30323 7040 30331 7104
rect 30395 7040 30411 7104
rect 30475 7040 30491 7104
rect 30555 7040 30571 7104
rect 30635 7040 30643 7104
rect 30323 6016 30643 7040
rect 30323 5952 30331 6016
rect 30395 5952 30411 6016
rect 30475 5952 30491 6016
rect 30555 5952 30571 6016
rect 30635 5952 30643 6016
rect 30323 4928 30643 5952
rect 30323 4864 30331 4928
rect 30395 4864 30411 4928
rect 30475 4864 30491 4928
rect 30555 4864 30571 4928
rect 30635 4864 30643 4928
rect 30323 3840 30643 4864
rect 30323 3776 30331 3840
rect 30395 3776 30411 3840
rect 30475 3776 30491 3840
rect 30555 3776 30571 3840
rect 30635 3776 30643 3840
rect 30323 2752 30643 3776
rect 30323 2688 30331 2752
rect 30395 2688 30411 2752
rect 30475 2688 30491 2752
rect 30555 2688 30571 2752
rect 30635 2688 30643 2752
rect 30323 2128 30643 2688
rect 34520 34848 34840 35408
rect 34520 34784 34528 34848
rect 34592 34784 34608 34848
rect 34672 34784 34688 34848
rect 34752 34784 34768 34848
rect 34832 34784 34840 34848
rect 34520 33760 34840 34784
rect 34520 33696 34528 33760
rect 34592 33696 34608 33760
rect 34672 33696 34688 33760
rect 34752 33696 34768 33760
rect 34832 33696 34840 33760
rect 34520 32672 34840 33696
rect 34520 32608 34528 32672
rect 34592 32608 34608 32672
rect 34672 32608 34688 32672
rect 34752 32608 34768 32672
rect 34832 32608 34840 32672
rect 34520 31584 34840 32608
rect 34520 31520 34528 31584
rect 34592 31520 34608 31584
rect 34672 31520 34688 31584
rect 34752 31520 34768 31584
rect 34832 31520 34840 31584
rect 34520 30496 34840 31520
rect 34520 30432 34528 30496
rect 34592 30432 34608 30496
rect 34672 30432 34688 30496
rect 34752 30432 34768 30496
rect 34832 30432 34840 30496
rect 34520 29408 34840 30432
rect 34520 29344 34528 29408
rect 34592 29344 34608 29408
rect 34672 29344 34688 29408
rect 34752 29344 34768 29408
rect 34832 29344 34840 29408
rect 34520 28320 34840 29344
rect 34520 28256 34528 28320
rect 34592 28256 34608 28320
rect 34672 28256 34688 28320
rect 34752 28256 34768 28320
rect 34832 28256 34840 28320
rect 34520 27232 34840 28256
rect 34520 27168 34528 27232
rect 34592 27168 34608 27232
rect 34672 27168 34688 27232
rect 34752 27168 34768 27232
rect 34832 27168 34840 27232
rect 34520 26144 34840 27168
rect 34520 26080 34528 26144
rect 34592 26080 34608 26144
rect 34672 26080 34688 26144
rect 34752 26080 34768 26144
rect 34832 26080 34840 26144
rect 34520 25056 34840 26080
rect 34520 24992 34528 25056
rect 34592 24992 34608 25056
rect 34672 24992 34688 25056
rect 34752 24992 34768 25056
rect 34832 24992 34840 25056
rect 34520 23968 34840 24992
rect 34520 23904 34528 23968
rect 34592 23904 34608 23968
rect 34672 23904 34688 23968
rect 34752 23904 34768 23968
rect 34832 23904 34840 23968
rect 34520 22880 34840 23904
rect 34520 22816 34528 22880
rect 34592 22816 34608 22880
rect 34672 22816 34688 22880
rect 34752 22816 34768 22880
rect 34832 22816 34840 22880
rect 34520 21792 34840 22816
rect 34520 21728 34528 21792
rect 34592 21728 34608 21792
rect 34672 21728 34688 21792
rect 34752 21728 34768 21792
rect 34832 21728 34840 21792
rect 34520 20704 34840 21728
rect 34520 20640 34528 20704
rect 34592 20640 34608 20704
rect 34672 20640 34688 20704
rect 34752 20640 34768 20704
rect 34832 20640 34840 20704
rect 34520 19616 34840 20640
rect 34520 19552 34528 19616
rect 34592 19552 34608 19616
rect 34672 19552 34688 19616
rect 34752 19552 34768 19616
rect 34832 19552 34840 19616
rect 34520 18528 34840 19552
rect 34520 18464 34528 18528
rect 34592 18464 34608 18528
rect 34672 18464 34688 18528
rect 34752 18464 34768 18528
rect 34832 18464 34840 18528
rect 34520 17440 34840 18464
rect 34520 17376 34528 17440
rect 34592 17376 34608 17440
rect 34672 17376 34688 17440
rect 34752 17376 34768 17440
rect 34832 17376 34840 17440
rect 34520 16352 34840 17376
rect 34520 16288 34528 16352
rect 34592 16288 34608 16352
rect 34672 16288 34688 16352
rect 34752 16288 34768 16352
rect 34832 16288 34840 16352
rect 34520 15264 34840 16288
rect 34520 15200 34528 15264
rect 34592 15200 34608 15264
rect 34672 15200 34688 15264
rect 34752 15200 34768 15264
rect 34832 15200 34840 15264
rect 34520 14176 34840 15200
rect 34520 14112 34528 14176
rect 34592 14112 34608 14176
rect 34672 14112 34688 14176
rect 34752 14112 34768 14176
rect 34832 14112 34840 14176
rect 34520 13088 34840 14112
rect 34520 13024 34528 13088
rect 34592 13024 34608 13088
rect 34672 13024 34688 13088
rect 34752 13024 34768 13088
rect 34832 13024 34840 13088
rect 34520 12000 34840 13024
rect 34520 11936 34528 12000
rect 34592 11936 34608 12000
rect 34672 11936 34688 12000
rect 34752 11936 34768 12000
rect 34832 11936 34840 12000
rect 34520 10912 34840 11936
rect 34520 10848 34528 10912
rect 34592 10848 34608 10912
rect 34672 10848 34688 10912
rect 34752 10848 34768 10912
rect 34832 10848 34840 10912
rect 34520 9824 34840 10848
rect 34520 9760 34528 9824
rect 34592 9760 34608 9824
rect 34672 9760 34688 9824
rect 34752 9760 34768 9824
rect 34832 9760 34840 9824
rect 34520 8736 34840 9760
rect 34520 8672 34528 8736
rect 34592 8672 34608 8736
rect 34672 8672 34688 8736
rect 34752 8672 34768 8736
rect 34832 8672 34840 8736
rect 34520 7648 34840 8672
rect 34520 7584 34528 7648
rect 34592 7584 34608 7648
rect 34672 7584 34688 7648
rect 34752 7584 34768 7648
rect 34832 7584 34840 7648
rect 34520 6560 34840 7584
rect 34520 6496 34528 6560
rect 34592 6496 34608 6560
rect 34672 6496 34688 6560
rect 34752 6496 34768 6560
rect 34832 6496 34840 6560
rect 34520 5472 34840 6496
rect 34520 5408 34528 5472
rect 34592 5408 34608 5472
rect 34672 5408 34688 5472
rect 34752 5408 34768 5472
rect 34832 5408 34840 5472
rect 34520 4384 34840 5408
rect 34520 4320 34528 4384
rect 34592 4320 34608 4384
rect 34672 4320 34688 4384
rect 34752 4320 34768 4384
rect 34832 4320 34840 4384
rect 34520 3296 34840 4320
rect 34520 3232 34528 3296
rect 34592 3232 34608 3296
rect 34672 3232 34688 3296
rect 34752 3232 34768 3296
rect 34832 3232 34840 3296
rect 34520 2208 34840 3232
rect 34520 2144 34528 2208
rect 34592 2144 34608 2208
rect 34672 2144 34688 2208
rect 34752 2144 34768 2208
rect 34832 2144 34840 2208
rect 34520 2128 34840 2144
use sky130_fd_sc_hd__inv_2  _0779_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0780_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _0781_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _0782_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_2  _0783_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6256 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _0784_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7728 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__or3_2  _0785_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3680 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0786_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4416 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0787_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _0788_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__o31a_2  _0789_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _0790_
timestamp 1688980957
transform 1 0 4416 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_2  _0791_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_4  _0792_
timestamp 1688980957
transform 1 0 11592 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0793_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9936 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1688980957
transform -1 0 11040 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0795_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10304 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0796_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10212 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0797_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0798_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0799_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_4  _0800_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_4  _0801_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 1688980957
transform 1 0 7176 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0803_
timestamp 1688980957
transform 1 0 7728 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0804_
timestamp 1688980957
transform 1 0 3404 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0805_
timestamp 1688980957
transform -1 0 9568 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0806_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0807_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _0808_
timestamp 1688980957
transform -1 0 8004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0810_
timestamp 1688980957
transform 1 0 4048 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _0811_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0812_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0813_
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0814_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0815_
timestamp 1688980957
transform 1 0 5520 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0816_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9844 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0817_
timestamp 1688980957
transform 1 0 12144 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1688980957
transform 1 0 3956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0819_
timestamp 1688980957
transform 1 0 6440 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0820_
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1688980957
transform 1 0 4232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0822_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0823_
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0824_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4048 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0825_
timestamp 1688980957
transform -1 0 5520 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0826_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12512 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1688980957
transform -1 0 13800 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0828_
timestamp 1688980957
transform -1 0 13524 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0829_
timestamp 1688980957
transform 1 0 12880 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1688980957
transform 1 0 6256 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0831_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11960 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0832_
timestamp 1688980957
transform -1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0833_
timestamp 1688980957
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0834_
timestamp 1688980957
transform 1 0 8004 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0835_
timestamp 1688980957
transform 1 0 4508 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0836_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0838_
timestamp 1688980957
transform -1 0 11500 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0839_
timestamp 1688980957
transform -1 0 11868 0 1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__a41o_1  _0840_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0841_
timestamp 1688980957
transform -1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0842_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0843_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0844_
timestamp 1688980957
transform -1 0 3496 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0845_
timestamp 1688980957
transform -1 0 9476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 1688980957
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0847_
timestamp 1688980957
transform 1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0848_
timestamp 1688980957
transform -1 0 5520 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0849_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0850_
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0851_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9844 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0852_
timestamp 1688980957
transform -1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _0853_
timestamp 1688980957
transform 1 0 4968 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__o31a_1  _0854_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10212 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0855_
timestamp 1688980957
transform -1 0 9936 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _0856_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10304 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0857_
timestamp 1688980957
transform -1 0 10212 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0858_
timestamp 1688980957
transform 1 0 10304 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0859_
timestamp 1688980957
transform 1 0 9016 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0860_
timestamp 1688980957
transform 1 0 9752 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1688980957
transform -1 0 8096 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0862_
timestamp 1688980957
transform 1 0 5428 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0863_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0864_
timestamp 1688980957
transform 1 0 13800 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1688980957
transform 1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0866_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13800 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0867_
timestamp 1688980957
transform -1 0 13800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1688980957
transform -1 0 12420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0869_
timestamp 1688980957
transform -1 0 13800 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0870_
timestamp 1688980957
transform -1 0 5244 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0871_
timestamp 1688980957
transform -1 0 11316 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0872_
timestamp 1688980957
transform -1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0873_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13248 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0874_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10488 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0875_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0876_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0877_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0878_
timestamp 1688980957
transform 1 0 9200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0879_
timestamp 1688980957
transform -1 0 7176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0880_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0881_
timestamp 1688980957
transform -1 0 5704 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0882_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6716 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0883_
timestamp 1688980957
transform -1 0 6992 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0884_
timestamp 1688980957
transform -1 0 6440 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0885_
timestamp 1688980957
transform -1 0 9200 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0886_
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1688980957
transform 1 0 8280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1688980957
transform 1 0 7820 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0889_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0890_
timestamp 1688980957
transform -1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0891_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8832 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _0892_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7176 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a311oi_1  _0893_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0894_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0895_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6348 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0896_
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0897_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9752 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0898_
timestamp 1688980957
transform 1 0 8740 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0899_
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_2  _0900_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0901_
timestamp 1688980957
transform -1 0 12512 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0902_
timestamp 1688980957
transform 1 0 6992 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0903_
timestamp 1688980957
transform 1 0 7452 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0904_
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0905_
timestamp 1688980957
transform -1 0 6808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0906_
timestamp 1688980957
transform -1 0 7452 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0907_
timestamp 1688980957
transform -1 0 11960 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _0908_
timestamp 1688980957
transform -1 0 13340 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _0909_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0910_
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0911_
timestamp 1688980957
transform -1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0912_
timestamp 1688980957
transform 1 0 6992 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0913_
timestamp 1688980957
transform 1 0 13156 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0914_
timestamp 1688980957
transform -1 0 12972 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1688980957
transform 1 0 7544 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0916_
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0917_
timestamp 1688980957
transform -1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0918_
timestamp 1688980957
transform -1 0 9752 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0919_
timestamp 1688980957
transform -1 0 7360 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0920_
timestamp 1688980957
transform -1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0921_
timestamp 1688980957
transform -1 0 14076 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _0922_
timestamp 1688980957
transform -1 0 13432 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0923_
timestamp 1688980957
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_4  _0924_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_4  _0925_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13800 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0926_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1688980957
transform 1 0 7452 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 1688980957
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1688980957
transform 1 0 8188 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0930_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8924 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0931_
timestamp 1688980957
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_4  _0932_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_1  _0933_
timestamp 1688980957
transform 1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0934_
timestamp 1688980957
transform 1 0 10396 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0935_
timestamp 1688980957
transform 1 0 9936 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0936_
timestamp 1688980957
transform -1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0937_
timestamp 1688980957
transform -1 0 11408 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1688980957
transform -1 0 13616 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0939_
timestamp 1688980957
transform -1 0 12052 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0940_
timestamp 1688980957
transform 1 0 12052 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0941_
timestamp 1688980957
transform 1 0 13524 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1688980957
transform -1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0943_
timestamp 1688980957
transform -1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0944_
timestamp 1688980957
transform -1 0 8648 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0945_
timestamp 1688980957
transform -1 0 12788 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0946_
timestamp 1688980957
transform -1 0 11684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0947_
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0948_
timestamp 1688980957
transform -1 0 11684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0949_
timestamp 1688980957
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1688980957
transform 1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0951_
timestamp 1688980957
transform -1 0 10672 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0952_
timestamp 1688980957
transform -1 0 11132 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0953_
timestamp 1688980957
transform 1 0 11040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0954_
timestamp 1688980957
transform 1 0 10672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0955_
timestamp 1688980957
transform -1 0 13616 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0956_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9752 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0957_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0958_
timestamp 1688980957
transform 1 0 14444 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0959_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0960_
timestamp 1688980957
transform 1 0 12052 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0961_
timestamp 1688980957
transform -1 0 16284 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0962_
timestamp 1688980957
transform 1 0 14536 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 1688980957
transform 1 0 15640 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0964_
timestamp 1688980957
transform -1 0 15364 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0965_
timestamp 1688980957
transform 1 0 14904 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0966_
timestamp 1688980957
transform -1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1688980957
transform 1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0968_
timestamp 1688980957
transform 1 0 15088 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0969_
timestamp 1688980957
transform -1 0 16008 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0970_
timestamp 1688980957
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0972_
timestamp 1688980957
transform 1 0 15180 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _0973_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15088 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0974_
timestamp 1688980957
transform 1 0 12512 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_4  _0975_
timestamp 1688980957
transform 1 0 12880 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__or2b_1  _0976_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15088 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _0977_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16284 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0978_
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_8  _0979_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0980_
timestamp 1688980957
transform -1 0 16376 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0981_
timestamp 1688980957
transform 1 0 16100 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0982_
timestamp 1688980957
transform 1 0 14720 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0985_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_1  _0986_
timestamp 1688980957
transform 1 0 16008 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0987_
timestamp 1688980957
transform 1 0 15272 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0988_
timestamp 1688980957
transform -1 0 16928 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 1688980957
transform -1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0990_
timestamp 1688980957
transform 1 0 17572 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0991_
timestamp 1688980957
transform 1 0 16928 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1688980957
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1688980957
transform -1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0994_
timestamp 1688980957
transform -1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0995_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0996_
timestamp 1688980957
transform -1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0997_
timestamp 1688980957
transform -1 0 16468 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0998_
timestamp 1688980957
transform -1 0 17296 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0999_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18584 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1000_
timestamp 1688980957
transform -1 0 14904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1001_
timestamp 1688980957
transform -1 0 15548 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1002_
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1003_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1004_
timestamp 1688980957
transform -1 0 17572 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1005_
timestamp 1688980957
transform -1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1006_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18676 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1007_
timestamp 1688980957
transform 1 0 20332 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1009_
timestamp 1688980957
transform 1 0 21712 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1010_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1011_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _1012_
timestamp 1688980957
transform 1 0 23276 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1013_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1014_
timestamp 1688980957
transform -1 0 21896 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1015_
timestamp 1688980957
transform 1 0 20976 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1017_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22264 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1018_
timestamp 1688980957
transform -1 0 23184 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 1688980957
transform 1 0 23552 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1020_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1021_
timestamp 1688980957
transform 1 0 22724 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1022_
timestamp 1688980957
transform 1 0 23000 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1024_
timestamp 1688980957
transform -1 0 23552 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1025_
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1026_
timestamp 1688980957
transform 1 0 19964 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1688980957
transform -1 0 20792 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1028_
timestamp 1688980957
transform 1 0 20424 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1029_
timestamp 1688980957
transform -1 0 20424 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1688980957
transform -1 0 22264 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_4  _1031_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24196 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_1  _1032_
timestamp 1688980957
transform 1 0 20608 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1033_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _1034_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_2  _1035_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19780 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1036_
timestamp 1688980957
transform -1 0 20056 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1037_
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1038_
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 1688980957
transform -1 0 21712 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1040_
timestamp 1688980957
transform -1 0 21436 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1041_
timestamp 1688980957
transform 1 0 23368 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1042_
timestamp 1688980957
transform 1 0 22172 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1043_
timestamp 1688980957
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1044_
timestamp 1688980957
transform 1 0 22540 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1045_
timestamp 1688980957
transform 1 0 20332 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_4  _1046_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1688980957
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _1048_
timestamp 1688980957
transform -1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _1049_
timestamp 1688980957
transform -1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1050_
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1051_
timestamp 1688980957
transform -1 0 21160 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1052_
timestamp 1688980957
transform -1 0 21528 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1053_
timestamp 1688980957
transform 1 0 20700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1054_
timestamp 1688980957
transform -1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1055_
timestamp 1688980957
transform -1 0 18308 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1056_
timestamp 1688980957
transform -1 0 18952 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1057_
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1058_
timestamp 1688980957
transform 1 0 20608 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_2  _1059_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21160 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o22ai_1  _1060_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _1061_
timestamp 1688980957
transform 1 0 21620 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1062_
timestamp 1688980957
transform -1 0 21712 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1063_
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_4  _1064_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__a32o_1  _1065_
timestamp 1688980957
transform 1 0 22540 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1066_
timestamp 1688980957
transform -1 0 20332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1067_
timestamp 1688980957
transform -1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1688980957
transform -1 0 24104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1069_
timestamp 1688980957
transform 1 0 22540 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1070_
timestamp 1688980957
transform 1 0 21988 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1071_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20884 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1072_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1073_
timestamp 1688980957
transform -1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1074_
timestamp 1688980957
transform 1 0 21344 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1075_
timestamp 1688980957
transform 1 0 23276 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1076_
timestamp 1688980957
transform 1 0 22816 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_4  _1077_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23368 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__nand4_1  _1078_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17112 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1079_
timestamp 1688980957
transform -1 0 19044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1081_
timestamp 1688980957
transform -1 0 19872 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1688980957
transform -1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1083_
timestamp 1688980957
transform -1 0 19780 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1084_
timestamp 1688980957
transform 1 0 20240 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1085_
timestamp 1688980957
transform 1 0 19504 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1688980957
transform -1 0 19872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1087_
timestamp 1688980957
transform -1 0 17940 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1088_
timestamp 1688980957
transform -1 0 18308 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1089_
timestamp 1688980957
transform 1 0 17112 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1688980957
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 1688980957
transform -1 0 17848 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1092_
timestamp 1688980957
transform 1 0 17020 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1093_
timestamp 1688980957
transform 1 0 17480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1688980957
transform -1 0 18492 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1095_
timestamp 1688980957
transform -1 0 18400 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1688980957
transform 1 0 17480 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1097_
timestamp 1688980957
transform 1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1688980957
transform -1 0 18400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1099_
timestamp 1688980957
transform 1 0 16100 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1688980957
transform -1 0 17940 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1101_
timestamp 1688980957
transform -1 0 17204 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1688980957
transform 1 0 15364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1103_
timestamp 1688980957
transform -1 0 18400 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1104_
timestamp 1688980957
transform 1 0 17112 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1105_
timestamp 1688980957
transform 1 0 17204 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1688980957
transform 1 0 18400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1688980957
transform 1 0 17204 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1108_
timestamp 1688980957
transform 1 0 18400 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1109_
timestamp 1688980957
transform 1 0 17664 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1110_
timestamp 1688980957
transform -1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1111_
timestamp 1688980957
transform -1 0 18584 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1113_
timestamp 1688980957
transform 1 0 17572 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1688980957
transform -1 0 18952 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1115_
timestamp 1688980957
transform -1 0 17940 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1688980957
transform 1 0 17020 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1117_
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1118_
timestamp 1688980957
transform -1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1119_
timestamp 1688980957
transform 1 0 16928 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1120_
timestamp 1688980957
transform 1 0 17112 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1121_
timestamp 1688980957
transform -1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1688980957
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1123_
timestamp 1688980957
transform -1 0 18584 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1124_
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1125_
timestamp 1688980957
transform 1 0 17572 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1126_
timestamp 1688980957
transform 1 0 18768 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1127_
timestamp 1688980957
transform -1 0 19688 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1688980957
transform -1 0 19228 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1129_
timestamp 1688980957
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1130_
timestamp 1688980957
transform -1 0 19872 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1688980957
transform 1 0 19412 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1132_
timestamp 1688980957
transform 1 0 18952 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1133_
timestamp 1688980957
transform -1 0 19872 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1134_
timestamp 1688980957
transform -1 0 19596 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1135_
timestamp 1688980957
transform -1 0 18952 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1136_
timestamp 1688980957
transform 1 0 17204 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1137_
timestamp 1688980957
transform 1 0 18216 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1138_
timestamp 1688980957
transform -1 0 11408 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1139_
timestamp 1688980957
transform -1 0 12604 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1140_
timestamp 1688980957
transform -1 0 12696 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1141_
timestamp 1688980957
transform -1 0 11960 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 1688980957
transform 1 0 11040 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1143_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10948 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1144_
timestamp 1688980957
transform 1 0 10120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1145_
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1146_
timestamp 1688980957
transform 1 0 11868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1147_
timestamp 1688980957
transform 1 0 10212 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1148_
timestamp 1688980957
transform 1 0 11776 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1149_
timestamp 1688980957
transform 1 0 11224 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1150_
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1151_
timestamp 1688980957
transform -1 0 12144 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1152_
timestamp 1688980957
transform -1 0 12788 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1688980957
transform -1 0 12972 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1154_
timestamp 1688980957
transform 1 0 14168 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1155_
timestamp 1688980957
transform 1 0 14720 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1156_
timestamp 1688980957
transform -1 0 14720 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1157_
timestamp 1688980957
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1158_
timestamp 1688980957
transform 1 0 15364 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1159_
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1160_
timestamp 1688980957
transform -1 0 16284 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1161_
timestamp 1688980957
transform 1 0 15456 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1162_
timestamp 1688980957
transform -1 0 18032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1163_
timestamp 1688980957
transform -1 0 17020 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1164_
timestamp 1688980957
transform 1 0 16008 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1165_
timestamp 1688980957
transform -1 0 17112 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1166_
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1167_
timestamp 1688980957
transform -1 0 16100 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1168_
timestamp 1688980957
transform -1 0 15364 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1169_
timestamp 1688980957
transform 1 0 13524 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1170_
timestamp 1688980957
transform 1 0 13800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1171_
timestamp 1688980957
transform 1 0 14168 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1172_
timestamp 1688980957
transform -1 0 14260 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1173_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1174_
timestamp 1688980957
transform -1 0 15272 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1175_
timestamp 1688980957
transform 1 0 15180 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1176_
timestamp 1688980957
transform 1 0 14720 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1688980957
transform -1 0 15640 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1178_
timestamp 1688980957
transform -1 0 15364 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1179_
timestamp 1688980957
transform -1 0 14536 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1180_
timestamp 1688980957
transform -1 0 14904 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1182_
timestamp 1688980957
transform -1 0 15732 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1183_
timestamp 1688980957
transform -1 0 15088 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1184_
timestamp 1688980957
transform 1 0 5336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1185_
timestamp 1688980957
transform -1 0 9476 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1186_
timestamp 1688980957
transform 1 0 5336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1187_
timestamp 1688980957
transform -1 0 7268 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1188_
timestamp 1688980957
transform 1 0 5428 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1189_
timestamp 1688980957
transform -1 0 7084 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1190_
timestamp 1688980957
transform -1 0 7084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1191_
timestamp 1688980957
transform 1 0 5796 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1192_
timestamp 1688980957
transform 1 0 6256 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1193_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6992 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1194_
timestamp 1688980957
transform 1 0 7360 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1195_
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1196_
timestamp 1688980957
transform -1 0 7912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1197_
timestamp 1688980957
transform -1 0 7452 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1198_
timestamp 1688980957
transform 1 0 6440 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1199_
timestamp 1688980957
transform -1 0 6992 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1200_
timestamp 1688980957
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1201_
timestamp 1688980957
transform -1 0 5244 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1202_
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1203_
timestamp 1688980957
transform 1 0 4324 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1204_
timestamp 1688980957
transform -1 0 4140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1205_
timestamp 1688980957
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1206_
timestamp 1688980957
transform -1 0 5060 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1207_
timestamp 1688980957
transform 1 0 4508 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1208_
timestamp 1688980957
transform -1 0 4416 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1688980957
transform -1 0 3680 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1210_
timestamp 1688980957
transform -1 0 3680 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1211_
timestamp 1688980957
transform 1 0 3496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1212_
timestamp 1688980957
transform 1 0 2944 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1213_
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1214_
timestamp 1688980957
transform -1 0 4140 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1215_
timestamp 1688980957
transform 1 0 4416 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1216_
timestamp 1688980957
transform 1 0 5520 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1217_
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1218_
timestamp 1688980957
transform 1 0 5336 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1219_
timestamp 1688980957
transform 1 0 6900 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1688980957
transform -1 0 7820 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1221_
timestamp 1688980957
transform 1 0 6900 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1222_
timestamp 1688980957
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1223_
timestamp 1688980957
transform 1 0 9568 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1224_
timestamp 1688980957
transform 1 0 8832 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1225_
timestamp 1688980957
transform 1 0 9016 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1226_
timestamp 1688980957
transform -1 0 8832 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1227_
timestamp 1688980957
transform 1 0 9476 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1228_
timestamp 1688980957
transform -1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1229_
timestamp 1688980957
transform 1 0 9108 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1230_
timestamp 1688980957
transform 1 0 9752 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1231_
timestamp 1688980957
transform 1 0 9568 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1232_
timestamp 1688980957
transform -1 0 10672 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1233_
timestamp 1688980957
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1234_
timestamp 1688980957
transform 1 0 7728 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1235_
timestamp 1688980957
transform -1 0 8464 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1236_
timestamp 1688980957
transform 1 0 8924 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1237_
timestamp 1688980957
transform 1 0 8096 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1238_
timestamp 1688980957
transform -1 0 9108 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1239_
timestamp 1688980957
transform -1 0 7544 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1688980957
transform 1 0 8096 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1241_
timestamp 1688980957
transform 1 0 7452 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1242_
timestamp 1688980957
transform 1 0 7912 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1243_
timestamp 1688980957
transform -1 0 6716 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1244_
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1245_
timestamp 1688980957
transform -1 0 5612 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1246_
timestamp 1688980957
transform 1 0 5612 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1247_
timestamp 1688980957
transform 1 0 3956 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1248_
timestamp 1688980957
transform 1 0 4600 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1249_
timestamp 1688980957
transform -1 0 4324 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1250_
timestamp 1688980957
transform -1 0 4324 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1251_
timestamp 1688980957
transform -1 0 4324 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1252_
timestamp 1688980957
transform 1 0 2300 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1253_
timestamp 1688980957
transform 1 0 4324 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 1688980957
transform 1 0 4416 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1255_
timestamp 1688980957
transform -1 0 5428 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1688980957
transform 1 0 3220 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1257_
timestamp 1688980957
transform -1 0 6440 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1258_
timestamp 1688980957
transform -1 0 6072 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1259_
timestamp 1688980957
transform -1 0 15364 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1260_
timestamp 1688980957
transform -1 0 13064 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1261_
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1262_
timestamp 1688980957
transform -1 0 13156 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1263_
timestamp 1688980957
transform -1 0 12236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1264_
timestamp 1688980957
transform 1 0 12144 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1688980957
transform 1 0 20516 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1266_
timestamp 1688980957
transform 1 0 20792 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1267_
timestamp 1688980957
transform -1 0 19964 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1268_
timestamp 1688980957
transform 1 0 19136 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1269_
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1270_
timestamp 1688980957
transform 1 0 18308 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1271_
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1272_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19596 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1273_
timestamp 1688980957
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1274_
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _1275_
timestamp 1688980957
transform -1 0 20792 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1276_
timestamp 1688980957
transform -1 0 19504 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1277_
timestamp 1688980957
transform 1 0 18308 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1278_
timestamp 1688980957
transform -1 0 21712 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1279_
timestamp 1688980957
transform 1 0 20332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1280_
timestamp 1688980957
transform 1 0 20608 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1688980957
transform 1 0 19780 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1282_
timestamp 1688980957
transform -1 0 21344 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1283_
timestamp 1688980957
transform -1 0 21620 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1284_
timestamp 1688980957
transform 1 0 20792 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1285_
timestamp 1688980957
transform 1 0 20148 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1286_
timestamp 1688980957
transform -1 0 21252 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1287_
timestamp 1688980957
transform -1 0 21620 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1288_
timestamp 1688980957
transform 1 0 20700 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1289_
timestamp 1688980957
transform -1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1290_
timestamp 1688980957
transform 1 0 20424 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1688980957
transform -1 0 21160 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1292_
timestamp 1688980957
transform 1 0 20424 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1293_
timestamp 1688980957
transform -1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1294_
timestamp 1688980957
transform -1 0 18952 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1295_
timestamp 1688980957
transform 1 0 19320 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1296_
timestamp 1688980957
transform -1 0 20056 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1297_
timestamp 1688980957
transform 1 0 19320 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1298_
timestamp 1688980957
transform -1 0 19228 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1299_
timestamp 1688980957
transform -1 0 18860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1300_
timestamp 1688980957
transform 1 0 18216 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1301_
timestamp 1688980957
transform -1 0 18216 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1302_
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1303_
timestamp 1688980957
transform -1 0 18032 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1304_
timestamp 1688980957
transform -1 0 17940 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1305_
timestamp 1688980957
transform 1 0 17112 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1306_
timestamp 1688980957
transform -1 0 17848 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _1307_
timestamp 1688980957
transform 1 0 17388 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1688980957
transform 1 0 27784 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1309_
timestamp 1688980957
transform 1 0 26404 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1310_
timestamp 1688980957
transform 1 0 27324 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1311_
timestamp 1688980957
transform 1 0 29900 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1312_
timestamp 1688980957
transform -1 0 27324 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1313_
timestamp 1688980957
transform 1 0 28980 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1314_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28152 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__a21oi_1  _1315_
timestamp 1688980957
transform 1 0 30360 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1316_
timestamp 1688980957
transform -1 0 29440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1317_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29624 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1688980957
transform 1 0 26036 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1319_
timestamp 1688980957
transform 1 0 27324 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _1320_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1321_
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1322_
timestamp 1688980957
transform 1 0 27232 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__or2b_1  _1323_
timestamp 1688980957
transform 1 0 29992 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1324_
timestamp 1688980957
transform 1 0 29992 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1325_
timestamp 1688980957
transform 1 0 30084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1326_
timestamp 1688980957
transform 1 0 30176 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1688980957
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1328_
timestamp 1688980957
transform 1 0 30176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1329_
timestamp 1688980957
transform -1 0 31556 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1330_
timestamp 1688980957
transform 1 0 27968 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1331_
timestamp 1688980957
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1332_
timestamp 1688980957
transform 1 0 30360 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1333_
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1334_
timestamp 1688980957
transform 1 0 29716 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1335_
timestamp 1688980957
transform -1 0 31924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1336_
timestamp 1688980957
transform 1 0 29808 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1337_
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1338_
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1339_
timestamp 1688980957
transform -1 0 31372 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1340_
timestamp 1688980957
transform 1 0 31096 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1341_
timestamp 1688980957
transform 1 0 33488 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1342_
timestamp 1688980957
transform 1 0 30268 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1343_
timestamp 1688980957
transform 1 0 30728 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1344_
timestamp 1688980957
transform -1 0 32384 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1345_
timestamp 1688980957
transform 1 0 31096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1346_
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1347_
timestamp 1688980957
transform 1 0 29716 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1348_
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1349_
timestamp 1688980957
transform 1 0 30544 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1350_
timestamp 1688980957
transform -1 0 31648 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1351_
timestamp 1688980957
transform 1 0 29900 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1352_
timestamp 1688980957
transform 1 0 31556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1353_
timestamp 1688980957
transform 1 0 31188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1354_
timestamp 1688980957
transform 1 0 29900 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1355_
timestamp 1688980957
transform -1 0 31096 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1356_
timestamp 1688980957
transform -1 0 31556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1357_
timestamp 1688980957
transform -1 0 32108 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 1688980957
transform 1 0 31464 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1359_
timestamp 1688980957
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1360_
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1361_
timestamp 1688980957
transform 1 0 28704 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1362_
timestamp 1688980957
transform 1 0 30084 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1363_
timestamp 1688980957
transform 1 0 30452 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1364_
timestamp 1688980957
transform 1 0 30084 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1365_
timestamp 1688980957
transform 1 0 30452 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1366_
timestamp 1688980957
transform 1 0 29256 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1367_
timestamp 1688980957
transform 1 0 28796 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1368_
timestamp 1688980957
transform -1 0 30360 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1369_
timestamp 1688980957
transform -1 0 31372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1370_
timestamp 1688980957
transform -1 0 30176 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1371_
timestamp 1688980957
transform 1 0 31188 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1372_
timestamp 1688980957
transform 1 0 30912 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1373_
timestamp 1688980957
transform 1 0 30084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1374_
timestamp 1688980957
transform 1 0 30636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1375_
timestamp 1688980957
transform 1 0 31188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1376_
timestamp 1688980957
transform 1 0 31464 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1377_
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1378_
timestamp 1688980957
transform 1 0 33120 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1379_
timestamp 1688980957
transform 1 0 31556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1380_
timestamp 1688980957
transform 1 0 31280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1381_
timestamp 1688980957
transform -1 0 32660 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1382_
timestamp 1688980957
transform 1 0 28520 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1383_
timestamp 1688980957
transform 1 0 29072 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1384_
timestamp 1688980957
transform 1 0 29624 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1385_
timestamp 1688980957
transform 1 0 30176 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1386_
timestamp 1688980957
transform 1 0 32936 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1387_
timestamp 1688980957
transform -1 0 34224 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1388_
timestamp 1688980957
transform -1 0 31740 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1389_
timestamp 1688980957
transform -1 0 31372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1390_
timestamp 1688980957
transform 1 0 28428 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1391_
timestamp 1688980957
transform 1 0 30728 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1392_
timestamp 1688980957
transform -1 0 32016 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1393_
timestamp 1688980957
transform 1 0 30360 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1394_
timestamp 1688980957
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _1395_
timestamp 1688980957
transform 1 0 33120 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1396_
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1397_
timestamp 1688980957
transform 1 0 24748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1398_
timestamp 1688980957
transform 1 0 27324 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1399_
timestamp 1688980957
transform 1 0 27416 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1400_
timestamp 1688980957
transform -1 0 27600 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1401_
timestamp 1688980957
transform -1 0 26864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1402_
timestamp 1688980957
transform -1 0 27324 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1403_
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1404_
timestamp 1688980957
transform -1 0 30084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1405_
timestamp 1688980957
transform -1 0 30636 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1406_
timestamp 1688980957
transform 1 0 28428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _1407_
timestamp 1688980957
transform 1 0 27876 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1408_
timestamp 1688980957
transform 1 0 28336 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1409_
timestamp 1688980957
transform -1 0 28796 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1410_
timestamp 1688980957
transform -1 0 30912 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1411_
timestamp 1688980957
transform 1 0 31464 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1412_
timestamp 1688980957
transform -1 0 33120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1413_
timestamp 1688980957
transform 1 0 31464 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1414_
timestamp 1688980957
transform 1 0 32200 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1415_
timestamp 1688980957
transform -1 0 31096 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1416_
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1417_
timestamp 1688980957
transform 1 0 32660 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1418_
timestamp 1688980957
transform 1 0 27968 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1419_
timestamp 1688980957
transform 1 0 28428 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1420_
timestamp 1688980957
transform -1 0 32292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1421_
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1422_
timestamp 1688980957
transform 1 0 32660 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1423_
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1424_
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1425_
timestamp 1688980957
transform -1 0 31740 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1426_
timestamp 1688980957
transform 1 0 32476 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1427_
timestamp 1688980957
transform 1 0 33120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1428_
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1429_
timestamp 1688980957
transform 1 0 30176 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1430_
timestamp 1688980957
transform -1 0 31556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1431_
timestamp 1688980957
transform -1 0 32016 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1432_
timestamp 1688980957
transform -1 0 32568 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1433_
timestamp 1688980957
transform -1 0 32568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1688980957
transform -1 0 32200 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1435_
timestamp 1688980957
transform 1 0 28244 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1436_
timestamp 1688980957
transform -1 0 28704 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1437_
timestamp 1688980957
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1438_
timestamp 1688980957
transform -1 0 32568 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1439_
timestamp 1688980957
transform -1 0 32936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1440_
timestamp 1688980957
transform -1 0 30176 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1441_
timestamp 1688980957
transform -1 0 28520 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1442_
timestamp 1688980957
transform -1 0 34132 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1443_
timestamp 1688980957
transform 1 0 33212 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1688980957
transform 1 0 33672 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1445_
timestamp 1688980957
transform 1 0 28244 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1446_
timestamp 1688980957
transform 1 0 27968 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1447_
timestamp 1688980957
transform -1 0 32936 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1448_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32660 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 1688980957
transform 1 0 33304 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1450_
timestamp 1688980957
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1451_
timestamp 1688980957
transform -1 0 30636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1452_
timestamp 1688980957
transform -1 0 28888 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1453_
timestamp 1688980957
transform 1 0 32752 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1454_
timestamp 1688980957
transform 1 0 32568 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1455_
timestamp 1688980957
transform 1 0 32752 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1688980957
transform 1 0 31280 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1457_
timestamp 1688980957
transform 1 0 32200 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1458_
timestamp 1688980957
transform 1 0 31004 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1459_
timestamp 1688980957
transform -1 0 33120 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1460_
timestamp 1688980957
transform 1 0 31648 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1461_
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1462_
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1463_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1464_
timestamp 1688980957
transform -1 0 33304 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1465_
timestamp 1688980957
transform -1 0 31924 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1466_
timestamp 1688980957
transform 1 0 31924 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1688980957
transform 1 0 32752 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 1688980957
transform 1 0 31188 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1469_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1470_
timestamp 1688980957
transform 1 0 30912 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1471_
timestamp 1688980957
transform 1 0 29808 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1472_
timestamp 1688980957
transform 1 0 30084 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1473_
timestamp 1688980957
transform 1 0 28152 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1474_
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1475_
timestamp 1688980957
transform 1 0 30452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1476_
timestamp 1688980957
transform -1 0 30176 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1477_
timestamp 1688980957
transform 1 0 28336 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1478_
timestamp 1688980957
transform -1 0 27232 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1479_
timestamp 1688980957
transform 1 0 27232 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1480_
timestamp 1688980957
transform -1 0 27784 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1481_
timestamp 1688980957
transform 1 0 22080 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1482_
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1483_
timestamp 1688980957
transform 1 0 22632 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 1688980957
transform 1 0 22264 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1485_
timestamp 1688980957
transform 1 0 23000 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1486_
timestamp 1688980957
transform 1 0 22632 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1487_
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1488_
timestamp 1688980957
transform 1 0 24748 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1489_
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1688980957
transform -1 0 26772 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1491_
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1688980957
transform 1 0 22540 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 1688980957
transform 1 0 22448 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1688980957
transform 1 0 21988 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1495_
timestamp 1688980957
transform 1 0 23368 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1688980957
transform 1 0 22908 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1497_
timestamp 1688980957
transform -1 0 25576 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1498_
timestamp 1688980957
transform 1 0 23552 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1499_
timestamp 1688980957
transform 1 0 24288 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1500_
timestamp 1688980957
transform 1 0 25944 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1501_
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1502_
timestamp 1688980957
transform 1 0 28336 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1503_
timestamp 1688980957
transform 1 0 23552 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1504_
timestamp 1688980957
transform 1 0 24748 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1505_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1506_
timestamp 1688980957
transform 1 0 23460 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1507_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 1688980957
transform -1 0 27048 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1509_
timestamp 1688980957
transform 1 0 27048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1510_
timestamp 1688980957
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1511_
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 1688980957
transform -1 0 24196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1513_
timestamp 1688980957
transform 1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1514_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1515_
timestamp 1688980957
transform -1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1516_
timestamp 1688980957
transform 1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1517_
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1518_
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1519_
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1520_
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1521_
timestamp 1688980957
transform -1 0 26956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1522_
timestamp 1688980957
transform -1 0 23828 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1523_
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1688980957
transform -1 0 26680 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1688980957
transform -1 0 27232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1526_
timestamp 1688980957
transform -1 0 23736 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1527_
timestamp 1688980957
transform 1 0 25760 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1528_
timestamp 1688980957
transform -1 0 25760 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1529_
timestamp 1688980957
transform 1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1530_
timestamp 1688980957
transform -1 0 26680 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1688980957
transform 1 0 26680 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1532_
timestamp 1688980957
transform 1 0 23552 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1533_
timestamp 1688980957
transform 1 0 26312 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1534_
timestamp 1688980957
transform -1 0 26772 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1535_
timestamp 1688980957
transform 1 0 24656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1536_
timestamp 1688980957
transform 1 0 25300 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1537_
timestamp 1688980957
transform 1 0 25392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1538_
timestamp 1688980957
transform 1 0 23184 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1539_
timestamp 1688980957
transform 1 0 26680 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1540_
timestamp 1688980957
transform -1 0 26864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1541_
timestamp 1688980957
transform 1 0 22172 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1542_
timestamp 1688980957
transform -1 0 25208 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1543_
timestamp 1688980957
transform 1 0 24748 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1544_
timestamp 1688980957
transform 1 0 23920 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1545_
timestamp 1688980957
transform 1 0 23644 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1546_
timestamp 1688980957
transform 1 0 20792 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1547_
timestamp 1688980957
transform 1 0 24932 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1548_
timestamp 1688980957
transform -1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1549_
timestamp 1688980957
transform -1 0 5336 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1550_
timestamp 1688980957
transform 1 0 4692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1551_
timestamp 1688980957
transform 1 0 5060 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1552_
timestamp 1688980957
transform 1 0 4784 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1553_
timestamp 1688980957
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1554_
timestamp 1688980957
transform -1 0 4692 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1555_
timestamp 1688980957
transform -1 0 4416 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1556_
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o41ai_1  _1557_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6992 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1558_
timestamp 1688980957
transform 1 0 3956 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 1688980957
transform -1 0 5428 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1560_
timestamp 1688980957
transform -1 0 5152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1561_
timestamp 1688980957
transform 1 0 4140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1688980957
transform 1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1563_
timestamp 1688980957
transform 1 0 4416 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1564_
timestamp 1688980957
transform -1 0 4048 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1565_
timestamp 1688980957
transform 1 0 5520 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1566_
timestamp 1688980957
transform 1 0 5060 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1567_
timestamp 1688980957
transform 1 0 4784 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1568_
timestamp 1688980957
transform 1 0 7820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1569_
timestamp 1688980957
transform 1 0 7176 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1570_
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1571_
timestamp 1688980957
transform -1 0 9660 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1572_
timestamp 1688980957
transform 1 0 9936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1573_
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1574_
timestamp 1688980957
transform 1 0 6716 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1575_
timestamp 1688980957
transform 1 0 6164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_8  _1576_
timestamp 1688980957
transform -1 0 18216 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1577_
timestamp 1688980957
transform 1 0 21344 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1578_
timestamp 1688980957
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1579_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1580_
timestamp 1688980957
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1581_
timestamp 1688980957
transform -1 0 22908 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1582_
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1583_
timestamp 1688980957
transform -1 0 23368 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1584_
timestamp 1688980957
transform 1 0 23368 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1585_
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1586_
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1587_
timestamp 1688980957
transform 1 0 24932 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1588_
timestamp 1688980957
transform -1 0 24748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1589_
timestamp 1688980957
transform 1 0 24564 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1590_
timestamp 1688980957
transform 1 0 24656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1591_
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1592_
timestamp 1688980957
transform -1 0 23920 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1593_
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1594_
timestamp 1688980957
transform -1 0 24104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1595_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1596_
timestamp 1688980957
transform -1 0 24656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1597_
timestamp 1688980957
transform -1 0 24288 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1598_
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1599_
timestamp 1688980957
transform -1 0 23828 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1600_
timestamp 1688980957
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1601_
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1602_
timestamp 1688980957
transform -1 0 22356 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1603_
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1604_
timestamp 1688980957
transform -1 0 21252 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1605_
timestamp 1688980957
transform 1 0 19320 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1606_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1607_
timestamp 1688980957
transform -1 0 21620 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1608_
timestamp 1688980957
transform -1 0 21344 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1609_
timestamp 1688980957
transform 1 0 26128 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1610_
timestamp 1688980957
transform 1 0 28336 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1611_
timestamp 1688980957
transform 1 0 26312 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1612_
timestamp 1688980957
transform -1 0 25392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1613_
timestamp 1688980957
transform 1 0 16744 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1614_
timestamp 1688980957
transform 1 0 18216 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1615_
timestamp 1688980957
transform 1 0 17848 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1616_
timestamp 1688980957
transform 1 0 19688 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1617_
timestamp 1688980957
transform -1 0 19872 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1618_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32568 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1619_
timestamp 1688980957
transform -1 0 31464 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1620_
timestamp 1688980957
transform 1 0 27140 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1621_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1622_
timestamp 1688980957
transform -1 0 13984 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1623_
timestamp 1688980957
transform 1 0 24932 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1624_
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1625_
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1626_
timestamp 1688980957
transform -1 0 34408 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1627_
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1628_
timestamp 1688980957
transform 1 0 32568 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1629_
timestamp 1688980957
transform -1 0 30452 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1630_
timestamp 1688980957
transform 1 0 27600 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1631_
timestamp 1688980957
transform 1 0 27140 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1632_
timestamp 1688980957
transform -1 0 29808 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1633_
timestamp 1688980957
transform 1 0 27876 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1634_
timestamp 1688980957
transform -1 0 34316 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1635_
timestamp 1688980957
transform -1 0 34408 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1636_
timestamp 1688980957
transform -1 0 33672 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1637_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28244 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1638_
timestamp 1688980957
transform 1 0 26496 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _1639_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16008 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1640_
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1641_
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1642_
timestamp 1688980957
transform 1 0 17020 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1643_
timestamp 1688980957
transform 1 0 18400 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1644_
timestamp 1688980957
transform 1 0 18400 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1645_
timestamp 1688980957
transform 1 0 14812 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1646_
timestamp 1688980957
transform 1 0 17940 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1647_
timestamp 1688980957
transform 1 0 18216 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1648_
timestamp 1688980957
transform 1 0 18492 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1649_
timestamp 1688980957
transform -1 0 21160 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1650_
timestamp 1688980957
transform 1 0 15548 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1651_
timestamp 1688980957
transform 1 0 18308 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1652_
timestamp 1688980957
transform 1 0 19872 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1653_
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1654_
timestamp 1688980957
transform 1 0 17296 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1655_
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1656_
timestamp 1688980957
transform -1 0 13708 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1657_
timestamp 1688980957
transform 1 0 9568 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1658_
timestamp 1688980957
transform 1 0 9292 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1659_
timestamp 1688980957
transform 1 0 10580 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1660_
timestamp 1688980957
transform -1 0 13984 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1661_
timestamp 1688980957
transform 1 0 13800 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1662_
timestamp 1688980957
transform 1 0 14720 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1663_
timestamp 1688980957
transform 1 0 20516 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1664_
timestamp 1688980957
transform 1 0 21712 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1665_
timestamp 1688980957
transform 1 0 22080 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1666_
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1667_
timestamp 1688980957
transform -1 0 28796 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1668_
timestamp 1688980957
transform 1 0 21988 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1669_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1670_
timestamp 1688980957
transform 1 0 22356 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1671_
timestamp 1688980957
transform -1 0 24840 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1672_
timestamp 1688980957
transform -1 0 25668 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1673_
timestamp 1688980957
transform -1 0 26404 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1674_
timestamp 1688980957
transform 1 0 26220 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1675_
timestamp 1688980957
transform 1 0 27968 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1676_
timestamp 1688980957
transform -1 0 30636 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1677_
timestamp 1688980957
transform -1 0 26036 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1678_
timestamp 1688980957
transform -1 0 26864 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1679_
timestamp 1688980957
transform 1 0 23460 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1680_
timestamp 1688980957
transform 1 0 26036 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1681_
timestamp 1688980957
transform 1 0 24196 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1682_
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1683_
timestamp 1688980957
transform 1 0 26036 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1684_
timestamp 1688980957
transform 1 0 26956 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1685_
timestamp 1688980957
transform 1 0 26496 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1686_
timestamp 1688980957
transform -1 0 27692 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1687_
timestamp 1688980957
transform 1 0 25760 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1688_
timestamp 1688980957
transform 1 0 25852 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1689_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1690_
timestamp 1688980957
transform 1 0 25024 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1691_
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1692_
timestamp 1688980957
transform 1 0 24564 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1693_
timestamp 1688980957
transform 1 0 23092 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1694_
timestamp 1688980957
transform 1 0 24840 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1695_
timestamp 1688980957
transform -1 0 3588 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1696_
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_4  _1697_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 -1 20672
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_4  _1698_
timestamp 1688980957
transform 1 0 1564 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1699_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1700_
timestamp 1688980957
transform 1 0 6992 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1701_
timestamp 1688980957
transform 1 0 9292 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1702_
timestamp 1688980957
transform 1 0 8464 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1703_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1704_
timestamp 1688980957
transform 1 0 19872 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1705_
timestamp 1688980957
transform 1 0 21896 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1706_
timestamp 1688980957
transform 1 0 21896 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1707_
timestamp 1688980957
transform 1 0 22448 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1708_
timestamp 1688980957
transform 1 0 22448 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1709_
timestamp 1688980957
transform 1 0 24748 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1710_
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1711_
timestamp 1688980957
transform 1 0 23920 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1712_
timestamp 1688980957
transform 1 0 24104 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1713_
timestamp 1688980957
transform 1 0 24196 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1714_
timestamp 1688980957
transform 1 0 23460 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1715_
timestamp 1688980957
transform 1 0 23092 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1716_
timestamp 1688980957
transform 1 0 22356 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1717_
timestamp 1688980957
transform 1 0 21252 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1718_
timestamp 1688980957
transform 1 0 19044 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1719_
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1720_
timestamp 1688980957
transform -1 0 27968 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1721_
timestamp 1688980957
transform 1 0 25208 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1722_
timestamp 1688980957
transform 1 0 24288 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1723_
timestamp 1688980957
transform 1 0 17112 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1724_
timestamp 1688980957
transform 1 0 15824 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1725_
timestamp 1688980957
transform 1 0 15548 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1726_
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1727_
timestamp 1688980957
transform 1 0 12052 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1728_
timestamp 1688980957
transform 1 0 15272 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1729_
timestamp 1688980957
transform 1 0 12420 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1730_
timestamp 1688980957
transform 1 0 15088 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1731_
timestamp 1688980957
transform 1 0 6900 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1732_
timestamp 1688980957
transform -1 0 9568 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1733_
timestamp 1688980957
transform 1 0 6256 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1734_
timestamp 1688980957
transform 1 0 3772 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1735_
timestamp 1688980957
transform 1 0 1840 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1736_
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1737_
timestamp 1688980957
transform 1 0 1564 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1738_
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1739_
timestamp 1688980957
transform 1 0 5152 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1740_
timestamp 1688980957
transform -1 0 8924 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1741_
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1742_
timestamp 1688980957
transform -1 0 12052 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1743_
timestamp 1688980957
transform -1 0 12052 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1744_
timestamp 1688980957
transform 1 0 6992 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1745_
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1746_
timestamp 1688980957
transform 1 0 7636 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1747_
timestamp 1688980957
transform -1 0 7176 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1748_
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1749_
timestamp 1688980957
transform 1 0 1840 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1750_
timestamp 1688980957
transform 1 0 2760 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1751_
timestamp 1688980957
transform 1 0 5152 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1752_
timestamp 1688980957
transform -1 0 17756 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1753_
timestamp 1688980957
transform 1 0 14536 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1754_
timestamp 1688980957
transform -1 0 19780 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1755_
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1756_
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1757_
timestamp 1688980957
transform 1 0 2668 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1758_
timestamp 1688980957
transform -1 0 16560 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1759_
timestamp 1688980957
transform 1 0 12880 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1760_
timestamp 1688980957
transform -1 0 16192 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1761_
timestamp 1688980957
transform -1 0 16008 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1762_
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1763_
timestamp 1688980957
transform 1 0 13432 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1764_
timestamp 1688980957
transform 1 0 12880 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1765_
timestamp 1688980957
transform 1 0 14168 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1766_
timestamp 1688980957
transform -1 0 34408 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1767_
timestamp 1688980957
transform -1 0 32016 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1768_
timestamp 1688980957
transform -1 0 34408 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1769_
timestamp 1688980957
transform -1 0 18584 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1770_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1771_
timestamp 1688980957
transform 1 0 7176 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1772_
timestamp 1688980957
transform 1 0 17296 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1773_
timestamp 1688980957
transform 1 0 19872 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1774_
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1775_
timestamp 1688980957
transform -1 0 16008 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1776_
timestamp 1688980957
transform 1 0 11868 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1777_
timestamp 1688980957
transform -1 0 34408 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1778_
timestamp 1688980957
transform -1 0 34408 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1779_
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1780_
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1781_
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1782_
timestamp 1688980957
transform 1 0 12328 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1783_
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1784_
timestamp 1688980957
transform 1 0 15272 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1785_
timestamp 1688980957
transform -1 0 15916 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19780 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1688980957
transform -1 0 8832 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform -1 0 9016 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform -1 0 13432 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform -1 0 13984 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform -1 0 8556 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform 1 0 7820 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform -1 0 15456 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform -1 0 15088 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform -1 0 24656 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 23276 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform -1 0 28796 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 25852 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 24656 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform -1 0 26404 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 29440 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout28
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout29
timestamp 1688980957
transform -1 0 9936 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout30
timestamp 1688980957
transform -1 0 16008 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout31
timestamp 1688980957
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout32
timestamp 1688980957
transform -1 0 17204 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout33
timestamp 1688980957
transform -1 0 20700 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout34
timestamp 1688980957
transform 1 0 29808 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout35
timestamp 1688980957
transform 1 0 23920 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout36
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout37
timestamp 1688980957
transform -1 0 27876 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp 1688980957
transform 1 0 21804 0 1 34816
box -38 -48 866 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_203
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_258
timestamp 1688980957
transform 1 0 24840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_270
timestamp 1688980957
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_278
timestamp 1688980957
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_321 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_328
timestamp 1688980957
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_357
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_169
timestamp 1688980957
transform 1 0 16652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_190
timestamp 1688980957
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_361
timestamp 1688980957
transform 1 0 34316 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_141
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_162
timestamp 1688980957
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_203
timestamp 1688980957
transform 1 0 19780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_215
timestamp 1688980957
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_231
timestamp 1688980957
transform 1 0 22356 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_243
timestamp 1688980957
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_247
timestamp 1688980957
transform 1 0 23828 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_271
timestamp 1688980957
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_301
timestamp 1688980957
transform 1 0 28796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_313
timestamp 1688980957
transform 1 0 29900 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_129
timestamp 1688980957
transform 1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_155
timestamp 1688980957
transform 1 0 15364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_167
timestamp 1688980957
transform 1 0 16468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_179
timestamp 1688980957
transform 1 0 17572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_246
timestamp 1688980957
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_262
timestamp 1688980957
transform 1 0 25208 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_274
timestamp 1688980957
transform 1 0 26312 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_286
timestamp 1688980957
transform 1 0 27416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_298
timestamp 1688980957
transform 1 0 28520 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_318
timestamp 1688980957
transform 1 0 30360 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_330
timestamp 1688980957
transform 1 0 31464 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_342
timestamp 1688980957
transform 1 0 32568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_354
timestamp 1688980957
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_201
timestamp 1688980957
transform 1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_234
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_246
timestamp 1688980957
transform 1 0 23736 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_255
timestamp 1688980957
transform 1 0 24564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_288
timestamp 1688980957
transform 1 0 27600 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_296
timestamp 1688980957
transform 1 0 28336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_306
timestamp 1688980957
transform 1 0 29256 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_324
timestamp 1688980957
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_149
timestamp 1688980957
transform 1 0 14812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_181
timestamp 1688980957
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_193
timestamp 1688980957
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_229
timestamp 1688980957
transform 1 0 22172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_279
timestamp 1688980957
transform 1 0 26772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_285
timestamp 1688980957
transform 1 0 27324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_295
timestamp 1688980957
transform 1 0 28244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_315
timestamp 1688980957
transform 1 0 30084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_327
timestamp 1688980957
transform 1 0 31188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_337
timestamp 1688980957
transform 1 0 32108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_344
timestamp 1688980957
transform 1 0 32752 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_356
timestamp 1688980957
transform 1 0 33856 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_6
timestamp 1688980957
transform 1 0 1656 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_18
timestamp 1688980957
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_30
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_42
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_86
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_133
timestamp 1688980957
transform 1 0 13340 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_154
timestamp 1688980957
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_201
timestamp 1688980957
transform 1 0 19596 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_212
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_242
timestamp 1688980957
transform 1 0 23368 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_251
timestamp 1688980957
transform 1 0 24196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_259
timestamp 1688980957
transform 1 0 24932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_271
timestamp 1688980957
transform 1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_310
timestamp 1688980957
transform 1 0 29624 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_324
timestamp 1688980957
transform 1 0 30912 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_341
timestamp 1688980957
transform 1 0 32476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 1688980957
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1688980957
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1688980957
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_204
timestamp 1688980957
transform 1 0 19872 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_216
timestamp 1688980957
transform 1 0 20976 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_228
timestamp 1688980957
transform 1 0 22080 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_240
timestamp 1688980957
transform 1 0 23184 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_291
timestamp 1688980957
transform 1 0 27876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_303
timestamp 1688980957
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_312
timestamp 1688980957
transform 1 0 29808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_320
timestamp 1688980957
transform 1 0 30544 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_326
timestamp 1688980957
transform 1 0 31096 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_337
timestamp 1688980957
transform 1 0 32108 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_348
timestamp 1688980957
transform 1 0 33120 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_360
timestamp 1688980957
transform 1 0 34224 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_73
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_82
timestamp 1688980957
transform 1 0 8648 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_94
timestamp 1688980957
transform 1 0 9752 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_102
timestamp 1688980957
transform 1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_121
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_142
timestamp 1688980957
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_172
timestamp 1688980957
transform 1 0 16928 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_176
timestamp 1688980957
transform 1 0 17296 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_180
timestamp 1688980957
transform 1 0 17664 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_195
timestamp 1688980957
transform 1 0 19044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_246
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_311
timestamp 1688980957
transform 1 0 29716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_117
timestamp 1688980957
transform 1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_164
timestamp 1688980957
transform 1 0 16192 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_172
timestamp 1688980957
transform 1 0 16928 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_187
timestamp 1688980957
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_214
timestamp 1688980957
transform 1 0 20792 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_226
timestamp 1688980957
transform 1 0 21896 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_237
timestamp 1688980957
transform 1 0 22908 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_247
timestamp 1688980957
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_270
timestamp 1688980957
transform 1 0 25944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_285
timestamp 1688980957
transform 1 0 27324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_291
timestamp 1688980957
transform 1 0 27876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_326
timestamp 1688980957
transform 1 0 31096 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_338
timestamp 1688980957
transform 1 0 32200 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_183
timestamp 1688980957
transform 1 0 17940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_195
timestamp 1688980957
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_203
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_215
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_221
timestamp 1688980957
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_264
timestamp 1688980957
transform 1 0 25392 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1688980957
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_284
timestamp 1688980957
transform 1 0 27232 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_292
timestamp 1688980957
transform 1 0 27968 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_313
timestamp 1688980957
transform 1 0 29900 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_325
timestamp 1688980957
transform 1 0 31004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_330
timestamp 1688980957
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_344
timestamp 1688980957
transform 1 0 32752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_356
timestamp 1688980957
transform 1 0 33856 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_89
timestamp 1688980957
transform 1 0 9292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_100
timestamp 1688980957
transform 1 0 10304 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_108
timestamp 1688980957
transform 1 0 11040 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_115
timestamp 1688980957
transform 1 0 11684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_127
timestamp 1688980957
transform 1 0 12788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_145
timestamp 1688980957
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_169
timestamp 1688980957
transform 1 0 16652 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_182
timestamp 1688980957
transform 1 0 17848 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_222
timestamp 1688980957
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_228
timestamp 1688980957
transform 1 0 22080 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_240
timestamp 1688980957
transform 1 0 23184 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_247
timestamp 1688980957
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_256
timestamp 1688980957
transform 1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_267
timestamp 1688980957
transform 1 0 25668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_339
timestamp 1688980957
transform 1 0 32292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_352
timestamp 1688980957
transform 1 0 33488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_360
timestamp 1688980957
transform 1 0 34224 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_38
timestamp 1688980957
transform 1 0 4600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_75
timestamp 1688980957
transform 1 0 8004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_102
timestamp 1688980957
transform 1 0 10488 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_127
timestamp 1688980957
transform 1 0 12788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_138
timestamp 1688980957
transform 1 0 13800 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_186
timestamp 1688980957
transform 1 0 18216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_209
timestamp 1688980957
transform 1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_230
timestamp 1688980957
transform 1 0 22264 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_236
timestamp 1688980957
transform 1 0 22816 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_246
timestamp 1688980957
transform 1 0 23736 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_255
timestamp 1688980957
transform 1 0 24564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_267
timestamp 1688980957
transform 1 0 25668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_276
timestamp 1688980957
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_290
timestamp 1688980957
transform 1 0 27784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_302
timestamp 1688980957
transform 1 0 28888 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_325
timestamp 1688980957
transform 1 0 31004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_333
timestamp 1688980957
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_45
timestamp 1688980957
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_50
timestamp 1688980957
transform 1 0 5704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_64
timestamp 1688980957
transform 1 0 6992 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_79
timestamp 1688980957
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_91
timestamp 1688980957
transform 1 0 9476 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_115
timestamp 1688980957
transform 1 0 11684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_119
timestamp 1688980957
transform 1 0 12052 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_188
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_229
timestamp 1688980957
transform 1 0 22172 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_268
timestamp 1688980957
transform 1 0 25760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_286
timestamp 1688980957
transform 1 0 27416 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_306
timestamp 1688980957
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_329
timestamp 1688980957
transform 1 0 31372 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_341
timestamp 1688980957
transform 1 0 32476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_29
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_37
timestamp 1688980957
transform 1 0 4508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_65
timestamp 1688980957
transform 1 0 7084 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_77
timestamp 1688980957
transform 1 0 8188 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_89
timestamp 1688980957
transform 1 0 9292 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_101
timestamp 1688980957
transform 1 0 10396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1688980957
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_208
timestamp 1688980957
transform 1 0 20240 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_220
timestamp 1688980957
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_240
timestamp 1688980957
transform 1 0 23184 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_252
timestamp 1688980957
transform 1 0 24288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_277
timestamp 1688980957
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_290
timestamp 1688980957
transform 1 0 27784 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_301
timestamp 1688980957
transform 1 0 28796 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_313
timestamp 1688980957
transform 1 0 29900 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_323
timestamp 1688980957
transform 1 0 30820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_352
timestamp 1688980957
transform 1 0 33488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_360
timestamp 1688980957
transform 1 0 34224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_23
timestamp 1688980957
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_37
timestamp 1688980957
transform 1 0 4508 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_49
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_63
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_94
timestamp 1688980957
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_102
timestamp 1688980957
transform 1 0 10488 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_114
timestamp 1688980957
transform 1 0 11592 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_122
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1688980957
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_170
timestamp 1688980957
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_182
timestamp 1688980957
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_218
timestamp 1688980957
transform 1 0 21160 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_230
timestamp 1688980957
transform 1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_237
timestamp 1688980957
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_242
timestamp 1688980957
transform 1 0 23368 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_248
timestamp 1688980957
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_323
timestamp 1688980957
transform 1 0 30820 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_340
timestamp 1688980957
transform 1 0 32384 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_352
timestamp 1688980957
transform 1 0 33488 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_360
timestamp 1688980957
transform 1 0 34224 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_32
timestamp 1688980957
transform 1 0 4048 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_44
timestamp 1688980957
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_141
timestamp 1688980957
transform 1 0 14076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_153
timestamp 1688980957
transform 1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_158
timestamp 1688980957
transform 1 0 15640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_162
timestamp 1688980957
transform 1 0 16008 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_203
timestamp 1688980957
transform 1 0 19780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_214
timestamp 1688980957
transform 1 0 20792 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_241
timestamp 1688980957
transform 1 0 23276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_253
timestamp 1688980957
transform 1 0 24380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_264
timestamp 1688980957
transform 1 0 25392 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_276
timestamp 1688980957
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_319
timestamp 1688980957
transform 1 0 30452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_333
timestamp 1688980957
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_21
timestamp 1688980957
transform 1 0 3036 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_48
timestamp 1688980957
transform 1 0 5520 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp 1688980957
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_92
timestamp 1688980957
transform 1 0 9568 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_104
timestamp 1688980957
transform 1 0 10672 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_113
timestamp 1688980957
transform 1 0 11500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_191
timestamp 1688980957
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_205
timestamp 1688980957
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_217
timestamp 1688980957
transform 1 0 21068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_236
timestamp 1688980957
transform 1 0 22816 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_273
timestamp 1688980957
transform 1 0 26220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_304
timestamp 1688980957
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_322
timestamp 1688980957
transform 1 0 30728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_340
timestamp 1688980957
transform 1 0 32384 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_358
timestamp 1688980957
transform 1 0 34040 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_85
timestamp 1688980957
transform 1 0 8924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_89
timestamp 1688980957
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_101
timestamp 1688980957
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_163
timestamp 1688980957
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_173
timestamp 1688980957
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_179
timestamp 1688980957
transform 1 0 17572 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_191
timestamp 1688980957
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_203
timestamp 1688980957
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_215
timestamp 1688980957
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_240
timestamp 1688980957
transform 1 0 23184 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_244
timestamp 1688980957
transform 1 0 23552 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_259
timestamp 1688980957
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_271
timestamp 1688980957
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_287
timestamp 1688980957
transform 1 0 27508 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_301
timestamp 1688980957
transform 1 0 28796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_313
timestamp 1688980957
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_325
timestamp 1688980957
transform 1 0 31004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_329
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_360
timestamp 1688980957
transform 1 0 34224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_6
timestamp 1688980957
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_18
timestamp 1688980957
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_35
timestamp 1688980957
transform 1 0 4324 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_43
timestamp 1688980957
transform 1 0 5060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_49
timestamp 1688980957
transform 1 0 5612 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_62
timestamp 1688980957
transform 1 0 6808 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_70
timestamp 1688980957
transform 1 0 7544 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_101
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_262
timestamp 1688980957
transform 1 0 25208 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_268
timestamp 1688980957
transform 1 0 25760 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_289
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_299
timestamp 1688980957
transform 1 0 28612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_315
timestamp 1688980957
transform 1 0 30084 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_361
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_23
timestamp 1688980957
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_66
timestamp 1688980957
transform 1 0 7176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_74
timestamp 1688980957
transform 1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_90
timestamp 1688980957
transform 1 0 9384 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_99
timestamp 1688980957
transform 1 0 10212 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1688980957
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_118
timestamp 1688980957
transform 1 0 11960 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_126
timestamp 1688980957
transform 1 0 12696 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_142
timestamp 1688980957
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1688980957
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_198
timestamp 1688980957
transform 1 0 19320 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_206
timestamp 1688980957
transform 1 0 20056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_214
timestamp 1688980957
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_268
timestamp 1688980957
transform 1 0 25760 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_284
timestamp 1688980957
transform 1 0 27232 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_290
timestamp 1688980957
transform 1 0 27784 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_300
timestamp 1688980957
transform 1 0 28704 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_312
timestamp 1688980957
transform 1 0 29808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_322
timestamp 1688980957
transform 1 0 30728 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_331
timestamp 1688980957
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_342
timestamp 1688980957
transform 1 0 32568 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_354
timestamp 1688980957
transform 1 0 33672 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_35
timestamp 1688980957
transform 1 0 4324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_57
timestamp 1688980957
transform 1 0 6348 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_63
timestamp 1688980957
transform 1 0 6900 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_105
timestamp 1688980957
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_115
timestamp 1688980957
transform 1 0 11684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_123
timestamp 1688980957
transform 1 0 12420 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1688980957
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_149
timestamp 1688980957
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_167
timestamp 1688980957
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_171
timestamp 1688980957
transform 1 0 16836 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_178
timestamp 1688980957
transform 1 0 17480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_191
timestamp 1688980957
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_211
timestamp 1688980957
transform 1 0 20516 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_217
timestamp 1688980957
transform 1 0 21068 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_228
timestamp 1688980957
transform 1 0 22080 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_232
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_246
timestamp 1688980957
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_278
timestamp 1688980957
transform 1 0 26680 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_342
timestamp 1688980957
transform 1 0 32568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_354
timestamp 1688980957
transform 1 0 33672 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 1688980957
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_61
timestamp 1688980957
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_71
timestamp 1688980957
transform 1 0 7636 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_77
timestamp 1688980957
transform 1 0 8188 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_85
timestamp 1688980957
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_95
timestamp 1688980957
transform 1 0 9844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_103
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_124
timestamp 1688980957
transform 1 0 12512 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_145
timestamp 1688980957
transform 1 0 14444 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_153
timestamp 1688980957
transform 1 0 15180 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_159
timestamp 1688980957
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_176
timestamp 1688980957
transform 1 0 17296 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_190
timestamp 1688980957
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_194
timestamp 1688980957
transform 1 0 18952 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_233
timestamp 1688980957
transform 1 0 22540 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_251
timestamp 1688980957
transform 1 0 24196 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_263
timestamp 1688980957
transform 1 0 25300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_267
timestamp 1688980957
transform 1 0 25668 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_300
timestamp 1688980957
transform 1 0 28704 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_312
timestamp 1688980957
transform 1 0 29808 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_320
timestamp 1688980957
transform 1 0 30544 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_345
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_357
timestamp 1688980957
transform 1 0 33948 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_72
timestamp 1688980957
transform 1 0 7728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_96
timestamp 1688980957
transform 1 0 9936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_118
timestamp 1688980957
transform 1 0 11960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_147
timestamp 1688980957
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_178
timestamp 1688980957
transform 1 0 17480 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_185
timestamp 1688980957
transform 1 0 18124 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_206
timestamp 1688980957
transform 1 0 20056 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_214
timestamp 1688980957
transform 1 0 20792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_229
timestamp 1688980957
transform 1 0 22172 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_246
timestamp 1688980957
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_288
timestamp 1688980957
transform 1 0 27600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_298
timestamp 1688980957
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_361
timestamp 1688980957
transform 1 0 34316 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_24
timestamp 1688980957
transform 1 0 3312 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_32
timestamp 1688980957
transform 1 0 4048 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_82
timestamp 1688980957
transform 1 0 8648 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_96
timestamp 1688980957
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1688980957
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_134
timestamp 1688980957
transform 1 0 13432 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_146
timestamp 1688980957
transform 1 0 14536 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_152
timestamp 1688980957
transform 1 0 15088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_159
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_185
timestamp 1688980957
transform 1 0 18124 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_207
timestamp 1688980957
transform 1 0 20148 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_219
timestamp 1688980957
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_234
timestamp 1688980957
transform 1 0 22632 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_270
timestamp 1688980957
transform 1 0 25944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_303
timestamp 1688980957
transform 1 0 28980 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_307
timestamp 1688980957
transform 1 0 29348 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_316
timestamp 1688980957
transform 1 0 30176 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_331
timestamp 1688980957
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_346
timestamp 1688980957
transform 1 0 32936 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_358
timestamp 1688980957
transform 1 0 34040 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_25
timestamp 1688980957
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1688980957
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_183
timestamp 1688980957
transform 1 0 17940 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_187
timestamp 1688980957
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_211
timestamp 1688980957
transform 1 0 20516 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_219
timestamp 1688980957
transform 1 0 21252 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_226
timestamp 1688980957
transform 1 0 21896 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_232
timestamp 1688980957
transform 1 0 22448 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_238
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_250
timestamp 1688980957
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_262
timestamp 1688980957
transform 1 0 25208 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_268
timestamp 1688980957
transform 1 0 25760 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_297
timestamp 1688980957
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_317
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_334
timestamp 1688980957
transform 1 0 31832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_343
timestamp 1688980957
transform 1 0 32660 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_359
timestamp 1688980957
transform 1 0 34132 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_31
timestamp 1688980957
transform 1 0 3956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_48
timestamp 1688980957
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_65
timestamp 1688980957
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_87
timestamp 1688980957
transform 1 0 9108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_95
timestamp 1688980957
transform 1 0 9844 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_103
timestamp 1688980957
transform 1 0 10580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_140
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_148
timestamp 1688980957
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_160
timestamp 1688980957
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_213
timestamp 1688980957
transform 1 0 20700 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_219
timestamp 1688980957
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_302
timestamp 1688980957
transform 1 0 28888 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_310
timestamp 1688980957
transform 1 0 29624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_319
timestamp 1688980957
transform 1 0 30452 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_332
timestamp 1688980957
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_353
timestamp 1688980957
transform 1 0 33580 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_357
timestamp 1688980957
transform 1 0 33948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_23
timestamp 1688980957
transform 1 0 3220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_39
timestamp 1688980957
transform 1 0 4692 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_59
timestamp 1688980957
transform 1 0 6532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_94
timestamp 1688980957
transform 1 0 9752 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_102
timestamp 1688980957
transform 1 0 10488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_120
timestamp 1688980957
transform 1 0 12144 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_128
timestamp 1688980957
transform 1 0 12880 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_145
timestamp 1688980957
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_150
timestamp 1688980957
transform 1 0 14904 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_158
timestamp 1688980957
transform 1 0 15640 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_179
timestamp 1688980957
transform 1 0 17572 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_190
timestamp 1688980957
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_210
timestamp 1688980957
transform 1 0 20424 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_214
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_224
timestamp 1688980957
transform 1 0 21712 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_232
timestamp 1688980957
transform 1 0 22448 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_245
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_262
timestamp 1688980957
transform 1 0 25208 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_268
timestamp 1688980957
transform 1 0 25760 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_281
timestamp 1688980957
transform 1 0 26956 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_289
timestamp 1688980957
transform 1 0 27692 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1688980957
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_329
timestamp 1688980957
transform 1 0 31372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_353
timestamp 1688980957
transform 1 0 33580 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_361
timestamp 1688980957
transform 1 0 34316 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_23
timestamp 1688980957
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_32
timestamp 1688980957
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_96
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_108
timestamp 1688980957
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_117
timestamp 1688980957
transform 1 0 11868 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_123
timestamp 1688980957
transform 1 0 12420 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_157
timestamp 1688980957
transform 1 0 15548 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1688980957
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_177
timestamp 1688980957
transform 1 0 17388 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_187
timestamp 1688980957
transform 1 0 18308 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_209
timestamp 1688980957
transform 1 0 20332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1688980957
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_271
timestamp 1688980957
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_291
timestamp 1688980957
transform 1 0 27876 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_321
timestamp 1688980957
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_333
timestamp 1688980957
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_346
timestamp 1688980957
transform 1 0 32936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_358
timestamp 1688980957
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_82
timestamp 1688980957
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_99
timestamp 1688980957
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1688980957
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_183
timestamp 1688980957
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_187
timestamp 1688980957
transform 1 0 18308 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1688980957
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_203
timestamp 1688980957
transform 1 0 19780 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_213
timestamp 1688980957
transform 1 0 20700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_243
timestamp 1688980957
transform 1 0 23460 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_247
timestamp 1688980957
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_256
timestamp 1688980957
transform 1 0 24656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_268
timestamp 1688980957
transform 1 0 25760 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_283
timestamp 1688980957
transform 1 0 27140 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_306
timestamp 1688980957
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_336
timestamp 1688980957
transform 1 0 32016 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_355
timestamp 1688980957
transform 1 0 33764 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_361
timestamp 1688980957
transform 1 0 34316 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_23
timestamp 1688980957
transform 1 0 3220 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_31
timestamp 1688980957
transform 1 0 3956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_48
timestamp 1688980957
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_71
timestamp 1688980957
transform 1 0 7636 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_79
timestamp 1688980957
transform 1 0 8372 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_88
timestamp 1688980957
transform 1 0 9200 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_100
timestamp 1688980957
transform 1 0 10304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_133
timestamp 1688980957
transform 1 0 13340 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_154
timestamp 1688980957
transform 1 0 15272 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1688980957
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_203
timestamp 1688980957
transform 1 0 19780 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_263
timestamp 1688980957
transform 1 0 25300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_275
timestamp 1688980957
transform 1 0 26404 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_301
timestamp 1688980957
transform 1 0 28796 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_313
timestamp 1688980957
transform 1 0 29900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_320
timestamp 1688980957
transform 1 0 30544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_324
timestamp 1688980957
transform 1 0 30912 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_334
timestamp 1688980957
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_341
timestamp 1688980957
transform 1 0 32476 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_6
timestamp 1688980957
transform 1 0 1656 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_14
timestamp 1688980957
transform 1 0 2392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_20
timestamp 1688980957
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_38
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_42
timestamp 1688980957
transform 1 0 4968 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_54
timestamp 1688980957
transform 1 0 6072 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_62
timestamp 1688980957
transform 1 0 6808 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_71
timestamp 1688980957
transform 1 0 7636 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_79
timestamp 1688980957
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_92
timestamp 1688980957
transform 1 0 9568 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_99
timestamp 1688980957
transform 1 0 10212 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_103
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_108
timestamp 1688980957
transform 1 0 11040 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_120
timestamp 1688980957
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_135
timestamp 1688980957
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_171
timestamp 1688980957
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_185
timestamp 1688980957
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_218
timestamp 1688980957
transform 1 0 21160 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_230
timestamp 1688980957
transform 1 0 22264 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_236
timestamp 1688980957
transform 1 0 22816 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_242
timestamp 1688980957
transform 1 0 23368 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_259
timestamp 1688980957
transform 1 0 24932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_272
timestamp 1688980957
transform 1 0 26128 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_278
timestamp 1688980957
transform 1 0 26680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_287
timestamp 1688980957
transform 1 0 27508 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_302
timestamp 1688980957
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_319
timestamp 1688980957
transform 1 0 30452 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_331
timestamp 1688980957
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_343
timestamp 1688980957
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_355
timestamp 1688980957
transform 1 0 33764 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_361
timestamp 1688980957
transform 1 0 34316 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_52
timestamp 1688980957
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_76
timestamp 1688980957
transform 1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_92
timestamp 1688980957
transform 1 0 9568 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_117
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_124
timestamp 1688980957
transform 1 0 12512 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_136
timestamp 1688980957
transform 1 0 13616 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_164
timestamp 1688980957
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_173
timestamp 1688980957
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_179
timestamp 1688980957
transform 1 0 17572 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_190
timestamp 1688980957
transform 1 0 18584 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_202
timestamp 1688980957
transform 1 0 19688 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_214
timestamp 1688980957
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1688980957
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_236
timestamp 1688980957
transform 1 0 22816 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_248
timestamp 1688980957
transform 1 0 23920 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_289
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_311
timestamp 1688980957
transform 1 0 29716 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_320
timestamp 1688980957
transform 1 0 30544 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_332
timestamp 1688980957
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_343
timestamp 1688980957
transform 1 0 32660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_353
timestamp 1688980957
transform 1 0 33580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_37
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_56
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_64
timestamp 1688980957
transform 1 0 6992 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_68
timestamp 1688980957
transform 1 0 7360 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_80
timestamp 1688980957
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_93
timestamp 1688980957
transform 1 0 9660 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_186
timestamp 1688980957
transform 1 0 18216 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_205
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_213
timestamp 1688980957
transform 1 0 20700 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_243
timestamp 1688980957
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_261
timestamp 1688980957
transform 1 0 25116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_267
timestamp 1688980957
transform 1 0 25668 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_275
timestamp 1688980957
transform 1 0 26404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_287
timestamp 1688980957
transform 1 0 27508 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_293
timestamp 1688980957
transform 1 0 28060 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_302
timestamp 1688980957
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_329
timestamp 1688980957
transform 1 0 31372 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_341
timestamp 1688980957
transform 1 0 32476 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_47
timestamp 1688980957
transform 1 0 5428 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_65
timestamp 1688980957
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_76
timestamp 1688980957
transform 1 0 8096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_84
timestamp 1688980957
transform 1 0 8832 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_99
timestamp 1688980957
transform 1 0 10212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_119
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_130
timestamp 1688980957
transform 1 0 13064 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_142
timestamp 1688980957
transform 1 0 14168 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_148
timestamp 1688980957
transform 1 0 14720 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_155
timestamp 1688980957
transform 1 0 15364 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1688980957
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_177
timestamp 1688980957
transform 1 0 17388 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_207
timestamp 1688980957
transform 1 0 20148 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_230
timestamp 1688980957
transform 1 0 22264 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_238
timestamp 1688980957
transform 1 0 23000 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_268
timestamp 1688980957
transform 1 0 25760 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_276
timestamp 1688980957
transform 1 0 26496 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_309
timestamp 1688980957
transform 1 0 29532 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_326
timestamp 1688980957
transform 1 0 31096 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_344
timestamp 1688980957
transform 1 0 32752 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_356
timestamp 1688980957
transform 1 0 33856 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_52
timestamp 1688980957
transform 1 0 5888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_61
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_73
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_112
timestamp 1688980957
transform 1 0 11408 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_131
timestamp 1688980957
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_161
timestamp 1688980957
transform 1 0 15916 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_173
timestamp 1688980957
transform 1 0 17020 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_185
timestamp 1688980957
transform 1 0 18124 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_191
timestamp 1688980957
transform 1 0 18676 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_237
timestamp 1688980957
transform 1 0 22908 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1688980957
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_278
timestamp 1688980957
transform 1 0 26680 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_290
timestamp 1688980957
transform 1 0 27784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_294
timestamp 1688980957
transform 1 0 28152 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_303
timestamp 1688980957
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_327
timestamp 1688980957
transform 1 0 31188 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_335
timestamp 1688980957
transform 1 0 31924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_344
timestamp 1688980957
transform 1 0 32752 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_354
timestamp 1688980957
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_63
timestamp 1688980957
transform 1 0 6900 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_87
timestamp 1688980957
transform 1 0 9108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_99
timestamp 1688980957
transform 1 0 10212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_117
timestamp 1688980957
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_141
timestamp 1688980957
transform 1 0 14076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_153
timestamp 1688980957
transform 1 0 15180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_165
timestamp 1688980957
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_174
timestamp 1688980957
transform 1 0 17112 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_185
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_191
timestamp 1688980957
transform 1 0 18676 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_202
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_210
timestamp 1688980957
transform 1 0 20424 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_219
timestamp 1688980957
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_258
timestamp 1688980957
transform 1 0 24840 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_270
timestamp 1688980957
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_278
timestamp 1688980957
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_304
timestamp 1688980957
transform 1 0 29072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_309
timestamp 1688980957
transform 1 0 29532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_316
timestamp 1688980957
transform 1 0 30176 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_324
timestamp 1688980957
transform 1 0 30912 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_330
timestamp 1688980957
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_46
timestamp 1688980957
transform 1 0 5336 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_70
timestamp 1688980957
transform 1 0 7544 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 1688980957
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_99
timestamp 1688980957
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_123
timestamp 1688980957
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_135
timestamp 1688980957
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_183
timestamp 1688980957
transform 1 0 17940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_187
timestamp 1688980957
transform 1 0 18308 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_224
timestamp 1688980957
transform 1 0 21712 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_228
timestamp 1688980957
transform 1 0 22080 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_241
timestamp 1688980957
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_249
timestamp 1688980957
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_260
timestamp 1688980957
transform 1 0 25024 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_272
timestamp 1688980957
transform 1 0 26128 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_305
timestamp 1688980957
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_316
timestamp 1688980957
transform 1 0 30176 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_329
timestamp 1688980957
transform 1 0 31372 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_341
timestamp 1688980957
transform 1 0 32476 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_353
timestamp 1688980957
transform 1 0 33580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_361
timestamp 1688980957
transform 1 0 34316 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_49
timestamp 1688980957
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_62
timestamp 1688980957
transform 1 0 6808 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_74
timestamp 1688980957
transform 1 0 7912 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_100
timestamp 1688980957
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_127
timestamp 1688980957
transform 1 0 12788 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_148
timestamp 1688980957
transform 1 0 14720 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_160
timestamp 1688980957
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_202
timestamp 1688980957
transform 1 0 19688 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_214
timestamp 1688980957
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1688980957
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_251
timestamp 1688980957
transform 1 0 24196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_271
timestamp 1688980957
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_290
timestamp 1688980957
transform 1 0 27784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_299
timestamp 1688980957
transform 1 0 28612 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_307
timestamp 1688980957
transform 1 0 29348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_318
timestamp 1688980957
transform 1 0 30360 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_330
timestamp 1688980957
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_350
timestamp 1688980957
transform 1 0 33304 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_44
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_76
timestamp 1688980957
transform 1 0 8096 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_120
timestamp 1688980957
transform 1 0 12144 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_132
timestamp 1688980957
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_159
timestamp 1688980957
transform 1 0 15732 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_171
timestamp 1688980957
transform 1 0 16836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_182
timestamp 1688980957
transform 1 0 17848 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_186
timestamp 1688980957
transform 1 0 18216 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_194
timestamp 1688980957
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_204
timestamp 1688980957
transform 1 0 19872 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_216
timestamp 1688980957
transform 1 0 20976 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_220
timestamp 1688980957
transform 1 0 21344 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_232
timestamp 1688980957
transform 1 0 22448 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_244
timestamp 1688980957
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_275
timestamp 1688980957
transform 1 0 26404 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_292
timestamp 1688980957
transform 1 0 27968 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_304
timestamp 1688980957
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_320
timestamp 1688980957
transform 1 0 30544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_324
timestamp 1688980957
transform 1 0 30912 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_337
timestamp 1688980957
transform 1 0 32108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_341
timestamp 1688980957
transform 1 0 32476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_7
timestamp 1688980957
transform 1 0 1748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_28
timestamp 1688980957
transform 1 0 3680 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_33
timestamp 1688980957
transform 1 0 4140 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_45
timestamp 1688980957
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_64
timestamp 1688980957
transform 1 0 6992 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_92
timestamp 1688980957
transform 1 0 9568 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_98
timestamp 1688980957
transform 1 0 10120 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_129
timestamp 1688980957
transform 1 0 12972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_141
timestamp 1688980957
transform 1 0 14076 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_147
timestamp 1688980957
transform 1 0 14628 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_189
timestamp 1688980957
transform 1 0 18492 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_197
timestamp 1688980957
transform 1 0 19228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_201
timestamp 1688980957
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_213
timestamp 1688980957
transform 1 0 20700 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_257
timestamp 1688980957
transform 1 0 24748 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_269
timestamp 1688980957
transform 1 0 25852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 1688980957
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_295
timestamp 1688980957
transform 1 0 28244 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_307
timestamp 1688980957
transform 1 0 29348 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_323
timestamp 1688980957
transform 1 0 30820 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_37
timestamp 1688980957
transform 1 0 4508 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_43
timestamp 1688980957
transform 1 0 5060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_55
timestamp 1688980957
transform 1 0 6164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_69
timestamp 1688980957
transform 1 0 7452 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_82
timestamp 1688980957
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_170
timestamp 1688980957
transform 1 0 16744 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_218
timestamp 1688980957
transform 1 0 21160 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_230
timestamp 1688980957
transform 1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_242
timestamp 1688980957
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 1688980957
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_267
timestamp 1688980957
transform 1 0 25668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_291
timestamp 1688980957
transform 1 0 27876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_299
timestamp 1688980957
transform 1 0 28612 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_306
timestamp 1688980957
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_318
timestamp 1688980957
transform 1 0 30360 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_324
timestamp 1688980957
transform 1 0 30912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_332
timestamp 1688980957
transform 1 0 31648 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_342
timestamp 1688980957
transform 1 0 32568 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_353
timestamp 1688980957
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_361
timestamp 1688980957
transform 1 0 34316 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_36
timestamp 1688980957
transform 1 0 4416 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_44
timestamp 1688980957
transform 1 0 5152 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_54
timestamp 1688980957
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_65
timestamp 1688980957
transform 1 0 7084 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_71
timestamp 1688980957
transform 1 0 7636 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_91
timestamp 1688980957
transform 1 0 9476 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_103
timestamp 1688980957
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_119
timestamp 1688980957
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_127
timestamp 1688980957
transform 1 0 12788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_139
timestamp 1688980957
transform 1 0 13892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_147
timestamp 1688980957
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_159
timestamp 1688980957
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_234
timestamp 1688980957
transform 1 0 22632 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_238
timestamp 1688980957
transform 1 0 23000 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_259
timestamp 1688980957
transform 1 0 24932 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_291
timestamp 1688980957
transform 1 0 27876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_303
timestamp 1688980957
transform 1 0 28980 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_311
timestamp 1688980957
transform 1 0 29716 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_319
timestamp 1688980957
transform 1 0 30452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_331
timestamp 1688980957
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_343
timestamp 1688980957
transform 1 0 32660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_355
timestamp 1688980957
transform 1 0 33764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_9
timestamp 1688980957
transform 1 0 1932 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_21
timestamp 1688980957
transform 1 0 3036 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_49
timestamp 1688980957
transform 1 0 5612 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_60
timestamp 1688980957
transform 1 0 6624 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_107
timestamp 1688980957
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_119
timestamp 1688980957
transform 1 0 12052 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_126
timestamp 1688980957
transform 1 0 12696 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_138
timestamp 1688980957
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_159
timestamp 1688980957
transform 1 0 15732 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_180
timestamp 1688980957
transform 1 0 17664 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_192
timestamp 1688980957
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_207
timestamp 1688980957
transform 1 0 20148 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_215
timestamp 1688980957
transform 1 0 20884 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_247
timestamp 1688980957
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_261
timestamp 1688980957
transform 1 0 25116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_283
timestamp 1688980957
transform 1 0 27140 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_293
timestamp 1688980957
transform 1 0 28060 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_324
timestamp 1688980957
transform 1 0 30912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_354
timestamp 1688980957
transform 1 0 33672 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_63
timestamp 1688980957
transform 1 0 6900 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_70
timestamp 1688980957
transform 1 0 7544 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_82
timestamp 1688980957
transform 1 0 8648 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_90
timestamp 1688980957
transform 1 0 9384 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_118
timestamp 1688980957
transform 1 0 11960 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_127
timestamp 1688980957
transform 1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_158
timestamp 1688980957
transform 1 0 15640 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_173
timestamp 1688980957
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_228
timestamp 1688980957
transform 1 0 22080 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_236
timestamp 1688980957
transform 1 0 22816 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_266
timestamp 1688980957
transform 1 0 25576 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 1688980957
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_316
timestamp 1688980957
transform 1 0 30176 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_328
timestamp 1688980957
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_64
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_76
timestamp 1688980957
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_101
timestamp 1688980957
transform 1 0 10396 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_107
timestamp 1688980957
transform 1 0 10948 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_114
timestamp 1688980957
transform 1 0 11592 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_146
timestamp 1688980957
transform 1 0 14536 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_152
timestamp 1688980957
transform 1 0 15088 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_166
timestamp 1688980957
transform 1 0 16376 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_172
timestamp 1688980957
transform 1 0 16928 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_184
timestamp 1688980957
transform 1 0 18032 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1688980957
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_200
timestamp 1688980957
transform 1 0 19504 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_208
timestamp 1688980957
transform 1 0 20240 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_231
timestamp 1688980957
transform 1 0 22356 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_239
timestamp 1688980957
transform 1 0 23092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_264
timestamp 1688980957
transform 1 0 25392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_268
timestamp 1688980957
transform 1 0 25760 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_292
timestamp 1688980957
transform 1 0 27968 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_305
timestamp 1688980957
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_25
timestamp 1688980957
transform 1 0 3404 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_30
timestamp 1688980957
transform 1 0 3864 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_42
timestamp 1688980957
transform 1 0 4968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_49
timestamp 1688980957
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_85
timestamp 1688980957
transform 1 0 8924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_97
timestamp 1688980957
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_109
timestamp 1688980957
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_245
timestamp 1688980957
transform 1 0 23644 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_275
timestamp 1688980957
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_297
timestamp 1688980957
transform 1 0 28428 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_309
timestamp 1688980957
transform 1 0 29532 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_328
timestamp 1688980957
transform 1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_357
timestamp 1688980957
transform 1 0 33948 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_19
timestamp 1688980957
transform 1 0 2852 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_55
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_105
timestamp 1688980957
transform 1 0 10764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_117
timestamp 1688980957
transform 1 0 11868 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_129
timestamp 1688980957
transform 1 0 12972 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_137
timestamp 1688980957
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_162
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_168
timestamp 1688980957
transform 1 0 16560 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_174
timestamp 1688980957
transform 1 0 17112 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_186
timestamp 1688980957
transform 1 0 18216 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_193
timestamp 1688980957
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_206
timestamp 1688980957
transform 1 0 20056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_218
timestamp 1688980957
transform 1 0 21160 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_261
timestamp 1688980957
transform 1 0 25116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_273
timestamp 1688980957
transform 1 0 26220 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_280
timestamp 1688980957
transform 1 0 26864 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_292
timestamp 1688980957
transform 1 0 27968 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_322
timestamp 1688980957
transform 1 0 30728 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_334
timestamp 1688980957
transform 1 0 31832 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_346
timestamp 1688980957
transform 1 0 32936 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_358
timestamp 1688980957
transform 1 0 34040 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_23
timestamp 1688980957
transform 1 0 3220 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_33
timestamp 1688980957
transform 1 0 4140 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_45
timestamp 1688980957
transform 1 0 5244 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_54
timestamp 1688980957
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_92
timestamp 1688980957
transform 1 0 9568 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_106
timestamp 1688980957
transform 1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_133
timestamp 1688980957
transform 1 0 13340 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_163
timestamp 1688980957
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_175
timestamp 1688980957
transform 1 0 17204 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_197
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_209
timestamp 1688980957
transform 1 0 20332 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_229
timestamp 1688980957
transform 1 0 22172 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_233
timestamp 1688980957
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_243
timestamp 1688980957
transform 1 0 23460 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_251
timestamp 1688980957
transform 1 0 24196 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_275
timestamp 1688980957
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_330
timestamp 1688980957
transform 1 0 31464 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_49
timestamp 1688980957
transform 1 0 5612 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_61
timestamp 1688980957
transform 1 0 6716 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_73
timestamp 1688980957
transform 1 0 7820 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_91
timestamp 1688980957
transform 1 0 9476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_119
timestamp 1688980957
transform 1 0 12052 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_130
timestamp 1688980957
transform 1 0 13064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_134
timestamp 1688980957
transform 1 0 13432 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_155
timestamp 1688980957
transform 1 0 15364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_186
timestamp 1688980957
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_190
timestamp 1688980957
transform 1 0 18584 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_194
timestamp 1688980957
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_203
timestamp 1688980957
transform 1 0 19780 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_208
timestamp 1688980957
transform 1 0 20240 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_219
timestamp 1688980957
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_231
timestamp 1688980957
transform 1 0 22356 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_237
timestamp 1688980957
transform 1 0 22908 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_247
timestamp 1688980957
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_275
timestamp 1688980957
transform 1 0 26404 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_287
timestamp 1688980957
transform 1 0 27508 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_299
timestamp 1688980957
transform 1 0 28612 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_325
timestamp 1688980957
transform 1 0 31004 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_337
timestamp 1688980957
transform 1 0 32108 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_349
timestamp 1688980957
transform 1 0 33212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_361
timestamp 1688980957
transform 1 0 34316 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_77
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_98
timestamp 1688980957
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_110
timestamp 1688980957
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_133
timestamp 1688980957
transform 1 0 13340 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_143
timestamp 1688980957
transform 1 0 14260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_151
timestamp 1688980957
transform 1 0 14996 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_160
timestamp 1688980957
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_209
timestamp 1688980957
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_257
timestamp 1688980957
transform 1 0 24748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_277
timestamp 1688980957
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_289
timestamp 1688980957
transform 1 0 27692 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_312
timestamp 1688980957
transform 1 0 29808 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_324
timestamp 1688980957
transform 1 0 30912 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_96
timestamp 1688980957
transform 1 0 9936 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_108
timestamp 1688980957
transform 1 0 11040 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_116
timestamp 1688980957
transform 1 0 11776 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_174
timestamp 1688980957
transform 1 0 17112 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_184
timestamp 1688980957
transform 1 0 18032 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_200
timestamp 1688980957
transform 1 0 19504 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_212
timestamp 1688980957
transform 1 0 20608 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_223
timestamp 1688980957
transform 1 0 21620 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_235
timestamp 1688980957
transform 1 0 22724 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_247
timestamp 1688980957
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_361
timestamp 1688980957
transform 1 0 34316 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_38
timestamp 1688980957
transform 1 0 4600 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_54
timestamp 1688980957
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_66
timestamp 1688980957
transform 1 0 7176 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_78
timestamp 1688980957
transform 1 0 8280 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_89
timestamp 1688980957
transform 1 0 9292 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_99
timestamp 1688980957
transform 1 0 10212 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_104
timestamp 1688980957
transform 1 0 10672 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_145
timestamp 1688980957
transform 1 0 14444 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_158
timestamp 1688980957
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_166
timestamp 1688980957
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_173
timestamp 1688980957
transform 1 0 17020 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_183
timestamp 1688980957
transform 1 0 17940 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_195
timestamp 1688980957
transform 1 0 19044 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_200
timestamp 1688980957
transform 1 0 19504 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_206
timestamp 1688980957
transform 1 0 20056 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_211
timestamp 1688980957
transform 1 0 20516 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_221
timestamp 1688980957
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_236
timestamp 1688980957
transform 1 0 22816 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_246
timestamp 1688980957
transform 1 0 23736 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_254
timestamp 1688980957
transform 1 0 24472 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_260
timestamp 1688980957
transform 1 0 25024 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_272
timestamp 1688980957
transform 1 0 26128 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_11
timestamp 1688980957
transform 1 0 2116 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_16
timestamp 1688980957
transform 1 0 2576 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_58
timestamp 1688980957
transform 1 0 6440 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_70
timestamp 1688980957
transform 1 0 7544 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_125
timestamp 1688980957
transform 1 0 12604 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_129
timestamp 1688980957
transform 1 0 12972 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_146
timestamp 1688980957
transform 1 0 14536 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_158
timestamp 1688980957
transform 1 0 15640 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_170
timestamp 1688980957
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_182
timestamp 1688980957
transform 1 0 17848 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_186
timestamp 1688980957
transform 1 0 18216 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_207
timestamp 1688980957
transform 1 0 20148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_219
timestamp 1688980957
transform 1 0 21252 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_247
timestamp 1688980957
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_261
timestamp 1688980957
transform 1 0 25116 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_273
timestamp 1688980957
transform 1 0 26220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_286
timestamp 1688980957
transform 1 0 27416 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_303
timestamp 1688980957
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_357
timestamp 1688980957
transform 1 0 33948 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_361
timestamp 1688980957
transform 1 0 34316 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_7
timestamp 1688980957
transform 1 0 1748 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_35
timestamp 1688980957
transform 1 0 4324 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_41
timestamp 1688980957
transform 1 0 4876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_53
timestamp 1688980957
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_67
timestamp 1688980957
transform 1 0 7268 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_80
timestamp 1688980957
transform 1 0 8464 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_84
timestamp 1688980957
transform 1 0 8832 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_92
timestamp 1688980957
transform 1 0 9568 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_104
timestamp 1688980957
transform 1 0 10672 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_121
timestamp 1688980957
transform 1 0 12236 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_159
timestamp 1688980957
transform 1 0 15732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_182
timestamp 1688980957
transform 1 0 17848 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_194
timestamp 1688980957
transform 1 0 18952 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_201
timestamp 1688980957
transform 1 0 19596 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_243
timestamp 1688980957
transform 1 0 23460 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_271
timestamp 1688980957
transform 1 0 26036 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_275
timestamp 1688980957
transform 1 0 26404 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_321
timestamp 1688980957
transform 1 0 30636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_333
timestamp 1688980957
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_9
timestamp 1688980957
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_21
timestamp 1688980957
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_35
timestamp 1688980957
transform 1 0 4324 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_47
timestamp 1688980957
transform 1 0 5428 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_61
timestamp 1688980957
transform 1 0 6716 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_73
timestamp 1688980957
transform 1 0 7820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_105
timestamp 1688980957
transform 1 0 10764 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_117
timestamp 1688980957
transform 1 0 11868 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_131
timestamp 1688980957
transform 1 0 13156 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_147
timestamp 1688980957
transform 1 0 14628 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_172
timestamp 1688980957
transform 1 0 16928 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_183
timestamp 1688980957
transform 1 0 17940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_205
timestamp 1688980957
transform 1 0 19964 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_217
timestamp 1688980957
transform 1 0 21068 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_225
timestamp 1688980957
transform 1 0 21804 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_230
timestamp 1688980957
transform 1 0 22264 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_241
timestamp 1688980957
transform 1 0 23276 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_249
timestamp 1688980957
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_264
timestamp 1688980957
transform 1 0 25392 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_272
timestamp 1688980957
transform 1 0 26128 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_282
timestamp 1688980957
transform 1 0 27048 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_294
timestamp 1688980957
transform 1 0 28152 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_306
timestamp 1688980957
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_341
timestamp 1688980957
transform 1 0 32476 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_43
timestamp 1688980957
transform 1 0 5060 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_70
timestamp 1688980957
transform 1 0 7544 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_82
timestamp 1688980957
transform 1 0 8648 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_87
timestamp 1688980957
transform 1 0 9108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_99
timestamp 1688980957
transform 1 0 10212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_183
timestamp 1688980957
transform 1 0 17940 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_202
timestamp 1688980957
transform 1 0 19688 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_220
timestamp 1688980957
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_245
timestamp 1688980957
transform 1 0 23644 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_257
timestamp 1688980957
transform 1 0 24748 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_267
timestamp 1688980957
transform 1 0 25668 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_278
timestamp 1688980957
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_45
timestamp 1688980957
transform 1 0 5244 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_66
timestamp 1688980957
transform 1 0 7176 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_81
timestamp 1688980957
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_151
timestamp 1688980957
transform 1 0 14996 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_174
timestamp 1688980957
transform 1 0 17112 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_185
timestamp 1688980957
transform 1 0 18124 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_201
timestamp 1688980957
transform 1 0 19596 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_214
timestamp 1688980957
transform 1 0 20792 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_226
timestamp 1688980957
transform 1 0 21896 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_234
timestamp 1688980957
transform 1 0 22632 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_240
timestamp 1688980957
transform 1 0 23184 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_259
timestamp 1688980957
transform 1 0 24932 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_291
timestamp 1688980957
transform 1 0 27876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_303
timestamp 1688980957
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_353
timestamp 1688980957
transform 1 0 33580 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_47
timestamp 1688980957
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_65
timestamp 1688980957
transform 1 0 7084 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_91
timestamp 1688980957
transform 1 0 9476 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_121
timestamp 1688980957
transform 1 0 12236 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_197
timestamp 1688980957
transform 1 0 19228 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_251
timestamp 1688980957
transform 1 0 24196 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_272
timestamp 1688980957
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_357
timestamp 1688980957
transform 1 0 33948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_9
timestamp 1688980957
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_21
timestamp 1688980957
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_57
timestamp 1688980957
transform 1 0 6348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_69
timestamp 1688980957
transform 1 0 7452 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_73
timestamp 1688980957
transform 1 0 7820 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_80
timestamp 1688980957
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_113
timestamp 1688980957
transform 1 0 11500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_125
timestamp 1688980957
transform 1 0 12604 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_167
timestamp 1688980957
transform 1 0 16468 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_175
timestamp 1688980957
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_187
timestamp 1688980957
transform 1 0 18308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_205
timestamp 1688980957
transform 1 0 19964 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_210
timestamp 1688980957
transform 1 0 20424 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_222
timestamp 1688980957
transform 1 0 21528 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_234
timestamp 1688980957
transform 1 0 22632 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_246
timestamp 1688980957
transform 1 0 23736 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_287
timestamp 1688980957
transform 1 0 27508 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_299
timestamp 1688980957
transform 1 0 28612 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_337
timestamp 1688980957
transform 1 0 32108 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_349
timestamp 1688980957
transform 1 0 33212 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_361
timestamp 1688980957
transform 1 0 34316 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 7912 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 14260 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 13984 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 14628 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 33672 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 8464 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 24564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 16468 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 25116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 25944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 25116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 7176 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 30268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 18860 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 25668 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 25944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 17388 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27048 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 7912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 8740 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 17204 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 11868 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 17756 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 28428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 28796 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform -1 0 27692 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 29164 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 28336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 26404 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 24932 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 23276 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 26404 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 26680 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 29624 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 31004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 28612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 27140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform -1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 26772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 28888 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 12788 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 12052 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 13064 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 26864 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 9292 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 8280 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 25668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform -1 0 28612 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 27232 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform -1 0 10580 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 24656 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 10212 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 25484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 27324 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 29532 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 28244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 28796 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 23644 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 28428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 27692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform -1 0 22540 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 24564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 24840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 23736 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 26680 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 23828 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 23828 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 21620 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 8464 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 13616 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 32936 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 34132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 6164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 34408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 34132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 34132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1688980957
transform 1 0 20056 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap23
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap24
timestamp 1688980957
transform -1 0 11868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap25
timestamp 1688980957
transform 1 0 8280 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap26
timestamp 1688980957
transform -1 0 5980 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap27
timestamp 1688980957
transform 1 0 4600 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 26956 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1688980957
transform -1 0 1932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform -1 0 1932 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1688980957
transform 1 0 34040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 34684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 34684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 34684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 34684 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 34684 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 34684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 34684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 34684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 34684 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 34684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 34684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 34684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 34684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 34684 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 34684 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 34684 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 34684 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 34684 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 34684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 34684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 34684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 34684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 34684 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 34684 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 34684 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 34684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 34684 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 34684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 34684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 34684 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 34684 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 34684 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 34684 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 34684 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 34684 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 6256 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 16560 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 21712 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 26864 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 32016 0 1 34816
box -38 -48 130 592
<< labels >>
flabel metal3 s 35073 34688 35873 34808 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 en
port 1 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 keypad_i[0]
port 2 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 keypad_i[10]
port 3 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 keypad_i[11]
port 4 nsew signal input
flabel metal2 s 7746 37217 7802 38017 0 FreeSans 224 90 0 0 keypad_i[12]
port 5 nsew signal input
flabel metal2 s 13542 37217 13598 38017 0 FreeSans 224 90 0 0 keypad_i[13]
port 6 nsew signal input
flabel metal2 s 32862 37217 32918 38017 0 FreeSans 224 90 0 0 keypad_i[14]
port 7 nsew signal input
flabel metal3 s 35073 8168 35873 8288 0 FreeSans 480 0 0 0 keypad_i[1]
port 8 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 keypad_i[2]
port 9 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 keypad_i[3]
port 10 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 keypad_i[4]
port 11 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 keypad_i[5]
port 12 nsew signal input
flabel metal3 s 35073 1368 35873 1488 0 FreeSans 480 0 0 0 keypad_i[6]
port 13 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 keypad_i[7]
port 14 nsew signal input
flabel metal3 s 35073 21088 35873 21208 0 FreeSans 480 0 0 0 keypad_i[8]
port 15 nsew signal input
flabel metal3 s 35073 27888 35873 28008 0 FreeSans 480 0 0 0 keypad_i[9]
port 16 nsew signal input
flabel metal2 s 19982 37217 20038 38017 0 FreeSans 224 90 0 0 n_rst
port 17 nsew signal input
flabel metal2 s 26422 37217 26478 38017 0 FreeSans 224 90 0 0 pwm_o
port 18 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 sound_series[0]
port 19 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 sound_series[1]
port 20 nsew signal tristate
flabel metal2 s 1306 37217 1362 38017 0 FreeSans 224 90 0 0 sound_series[2]
port 21 nsew signal tristate
flabel metal3 s 35073 14288 35873 14408 0 FreeSans 480 0 0 0 sound_series[3]
port 22 nsew signal tristate
flabel metal4 s 5141 2128 5461 35408 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 13535 2128 13855 35408 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 21929 2128 22249 35408 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 30323 2128 30643 35408 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 9338 2128 9658 35408 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
flabel metal4 s 17732 2128 18052 35408 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
flabel metal4 s 26126 2128 26446 35408 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
flabel metal4 s 34520 2128 34840 35408 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
rlabel metal1 17894 35360 17894 35360 0 vccd1
rlabel via1 17972 34816 17972 34816 0 vssd1
rlabel metal2 4094 15810 4094 15810 0 SS_FSM.count\[0\]
rlabel metal1 3266 16558 3266 16558 0 SS_FSM.count\[1\]
rlabel metal1 4324 20434 4324 20434 0 SS_FSM.count\[2\]
rlabel metal1 3726 18326 3726 18326 0 SS_FSM.count\[3\]
rlabel metal1 5750 18258 5750 18258 0 SS_FSM.count\[4\]
rlabel metal1 7452 20230 7452 20230 0 SS_FSM.count\[5\]
rlabel metal2 11362 21420 11362 21420 0 SS_FSM.count\[6\]
rlabel metal1 10120 20502 10120 20502 0 SS_FSM.count\[7\]
rlabel metal1 7406 20468 7406 20468 0 SS_FSM.count\[8\]
rlabel metal1 12236 22202 12236 22202 0 SS_FSM.next_sound\[0\]
rlabel metal1 13484 21114 13484 21114 0 SS_FSM.next_sound\[1\]
rlabel metal1 13386 19822 13386 19822 0 SS_FSM.sound\[0\]
rlabel metal1 8004 19822 8004 19822 0 SS_FSM.sound\[1\]
rlabel metal2 30958 27778 30958 27778 0 _0000_
rlabel metal2 31142 29478 31142 29478 0 _0001_
rlabel metal1 28244 29070 28244 29070 0 _0002_
rlabel metal1 25668 5338 25668 5338 0 _0003_
rlabel metal1 27048 4182 27048 4182 0 _0004_
rlabel metal1 28198 8058 28198 8058 0 _0005_
rlabel metal1 33166 5882 33166 5882 0 _0006_
rlabel metal1 29532 9962 29532 9962 0 _0007_
rlabel metal1 32512 10234 32512 10234 0 _0008_
rlabel metal1 30176 11798 30176 11798 0 _0009_
rlabel metal2 27922 14178 27922 14178 0 _0010_
rlabel metal1 28014 15674 28014 15674 0 _0011_
rlabel metal1 28704 17850 28704 17850 0 _0012_
rlabel metal1 28428 20026 28428 20026 0 _0013_
rlabel metal2 32246 22372 32246 22372 0 _0014_
rlabel metal1 33672 23834 33672 23834 0 _0015_
rlabel metal1 32614 26010 32614 26010 0 _0016_
rlabel metal1 28704 26554 28704 26554 0 _0017_
rlabel metal1 27048 23154 27048 23154 0 _0018_
rlabel metal1 21344 27098 21344 27098 0 _0019_
rlabel metal2 22310 28696 22310 28696 0 _0020_
rlabel metal1 22540 29818 22540 29818 0 _0021_
rlabel metal1 24741 30906 24741 30906 0 _0022_
rlabel metal1 28474 32504 28474 32504 0 _0023_
rlabel metal1 22448 31450 22448 31450 0 _0024_
rlabel metal2 22310 33235 22310 33235 0 _0025_
rlabel metal1 22816 34170 22816 34170 0 _0026_
rlabel metal1 24518 27064 24518 27064 0 _0027_
rlabel metal1 26036 27982 26036 27982 0 _0028_
rlabel metal1 24932 29070 24932 29070 0 _0029_
rlabel metal1 27048 30158 27048 30158 0 _0030_
rlabel metal1 28336 31654 28336 31654 0 _0031_
rlabel metal2 28934 32164 28934 32164 0 _0032_
rlabel metal1 24288 31858 24288 31858 0 _0033_
rlabel metal1 25668 33082 25668 33082 0 _0034_
rlabel metal2 23782 8602 23782 8602 0 _0035_
rlabel metal1 26719 6970 26719 6970 0 _0036_
rlabel metal1 24334 4046 24334 4046 0 _0037_
rlabel metal1 24518 7310 24518 7310 0 _0038_
rlabel metal2 26358 9180 26358 9180 0 _0039_
rlabel metal1 27094 11050 27094 11050 0 _0040_
rlabel metal2 27002 12517 27002 12517 0 _0041_
rlabel metal1 27324 13362 27324 13362 0 _0042_
rlabel metal1 25898 15402 25898 15402 0 _0043_
rlabel metal1 26443 16762 26443 16762 0 _0044_
rlabel metal1 27002 19278 27002 19278 0 _0045_
rlabel metal1 25392 20502 25392 20502 0 _0046_
rlabel metal1 27048 21454 27048 21454 0 _0047_
rlabel metal1 24840 23290 24840 23290 0 _0048_
rlabel metal2 23690 25432 23690 25432 0 _0049_
rlabel metal1 24794 21896 24794 21896 0 _0050_
rlabel metal1 3551 15674 3551 15674 0 _0051_
rlabel metal1 2484 17102 2484 17102 0 _0052_
rlabel metal1 2530 20026 2530 20026 0 _0053_
rlabel metal2 1886 18530 1886 18530 0 _0054_
rlabel metal1 4600 21658 4600 21658 0 _0055_
rlabel metal1 7268 21658 7268 21658 0 _0056_
rlabel metal1 9430 21658 9430 21658 0 _0057_
rlabel metal1 8510 23630 8510 23630 0 _0058_
rlabel metal1 6118 22202 6118 22202 0 _0059_
rlabel metal1 20240 5270 20240 5270 0 _0060_
rlabel metal1 21965 4454 21965 4454 0 _0061_
rlabel metal1 22218 7480 22218 7480 0 _0062_
rlabel metal1 23085 5882 23085 5882 0 _0063_
rlabel metal1 22855 10234 22855 10234 0 _0064_
rlabel metal1 24886 10710 24886 10710 0 _0065_
rlabel metal2 24702 12376 24702 12376 0 _0066_
rlabel metal1 24058 13838 24058 13838 0 _0067_
rlabel metal1 24242 16014 24242 16014 0 _0068_
rlabel metal1 24518 18360 24518 18360 0 _0069_
rlabel metal1 24104 19278 24104 19278 0 _0070_
rlabel metal1 23644 21454 23644 21454 0 _0071_
rlabel metal1 22494 23630 22494 23630 0 _0072_
rlabel metal1 21482 26418 21482 26418 0 _0073_
rlabel metal1 19366 27064 19366 27064 0 _0074_
rlabel metal2 21298 24582 21298 24582 0 _0075_
rlabel metal1 27002 28118 27002 28118 0 _0076_
rlabel metal1 25300 26010 25300 26010 0 _0077_
rlabel metal1 17756 34170 17756 34170 0 _0078_
rlabel metal1 20010 34510 20010 34510 0 _0079_
rlabel metal1 22954 29614 22954 29614 0 _0080_
rlabel metal1 25070 30362 25070 30362 0 _0081_
rlabel metal1 26588 31994 26588 31994 0 _0082_
rlabel metal1 22862 31314 22862 31314 0 _0083_
rlabel metal1 22356 32878 22356 32878 0 _0084_
rlabel metal1 23276 33966 23276 33966 0 _0085_
rlabel metal1 24150 9010 24150 9010 0 _0086_
rlabel metal1 26818 7922 26818 7922 0 _0087_
rlabel via1 27274 7854 27274 7854 0 _0088_
rlabel metal1 22862 4114 22862 4114 0 _0089_
rlabel metal1 23966 4148 23966 4148 0 _0090_
rlabel metal1 24196 7922 24196 7922 0 _0091_
rlabel metal1 24150 7412 24150 7412 0 _0092_
rlabel metal1 27002 9622 27002 9622 0 _0093_
rlabel metal1 26726 9554 26726 9554 0 _0094_
rlabel metal1 26910 10710 26910 10710 0 _0095_
rlabel metal1 26864 10778 26864 10778 0 _0096_
rlabel metal1 26128 12818 26128 12818 0 _0097_
rlabel metal1 27002 13974 27002 13974 0 _0098_
rlabel metal1 25622 15062 25622 15062 0 _0099_
rlabel metal1 25668 15130 25668 15130 0 _0100_
rlabel metal1 25070 17578 25070 17578 0 _0101_
rlabel metal1 26772 17646 26772 17646 0 _0102_
rlabel metal1 25254 18802 25254 18802 0 _0103_
rlabel metal1 26450 18938 26450 18938 0 _0104_
rlabel metal1 25300 19754 25300 19754 0 _0105_
rlabel metal1 25484 20026 25484 20026 0 _0106_
rlabel metal1 26450 20842 26450 20842 0 _0107_
rlabel metal1 26680 21114 26680 21114 0 _0108_
rlabel metal1 23506 23018 23506 23018 0 _0109_
rlabel metal1 25070 23086 25070 23086 0 _0110_
rlabel metal1 23920 24786 23920 24786 0 _0111_
rlabel metal2 25162 20366 25162 20366 0 _0112_
rlabel metal1 24794 21386 24794 21386 0 _0113_
rlabel metal1 5152 20502 5152 20502 0 _0114_
rlabel metal1 4922 19686 4922 19686 0 _0115_
rlabel metal2 5474 14144 5474 14144 0 _0116_
rlabel metal1 4094 19822 4094 19822 0 _0117_
rlabel metal1 4186 17680 4186 17680 0 _0118_
rlabel metal1 3864 18326 3864 18326 0 _0119_
rlabel metal1 7176 20434 7176 20434 0 _0120_
rlabel metal1 4600 20026 4600 20026 0 _0121_
rlabel metal2 5014 20706 5014 20706 0 _0122_
rlabel metal1 4876 20774 4876 20774 0 _0123_
rlabel metal1 2898 19856 2898 19856 0 _0124_
rlabel metal2 4002 18054 4002 18054 0 _0125_
rlabel metal1 5014 21488 5014 21488 0 _0126_
rlabel metal1 5106 21556 5106 21556 0 _0127_
rlabel metal1 7498 21556 7498 21556 0 _0128_
rlabel metal1 9338 21556 9338 21556 0 _0129_
rlabel metal1 10028 21658 10028 21658 0 _0130_
rlabel metal1 6578 20570 6578 20570 0 _0131_
rlabel metal1 18078 24888 18078 24888 0 _0132_
rlabel metal1 20976 5882 20976 5882 0 _0133_
rlabel metal1 21758 4590 21758 4590 0 _0134_
rlabel metal1 23000 8058 23000 8058 0 _0135_
rlabel metal1 23460 6426 23460 6426 0 _0136_
rlabel metal1 23046 9690 23046 9690 0 _0137_
rlabel metal1 24748 10234 24748 10234 0 _0138_
rlabel metal1 24748 11866 24748 11866 0 _0139_
rlabel metal1 24058 13498 24058 13498 0 _0140_
rlabel metal1 23874 16116 23874 16116 0 _0141_
rlabel metal2 24426 18292 24426 18292 0 _0142_
rlabel metal1 24426 19822 24426 19822 0 _0143_
rlabel metal1 23782 21896 23782 21896 0 _0144_
rlabel metal1 22402 23290 22402 23290 0 _0145_
rlabel metal1 21436 26010 21436 26010 0 _0146_
rlabel metal1 19412 26554 19412 26554 0 _0147_
rlabel metal1 21344 24174 21344 24174 0 _0148_
rlabel metal1 26680 27098 26680 27098 0 _0149_
rlabel metal1 26542 28560 26542 28560 0 _0150_
rlabel metal2 18814 34204 18814 34204 0 _0151_
rlabel metal1 18170 33966 18170 33966 0 _0152_
rlabel metal1 19688 34170 19688 34170 0 _0153_
rlabel metal1 8188 13294 8188 13294 0 _0154_
rlabel metal1 3036 16014 3036 16014 0 _0155_
rlabel metal1 5888 16762 5888 16762 0 _0156_
rlabel metal2 7406 18258 7406 18258 0 _0157_
rlabel metal1 6900 18734 6900 18734 0 _0158_
rlabel metal1 7222 15079 7222 15079 0 _0159_
rlabel metal1 3266 11798 3266 11798 0 _0160_
rlabel metal1 4416 12342 4416 12342 0 _0161_
rlabel metal2 9936 13770 9936 13770 0 _0162_
rlabel metal1 4968 14858 4968 14858 0 _0163_
rlabel metal1 4968 16014 4968 16014 0 _0164_
rlabel metal2 4554 12104 4554 12104 0 _0165_
rlabel metal1 11086 17204 11086 17204 0 _0166_
rlabel metal1 6164 20910 6164 20910 0 _0167_
rlabel metal1 13570 14960 13570 14960 0 _0168_
rlabel metal1 10994 19686 10994 19686 0 _0169_
rlabel metal1 10902 20400 10902 20400 0 _0170_
rlabel metal1 9614 20366 9614 20366 0 _0171_
rlabel metal2 5382 19788 5382 19788 0 _0172_
rlabel metal1 5106 19482 5106 19482 0 _0173_
rlabel metal2 8970 19703 8970 19703 0 _0174_
rlabel metal1 8740 20298 8740 20298 0 _0175_
rlabel metal1 12006 13294 12006 13294 0 _0176_
rlabel metal1 7682 18734 7682 18734 0 _0177_
rlabel metal1 8924 18258 8924 18258 0 _0178_
rlabel metal2 7682 16660 7682 16660 0 _0179_
rlabel metal1 7461 19822 7461 19822 0 _0180_
rlabel metal1 7544 20026 7544 20026 0 _0181_
rlabel via2 3634 17187 3634 17187 0 _0182_
rlabel metal1 7820 11730 7820 11730 0 _0183_
rlabel metal1 7222 15640 7222 15640 0 _0184_
rlabel metal1 7498 12614 7498 12614 0 _0185_
rlabel metal2 12466 9197 12466 9197 0 _0186_
rlabel metal1 13110 13838 13110 13838 0 _0187_
rlabel metal1 5014 15062 5014 15062 0 _0188_
rlabel metal1 5796 15130 5796 15130 0 _0189_
rlabel metal1 6302 14280 6302 14280 0 _0190_
rlabel metal1 8694 16490 8694 16490 0 _0191_
rlabel metal1 13156 15470 13156 15470 0 _0192_
rlabel metal1 7005 14042 7005 14042 0 _0193_
rlabel metal1 13202 13328 13202 13328 0 _0194_
rlabel metal2 10074 11441 10074 11441 0 _0195_
rlabel metal1 5198 13940 5198 13940 0 _0196_
rlabel metal1 12742 11084 12742 11084 0 _0197_
rlabel metal1 6854 10676 6854 10676 0 _0198_
rlabel metal1 4048 11866 4048 11866 0 _0199_
rlabel via2 12742 12189 12742 12189 0 _0200_
rlabel metal1 12512 13226 12512 13226 0 _0201_
rlabel metal1 12972 13294 12972 13294 0 _0202_
rlabel metal1 13432 13498 13432 13498 0 _0203_
rlabel metal1 13018 14042 13018 14042 0 _0204_
rlabel metal2 6394 16150 6394 16150 0 _0205_
rlabel metal1 12144 14994 12144 14994 0 _0206_
rlabel metal1 13524 14382 13524 14382 0 _0207_
rlabel metal1 12926 14348 12926 14348 0 _0208_
rlabel metal1 9338 16218 9338 16218 0 _0209_
rlabel metal1 4784 14042 4784 14042 0 _0210_
rlabel metal1 6716 16218 6716 16218 0 _0211_
rlabel via2 5106 11747 5106 11747 0 _0212_
rlabel metal1 11040 14382 11040 14382 0 _0213_
rlabel metal1 9798 21114 9798 21114 0 _0214_
rlabel metal1 12328 14450 12328 14450 0 _0215_
rlabel metal1 10442 20468 10442 20468 0 _0216_
rlabel metal1 10810 20230 10810 20230 0 _0217_
rlabel metal1 13800 14586 13800 14586 0 _0218_
rlabel metal1 4508 19822 4508 19822 0 _0219_
rlabel metal1 9476 17646 9476 17646 0 _0220_
rlabel metal1 9292 16966 9292 16966 0 _0221_
rlabel metal1 4462 13498 4462 13498 0 _0222_
rlabel metal1 5244 16966 5244 16966 0 _0223_
rlabel metal1 5520 10030 5520 10030 0 _0224_
rlabel via1 9522 11658 9522 11658 0 _0225_
rlabel metal1 9660 16558 9660 16558 0 _0226_
rlabel metal2 10718 16252 10718 16252 0 _0227_
rlabel metal1 8050 9520 8050 9520 0 _0228_
rlabel metal1 10580 11730 10580 11730 0 _0229_
rlabel metal1 10258 15470 10258 15470 0 _0230_
rlabel metal1 10442 15674 10442 15674 0 _0231_
rlabel metal2 9154 14042 9154 14042 0 _0232_
rlabel metal1 14214 15062 14214 15062 0 _0233_
rlabel metal1 8510 18394 8510 18394 0 _0234_
rlabel metal1 10028 18258 10028 18258 0 _0235_
rlabel metal1 5014 19244 5014 19244 0 _0236_
rlabel metal2 13110 17340 13110 17340 0 _0237_
rlabel metal2 13110 14688 13110 14688 0 _0238_
rlabel metal1 13202 15028 13202 15028 0 _0239_
rlabel metal2 12282 20230 12282 20230 0 _0240_
rlabel metal1 13340 9690 13340 9690 0 _0241_
rlabel metal1 13294 10098 13294 10098 0 _0242_
rlabel metal1 13478 9962 13478 9962 0 _0243_
rlabel metal1 9844 9690 9844 9690 0 _0244_
rlabel metal1 13202 10234 13202 10234 0 _0245_
rlabel metal1 12788 9894 12788 9894 0 _0246_
rlabel metal1 9430 9996 9430 9996 0 _0247_
rlabel metal1 9936 9486 9936 9486 0 _0248_
rlabel metal1 9200 12818 9200 12818 0 _0249_
rlabel metal1 9706 13702 9706 13702 0 _0250_
rlabel metal1 9384 9146 9384 9146 0 _0251_
rlabel metal1 8970 9486 8970 9486 0 _0252_
rlabel metal2 7038 13129 7038 13129 0 _0253_
rlabel metal1 6256 10166 6256 10166 0 _0254_
rlabel metal1 5842 10166 5842 10166 0 _0255_
rlabel metal1 6624 10234 6624 10234 0 _0256_
rlabel metal1 12673 13294 12673 13294 0 _0257_
rlabel metal1 7912 9350 7912 9350 0 _0258_
rlabel metal1 9200 9690 9200 9690 0 _0259_
rlabel metal1 8832 10234 8832 10234 0 _0260_
rlabel metal2 8142 11696 8142 11696 0 _0261_
rlabel metal1 8280 11118 8280 11118 0 _0262_
rlabel metal1 8878 11322 8878 11322 0 _0263_
rlabel metal1 9200 12954 9200 12954 0 _0264_
rlabel metal1 8970 11866 8970 11866 0 _0265_
rlabel metal1 7360 11526 7360 11526 0 _0266_
rlabel metal1 8096 11866 8096 11866 0 _0267_
rlabel metal1 9016 12410 9016 12410 0 _0268_
rlabel metal1 7498 14348 7498 14348 0 _0269_
rlabel metal1 8648 13226 8648 13226 0 _0270_
rlabel metal1 9614 13498 9614 13498 0 _0271_
rlabel metal1 8694 13906 8694 13906 0 _0272_
rlabel metal1 7820 14042 7820 14042 0 _0273_
rlabel metal1 12558 20230 12558 20230 0 _0274_
rlabel metal1 7498 15674 7498 15674 0 _0275_
rlabel metal1 7222 16762 7222 16762 0 _0276_
rlabel metal1 7222 16592 7222 16592 0 _0277_
rlabel metal1 7130 16592 7130 16592 0 _0278_
rlabel metal1 8648 16694 8648 16694 0 _0279_
rlabel metal1 12742 15504 12742 15504 0 _0280_
rlabel metal2 13294 15810 13294 15810 0 _0281_
rlabel metal2 13938 16898 13938 16898 0 _0282_
rlabel metal1 12006 17102 12006 17102 0 _0283_
rlabel metal1 11864 17306 11864 17306 0 _0284_
rlabel metal2 12834 15487 12834 15487 0 _0285_
rlabel metal1 12926 16218 12926 16218 0 _0286_
rlabel metal1 13938 17204 13938 17204 0 _0287_
rlabel metal1 11822 9078 11822 9078 0 _0288_
rlabel metal2 12374 11526 12374 11526 0 _0289_
rlabel metal1 13110 11560 13110 11560 0 _0290_
rlabel metal1 10028 11254 10028 11254 0 _0291_
rlabel metal2 9614 12580 9614 12580 0 _0292_
rlabel metal1 13478 11798 13478 11798 0 _0293_
rlabel metal1 12926 11696 12926 11696 0 _0294_
rlabel metal1 13340 11866 13340 11866 0 _0295_
rlabel metal1 13570 17034 13570 17034 0 _0296_
rlabel metal2 8556 18734 8556 18734 0 _0297_
rlabel metal1 12972 18666 12972 18666 0 _0298_
rlabel metal2 12006 18768 12006 18768 0 _0299_
rlabel metal1 8328 15470 8328 15470 0 _0300_
rlabel metal2 8234 15351 8234 15351 0 _0301_
rlabel metal2 8602 17408 8602 17408 0 _0302_
rlabel metal1 8096 15130 8096 15130 0 _0303_
rlabel metal2 8602 15895 8602 15895 0 _0304_
rlabel metal1 13386 9622 13386 9622 0 _0305_
rlabel metal2 11178 11628 11178 11628 0 _0306_
rlabel metal1 10856 11322 10856 11322 0 _0307_
rlabel metal1 10955 11730 10955 11730 0 _0308_
rlabel metal1 13110 11152 13110 11152 0 _0309_
rlabel metal2 13892 13770 13892 13770 0 _0310_
rlabel metal1 12190 13226 12190 13226 0 _0311_
rlabel metal2 12742 13634 12742 13634 0 _0312_
rlabel metal2 13248 17170 13248 17170 0 _0313_
rlabel metal1 10626 9146 10626 9146 0 _0314_
rlabel metal2 8234 9860 8234 9860 0 _0315_
rlabel metal2 9430 9520 9430 9520 0 _0316_
rlabel metal1 12742 9656 12742 9656 0 _0317_
rlabel metal1 11592 9146 11592 9146 0 _0318_
rlabel metal1 11500 9690 11500 9690 0 _0319_
rlabel metal1 11178 9588 11178 9588 0 _0320_
rlabel metal2 10672 16524 10672 16524 0 _0321_
rlabel metal1 10626 13940 10626 13940 0 _0322_
rlabel metal1 10396 14042 10396 14042 0 _0323_
rlabel metal1 11270 14790 11270 14790 0 _0324_
rlabel metal1 10948 17646 10948 17646 0 _0325_
rlabel metal1 12742 17782 12742 17782 0 _0326_
rlabel metal2 14674 17408 14674 17408 0 _0327_
rlabel metal1 10672 18190 10672 18190 0 _0328_
rlabel metal1 14490 18258 14490 18258 0 _0329_
rlabel metal1 16238 14824 16238 14824 0 _0330_
rlabel metal1 14950 32198 14950 32198 0 _0331_
rlabel metal1 15456 12614 15456 12614 0 _0332_
rlabel metal1 15088 12818 15088 12818 0 _0333_
rlabel metal1 15962 16082 15962 16082 0 _0334_
rlabel metal1 15042 16422 15042 16422 0 _0335_
rlabel metal1 15456 16558 15456 16558 0 _0336_
rlabel metal2 15410 15130 15410 15130 0 _0337_
rlabel metal1 15870 13362 15870 13362 0 _0338_
rlabel metal2 15686 9078 15686 9078 0 _0339_
rlabel metal1 15456 13498 15456 13498 0 _0340_
rlabel metal1 15640 14382 15640 14382 0 _0341_
rlabel metal2 15410 16252 15410 16252 0 _0342_
rlabel metal2 15778 15198 15778 15198 0 _0343_
rlabel metal1 15916 18258 15916 18258 0 _0344_
rlabel metal1 13248 18122 13248 18122 0 _0345_
rlabel metal1 15318 18156 15318 18156 0 _0346_
rlabel metal1 15870 12954 15870 12954 0 _0347_
rlabel metal1 16376 17510 16376 17510 0 _0348_
rlabel metal1 16422 17646 16422 17646 0 _0349_
rlabel metal2 17020 20570 17020 20570 0 _0350_
rlabel metal1 20010 17748 20010 17748 0 _0351_
rlabel metal1 18078 14994 18078 14994 0 _0352_
rlabel metal1 16974 15436 16974 15436 0 _0353_
rlabel metal1 15916 13974 15916 13974 0 _0354_
rlabel metal1 16744 7514 16744 7514 0 _0355_
rlabel metal1 16054 8976 16054 8976 0 _0356_
rlabel metal1 16146 13838 16146 13838 0 _0357_
rlabel metal1 16008 14042 16008 14042 0 _0358_
rlabel metal1 17250 15504 17250 15504 0 _0359_
rlabel metal1 17526 15470 17526 15470 0 _0360_
rlabel metal1 18078 13974 18078 13974 0 _0361_
rlabel metal1 17342 14280 17342 14280 0 _0362_
rlabel metal1 15916 9078 15916 9078 0 _0363_
rlabel metal1 15870 7718 15870 7718 0 _0364_
rlabel metal1 15916 8942 15916 8942 0 _0365_
rlabel metal1 15548 9146 15548 9146 0 _0366_
rlabel metal1 15824 9622 15824 9622 0 _0367_
rlabel metal1 16790 14518 16790 14518 0 _0368_
rlabel metal1 18354 15028 18354 15028 0 _0369_
rlabel metal2 20286 16218 20286 16218 0 _0370_
rlabel metal1 14950 18190 14950 18190 0 _0371_
rlabel metal1 15778 18768 15778 18768 0 _0372_
rlabel metal1 18009 18666 18009 18666 0 _0373_
rlabel metal1 20884 16626 20884 16626 0 _0374_
rlabel metal1 18354 13974 18354 13974 0 _0375_
rlabel metal1 21344 16762 21344 16762 0 _0376_
rlabel metal1 20562 13940 20562 13940 0 _0377_
rlabel metal1 20792 14994 20792 14994 0 _0378_
rlabel metal1 21758 15504 21758 15504 0 _0379_
rlabel metal1 22172 13294 22172 13294 0 _0380_
rlabel metal1 23046 15368 23046 15368 0 _0381_
rlabel metal1 20424 19346 20424 19346 0 _0382_
rlabel metal1 23230 14416 23230 14416 0 _0383_
rlabel metal1 21574 15674 21574 15674 0 _0384_
rlabel metal1 22724 20910 22724 20910 0 _0385_
rlabel metal2 22770 14722 22770 14722 0 _0386_
rlabel metal1 22494 20808 22494 20808 0 _0387_
rlabel metal1 22954 20434 22954 20434 0 _0388_
rlabel metal1 22310 20264 22310 20264 0 _0389_
rlabel metal1 23230 16048 23230 16048 0 _0390_
rlabel metal1 20608 13294 20608 13294 0 _0391_
rlabel metal1 22954 13498 22954 13498 0 _0392_
rlabel metal1 23184 17510 23184 17510 0 _0393_
rlabel metal1 22908 16082 22908 16082 0 _0394_
rlabel metal2 22586 19074 22586 19074 0 _0395_
rlabel metal1 22540 20026 22540 20026 0 _0396_
rlabel metal1 20700 19346 20700 19346 0 _0397_
rlabel metal1 20378 20842 20378 20842 0 _0398_
rlabel metal1 20654 21386 20654 21386 0 _0399_
rlabel metal1 20838 21046 20838 21046 0 _0400_
rlabel metal1 21620 21522 21620 21522 0 _0401_
rlabel metal2 20746 18088 20746 18088 0 _0402_
rlabel metal1 21356 21590 21356 21590 0 _0403_
rlabel metal1 21850 20400 21850 20400 0 _0404_
rlabel metal1 21896 20570 21896 20570 0 _0405_
rlabel metal1 19734 15062 19734 15062 0 _0406_
rlabel metal1 23690 15436 23690 15436 0 _0407_
rlabel via1 23874 17647 23874 17647 0 _0408_
rlabel metal1 22034 18802 22034 18802 0 _0409_
rlabel metal1 21206 17714 21206 17714 0 _0410_
rlabel metal1 22356 18666 22356 18666 0 _0411_
rlabel metal1 22954 18734 22954 18734 0 _0412_
rlabel metal1 21965 18666 21965 18666 0 _0413_
rlabel metal1 21804 20910 21804 20910 0 _0414_
rlabel metal1 21206 20876 21206 20876 0 _0415_
rlabel metal1 20976 20978 20976 20978 0 _0416_
rlabel metal1 17618 19686 17618 19686 0 _0417_
rlabel metal1 22586 12206 22586 12206 0 _0418_
rlabel metal1 23552 14314 23552 14314 0 _0419_
rlabel metal1 19872 14246 19872 14246 0 _0420_
rlabel metal1 20838 13362 20838 13362 0 _0421_
rlabel metal2 21206 12750 21206 12750 0 _0422_
rlabel metal1 20976 9486 20976 9486 0 _0423_
rlabel metal1 21298 9622 21298 9622 0 _0424_
rlabel metal1 18768 13906 18768 13906 0 _0425_
rlabel metal1 18676 13838 18676 13838 0 _0426_
rlabel metal1 19826 14042 19826 14042 0 _0427_
rlabel metal2 21390 9078 21390 9078 0 _0428_
rlabel metal1 21068 14586 21068 14586 0 _0429_
rlabel metal1 21758 14450 21758 14450 0 _0430_
rlabel metal1 21920 9452 21920 9452 0 _0431_
rlabel metal2 21206 9350 21206 9350 0 _0432_
rlabel metal2 21666 10642 21666 10642 0 _0433_
rlabel metal2 21574 11526 21574 11526 0 _0434_
rlabel metal2 20102 11390 20102 11390 0 _0435_
rlabel metal1 21298 11118 21298 11118 0 _0436_
rlabel metal1 20286 11730 20286 11730 0 _0437_
rlabel metal1 20884 11662 20884 11662 0 _0438_
rlabel metal1 23276 12750 23276 12750 0 _0439_
rlabel metal1 22448 12614 22448 12614 0 _0440_
rlabel metal1 21574 12240 21574 12240 0 _0441_
rlabel metal1 21758 11730 21758 11730 0 _0442_
rlabel metal2 22494 15062 22494 15062 0 _0443_
rlabel metal1 21206 12206 21206 12206 0 _0444_
rlabel metal1 22172 12410 22172 12410 0 _0445_
rlabel metal2 23230 18394 23230 18394 0 _0446_
rlabel metal1 23322 18326 23322 18326 0 _0447_
rlabel metal1 18308 17170 18308 17170 0 _0448_
rlabel metal2 19550 6970 19550 6970 0 _0449_
rlabel metal1 19228 6426 19228 6426 0 _0450_
rlabel metal1 19366 6358 19366 6358 0 _0451_
rlabel metal1 17664 8466 17664 8466 0 _0452_
rlabel metal1 20160 7786 20160 7786 0 _0453_
rlabel metal1 19688 7378 19688 7378 0 _0454_
rlabel metal1 17204 9622 17204 9622 0 _0455_
rlabel metal1 17768 7786 17768 7786 0 _0456_
rlabel metal1 17526 7378 17526 7378 0 _0457_
rlabel metal1 17480 9486 17480 9486 0 _0458_
rlabel metal1 17722 9622 17722 9622 0 _0459_
rlabel metal1 18216 8942 18216 8942 0 _0460_
rlabel metal1 17296 11798 17296 11798 0 _0461_
rlabel metal2 17894 10404 17894 10404 0 _0462_
rlabel metal1 18124 10642 18124 10642 0 _0463_
rlabel metal1 17020 12206 17020 12206 0 _0464_
rlabel metal1 17296 11866 17296 11866 0 _0465_
rlabel metal1 15594 11764 15594 11764 0 _0466_
rlabel metal1 18584 17238 18584 17238 0 _0467_
rlabel metal1 17630 12274 17630 12274 0 _0468_
rlabel metal1 18262 12206 18262 12206 0 _0469_
rlabel metal2 17618 17408 17618 17408 0 _0470_
rlabel metal1 18274 17102 18274 17102 0 _0471_
rlabel metal1 18124 16558 18124 16558 0 _0472_
rlabel via1 17166 19686 17166 19686 0 _0473_
rlabel metal2 18078 17918 18078 17918 0 _0474_
rlabel metal1 18492 18394 18492 18394 0 _0475_
rlabel metal1 17740 20502 17740 20502 0 _0476_
rlabel metal1 17526 19482 17526 19482 0 _0477_
rlabel metal1 18308 18734 18308 18734 0 _0478_
rlabel metal1 18216 20910 18216 20910 0 _0479_
rlabel metal2 17526 20740 17526 20740 0 _0480_
rlabel metal1 16928 21114 16928 21114 0 _0481_
rlabel metal1 17894 21522 17894 21522 0 _0482_
rlabel metal1 18538 21114 18538 21114 0 _0483_
rlabel metal1 18262 21488 18262 21488 0 _0484_
rlabel metal1 19366 23698 19366 23698 0 _0485_
rlabel metal1 18860 22746 18860 22746 0 _0486_
rlabel metal1 19366 23086 19366 23086 0 _0487_
rlabel metal1 19550 24208 19550 24208 0 _0488_
rlabel metal1 19412 23834 19412 23834 0 _0489_
rlabel metal1 19320 24378 19320 24378 0 _0490_
rlabel metal1 17986 24106 17986 24106 0 _0491_
rlabel metal1 18124 24378 18124 24378 0 _0492_
rlabel metal1 12512 26350 12512 26350 0 _0493_
rlabel metal1 11224 26486 11224 26486 0 _0494_
rlabel metal1 10810 26282 10810 26282 0 _0495_
rlabel metal2 10350 26996 10350 26996 0 _0496_
rlabel metal1 11500 24378 11500 24378 0 _0497_
rlabel metal1 10442 24718 10442 24718 0 _0498_
rlabel metal1 11454 24242 11454 24242 0 _0499_
rlabel metal2 12742 25330 12742 25330 0 _0500_
rlabel metal2 12098 25432 12098 25432 0 _0501_
rlabel metal2 12558 25262 12558 25262 0 _0502_
rlabel metal1 15548 25194 15548 25194 0 _0503_
rlabel metal1 14490 26282 14490 26282 0 _0504_
rlabel metal2 14122 26996 14122 26996 0 _0505_
rlabel metal1 15916 25466 15916 25466 0 _0506_
rlabel metal1 16836 25194 16836 25194 0 _0507_
rlabel metal1 15778 24174 15778 24174 0 _0508_
rlabel metal2 16698 27234 16698 27234 0 _0509_
rlabel metal1 16330 29002 16330 29002 0 _0510_
rlabel metal1 16192 28934 16192 28934 0 _0511_
rlabel metal2 15502 29444 15502 29444 0 _0512_
rlabel via1 14582 30703 14582 30703 0 _0513_
rlabel metal1 14168 29138 14168 29138 0 _0514_
rlabel metal1 14260 30362 14260 30362 0 _0515_
rlabel metal1 15088 32402 15088 32402 0 _0516_
rlabel metal2 15226 30872 15226 30872 0 _0517_
rlabel metal1 15364 31314 15364 31314 0 _0518_
rlabel metal1 14858 32470 14858 32470 0 _0519_
rlabel metal2 14122 32232 14122 32232 0 _0520_
rlabel metal1 13294 31824 13294 31824 0 _0521_
rlabel metal2 15410 32674 15410 32674 0 _0522_
rlabel metal1 6348 25806 6348 25806 0 _0523_
rlabel metal1 7038 30124 7038 30124 0 _0524_
rlabel metal1 6394 29274 6394 29274 0 _0525_
rlabel metal1 6624 30294 6624 30294 0 _0526_
rlabel metal1 6164 31926 6164 31926 0 _0527_
rlabel metal1 6992 25942 6992 25942 0 _0528_
rlabel metal1 6164 25670 6164 25670 0 _0529_
rlabel metal1 6256 26350 6256 26350 0 _0530_
rlabel metal1 5566 28730 5566 28730 0 _0531_
rlabel metal1 7544 25874 7544 25874 0 _0532_
rlabel metal1 8188 25194 8188 25194 0 _0533_
rlabel metal1 5014 24854 5014 24854 0 _0534_
rlabel metal1 6532 24922 6532 24922 0 _0535_
rlabel metal1 6578 23698 6578 23698 0 _0536_
rlabel metal1 3634 24786 3634 24786 0 _0537_
rlabel metal1 4554 24208 4554 24208 0 _0538_
rlabel metal1 4094 24684 4094 24684 0 _0539_
rlabel via1 4002 28509 4002 28509 0 _0540_
rlabel metal1 4278 25670 4278 25670 0 _0541_
rlabel metal1 3634 26010 3634 26010 0 _0542_
rlabel metal1 3964 28390 3964 28390 0 _0543_
rlabel metal1 3772 28186 3772 28186 0 _0544_
rlabel metal1 3864 28730 3864 28730 0 _0545_
rlabel metal1 7452 29138 7452 29138 0 _0546_
rlabel metal1 5428 28458 5428 28458 0 _0547_
rlabel metal1 5520 28050 5520 28050 0 _0548_
rlabel metal1 7268 28934 7268 28934 0 _0549_
rlabel metal1 7360 28458 7360 28458 0 _0550_
rlabel metal1 8142 28526 8142 28526 0 _0551_
rlabel metal1 9062 29172 9062 29172 0 _0552_
rlabel metal2 9200 32334 9200 32334 0 _0553_
rlabel metal1 8924 29818 8924 29818 0 _0554_
rlabel metal1 10350 29138 10350 29138 0 _0555_
rlabel metal1 8188 31994 8188 31994 0 _0556_
rlabel metal1 10074 31450 10074 31450 0 _0557_
rlabel metal1 10304 31654 10304 31654 0 _0558_
rlabel metal1 7958 31858 7958 31858 0 _0559_
rlabel metal1 6486 32844 6486 32844 0 _0560_
rlabel metal1 8740 32538 8740 32538 0 _0561_
rlabel metal1 8786 33082 8786 33082 0 _0562_
rlabel metal1 6854 33456 6854 33456 0 _0563_
rlabel metal1 7866 33932 7866 33932 0 _0564_
rlabel metal1 8096 34170 8096 34170 0 _0565_
rlabel metal1 6624 33082 6624 33082 0 _0566_
rlabel metal1 4140 32878 4140 32878 0 _0567_
rlabel metal1 5014 33626 5014 33626 0 _0568_
rlabel metal1 4692 33966 4692 33966 0 _0569_
rlabel metal1 4278 32266 4278 32266 0 _0570_
rlabel metal2 3910 32640 3910 32640 0 _0571_
rlabel metal1 2645 31790 2645 31790 0 _0572_
rlabel metal1 5474 31858 5474 31858 0 _0573_
rlabel metal1 4922 32198 4922 32198 0 _0574_
rlabel metal2 4830 31178 4830 31178 0 _0575_
rlabel metal1 6072 31382 6072 31382 0 _0576_
rlabel metal1 13018 21488 13018 21488 0 _0577_
rlabel metal1 12972 21658 12972 21658 0 _0578_
rlabel metal1 12788 21998 12788 21998 0 _0579_
rlabel metal1 12581 22066 12581 22066 0 _0580_
rlabel metal1 20424 33830 20424 33830 0 _0581_
rlabel metal2 21022 32810 21022 32810 0 _0582_
rlabel metal1 19780 33082 19780 33082 0 _0583_
rlabel metal1 18998 33490 18998 33490 0 _0584_
rlabel metal1 19136 33422 19136 33422 0 _0585_
rlabel metal1 17434 33592 17434 33592 0 _0586_
rlabel metal1 19458 32504 19458 32504 0 _0587_
rlabel metal1 20056 31994 20056 31994 0 _0588_
rlabel metal2 19458 31620 19458 31620 0 _0589_
rlabel metal1 19136 31790 19136 31790 0 _0590_
rlabel metal2 21114 32980 21114 32980 0 _0591_
rlabel metal1 19136 30906 19136 30906 0 _0592_
rlabel metal1 17434 31892 17434 31892 0 _0593_
rlabel metal1 21114 32402 21114 32402 0 _0594_
rlabel metal1 20654 32334 20654 32334 0 _0595_
rlabel metal1 20378 31858 20378 31858 0 _0596_
rlabel metal1 18814 32266 18814 32266 0 _0597_
rlabel metal1 21022 30906 21022 30906 0 _0598_
rlabel metal1 21436 30906 21436 30906 0 _0599_
rlabel metal1 20654 31246 20654 31246 0 _0600_
rlabel metal1 17526 31212 17526 31212 0 _0601_
rlabel metal1 20930 29818 20930 29818 0 _0602_
rlabel metal1 20930 30124 20930 30124 0 _0603_
rlabel metal1 20378 30158 20378 30158 0 _0604_
rlabel metal2 17618 29818 17618 29818 0 _0605_
rlabel metal1 20792 28730 20792 28730 0 _0606_
rlabel metal2 21022 28934 21022 28934 0 _0607_
rlabel metal1 20194 29274 20194 29274 0 _0608_
rlabel metal1 17802 29580 17802 29580 0 _0609_
rlabel metal2 18630 29308 18630 29308 0 _0610_
rlabel metal1 19688 28730 19688 28730 0 _0611_
rlabel metal1 19734 28662 19734 28662 0 _0612_
rlabel metal1 19136 29070 19136 29070 0 _0613_
rlabel via1 18814 29138 18814 29138 0 _0614_
rlabel metal1 18170 28730 18170 28730 0 _0615_
rlabel metal1 18216 29138 18216 29138 0 _0616_
rlabel metal1 17480 29274 17480 29274 0 _0617_
rlabel metal2 18170 30260 18170 30260 0 _0618_
rlabel metal1 17618 30906 17618 30906 0 _0619_
rlabel metal2 17158 31620 17158 31620 0 _0620_
rlabel metal2 17802 32198 17802 32198 0 _0621_
rlabel metal2 17066 32912 17066 32912 0 _0622_
rlabel metal1 27140 25874 27140 25874 0 _0623_
rlabel metal1 27462 25840 27462 25840 0 _0624_
rlabel via1 28842 17187 28842 17187 0 _0625_
rlabel metal1 28198 27506 28198 27506 0 _0626_
rlabel metal1 29302 29036 29302 29036 0 _0627_
rlabel metal1 32568 5678 32568 5678 0 _0628_
rlabel metal2 30866 29172 30866 29172 0 _0629_
rlabel metal1 26956 25194 26956 25194 0 _0630_
rlabel metal2 26910 18292 26910 18292 0 _0631_
rlabel metal1 32522 23596 32522 23596 0 _0632_
rlabel metal1 27186 24718 27186 24718 0 _0633_
rlabel metal2 31372 21420 31372 21420 0 _0634_
rlabel metal1 31786 19414 31786 19414 0 _0635_
rlabel metal1 31786 18700 31786 18700 0 _0636_
rlabel metal1 31464 16082 31464 16082 0 _0637_
rlabel metal1 31418 14280 31418 14280 0 _0638_
rlabel metal1 29532 17170 29532 17170 0 _0639_
rlabel metal1 31786 16592 31786 16592 0 _0640_
rlabel metal1 31188 16762 31188 16762 0 _0641_
rlabel metal1 28796 6222 28796 6222 0 _0642_
rlabel metal1 30820 5202 30820 5202 0 _0643_
rlabel metal1 30636 6698 30636 6698 0 _0644_
rlabel metal1 30314 6256 30314 6256 0 _0645_
rlabel metal2 29762 7106 29762 7106 0 _0646_
rlabel metal2 31418 8636 31418 8636 0 _0647_
rlabel metal1 30912 7378 30912 7378 0 _0648_
rlabel metal1 31188 7718 31188 7718 0 _0649_
rlabel metal1 31004 10438 31004 10438 0 _0650_
rlabel metal2 30866 9350 30866 9350 0 _0651_
rlabel metal1 31602 9418 31602 9418 0 _0652_
rlabel metal1 33120 12070 33120 12070 0 _0653_
rlabel metal1 31234 11764 31234 11764 0 _0654_
rlabel metal1 31326 13430 31326 13430 0 _0655_
rlabel metal1 31832 12410 31832 12410 0 _0656_
rlabel metal1 31280 15062 31280 15062 0 _0657_
rlabel metal1 33166 17680 33166 17680 0 _0658_
rlabel metal2 30958 16796 30958 16796 0 _0659_
rlabel metal2 32798 16218 32798 16218 0 _0660_
rlabel metal1 32752 17170 32752 17170 0 _0661_
rlabel metal1 31648 17306 31648 17306 0 _0662_
rlabel metal1 31050 19312 31050 19312 0 _0663_
rlabel metal1 32660 17646 32660 17646 0 _0664_
rlabel metal1 31050 18938 31050 18938 0 _0665_
rlabel metal1 31142 20944 31142 20944 0 _0666_
rlabel metal1 30728 21114 30728 21114 0 _0667_
rlabel metal1 31924 24786 31924 24786 0 _0668_
rlabel metal1 31510 24752 31510 24752 0 _0669_
rlabel metal1 31694 24786 31694 24786 0 _0670_
rlabel metal2 31878 25092 31878 25092 0 _0671_
rlabel metal1 30636 24786 30636 24786 0 _0672_
rlabel metal1 29946 25262 29946 25262 0 _0673_
rlabel metal1 30130 25466 30130 25466 0 _0674_
rlabel metal1 30498 21318 30498 21318 0 _0675_
rlabel metal1 30912 21522 30912 21522 0 _0676_
rlabel metal1 31142 21658 31142 21658 0 _0677_
rlabel metal1 29854 22610 29854 22610 0 _0678_
rlabel metal1 30498 24718 30498 24718 0 _0679_
rlabel metal2 31326 23290 31326 23290 0 _0680_
rlabel metal1 30958 23154 30958 23154 0 _0681_
rlabel metal1 30406 22746 30406 22746 0 _0682_
rlabel metal2 31648 13668 31648 13668 0 _0683_
rlabel metal1 31510 7310 31510 7310 0 _0684_
rlabel metal1 30452 4794 30452 4794 0 _0685_
rlabel metal1 31188 5338 31188 5338 0 _0686_
rlabel metal1 32246 8908 32246 8908 0 _0687_
rlabel metal2 31832 13294 31832 13294 0 _0688_
rlabel metal1 32292 18258 32292 18258 0 _0689_
rlabel metal1 32522 16660 32522 16660 0 _0690_
rlabel metal2 33166 16966 33166 16966 0 _0691_
rlabel metal1 32522 16150 32522 16150 0 _0692_
rlabel metal1 32062 16422 32062 16422 0 _0693_
rlabel metal1 29210 6154 29210 6154 0 _0694_
rlabel metal2 29578 7990 29578 7990 0 _0695_
rlabel metal2 31234 13707 31234 13707 0 _0696_
rlabel via1 31142 13362 31142 13362 0 _0697_
rlabel metal1 33810 12342 33810 12342 0 _0698_
rlabel metal1 33258 12818 33258 12818 0 _0699_
rlabel metal2 31326 14144 31326 14144 0 _0700_
rlabel metal1 32338 21556 32338 21556 0 _0701_
rlabel metal2 30084 20468 30084 20468 0 _0702_
rlabel metal1 31855 15062 31855 15062 0 _0703_
rlabel metal2 31510 16269 31510 16269 0 _0704_
rlabel metal1 31188 22678 31188 22678 0 _0705_
rlabel metal2 32154 22277 32154 22277 0 _0706_
rlabel metal1 32430 6766 32430 6766 0 _0707_
rlabel metal1 24794 5236 24794 5236 0 _0708_
rlabel metal2 27830 5814 27830 5814 0 _0709_
rlabel metal1 26358 5236 26358 5236 0 _0710_
rlabel metal1 26818 5202 26818 5202 0 _0711_
rlabel metal1 28152 19890 28152 19890 0 _0712_
rlabel metal1 29670 5780 29670 5780 0 _0713_
rlabel metal1 30130 5882 30130 5882 0 _0714_
rlabel metal1 29440 5338 29440 5338 0 _0715_
rlabel metal1 28520 5338 28520 5338 0 _0716_
rlabel metal2 28198 18700 28198 18700 0 _0717_
rlabel metal2 28750 8330 28750 8330 0 _0718_
rlabel metal1 30774 6800 30774 6800 0 _0719_
rlabel metal1 32384 6630 32384 6630 0 _0720_
rlabel metal2 33074 6154 33074 6154 0 _0721_
rlabel metal1 32246 5678 32246 5678 0 _0722_
rlabel metal2 31050 7684 31050 7684 0 _0723_
rlabel metal1 32890 8398 32890 8398 0 _0724_
rlabel metal1 32476 9146 32476 9146 0 _0725_
rlabel metal1 28428 10030 28428 10030 0 _0726_
rlabel metal2 32062 10166 32062 10166 0 _0727_
rlabel metal2 33074 10880 33074 10880 0 _0728_
rlabel metal1 32660 10642 32660 10642 0 _0729_
rlabel metal1 32154 10642 32154 10642 0 _0730_
rlabel metal2 31510 12546 31510 12546 0 _0731_
rlabel metal1 33304 12954 33304 12954 0 _0732_
rlabel metal1 32062 12104 32062 12104 0 _0733_
rlabel metal1 30268 12206 30268 12206 0 _0734_
rlabel metal2 32338 14110 32338 14110 0 _0735_
rlabel via1 32246 13906 32246 13906 0 _0736_
rlabel metal1 32062 14042 32062 14042 0 _0737_
rlabel metal1 32154 14416 32154 14416 0 _0738_
rlabel metal1 28474 13872 28474 13872 0 _0739_
rlabel metal2 28658 14348 28658 14348 0 _0740_
rlabel metal1 32384 16082 32384 16082 0 _0741_
rlabel metal2 32982 16524 32982 16524 0 _0742_
rlabel metal1 32890 15980 32890 15980 0 _0743_
rlabel metal1 28980 15470 28980 15470 0 _0744_
rlabel metal1 33764 16626 33764 16626 0 _0745_
rlabel metal1 33764 16762 33764 16762 0 _0746_
rlabel metal1 28750 17204 28750 17204 0 _0747_
rlabel metal1 28152 17306 28152 17306 0 _0748_
rlabel metal1 33350 18598 33350 18598 0 _0749_
rlabel viali 32704 18712 32704 18712 0 _0750_
rlabel metal1 33166 18870 33166 18870 0 _0751_
rlabel metal1 32430 18836 32430 18836 0 _0752_
rlabel metal1 29670 18938 29670 18938 0 _0753_
rlabel metal1 32752 18938 32752 18938 0 _0754_
rlabel metal1 33120 19482 33120 19482 0 _0755_
rlabel metal1 32752 20570 32752 20570 0 _0756_
rlabel metal1 32154 21862 32154 21862 0 _0757_
rlabel metal2 32154 18428 32154 18428 0 _0758_
rlabel metal1 32384 17646 32384 17646 0 _0759_
rlabel metal1 31993 21454 31993 21454 0 _0760_
rlabel metal1 32982 21454 32982 21454 0 _0761_
rlabel metal1 32844 21862 32844 21862 0 _0762_
rlabel metal1 33074 23732 33074 23732 0 _0763_
rlabel metal2 31418 25058 31418 25058 0 _0764_
rlabel metal1 32844 25126 32844 25126 0 _0765_
rlabel metal1 32706 25466 32706 25466 0 _0766_
rlabel metal1 32062 26214 32062 26214 0 _0767_
rlabel metal1 30774 24820 30774 24820 0 _0768_
rlabel metal1 30452 26010 30452 26010 0 _0769_
rlabel metal1 29486 26350 29486 26350 0 _0770_
rlabel metal1 28888 26350 28888 26350 0 _0771_
rlabel metal1 30084 23154 30084 23154 0 _0772_
rlabel metal1 29164 23018 29164 23018 0 _0773_
rlabel metal2 28382 23494 28382 23494 0 _0774_
rlabel metal1 27278 24276 27278 24276 0 _0775_
rlabel metal1 23276 32946 23276 32946 0 _0776_
rlabel metal2 22310 27404 22310 27404 0 _0777_
rlabel metal1 22586 29138 22586 29138 0 _0778_
rlabel metal3 35052 34680 35052 34680 0 clk
rlabel metal1 8878 25466 8878 25466 0 clk8.count\[0\]
rlabel metal1 10626 29070 10626 29070 0 clk8.count\[10\]
rlabel metal1 9108 29546 9108 29546 0 clk8.count\[11\]
rlabel metal1 9522 32334 9522 32334 0 clk8.count\[12\]
rlabel metal1 9246 32300 9246 32300 0 clk8.count\[13\]
rlabel metal1 10074 32402 10074 32402 0 clk8.count\[14\]
rlabel metal1 8878 33898 8878 33898 0 clk8.count\[15\]
rlabel metal2 6394 32572 6394 32572 0 clk8.count\[16\]
rlabel metal1 5520 33286 5520 33286 0 clk8.count\[17\]
rlabel metal1 4692 31994 4692 31994 0 clk8.count\[18\]
rlabel metal2 4554 32028 4554 32028 0 clk8.count\[19\]
rlabel metal1 6900 25126 6900 25126 0 clk8.count\[1\]
rlabel metal1 6992 31314 6992 31314 0 clk8.count\[20\]
rlabel via1 7214 25126 7214 25126 0 clk8.count\[2\]
rlabel metal1 5658 25874 5658 25874 0 clk8.count\[3\]
rlabel metal1 4830 25772 4830 25772 0 clk8.count\[4\]
rlabel metal1 5474 25942 5474 25942 0 clk8.count\[5\]
rlabel metal1 5842 28492 5842 28492 0 clk8.count\[6\]
rlabel metal1 5474 29138 5474 29138 0 clk8.count\[7\]
rlabel metal1 6256 28526 6256 28526 0 clk8.count\[8\]
rlabel metal1 8234 29614 8234 29614 0 clk8.count\[9\]
rlabel metal1 7314 26010 7314 26010 0 clk8.next_count\[0\]
rlabel metal1 9200 28458 9200 28458 0 clk8.next_count\[10\]
rlabel metal1 10810 29104 10810 29104 0 clk8.next_count\[11\]
rlabel metal1 11178 31450 11178 31450 0 clk8.next_count\[12\]
rlabel metal1 7958 31654 7958 31654 0 clk8.next_count\[13\]
rlabel metal1 9200 32810 9200 32810 0 clk8.next_count\[14\]
rlabel metal2 7958 34782 7958 34782 0 clk8.next_count\[15\]
rlabel metal1 6624 33626 6624 33626 0 clk8.next_count\[16\]
rlabel metal2 4646 34272 4646 34272 0 clk8.next_count\[17\]
rlabel metal1 2254 31994 2254 31994 0 clk8.next_count\[18\]
rlabel metal1 3174 30906 3174 30906 0 clk8.next_count\[19\]
rlabel metal1 8326 25806 8326 25806 0 clk8.next_count\[1\]
rlabel metal1 5743 30906 5743 30906 0 clk8.next_count\[20\]
rlabel metal2 6578 23970 6578 23970 0 clk8.next_count\[2\]
rlabel metal1 4094 23800 4094 23800 0 clk8.next_count\[3\]
rlabel metal2 2898 24922 2898 24922 0 clk8.next_count\[4\]
rlabel metal1 3864 26282 3864 26282 0 clk8.next_count\[5\]
rlabel metal1 1886 28152 1886 28152 0 clk8.next_count\[6\]
rlabel metal2 4094 29410 4094 29410 0 clk8.next_count\[7\]
rlabel metal1 5513 27642 5513 27642 0 clk8.next_count\[8\]
rlabel metal2 8602 28254 8602 28254 0 clk8.next_count\[9\]
rlabel metal1 13018 29546 13018 29546 0 clk_div.count\[0\]
rlabel metal1 11684 27302 11684 27302 0 clk_div.count\[1\]
rlabel metal1 11316 27098 11316 27098 0 clk_div.count\[2\]
rlabel metal2 11730 25024 11730 25024 0 clk_div.count\[3\]
rlabel metal1 12374 24684 12374 24684 0 clk_div.count\[4\]
rlabel metal2 12190 24990 12190 24990 0 clk_div.count\[5\]
rlabel metal1 14904 26350 14904 26350 0 clk_div.count\[6\]
rlabel metal1 16514 25296 16514 25296 0 clk_div.count\[7\]
rlabel metal1 11730 29070 11730 29070 0 clk_div.next_count\[0\]
rlabel metal1 12880 26554 12880 26554 0 clk_div.next_count\[1\]
rlabel metal1 9890 27064 9890 27064 0 clk_div.next_count\[2\]
rlabel metal1 10074 24922 10074 24922 0 clk_div.next_count\[3\]
rlabel metal1 11086 23154 11086 23154 0 clk_div.next_count\[4\]
rlabel metal1 13294 24922 13294 24922 0 clk_div.next_count\[5\]
rlabel metal1 14122 27064 14122 27064 0 clk_div.next_count\[6\]
rlabel metal1 15272 24378 15272 24378 0 clk_div.next_count\[7\]
rlabel metal1 15410 29240 15410 29240 0 clknet_0_clk
rlabel metal1 2070 6834 2070 6834 0 clknet_4_0_0_clk
rlabel metal2 34362 5202 34362 5202 0 clknet_4_10_0_clk
rlabel metal1 27048 16082 27048 16082 0 clknet_4_11_0_clk
rlabel metal1 21850 24650 21850 24650 0 clknet_4_12_0_clk
rlabel metal1 21804 28594 21804 28594 0 clknet_4_13_0_clk
rlabel metal2 27002 21046 27002 21046 0 clknet_4_14_0_clk
rlabel metal1 32292 34510 32292 34510 0 clknet_4_15_0_clk
rlabel metal2 1426 19074 1426 19074 0 clknet_4_1_0_clk
rlabel metal2 13800 16626 13800 16626 0 clknet_4_2_0_clk
rlabel metal1 18354 21590 18354 21590 0 clknet_4_3_0_clk
rlabel metal1 1886 24650 1886 24650 0 clknet_4_4_0_clk
rlabel metal1 1886 32266 1886 32266 0 clknet_4_5_0_clk
rlabel metal2 13938 24548 13938 24548 0 clknet_4_6_0_clk
rlabel metal1 17342 34646 17342 34646 0 clknet_4_7_0_clk
rlabel metal2 18446 10064 18446 10064 0 clknet_4_8_0_clk
rlabel metal1 18400 18190 18400 18190 0 clknet_4_9_0_clk
rlabel metal3 820 32708 820 32708 0 en
rlabel metal2 30958 1027 30958 1027 0 keypad_i[0]
rlabel metal3 820 6188 820 6188 0 keypad_i[10]
rlabel metal3 820 19788 820 19788 0 keypad_i[11]
rlabel metal1 8234 35020 8234 35020 0 keypad_i[12]
rlabel metal1 13892 35054 13892 35054 0 keypad_i[13]
rlabel metal1 33028 35054 33028 35054 0 keypad_i[14]
rlabel metal1 34592 8466 34592 8466 0 keypad_i[1]
rlabel metal2 24518 1588 24518 1588 0 keypad_i[2]
rlabel metal2 46 1588 46 1588 0 keypad_i[3]
rlabel metal2 5842 1027 5842 1027 0 keypad_i[4]
rlabel metal3 820 12988 820 12988 0 keypad_i[5]
rlabel metal1 34408 2414 34408 2414 0 keypad_i[6]
rlabel metal2 12282 1588 12282 1588 0 keypad_i[7]
rlabel metal1 34592 21522 34592 21522 0 keypad_i[8]
rlabel metal1 34362 28016 34362 28016 0 keypad_i[9]
rlabel metal1 16928 34170 16928 34170 0 kp_encoder.last_mk
rlabel metal1 15318 21624 15318 21624 0 kp_encoder.last_sk
rlabel metal2 30222 4624 30222 4624 0 kp_encoder.q\[0\]
rlabel metal1 5566 6834 5566 6834 0 kp_encoder.q\[10\]
rlabel metal2 8510 19329 8510 19329 0 kp_encoder.q\[11\]
rlabel metal1 11822 28594 11822 28594 0 kp_encoder.q\[12\]
rlabel metal1 14214 33966 14214 33966 0 kp_encoder.q\[13\]
rlabel metal1 33856 34034 33856 34034 0 kp_encoder.q\[14\]
rlabel metal1 32614 7956 32614 7956 0 kp_encoder.q\[1\]
rlabel metal1 17480 3706 17480 3706 0 kp_encoder.q\[2\]
rlabel metal1 13984 5746 13984 5746 0 kp_encoder.q\[3\]
rlabel metal1 9844 6426 9844 6426 0 kp_encoder.q\[4\]
rlabel metal1 3404 10642 3404 10642 0 kp_encoder.q\[5\]
rlabel metal1 14444 4250 14444 4250 0 kp_encoder.q\[6\]
rlabel metal1 13754 4046 13754 4046 0 kp_encoder.q\[7\]
rlabel metal1 32177 20774 32177 20774 0 kp_encoder.q\[8\]
rlabel metal2 32614 26877 32614 26877 0 kp_encoder.q\[9\]
rlabel metal2 15962 6324 15962 6324 0 kp_encoder.sync_out\[0\]
rlabel metal1 15594 13872 15594 13872 0 kp_encoder.sync_out\[10\]
rlabel metal2 15318 18224 15318 18224 0 kp_encoder.sync_out\[11\]
rlabel metal1 14812 23494 14812 23494 0 kp_encoder.sync_out\[12\]
rlabel metal1 16054 34510 16054 34510 0 kp_encoder.sync_out\[13\]
rlabel metal2 32614 30464 32614 30464 0 kp_encoder.sync_out\[14\]
rlabel metal1 16376 7514 16376 7514 0 kp_encoder.sync_out\[1\]
rlabel metal1 16882 7344 16882 7344 0 kp_encoder.sync_out\[2\]
rlabel metal1 15732 6698 15732 6698 0 kp_encoder.sync_out\[3\]
rlabel metal1 15042 8874 15042 8874 0 kp_encoder.sync_out\[4\]
rlabel metal1 4462 9010 4462 9010 0 kp_encoder.sync_out\[5\]
rlabel metal1 14812 8942 14812 8942 0 kp_encoder.sync_out\[6\]
rlabel metal1 14628 8874 14628 8874 0 kp_encoder.sync_out\[7\]
rlabel metal1 14720 16558 14720 16558 0 kp_encoder.sync_out\[8\]
rlabel metal1 15364 16762 15364 16762 0 kp_encoder.sync_out\[9\]
rlabel metal1 21344 33490 21344 33490 0 mode_FSM.mode\[0\]
rlabel metal1 19412 32810 19412 32810 0 mode_FSM.mode\[1\]
rlabel metal1 20056 35054 20056 35054 0 n_rst
rlabel metal1 16054 18700 16054 18700 0 net1
rlabel metal1 6716 2278 6716 2278 0 net10
rlabel metal1 27462 16184 27462 16184 0 net100
rlabel metal1 8418 31858 8418 31858 0 net101
rlabel metal1 7353 30906 7353 30906 0 net102
rlabel metal1 3680 25262 3680 25262 0 net103
rlabel metal1 24794 8942 24794 8942 0 net104
rlabel metal2 7038 33932 7038 33932 0 net105
rlabel metal1 3450 29172 3450 29172 0 net106
rlabel metal1 31326 10710 31326 10710 0 net107
rlabel metal1 27554 23630 27554 23630 0 net108
rlabel metal1 27462 23732 27462 23732 0 net109
rlabel metal1 6808 2618 6808 2618 0 net11
rlabel metal1 9706 29138 9706 29138 0 net110
rlabel metal2 28474 26826 28474 26826 0 net111
rlabel metal1 9154 22950 9154 22950 0 net112
rlabel metal1 27278 5168 27278 5168 0 net113
rlabel metal1 31418 26350 31418 26350 0 net114
rlabel metal1 27508 20910 27508 20910 0 net115
rlabel metal1 6900 21998 6900 21998 0 net116
rlabel metal1 31602 21896 31602 21896 0 net117
rlabel metal1 27738 10642 27738 10642 0 net118
rlabel metal1 27278 18666 27278 18666 0 net119
rlabel metal2 1702 12172 1702 12172 0 net12
rlabel metal1 22724 28050 22724 28050 0 net120
rlabel metal1 27370 31450 27370 31450 0 net121
rlabel metal1 25714 30226 25714 30226 0 net122
rlabel metal1 21804 5678 21804 5678 0 net123
rlabel metal1 23598 9554 23598 9554 0 net124
rlabel metal1 23552 21930 23552 21930 0 net125
rlabel metal1 22632 5202 22632 5202 0 net126
rlabel metal1 25668 9962 25668 9962 0 net127
rlabel metal1 22816 7786 22816 7786 0 net128
rlabel metal1 22678 26010 22678 26010 0 net129
rlabel metal1 20953 2482 20953 2482 0 net13
rlabel metal1 20332 26350 20332 26350 0 net130
rlabel metal1 12282 2618 12282 2618 0 net14
rlabel metal1 34178 20978 34178 20978 0 net15
rlabel metal1 34417 27642 34417 27642 0 net16
rlabel metal2 17388 17204 17388 17204 0 net17
rlabel metal1 26588 34714 26588 34714 0 net18
rlabel metal1 18170 2414 18170 2414 0 net19
rlabel metal1 31464 2618 31464 2618 0 net2
rlabel metal2 1932 20196 1932 20196 0 net20
rlabel metal2 1840 20060 1840 20060 0 net21
rlabel metal1 34132 14382 34132 14382 0 net22
rlabel metal1 4370 19992 4370 19992 0 net23
rlabel metal1 11592 20570 11592 20570 0 net24
rlabel metal1 10718 18802 10718 18802 0 net25
rlabel metal1 5934 15878 5934 15878 0 net26
rlabel metal1 4922 17714 4922 17714 0 net27
rlabel metal1 16659 11118 16659 11118 0 net28
rlabel metal1 8885 30634 8885 30634 0 net29
rlabel metal1 1656 6426 1656 6426 0 net3
rlabel metal2 14766 19924 14766 19924 0 net30
rlabel metal1 16567 32878 16567 32878 0 net31
rlabel metal1 15916 34578 15916 34578 0 net32
rlabel via1 19550 18309 19550 18309 0 net33
rlabel metal1 32561 6290 32561 6290 0 net34
rlabel metal2 19734 20672 19734 20672 0 net35
rlabel metal2 18998 27472 18998 27472 0 net36
rlabel metal1 32943 22610 32943 22610 0 net37
rlabel metal2 32982 30158 32982 30158 0 net38
rlabel metal2 12466 7650 12466 7650 0 net39
rlabel metal1 1656 19414 1656 19414 0 net4
rlabel metal2 14122 6052 14122 6052 0 net40
rlabel metal1 3036 9622 3036 9622 0 net41
rlabel metal1 10626 7446 10626 7446 0 net42
rlabel metal1 14720 34170 14720 34170 0 net43
rlabel metal1 13248 4794 13248 4794 0 net44
rlabel metal1 15778 4794 15778 4794 0 net45
rlabel metal1 34224 32810 34224 32810 0 net46
rlabel metal1 11454 19414 11454 19414 0 net47
rlabel metal2 19458 4250 19458 4250 0 net48
rlabel metal1 21758 5576 21758 5576 0 net49
rlabel metal1 9844 34646 9844 34646 0 net5
rlabel metal1 15640 33898 15640 33898 0 net50
rlabel metal2 13202 26078 13202 26078 0 net51
rlabel metal1 18998 20332 18998 20332 0 net52
rlabel metal2 19642 7582 19642 7582 0 net53
rlabel metal1 15686 22576 15686 22576 0 net54
rlabel metal2 24334 25296 24334 25296 0 net55
rlabel metal1 6440 31450 6440 31450 0 net56
rlabel metal1 29486 29138 29486 29138 0 net57
rlabel metal1 17986 27472 17986 27472 0 net58
rlabel metal1 24380 33626 24380 33626 0 net59
rlabel metal1 12650 34680 12650 34680 0 net6
rlabel metal1 26588 33626 26588 33626 0 net60
rlabel metal1 17112 33490 17112 33490 0 net61
rlabel metal1 27370 32742 27370 32742 0 net62
rlabel metal1 25392 31994 25392 31994 0 net63
rlabel metal1 12328 29478 12328 29478 0 net64
rlabel metal1 8142 25126 8142 25126 0 net65
rlabel metal1 9200 24718 9200 24718 0 net66
rlabel metal1 17526 32436 17526 32436 0 net67
rlabel metal1 25162 5304 25162 5304 0 net68
rlabel metal1 25300 5746 25300 5746 0 net69
rlabel metal1 32568 34646 32568 34646 0 net7
rlabel metal1 10902 24786 10902 24786 0 net70
rlabel metal1 16698 27438 16698 27438 0 net71
rlabel metal1 16323 26554 16323 26554 0 net72
rlabel metal2 27738 28356 27738 28356 0 net73
rlabel via1 27652 27642 27652 27642 0 net74
rlabel metal2 28106 30294 28106 30294 0 net75
rlabel metal1 26772 30362 26772 30362 0 net76
rlabel metal1 28428 31722 28428 31722 0 net77
rlabel metal1 28566 12138 28566 12138 0 net78
rlabel metal1 24334 29172 24334 29172 0 net79
rlabel metal2 34086 8092 34086 8092 0 net8
rlabel metal1 25852 29274 25852 29274 0 net80
rlabel metal1 23920 27642 23920 27642 0 net81
rlabel metal1 25530 27982 25530 27982 0 net82
rlabel metal1 29026 10098 29026 10098 0 net83
rlabel metal1 30360 28458 30360 28458 0 net84
rlabel metal1 29394 29580 29394 29580 0 net85
rlabel metal1 30360 28050 30360 28050 0 net86
rlabel metal1 27692 12818 27692 12818 0 net87
rlabel metal2 27830 17884 27830 17884 0 net88
rlabel metal1 29446 18054 29446 18054 0 net89
rlabel metal1 21436 3434 21436 3434 0 net9
rlabel metal1 4830 24140 4830 24140 0 net90
rlabel metal1 25668 19958 25668 19958 0 net91
rlabel via1 28191 20230 28191 20230 0 net92
rlabel metal1 12052 24038 12052 24038 0 net93
rlabel metal2 12374 27574 12374 27574 0 net94
rlabel metal1 13570 27098 13570 27098 0 net95
rlabel metal1 27968 7854 27968 7854 0 net96
rlabel metal1 17158 22746 17158 22746 0 net97
rlabel metal1 26818 14314 26818 14314 0 net98
rlabel metal1 25806 16218 25806 16218 0 net99
rlabel metal1 18998 8568 18998 8568 0 osc.count\[0\]
rlabel metal1 18630 19346 18630 19346 0 osc.count\[10\]
rlabel metal1 19780 20230 19780 20230 0 osc.count\[11\]
rlabel metal1 19044 20842 19044 20842 0 osc.count\[12\]
rlabel metal1 21850 21590 21850 21590 0 osc.count\[13\]
rlabel metal1 20562 21522 20562 21522 0 osc.count\[14\]
rlabel metal1 20654 20944 20654 20944 0 osc.count\[15\]
rlabel metal1 19136 7378 19136 7378 0 osc.count\[1\]
rlabel metal2 20470 8058 20470 8058 0 osc.count\[2\]
rlabel metal1 18446 7786 18446 7786 0 osc.count\[3\]
rlabel metal1 18630 10234 18630 10234 0 osc.count\[4\]
rlabel metal1 20286 11628 20286 11628 0 osc.count\[5\]
rlabel metal1 20562 11798 20562 11798 0 osc.count\[6\]
rlabel metal1 17848 12818 17848 12818 0 osc.count\[7\]
rlabel metal1 23460 17578 23460 17578 0 osc.count\[8\]
rlabel metal1 19412 17578 19412 17578 0 osc.count\[9\]
rlabel metal2 16422 22916 16422 22916 0 osc.next_count\[0\]
rlabel metal1 19136 18938 19136 18938 0 osc.next_count\[10\]
rlabel metal1 15909 21114 15909 21114 0 osc.next_count\[11\]
rlabel metal1 18722 21862 18722 21862 0 osc.next_count\[12\]
rlabel metal1 20010 23018 20010 23018 0 osc.next_count\[13\]
rlabel metal2 19550 25058 19550 25058 0 osc.next_count\[14\]
rlabel metal2 18262 25024 18262 25024 0 osc.next_count\[15\]
rlabel metal2 19550 5916 19550 5916 0 osc.next_count\[1\]
rlabel metal1 20010 7446 20010 7446 0 osc.next_count\[2\]
rlabel metal1 17381 6970 17381 6970 0 osc.next_count\[3\]
rlabel metal1 18584 9146 18584 9146 0 osc.next_count\[4\]
rlabel metal1 18538 10710 18538 10710 0 osc.next_count\[5\]
rlabel metal1 15180 11186 15180 11186 0 osc.next_count\[6\]
rlabel metal1 18446 11662 18446 11662 0 osc.next_count\[7\]
rlabel metal1 18538 16184 18538 16184 0 osc.next_count\[8\]
rlabel metal1 18814 18360 18814 18360 0 osc.next_count\[9\]
rlabel metal1 18860 27438 18860 27438 0 pwm.count\[0\]
rlabel metal1 17572 27438 17572 27438 0 pwm.count\[1\]
rlabel metal1 16882 29104 16882 29104 0 pwm.count\[2\]
rlabel metal1 17710 29580 17710 29580 0 pwm.count\[3\]
rlabel metal1 17820 30702 17820 30702 0 pwm.count\[4\]
rlabel metal1 17572 31314 17572 31314 0 pwm.count\[5\]
rlabel metal1 14306 31790 14306 31790 0 pwm.count\[6\]
rlabel metal2 17250 33184 17250 33184 0 pwm.count\[7\]
rlabel metal1 17434 27064 17434 27064 0 pwm.next_count\[0\]
rlabel metal1 16008 26962 16008 26962 0 pwm.next_count\[1\]
rlabel metal1 15594 29546 15594 29546 0 pwm.next_count\[2\]
rlabel metal1 14352 28458 14352 28458 0 pwm.next_count\[3\]
rlabel metal1 13241 30906 13241 30906 0 pwm.next_count\[4\]
rlabel metal2 15594 30940 15594 30940 0 pwm.next_count\[5\]
rlabel metal1 12926 31994 12926 31994 0 pwm.next_count\[6\]
rlabel metal1 15318 32946 15318 32946 0 pwm.next_count\[7\]
rlabel metal1 21758 34408 21758 34408 0 pwm.pwm
rlabel metal1 26818 35258 26818 35258 0 pwm_o
rlabel metal1 29762 6766 29762 6766 0 seq_div.D\[0\]
rlabel metal1 30176 19346 30176 19346 0 seq_div.D\[10\]
rlabel metal1 26266 20230 26266 20230 0 seq_div.D\[11\]
rlabel metal1 29072 21454 29072 21454 0 seq_div.D\[12\]
rlabel metal1 26680 24038 26680 24038 0 seq_div.D\[13\]
rlabel metal1 29279 25262 29279 25262 0 seq_div.D\[14\]
rlabel metal1 27646 21862 27646 21862 0 seq_div.D\[15\]
rlabel metal2 27830 7378 27830 7378 0 seq_div.D\[1\]
rlabel metal2 25990 4352 25990 4352 0 seq_div.D\[2\]
rlabel metal1 25484 7514 25484 7514 0 seq_div.D\[3\]
rlabel metal2 27830 9350 27830 9350 0 seq_div.D\[4\]
rlabel metal2 28750 10812 28750 10812 0 seq_div.D\[5\]
rlabel metal1 32338 12240 32338 12240 0 seq_div.D\[6\]
rlabel metal1 26404 14246 26404 14246 0 seq_div.D\[7\]
rlabel metal2 27554 15232 27554 15232 0 seq_div.D\[8\]
rlabel metal2 27646 17170 27646 17170 0 seq_div.D\[9\]
rlabel metal1 23460 27506 23460 27506 0 seq_div.Q\[0\]
rlabel metal1 23414 29138 23414 29138 0 seq_div.Q\[1\]
rlabel metal1 26450 29138 26450 29138 0 seq_div.Q\[2\]
rlabel metal1 27830 30906 27830 30906 0 seq_div.Q\[3\]
rlabel metal1 29440 31246 29440 31246 0 seq_div.Q\[4\]
rlabel metal1 27922 32334 27922 32334 0 seq_div.Q\[5\]
rlabel metal1 24656 32538 24656 32538 0 seq_div.Q\[6\]
rlabel metal1 25300 33490 25300 33490 0 seq_div.Q\[7\]
rlabel metal2 32614 7038 32614 7038 0 seq_div.R\[10\]
rlabel metal1 32200 6426 32200 6426 0 seq_div.R\[11\]
rlabel metal2 28198 10234 28198 10234 0 seq_div.R\[12\]
rlabel metal1 33856 12410 33856 12410 0 seq_div.R\[13\]
rlabel metal2 29578 11934 29578 11934 0 seq_div.R\[14\]
rlabel metal2 29394 14790 29394 14790 0 seq_div.R\[15\]
rlabel metal1 28566 15878 28566 15878 0 seq_div.R\[16\]
rlabel metal1 28152 18054 28152 18054 0 seq_div.R\[17\]
rlabel metal1 32499 20366 32499 20366 0 seq_div.R\[18\]
rlabel metal1 32936 22066 32936 22066 0 seq_div.R\[19\]
rlabel metal2 32614 24786 32614 24786 0 seq_div.R\[20\]
rlabel metal1 28750 25228 28750 25228 0 seq_div.R\[21\]
rlabel metal1 28152 26350 28152 26350 0 seq_div.R\[22\]
rlabel metal1 28658 23222 28658 23222 0 seq_div.R\[23\]
rlabel metal1 25760 5882 25760 5882 0 seq_div.R\[8\]
rlabel metal1 28244 5202 28244 5202 0 seq_div.R\[9\]
rlabel metal1 29808 28526 29808 28526 0 seq_div.count_div\[0\]
rlabel metal2 29670 28764 29670 28764 0 seq_div.count_div\[1\]
rlabel metal1 29072 29002 29072 29002 0 seq_div.count_div\[2\]
rlabel metal1 22586 6290 22586 6290 0 seq_div.dividend\[0\]
rlabel metal1 25254 19346 25254 19346 0 seq_div.dividend\[10\]
rlabel metal1 27255 22066 27255 22066 0 seq_div.dividend\[11\]
rlabel metal1 32430 23630 32430 23630 0 seq_div.dividend\[12\]
rlabel metal1 25576 26418 25576 26418 0 seq_div.dividend\[13\]
rlabel metal1 21574 26996 21574 26996 0 seq_div.dividend\[14\]
rlabel metal1 23506 24582 23506 24582 0 seq_div.dividend\[15\]
rlabel metal1 24104 5202 24104 5202 0 seq_div.dividend\[1\]
rlabel metal1 24380 7854 24380 7854 0 seq_div.dividend\[2\]
rlabel metal1 25392 5542 25392 5542 0 seq_div.dividend\[3\]
rlabel metal1 25484 10166 25484 10166 0 seq_div.dividend\[4\]
rlabel metal1 27554 10438 27554 10438 0 seq_div.dividend\[5\]
rlabel metal1 28382 12342 28382 12342 0 seq_div.dividend\[6\]
rlabel metal2 25714 14212 25714 14212 0 seq_div.dividend\[7\]
rlabel metal1 26036 16014 26036 16014 0 seq_div.dividend\[8\]
rlabel metal1 26588 18190 26588 18190 0 seq_div.dividend\[9\]
rlabel metal1 20056 28526 20056 28526 0 seq_div.q_out\[0\]
rlabel metal2 20470 28832 20470 28832 0 seq_div.q_out\[1\]
rlabel metal1 20700 29614 20700 29614 0 seq_div.q_out\[2\]
rlabel metal2 21298 30430 21298 30430 0 seq_div.q_out\[3\]
rlabel metal1 27048 31858 27048 31858 0 seq_div.q_out\[4\]
rlabel metal1 19780 31790 19780 31790 0 seq_div.q_out\[5\]
rlabel metal1 19642 32878 19642 32878 0 seq_div.q_out\[6\]
rlabel metal1 24334 33966 24334 33966 0 seq_div.q_out\[7\]
rlabel metal1 26036 27030 26036 27030 0 seq_div.state\[0\]
rlabel metal1 27830 26996 27830 26996 0 seq_div.state\[1\]
rlabel metal2 18722 823 18722 823 0 sound_series[0]
rlabel metal3 751 25908 751 25908 0 sound_series[1]
rlabel metal1 1426 35258 1426 35258 0 sound_series[2]
rlabel metal1 34500 14586 34500 14586 0 sound_series[3]
<< properties >>
string FIXED_BBOX 0 0 35873 38017
<< end >>
