magic
tech sky130A
magscale 1 2
timestamp 1694009784
<< obsli1 >>
rect 1104 2159 86112 87057
<< obsm1 >>
rect 14 2128 87018 87088
<< metal2 >>
rect 662 88604 718 89404
rect 18050 88604 18106 89404
rect 35438 88604 35494 89404
rect 52826 88604 52882 89404
rect 70214 88604 70270 89404
rect 86958 88604 87014 89404
rect 18 0 74 800
rect 16762 0 16818 800
rect 34150 0 34206 800
rect 51538 0 51594 800
rect 68926 0 68982 800
rect 86314 0 86370 800
<< obsm2 >>
rect 20 88548 606 88754
rect 774 88548 17994 88754
rect 18162 88548 35382 88754
rect 35550 88548 52770 88754
rect 52938 88548 70158 88754
rect 70326 88548 86902 88754
rect 20 856 87012 88548
rect 130 800 16706 856
rect 16874 800 34094 856
rect 34262 800 51482 856
rect 51650 800 68870 856
rect 69038 800 86258 856
rect 86426 800 87012 856
<< metal3 >>
rect 0 72768 800 72888
rect 86460 71408 87260 71528
rect 0 54408 800 54528
rect 86460 53048 87260 53168
rect 0 36048 800 36168
rect 86460 34688 87260 34808
rect 0 17688 800 17808
rect 86460 16328 87260 16448
<< obsm3 >>
rect 798 72968 86460 87073
rect 880 72688 86460 72968
rect 798 71608 86460 72688
rect 798 71328 86380 71608
rect 798 54608 86460 71328
rect 880 54328 86460 54608
rect 798 53248 86460 54328
rect 798 52968 86380 53248
rect 798 36248 86460 52968
rect 880 35968 86460 36248
rect 798 34888 86460 35968
rect 798 34608 86380 34888
rect 798 17888 86460 34608
rect 880 17608 86460 17888
rect 798 16528 86460 17608
rect 798 16248 86380 16528
rect 798 2143 86460 16248
<< metal4 >>
rect 4208 2128 4528 87088
rect 19568 2128 19888 87088
rect 34928 2128 35248 87088
rect 50288 2128 50608 87088
rect 65648 2128 65968 87088
rect 81008 2128 81328 87088
<< obsm4 >>
rect 10547 7379 19488 85645
rect 19968 7379 34848 85645
rect 35328 7379 50208 85645
rect 50688 7379 65568 85645
rect 66048 7379 80717 85645
<< labels >>
rlabel metal3 s 86460 16328 87260 16448 6 clk
port 1 nsew signal input
rlabel metal2 s 86958 88604 87014 89404 6 mode_out[0]
port 2 nsew signal output
rlabel metal2 s 52826 88604 52882 89404 6 mode_out[1]
port 3 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 pb[0]
port 4 nsew signal input
rlabel metal3 s 86460 71408 87260 71528 6 pb[10]
port 5 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 pb[11]
port 6 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 pb[12]
port 7 nsew signal input
rlabel metal2 s 35438 88604 35494 89404 6 pb[13]
port 8 nsew signal input
rlabel metal2 s 18 0 74 800 6 pb[14]
port 9 nsew signal input
rlabel metal2 s 18050 88604 18106 89404 6 pb[1]
port 10 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 pb[2]
port 11 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 pb[3]
port 12 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 pb[4]
port 13 nsew signal input
rlabel metal3 s 86460 53048 87260 53168 6 pb[5]
port 14 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 pb[6]
port 15 nsew signal input
rlabel metal2 s 70214 88604 70270 89404 6 pb[7]
port 16 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 pb[8]
port 17 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 pb[9]
port 18 nsew signal input
rlabel metal2 s 662 88604 718 89404 6 reset
port 19 nsew signal input
rlabel metal3 s 86460 34688 87260 34808 6 sigout
port 20 nsew signal output
rlabel metal4 s 4208 2128 4528 87088 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 87088 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 87088 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 87088 6 vssd1
port 22 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 87088 6 vssd1
port 22 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 87088 6 vssd1
port 22 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 87260 89404
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 25703472
string GDS_FILE /home/designer-25/CUP/openlane/tmnt/runs/23_09_06_06_59/results/signoff/top_asic.magic.gds
string GDS_START 1129380
<< end >>

