magic
tech sky130A
magscale 1 2
timestamp 1694412481
<< obsli1 >>
rect 1104 2159 53820 54417
<< obsm1 >>
rect 14 1776 54818 54936
<< metal2 >>
rect 662 56309 718 57109
rect 1950 56309 2006 57109
rect 3238 56309 3294 57109
rect 5170 56309 5226 57109
rect 6458 56309 6514 57109
rect 8390 56309 8446 57109
rect 9678 56309 9734 57109
rect 11610 56309 11666 57109
rect 12898 56309 12954 57109
rect 14186 56309 14242 57109
rect 16118 56309 16174 57109
rect 17406 56309 17462 57109
rect 19338 56309 19394 57109
rect 20626 56309 20682 57109
rect 22558 56309 22614 57109
rect 23846 56309 23902 57109
rect 25134 56309 25190 57109
rect 27066 56309 27122 57109
rect 28354 56309 28410 57109
rect 30286 56309 30342 57109
rect 31574 56309 31630 57109
rect 33506 56309 33562 57109
rect 34794 56309 34850 57109
rect 36082 56309 36138 57109
rect 38014 56309 38070 57109
rect 39302 56309 39358 57109
rect 41234 56309 41290 57109
rect 42522 56309 42578 57109
rect 44454 56309 44510 57109
rect 45742 56309 45798 57109
rect 47030 56309 47086 57109
rect 48962 56309 49018 57109
rect 50250 56309 50306 57109
rect 52182 56309 52238 57109
rect 53470 56309 53526 57109
rect 54758 56309 54814 57109
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 48318 0 48374 800
rect 49606 0 49662 800
rect 51538 0 51594 800
rect 52826 0 52882 800
rect 54758 0 54814 800
<< obsm2 >>
rect 20 56253 606 56309
rect 774 56253 1894 56309
rect 2062 56253 3182 56309
rect 3350 56253 5114 56309
rect 5282 56253 6402 56309
rect 6570 56253 8334 56309
rect 8502 56253 9622 56309
rect 9790 56253 11554 56309
rect 11722 56253 12842 56309
rect 13010 56253 14130 56309
rect 14298 56253 16062 56309
rect 16230 56253 17350 56309
rect 17518 56253 19282 56309
rect 19450 56253 20570 56309
rect 20738 56253 22502 56309
rect 22670 56253 23790 56309
rect 23958 56253 25078 56309
rect 25246 56253 27010 56309
rect 27178 56253 28298 56309
rect 28466 56253 30230 56309
rect 30398 56253 31518 56309
rect 31686 56253 33450 56309
rect 33618 56253 34738 56309
rect 34906 56253 36026 56309
rect 36194 56253 37958 56309
rect 38126 56253 39246 56309
rect 39414 56253 41178 56309
rect 41346 56253 42466 56309
rect 42634 56253 44398 56309
rect 44566 56253 45686 56309
rect 45854 56253 46974 56309
rect 47142 56253 48906 56309
rect 49074 56253 50194 56309
rect 50362 56253 52126 56309
rect 52294 56253 53414 56309
rect 53582 56253 54702 56309
rect 20 856 54812 56253
rect 130 711 1250 856
rect 1418 711 2538 856
rect 2706 711 4470 856
rect 4638 711 5758 856
rect 5926 711 7690 856
rect 7858 711 8978 856
rect 9146 711 10910 856
rect 11078 711 12198 856
rect 12366 711 13486 856
rect 13654 711 15418 856
rect 15586 711 16706 856
rect 16874 711 18638 856
rect 18806 711 19926 856
rect 20094 711 21858 856
rect 22026 711 23146 856
rect 23314 711 24434 856
rect 24602 711 26366 856
rect 26534 711 27654 856
rect 27822 711 29586 856
rect 29754 711 30874 856
rect 31042 711 32162 856
rect 32330 711 34094 856
rect 34262 711 35382 856
rect 35550 711 37314 856
rect 37482 711 38602 856
rect 38770 711 40534 856
rect 40702 711 41822 856
rect 41990 711 43754 856
rect 43922 711 45042 856
rect 45210 711 46330 856
rect 46498 711 48262 856
rect 48430 711 49550 856
rect 49718 711 51482 856
rect 51650 711 52770 856
rect 52938 711 54702 856
<< metal3 >>
rect 0 55768 800 55888
rect 54165 55088 54965 55208
rect 0 54408 800 54528
rect 54165 53728 54965 53848
rect 0 52368 800 52488
rect 54165 51688 54965 51808
rect 0 51008 800 51128
rect 54165 50328 54965 50448
rect 0 48968 800 49088
rect 54165 48288 54965 48408
rect 0 47608 800 47728
rect 54165 46928 54965 47048
rect 0 45568 800 45688
rect 54165 45568 54965 45688
rect 0 44208 800 44328
rect 54165 43528 54965 43648
rect 0 42848 800 42968
rect 54165 42168 54965 42288
rect 0 40808 800 40928
rect 54165 40128 54965 40248
rect 0 39448 800 39568
rect 54165 38768 54965 38888
rect 0 37408 800 37528
rect 54165 36728 54965 36848
rect 0 36048 800 36168
rect 54165 35368 54965 35488
rect 0 34008 800 34128
rect 54165 34008 54965 34128
rect 0 32648 800 32768
rect 54165 31968 54965 32088
rect 0 31288 800 31408
rect 54165 30608 54965 30728
rect 0 29248 800 29368
rect 54165 28568 54965 28688
rect 0 27888 800 28008
rect 54165 27208 54965 27328
rect 0 25848 800 25968
rect 54165 25168 54965 25288
rect 0 24488 800 24608
rect 54165 23808 54965 23928
rect 0 22448 800 22568
rect 54165 21768 54965 21888
rect 0 21088 800 21208
rect 54165 20408 54965 20528
rect 0 19728 800 19848
rect 54165 19048 54965 19168
rect 0 17688 800 17808
rect 54165 17008 54965 17128
rect 0 16328 800 16448
rect 54165 15648 54965 15768
rect 0 14288 800 14408
rect 54165 13608 54965 13728
rect 0 12928 800 13048
rect 54165 12248 54965 12368
rect 0 10888 800 11008
rect 54165 10208 54965 10328
rect 0 9528 800 9648
rect 54165 8848 54965 8968
rect 0 8168 800 8288
rect 54165 7488 54965 7608
rect 0 6128 800 6248
rect 54165 5448 54965 5568
rect 0 4768 800 4888
rect 54165 4088 54965 4208
rect 0 2728 800 2848
rect 54165 2048 54965 2168
rect 0 1368 800 1488
rect 54165 688 54965 808
<< obsm3 >>
rect 880 55688 54727 55861
rect 800 55288 54727 55688
rect 800 55008 54085 55288
rect 800 54608 54727 55008
rect 880 54328 54727 54608
rect 800 53928 54727 54328
rect 800 53648 54085 53928
rect 800 52568 54727 53648
rect 880 52288 54727 52568
rect 800 51888 54727 52288
rect 800 51608 54085 51888
rect 800 51208 54727 51608
rect 880 50928 54727 51208
rect 800 50528 54727 50928
rect 800 50248 54085 50528
rect 800 49168 54727 50248
rect 880 48888 54727 49168
rect 800 48488 54727 48888
rect 800 48208 54085 48488
rect 800 47808 54727 48208
rect 880 47528 54727 47808
rect 800 47128 54727 47528
rect 800 46848 54085 47128
rect 800 45768 54727 46848
rect 880 45488 54085 45768
rect 800 44408 54727 45488
rect 880 44128 54727 44408
rect 800 43728 54727 44128
rect 800 43448 54085 43728
rect 800 43048 54727 43448
rect 880 42768 54727 43048
rect 800 42368 54727 42768
rect 800 42088 54085 42368
rect 800 41008 54727 42088
rect 880 40728 54727 41008
rect 800 40328 54727 40728
rect 800 40048 54085 40328
rect 800 39648 54727 40048
rect 880 39368 54727 39648
rect 800 38968 54727 39368
rect 800 38688 54085 38968
rect 800 37608 54727 38688
rect 880 37328 54727 37608
rect 800 36928 54727 37328
rect 800 36648 54085 36928
rect 800 36248 54727 36648
rect 880 35968 54727 36248
rect 800 35568 54727 35968
rect 800 35288 54085 35568
rect 800 34208 54727 35288
rect 880 33928 54085 34208
rect 800 32848 54727 33928
rect 880 32568 54727 32848
rect 800 32168 54727 32568
rect 800 31888 54085 32168
rect 800 31488 54727 31888
rect 880 31208 54727 31488
rect 800 30808 54727 31208
rect 800 30528 54085 30808
rect 800 29448 54727 30528
rect 880 29168 54727 29448
rect 800 28768 54727 29168
rect 800 28488 54085 28768
rect 800 28088 54727 28488
rect 880 27808 54727 28088
rect 800 27408 54727 27808
rect 800 27128 54085 27408
rect 800 26048 54727 27128
rect 880 25768 54727 26048
rect 800 25368 54727 25768
rect 800 25088 54085 25368
rect 800 24688 54727 25088
rect 880 24408 54727 24688
rect 800 24008 54727 24408
rect 800 23728 54085 24008
rect 800 22648 54727 23728
rect 880 22368 54727 22648
rect 800 21968 54727 22368
rect 800 21688 54085 21968
rect 800 21288 54727 21688
rect 880 21008 54727 21288
rect 800 20608 54727 21008
rect 800 20328 54085 20608
rect 800 19928 54727 20328
rect 880 19648 54727 19928
rect 800 19248 54727 19648
rect 800 18968 54085 19248
rect 800 17888 54727 18968
rect 880 17608 54727 17888
rect 800 17208 54727 17608
rect 800 16928 54085 17208
rect 800 16528 54727 16928
rect 880 16248 54727 16528
rect 800 15848 54727 16248
rect 800 15568 54085 15848
rect 800 14488 54727 15568
rect 880 14208 54727 14488
rect 800 13808 54727 14208
rect 800 13528 54085 13808
rect 800 13128 54727 13528
rect 880 12848 54727 13128
rect 800 12448 54727 12848
rect 800 12168 54085 12448
rect 800 11088 54727 12168
rect 880 10808 54727 11088
rect 800 10408 54727 10808
rect 800 10128 54085 10408
rect 800 9728 54727 10128
rect 880 9448 54727 9728
rect 800 9048 54727 9448
rect 800 8768 54085 9048
rect 800 8368 54727 8768
rect 880 8088 54727 8368
rect 800 7688 54727 8088
rect 800 7408 54085 7688
rect 800 6328 54727 7408
rect 880 6048 54727 6328
rect 800 5648 54727 6048
rect 800 5368 54085 5648
rect 800 4968 54727 5368
rect 880 4688 54727 4968
rect 800 4288 54727 4688
rect 800 4008 54085 4288
rect 800 2928 54727 4008
rect 880 2648 54727 2928
rect 800 2248 54727 2648
rect 800 1968 54085 2248
rect 800 1568 54727 1968
rect 880 1288 54727 1568
rect 800 888 54727 1288
rect 800 715 54085 888
<< metal4 >>
rect 4208 2128 4528 54448
rect 19568 2128 19888 54448
rect 34928 2128 35248 54448
rect 50288 2128 50608 54448
<< obsm4 >>
rect 6683 2211 19488 54093
rect 19968 2211 34848 54093
rect 35328 2211 50208 54093
rect 50688 2211 52381 54093
<< labels >>
rlabel metal2 s 15474 0 15530 800 6 clk
port 1 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 interrupt_gpio_in
port 2 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 keypad_input[0]
port 3 nsew signal input
rlabel metal3 s 54165 688 54965 808 6 keypad_input[10]
port 4 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 keypad_input[11]
port 5 nsew signal input
rlabel metal2 s 52182 56309 52238 57109 6 keypad_input[12]
port 6 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 keypad_input[13]
port 7 nsew signal input
rlabel metal3 s 54165 15648 54965 15768 6 keypad_input[14]
port 8 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 keypad_input[15]
port 9 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 keypad_input[1]
port 10 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 keypad_input[2]
port 11 nsew signal input
rlabel metal2 s 38014 56309 38070 57109 6 keypad_input[3]
port 12 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 keypad_input[4]
port 13 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 keypad_input[5]
port 14 nsew signal input
rlabel metal2 s 23846 56309 23902 57109 6 keypad_input[6]
port 15 nsew signal input
rlabel metal3 s 54165 10208 54965 10328 6 keypad_input[7]
port 16 nsew signal input
rlabel metal3 s 54165 35368 54965 35488 6 keypad_input[8]
port 17 nsew signal input
rlabel metal2 s 47030 56309 47086 57109 6 keypad_input[9]
port 18 nsew signal input
rlabel metal2 s 53470 56309 53526 57109 6 memory_address_out[0]
port 19 nsew signal output
rlabel metal2 s 17406 56309 17462 57109 6 memory_address_out[10]
port 20 nsew signal output
rlabel metal2 s 28354 56309 28410 57109 6 memory_address_out[11]
port 21 nsew signal output
rlabel metal3 s 54165 40128 54965 40248 6 memory_address_out[12]
port 22 nsew signal output
rlabel metal2 s 50250 56309 50306 57109 6 memory_address_out[13]
port 23 nsew signal output
rlabel metal3 s 54165 7488 54965 7608 6 memory_address_out[14]
port 24 nsew signal output
rlabel metal2 s 45742 56309 45798 57109 6 memory_address_out[15]
port 25 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 memory_address_out[1]
port 26 nsew signal output
rlabel metal3 s 54165 43528 54965 43648 6 memory_address_out[2]
port 27 nsew signal output
rlabel metal2 s 5170 56309 5226 57109 6 memory_address_out[3]
port 28 nsew signal output
rlabel metal2 s 31574 56309 31630 57109 6 memory_address_out[4]
port 29 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 memory_address_out[5]
port 30 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 memory_address_out[6]
port 31 nsew signal output
rlabel metal3 s 54165 17008 54965 17128 6 memory_address_out[7]
port 32 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 memory_address_out[8]
port 33 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 memory_address_out[9]
port 34 nsew signal output
rlabel metal3 s 54165 25168 54965 25288 6 memory_data_in[0]
port 35 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 memory_data_in[1]
port 36 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 memory_data_in[2]
port 37 nsew signal input
rlabel metal2 s 6458 56309 6514 57109 6 memory_data_in[3]
port 38 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 memory_data_in[4]
port 39 nsew signal input
rlabel metal2 s 36082 56309 36138 57109 6 memory_data_in[5]
port 40 nsew signal input
rlabel metal2 s 27066 56309 27122 57109 6 memory_data_in[6]
port 41 nsew signal input
rlabel metal3 s 54165 38768 54965 38888 6 memory_data_in[7]
port 42 nsew signal input
rlabel metal3 s 54165 45568 54965 45688 6 memory_data_out[0]
port 43 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 memory_data_out[1]
port 44 nsew signal output
rlabel metal3 s 54165 23808 54965 23928 6 memory_data_out[2]
port 45 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 memory_data_out[3]
port 46 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 memory_data_out[4]
port 47 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 memory_data_out[5]
port 48 nsew signal output
rlabel metal3 s 54165 2048 54965 2168 6 memory_data_out[6]
port 49 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 memory_data_out[7]
port 50 nsew signal output
rlabel metal3 s 54165 30608 54965 30728 6 memory_wr
port 51 nsew signal output
rlabel metal2 s 44454 56309 44510 57109 6 nrst
port 52 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 programmable_gpio_in[0]
port 53 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 programmable_gpio_in[1]
port 54 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 programmable_gpio_in[2]
port 55 nsew signal input
rlabel metal3 s 54165 50328 54965 50448 6 programmable_gpio_in[3]
port 56 nsew signal input
rlabel metal3 s 54165 19048 54965 19168 6 programmable_gpio_in[4]
port 57 nsew signal input
rlabel metal2 s 16118 56309 16174 57109 6 programmable_gpio_in[5]
port 58 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 programmable_gpio_in[6]
port 59 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 programmable_gpio_in[7]
port 60 nsew signal input
rlabel metal2 s 22558 56309 22614 57109 6 programmable_gpio_out[0]
port 61 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 programmable_gpio_out[1]
port 62 nsew signal output
rlabel metal3 s 54165 46928 54965 47048 6 programmable_gpio_out[2]
port 63 nsew signal output
rlabel metal3 s 54165 12248 54965 12368 6 programmable_gpio_out[3]
port 64 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 programmable_gpio_out[4]
port 65 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 programmable_gpio_out[5]
port 66 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 programmable_gpio_out[6]
port 67 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 programmable_gpio_out[7]
port 68 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 programmable_gpio_wr[0]
port 69 nsew signal output
rlabel metal3 s 54165 34008 54965 34128 6 programmable_gpio_wr[1]
port 70 nsew signal output
rlabel metal2 s 11610 56309 11666 57109 6 programmable_gpio_wr[2]
port 71 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 programmable_gpio_wr[3]
port 72 nsew signal output
rlabel metal3 s 54165 53728 54965 53848 6 programmable_gpio_wr[4]
port 73 nsew signal output
rlabel metal2 s 25134 56309 25190 57109 6 programmable_gpio_wr[5]
port 74 nsew signal output
rlabel metal2 s 1950 56309 2006 57109 6 programmable_gpio_wr[6]
port 75 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 programmable_gpio_wr[7]
port 76 nsew signal output
rlabel metal2 s 19338 56309 19394 57109 6 ss0[0]
port 77 nsew signal output
rlabel metal2 s 12898 56309 12954 57109 6 ss0[1]
port 78 nsew signal output
rlabel metal2 s 8390 56309 8446 57109 6 ss0[2]
port 79 nsew signal output
rlabel metal3 s 54165 20408 54965 20528 6 ss0[3]
port 80 nsew signal output
rlabel metal3 s 54165 55088 54965 55208 6 ss0[4]
port 81 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 ss0[5]
port 82 nsew signal output
rlabel metal3 s 54165 4088 54965 4208 6 ss0[6]
port 83 nsew signal output
rlabel metal3 s 54165 21768 54965 21888 6 ss0[7]
port 84 nsew signal output
rlabel metal2 s 34794 56309 34850 57109 6 ss1[0]
port 85 nsew signal output
rlabel metal2 s 3238 56309 3294 57109 6 ss1[1]
port 86 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 ss1[2]
port 87 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 ss1[3]
port 88 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 ss1[4]
port 89 nsew signal output
rlabel metal2 s 54758 56309 54814 57109 6 ss1[5]
port 90 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 ss1[6]
port 91 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 ss1[7]
port 92 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 ss2[0]
port 93 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 ss2[1]
port 94 nsew signal output
rlabel metal2 s 20626 56309 20682 57109 6 ss2[2]
port 95 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 ss2[3]
port 96 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 ss2[4]
port 97 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 ss2[5]
port 98 nsew signal output
rlabel metal3 s 54165 5448 54965 5568 6 ss2[6]
port 99 nsew signal output
rlabel metal3 s 54165 42168 54965 42288 6 ss2[7]
port 100 nsew signal output
rlabel metal3 s 54165 28568 54965 28688 6 ss3[0]
port 101 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 ss3[1]
port 102 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 ss3[2]
port 103 nsew signal output
rlabel metal3 s 54165 13608 54965 13728 6 ss3[3]
port 104 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 ss3[4]
port 105 nsew signal output
rlabel metal3 s 54165 31968 54965 32088 6 ss3[5]
port 106 nsew signal output
rlabel metal3 s 54165 48288 54965 48408 6 ss3[6]
port 107 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 ss3[7]
port 108 nsew signal output
rlabel metal3 s 54165 51688 54965 51808 6 ss4[0]
port 109 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 ss4[1]
port 110 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 ss4[2]
port 111 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 ss4[3]
port 112 nsew signal output
rlabel metal2 s 18 0 74 800 6 ss4[4]
port 113 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 ss4[5]
port 114 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 ss4[6]
port 115 nsew signal output
rlabel metal2 s 14186 56309 14242 57109 6 ss4[7]
port 116 nsew signal output
rlabel metal2 s 33506 56309 33562 57109 6 ss5[0]
port 117 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 ss5[1]
port 118 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 ss5[2]
port 119 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 ss5[3]
port 120 nsew signal output
rlabel metal2 s 42522 56309 42578 57109 6 ss5[4]
port 121 nsew signal output
rlabel metal2 s 30286 56309 30342 57109 6 ss5[5]
port 122 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 ss5[6]
port 123 nsew signal output
rlabel metal2 s 48962 56309 49018 57109 6 ss5[7]
port 124 nsew signal output
rlabel metal3 s 54165 8848 54965 8968 6 ss6[0]
port 125 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 ss6[1]
port 126 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 ss6[2]
port 127 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 ss6[3]
port 128 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 ss6[4]
port 129 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 ss6[5]
port 130 nsew signal output
rlabel metal3 s 54165 36728 54965 36848 6 ss6[6]
port 131 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 ss6[7]
port 132 nsew signal output
rlabel metal2 s 41234 56309 41290 57109 6 ss7[0]
port 133 nsew signal output
rlabel metal2 s 39302 56309 39358 57109 6 ss7[1]
port 134 nsew signal output
rlabel metal2 s 662 56309 718 57109 6 ss7[2]
port 135 nsew signal output
rlabel metal2 s 9678 56309 9734 57109 6 ss7[3]
port 136 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 ss7[4]
port 137 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 ss7[5]
port 138 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 ss7[6]
port 139 nsew signal output
rlabel metal3 s 54165 27208 54965 27328 6 ss7[7]
port 140 nsew signal output
rlabel metal4 s 4208 2128 4528 54448 6 vccd1
port 141 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 54448 6 vccd1
port 141 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 54448 6 vssd1
port 142 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 54448 6 vssd1
port 142 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 54965 57109
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13456556
string GDS_FILE /home/designer-05/Caravel_STARS_2023/openlane/z23/runs/23_09_10_22_52/results/signoff/z23.magic.gds
string GDS_START 1306742
<< end >>

