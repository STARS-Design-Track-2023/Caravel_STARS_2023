magic
tech sky130A
magscale 1 2
timestamp 1691549598
<< viali >>
rect 6745 30345 6779 30379
rect 10241 30277 10275 30311
rect 22293 30277 22327 30311
rect 25697 30277 25731 30311
rect 1593 30209 1627 30243
rect 2789 30209 2823 30243
rect 6653 30209 6687 30243
rect 9873 30209 9907 30243
rect 14197 30209 14231 30243
rect 17601 30209 17635 30243
rect 21925 30209 21959 30243
rect 25329 30209 25363 30243
rect 28365 30209 28399 30243
rect 28733 30209 28767 30243
rect 29009 30141 29043 30175
rect 14381 30073 14415 30107
rect 17785 30073 17819 30107
rect 1409 30005 1443 30039
rect 2881 30005 2915 30039
rect 28549 30005 28583 30039
rect 23673 29801 23707 29835
rect 5549 29665 5583 29699
rect 16773 29665 16807 29699
rect 5089 29597 5123 29631
rect 5457 29597 5491 29631
rect 5641 29597 5675 29631
rect 5733 29597 5767 29631
rect 9045 29597 9079 29631
rect 11253 29597 11287 29631
rect 14749 29597 14783 29631
rect 16865 29597 16899 29631
rect 17509 29597 17543 29631
rect 20821 29597 20855 29631
rect 23857 29597 23891 29631
rect 7389 29529 7423 29563
rect 7573 29529 7607 29563
rect 9413 29529 9447 29563
rect 15117 29529 15151 29563
rect 4905 29461 4939 29495
rect 5273 29461 5307 29495
rect 7757 29461 7791 29495
rect 11805 29461 11839 29495
rect 17233 29461 17267 29495
rect 17325 29461 17359 29495
rect 20637 29461 20671 29495
rect 6653 29257 6687 29291
rect 13277 29257 13311 29291
rect 16497 29257 16531 29291
rect 19165 29257 19199 29291
rect 1685 29189 1719 29223
rect 7205 29189 7239 29223
rect 8953 29189 8987 29223
rect 11805 29189 11839 29223
rect 16957 29189 16991 29223
rect 20177 29189 20211 29223
rect 24041 29189 24075 29223
rect 6837 29121 6871 29155
rect 8773 29121 8807 29155
rect 9045 29121 9079 29155
rect 10701 29121 10735 29155
rect 11345 29121 11379 29155
rect 16221 29121 16255 29155
rect 16313 29121 16347 29155
rect 19901 29121 19935 29155
rect 22661 29121 22695 29155
rect 23121 29121 23155 29155
rect 23305 29121 23339 29155
rect 24409 29121 24443 29155
rect 1409 29053 1443 29087
rect 3249 29053 3283 29087
rect 3525 29053 3559 29087
rect 5089 29053 5123 29087
rect 6929 29053 6963 29087
rect 8677 29053 8711 29087
rect 10793 29053 10827 29087
rect 11529 29053 11563 29087
rect 13461 29053 13495 29087
rect 13737 29053 13771 29087
rect 15301 29053 15335 29087
rect 16681 29053 16715 29087
rect 18521 29053 18555 29087
rect 22569 29053 22603 29087
rect 23397 29053 23431 29087
rect 24685 29053 24719 29087
rect 3157 28985 3191 29019
rect 5733 28985 5767 29019
rect 11069 28985 11103 29019
rect 4997 28917 5031 28951
rect 8769 28917 8803 28951
rect 11161 28917 11195 28951
rect 15209 28917 15243 28951
rect 15945 28917 15979 28951
rect 18429 28917 18463 28951
rect 21649 28917 21683 28951
rect 23029 28917 23063 28951
rect 23121 28917 23155 28951
rect 6101 28713 6135 28747
rect 7389 28713 7423 28747
rect 7849 28713 7883 28747
rect 9781 28713 9815 28747
rect 10333 28713 10367 28747
rect 12449 28713 12483 28747
rect 12633 28713 12667 28747
rect 13461 28713 13495 28747
rect 14933 28713 14967 28747
rect 16129 28713 16163 28747
rect 16681 28713 16715 28747
rect 20361 28713 20395 28747
rect 20545 28713 20579 28747
rect 21741 28713 21775 28747
rect 22017 28713 22051 28747
rect 6745 28645 6779 28679
rect 7573 28645 7607 28679
rect 15853 28645 15887 28679
rect 18521 28645 18555 28679
rect 22201 28645 22235 28679
rect 24225 28645 24259 28679
rect 3341 28577 3375 28611
rect 8217 28577 8251 28611
rect 9137 28577 9171 28611
rect 10701 28577 10735 28611
rect 13645 28577 13679 28611
rect 15393 28577 15427 28611
rect 17049 28577 17083 28611
rect 19533 28577 19567 28611
rect 22753 28577 22787 28611
rect 24777 28577 24811 28611
rect 25237 28577 25271 28611
rect 3249 28509 3283 28543
rect 4353 28509 4387 28543
rect 6469 28509 6503 28543
rect 6561 28509 6595 28543
rect 6929 28509 6963 28543
rect 7113 28509 7147 28543
rect 10425 28509 10459 28543
rect 13185 28509 13219 28543
rect 13369 28509 13403 28543
rect 13737 28509 13771 28543
rect 14197 28509 14231 28543
rect 15117 28509 15151 28543
rect 15301 28509 15335 28543
rect 15485 28509 15519 28543
rect 15669 28509 15703 28543
rect 16037 28509 16071 28543
rect 16221 28509 16255 28543
rect 16497 28509 16531 28543
rect 16773 28509 16807 28543
rect 19257 28509 19291 28543
rect 19349 28509 19383 28543
rect 20821 28509 20855 28543
rect 20913 28509 20947 28543
rect 21005 28509 21039 28543
rect 21097 28509 21131 28543
rect 21373 28509 21407 28543
rect 21465 28509 21499 28543
rect 21833 28509 21867 28543
rect 22293 28509 22327 28543
rect 22385 28509 22419 28543
rect 22477 28509 22511 28543
rect 24501 28509 24535 28543
rect 12495 28475 12529 28509
rect 3893 28441 3927 28475
rect 4077 28441 4111 28475
rect 4629 28441 4663 28475
rect 6193 28441 6227 28475
rect 7205 28441 7239 28475
rect 7421 28441 7455 28475
rect 7665 28441 7699 28475
rect 7865 28441 7899 28475
rect 8769 28441 8803 28475
rect 9965 28441 9999 28475
rect 10149 28441 10183 28475
rect 12265 28441 12299 28475
rect 13461 28441 13495 28475
rect 16313 28441 16347 28475
rect 20177 28441 20211 28475
rect 20393 28441 20427 28475
rect 22109 28441 22143 28475
rect 3617 28373 3651 28407
rect 4261 28373 4295 28407
rect 6377 28373 6411 28407
rect 7021 28373 7055 28407
rect 8033 28373 8067 28407
rect 12173 28373 12207 28407
rect 13277 28373 13311 28407
rect 13921 28373 13955 28407
rect 14749 28373 14783 28407
rect 19533 28373 19567 28407
rect 20637 28373 20671 28407
rect 25881 28373 25915 28407
rect 3433 28169 3467 28203
rect 5457 28169 5491 28203
rect 6009 28169 6043 28203
rect 7297 28169 7331 28203
rect 9413 28169 9447 28203
rect 9873 28169 9907 28203
rect 10977 28169 11011 28203
rect 13369 28169 13403 28203
rect 17049 28169 17083 28203
rect 20729 28169 20763 28203
rect 24685 28169 24719 28203
rect 3985 28101 4019 28135
rect 11529 28101 11563 28135
rect 11713 28101 11747 28135
rect 11805 28101 11839 28135
rect 13001 28101 13035 28135
rect 13201 28101 13235 28135
rect 16681 28101 16715 28135
rect 23213 28101 23247 28135
rect 3617 28033 3651 28067
rect 6377 28033 6411 28067
rect 6653 28033 6687 28067
rect 6837 28033 6871 28067
rect 7113 28033 7147 28067
rect 7297 28033 7331 28067
rect 7665 28033 7699 28067
rect 9689 28033 9723 28067
rect 10425 28033 10459 28067
rect 10793 28033 10827 28067
rect 11069 28033 11103 28067
rect 11253 28033 11287 28067
rect 11897 28033 11931 28067
rect 13461 28033 13495 28067
rect 15945 28033 15979 28067
rect 16037 28033 16071 28067
rect 16221 28033 16255 28067
rect 16865 28033 16899 28067
rect 16957 28033 16991 28067
rect 17325 28033 17359 28067
rect 17785 28033 17819 28067
rect 18521 28033 18555 28067
rect 20821 28033 20855 28067
rect 22569 28033 22603 28067
rect 22937 28033 22971 28067
rect 3709 27965 3743 27999
rect 5549 27965 5583 27999
rect 7941 27965 7975 27999
rect 9505 27965 9539 27999
rect 10333 27965 10367 27999
rect 13737 27965 13771 27999
rect 15301 27965 15335 27999
rect 17601 27965 17635 27999
rect 18245 27965 18279 27999
rect 18337 27965 18371 27999
rect 18429 27965 18463 27999
rect 18981 27965 19015 27999
rect 19257 27965 19291 27999
rect 21833 27965 21867 27999
rect 22845 27965 22879 27999
rect 5825 27897 5859 27931
rect 16037 27897 16071 27931
rect 21465 27897 21499 27931
rect 22661 27897 22695 27931
rect 6469 27829 6503 27863
rect 7021 27829 7055 27863
rect 10793 27829 10827 27863
rect 11161 27829 11195 27863
rect 12081 27829 12115 27863
rect 13185 27829 13219 27863
rect 15209 27829 15243 27863
rect 17233 27829 17267 27863
rect 17785 27829 17819 27863
rect 17969 27829 18003 27863
rect 18061 27829 18095 27863
rect 22477 27829 22511 27863
rect 22569 27829 22603 27863
rect 14565 27625 14599 27659
rect 18245 27625 18279 27659
rect 19257 27625 19291 27659
rect 20164 27625 20198 27659
rect 4629 27557 4663 27591
rect 8125 27557 8159 27591
rect 12173 27557 12207 27591
rect 13921 27557 13955 27591
rect 14841 27557 14875 27591
rect 21741 27557 21775 27591
rect 2697 27489 2731 27523
rect 4261 27489 4295 27523
rect 4813 27489 4847 27523
rect 9321 27489 9355 27523
rect 9413 27489 9447 27523
rect 10241 27489 10275 27523
rect 11529 27489 11563 27523
rect 11713 27489 11747 27523
rect 11805 27489 11839 27523
rect 12725 27489 12759 27523
rect 13001 27489 13035 27523
rect 13277 27489 13311 27523
rect 14197 27489 14231 27523
rect 19901 27489 19935 27523
rect 22201 27489 22235 27523
rect 22753 27489 22787 27523
rect 4445 27421 4479 27455
rect 4721 27421 4755 27455
rect 4905 27421 4939 27455
rect 8493 27421 8527 27455
rect 9137 27421 9171 27455
rect 9689 27421 9723 27455
rect 10333 27421 10367 27455
rect 10517 27421 10551 27455
rect 11621 27421 11655 27455
rect 11989 27421 12023 27455
rect 12633 27421 12667 27455
rect 14289 27421 14323 27455
rect 14657 27421 14691 27455
rect 16405 27421 16439 27455
rect 16497 27421 16531 27455
rect 19533 27421 19567 27455
rect 21925 27421 21959 27455
rect 22017 27421 22051 27455
rect 22385 27421 22419 27455
rect 22661 27421 22695 27455
rect 22845 27421 22879 27455
rect 1501 27353 1535 27387
rect 7757 27353 7791 27387
rect 7941 27353 7975 27387
rect 10425 27353 10459 27387
rect 16773 27353 16807 27387
rect 19257 27353 19291 27387
rect 21741 27353 21775 27387
rect 1593 27285 1627 27319
rect 3341 27285 3375 27319
rect 8585 27285 8619 27319
rect 8953 27285 8987 27319
rect 11345 27285 11379 27319
rect 16221 27285 16255 27319
rect 19441 27285 19475 27319
rect 21649 27285 21683 27319
rect 22569 27285 22603 27319
rect 9689 27081 9723 27115
rect 14565 27081 14599 27115
rect 17601 27081 17635 27115
rect 21189 27081 21223 27115
rect 8217 27013 8251 27047
rect 14381 27013 14415 27047
rect 17141 27013 17175 27047
rect 20821 27013 20855 27047
rect 21021 27013 21055 27047
rect 11805 26945 11839 26979
rect 11897 26945 11931 26979
rect 12530 26945 12564 26979
rect 14657 26945 14691 26979
rect 28825 26945 28859 26979
rect 7941 26877 7975 26911
rect 11713 26877 11747 26911
rect 14289 26809 14323 26843
rect 14381 26809 14415 26843
rect 17509 26809 17543 26843
rect 11529 26741 11563 26775
rect 12804 26741 12838 26775
rect 21005 26741 21039 26775
rect 29009 26741 29043 26775
rect 2237 26537 2271 26571
rect 11056 26537 11090 26571
rect 12541 26537 12575 26571
rect 6837 26401 6871 26435
rect 10793 26401 10827 26435
rect 2421 26333 2455 26367
rect 5733 26333 5767 26367
rect 5917 26333 5951 26367
rect 6285 26333 6319 26367
rect 19625 26333 19659 26367
rect 19257 26265 19291 26299
rect 19441 26265 19475 26299
rect 5825 26197 5859 26231
rect 6193 25993 6227 26027
rect 19073 25925 19107 25959
rect 4997 25857 5031 25891
rect 5181 25857 5215 25891
rect 5273 25857 5307 25891
rect 5457 25857 5491 25891
rect 5733 25857 5767 25891
rect 6009 25857 6043 25891
rect 7113 25857 7147 25891
rect 7297 25857 7331 25891
rect 7389 25857 7423 25891
rect 8125 25857 8159 25891
rect 8217 25857 8251 25891
rect 8401 25857 8435 25891
rect 5917 25789 5951 25823
rect 6469 25789 6503 25823
rect 7573 25789 7607 25823
rect 18797 25789 18831 25823
rect 7113 25721 7147 25755
rect 8217 25721 8251 25755
rect 4997 25653 5031 25687
rect 5641 25653 5675 25687
rect 5733 25653 5767 25687
rect 7021 25653 7055 25687
rect 20545 25653 20579 25687
rect 3617 25449 3651 25483
rect 6745 25449 6779 25483
rect 6929 25449 6963 25483
rect 7284 25449 7318 25483
rect 8769 25449 8803 25483
rect 1869 25313 1903 25347
rect 4997 25313 5031 25347
rect 7021 25313 7055 25347
rect 15025 25313 15059 25347
rect 20361 25313 20395 25347
rect 20637 25313 20671 25347
rect 20913 25313 20947 25347
rect 4445 25245 4479 25279
rect 4629 25245 4663 25279
rect 4721 25245 4755 25279
rect 12081 25245 12115 25279
rect 18153 25245 18187 25279
rect 18613 25245 18647 25279
rect 18705 25245 18739 25279
rect 18797 25245 18831 25279
rect 18915 25245 18949 25279
rect 19073 25245 19107 25279
rect 19349 25245 19383 25279
rect 19533 25245 19567 25279
rect 2145 25177 2179 25211
rect 6561 25177 6595 25211
rect 15301 25177 15335 25211
rect 16957 25177 16991 25211
rect 17417 25177 17451 25211
rect 19625 25177 19659 25211
rect 22661 25177 22695 25211
rect 4629 25109 4663 25143
rect 6469 25109 6503 25143
rect 6771 25109 6805 25143
rect 11897 25109 11931 25143
rect 16773 25109 16807 25143
rect 17049 25109 17083 25143
rect 18429 25109 18463 25143
rect 19441 25109 19475 25143
rect 7389 24905 7423 24939
rect 14933 24905 14967 24939
rect 7113 24837 7147 24871
rect 7297 24837 7331 24871
rect 11805 24837 11839 24871
rect 14197 24837 14231 24871
rect 18061 24837 18095 24871
rect 18705 24837 18739 24871
rect 3157 24769 3191 24803
rect 5181 24769 5215 24803
rect 6377 24769 6411 24803
rect 7481 24769 7515 24803
rect 7665 24769 7699 24803
rect 9689 24769 9723 24803
rect 11529 24769 11563 24803
rect 15117 24769 15151 24803
rect 15209 24769 15243 24803
rect 15301 24769 15335 24803
rect 15419 24769 15453 24803
rect 15669 24769 15703 24803
rect 15853 24769 15887 24803
rect 16129 24769 16163 24803
rect 16313 24769 16347 24803
rect 16873 24769 16907 24803
rect 17877 24769 17911 24803
rect 17969 24769 18003 24803
rect 18179 24769 18213 24803
rect 20361 24769 20395 24803
rect 20821 24769 20855 24803
rect 3433 24701 3467 24735
rect 4905 24701 4939 24735
rect 4997 24701 5031 24735
rect 5549 24701 5583 24735
rect 7021 24701 7055 24735
rect 7849 24701 7883 24735
rect 8125 24701 8159 24735
rect 13553 24701 13587 24735
rect 14381 24701 14415 24735
rect 14473 24701 14507 24735
rect 14565 24701 14599 24735
rect 15577 24701 15611 24735
rect 18337 24701 18371 24735
rect 18429 24701 18463 24735
rect 20177 24701 20211 24735
rect 21005 24701 21039 24735
rect 6193 24633 6227 24667
rect 16037 24633 16071 24667
rect 17693 24633 17727 24667
rect 5365 24565 5399 24599
rect 9597 24565 9631 24599
rect 9781 24565 9815 24599
rect 10149 24565 10183 24599
rect 16221 24565 16255 24599
rect 16957 24565 16991 24599
rect 20453 24565 20487 24599
rect 4077 24361 4111 24395
rect 7021 24361 7055 24395
rect 16662 24361 16696 24395
rect 19257 24361 19291 24395
rect 19901 24361 19935 24395
rect 5273 24225 5307 24259
rect 11621 24225 11655 24259
rect 15301 24225 15335 24259
rect 16313 24225 16347 24259
rect 16405 24225 16439 24259
rect 4261 24157 4295 24191
rect 7113 24157 7147 24191
rect 7297 24157 7331 24191
rect 10057 24157 10091 24191
rect 15853 24157 15887 24191
rect 16175 24157 16209 24191
rect 19441 24157 19475 24191
rect 19717 24157 19751 24191
rect 19809 24157 19843 24191
rect 20085 24157 20119 24191
rect 5549 24089 5583 24123
rect 7205 24089 7239 24123
rect 11897 24089 11931 24123
rect 13645 24089 13679 24123
rect 14565 24089 14599 24123
rect 15945 24089 15979 24123
rect 16037 24089 16071 24123
rect 18429 24089 18463 24123
rect 19993 24089 20027 24123
rect 10609 24021 10643 24055
rect 15669 24021 15703 24055
rect 19625 24021 19659 24055
rect 13001 23817 13035 23851
rect 14749 23817 14783 23851
rect 17601 23817 17635 23851
rect 13369 23749 13403 23783
rect 15669 23749 15703 23783
rect 17509 23749 17543 23783
rect 1501 23681 1535 23715
rect 13461 23681 13495 23715
rect 14565 23681 14599 23715
rect 14841 23681 14875 23715
rect 15025 23681 15059 23715
rect 15301 23681 15335 23715
rect 15485 23681 15519 23715
rect 15577 23681 15611 23715
rect 17141 23681 17175 23715
rect 17233 23681 17267 23715
rect 17325 23681 17359 23715
rect 17785 23681 17819 23715
rect 9229 23613 9263 23647
rect 9505 23613 9539 23647
rect 11529 23613 11563 23647
rect 13645 23613 13679 23647
rect 14105 23613 14139 23647
rect 14473 23613 14507 23647
rect 15117 23613 15151 23647
rect 17877 23613 17911 23647
rect 17969 23613 18003 23647
rect 18061 23613 18095 23647
rect 15945 23545 15979 23579
rect 16957 23545 16991 23579
rect 1593 23477 1627 23511
rect 10977 23477 11011 23511
rect 12173 23477 12207 23511
rect 14841 23477 14875 23511
rect 16129 23477 16163 23511
rect 14657 23273 14691 23307
rect 15025 23273 15059 23307
rect 25237 23273 25271 23307
rect 10793 23205 10827 23239
rect 15209 23205 15243 23239
rect 15577 23205 15611 23239
rect 17601 23205 17635 23239
rect 6745 23137 6779 23171
rect 9045 23137 9079 23171
rect 11621 23137 11655 23171
rect 14841 23137 14875 23171
rect 16037 23137 16071 23171
rect 21005 23137 21039 23171
rect 4537 23069 4571 23103
rect 14105 23069 14139 23103
rect 14473 23069 14507 23103
rect 14749 23069 14783 23103
rect 15025 23069 15059 23103
rect 15301 23069 15335 23103
rect 15575 23047 15609 23081
rect 15761 23069 15795 23103
rect 15853 23069 15887 23103
rect 17601 23069 17635 23103
rect 17785 23069 17819 23103
rect 20729 23069 20763 23103
rect 20821 23069 20855 23103
rect 21097 23069 21131 23103
rect 24501 23069 24535 23103
rect 24593 23069 24627 23103
rect 24777 23069 24811 23103
rect 24869 23069 24903 23103
rect 6009 23001 6043 23035
rect 9321 23001 9355 23035
rect 10885 23001 10919 23035
rect 14381 23001 14415 23035
rect 15485 23001 15519 23035
rect 21189 23001 21223 23035
rect 25053 23001 25087 23035
rect 5089 22933 5123 22967
rect 14289 22933 14323 22967
rect 21005 22933 21039 22967
rect 9229 22729 9263 22763
rect 12817 22729 12851 22763
rect 20913 22729 20947 22763
rect 24409 22729 24443 22763
rect 25421 22729 25455 22763
rect 5273 22661 5307 22695
rect 8217 22661 8251 22695
rect 8953 22661 8987 22695
rect 12449 22661 12483 22695
rect 12541 22661 12575 22695
rect 15393 22661 15427 22695
rect 6745 22593 6779 22627
rect 6929 22593 6963 22627
rect 7021 22593 7055 22627
rect 7113 22593 7147 22627
rect 8677 22593 8711 22627
rect 8861 22593 8895 22627
rect 9045 22593 9079 22627
rect 9321 22593 9355 22627
rect 12265 22593 12299 22627
rect 12633 22593 12667 22627
rect 15025 22593 15059 22627
rect 15301 22593 15335 22627
rect 17325 22593 17359 22627
rect 20729 22593 20763 22627
rect 21281 22593 21315 22627
rect 21465 22593 21499 22627
rect 21557 22593 21591 22627
rect 21833 22593 21867 22627
rect 22017 22593 22051 22627
rect 22753 22593 22787 22627
rect 22937 22593 22971 22627
rect 23121 22593 23155 22627
rect 23305 22593 23339 22627
rect 23673 22593 23707 22627
rect 23765 22593 23799 22627
rect 23908 22593 23942 22627
rect 24041 22593 24075 22627
rect 24133 22593 24167 22627
rect 24317 22593 24351 22627
rect 24580 22593 24614 22627
rect 24685 22593 24719 22627
rect 24777 22593 24811 22627
rect 24869 22593 24903 22627
rect 25053 22593 25087 22627
rect 25237 22593 25271 22627
rect 28825 22593 28859 22627
rect 4537 22525 4571 22559
rect 6009 22525 6043 22559
rect 7665 22525 7699 22559
rect 9597 22525 9631 22559
rect 11069 22525 11103 22559
rect 11529 22525 11563 22559
rect 15209 22525 15243 22559
rect 16221 22525 16255 22559
rect 16681 22525 16715 22559
rect 20545 22525 20579 22559
rect 21373 22525 21407 22559
rect 24225 22525 24259 22559
rect 29009 22457 29043 22491
rect 5089 22389 5123 22423
rect 7297 22389 7331 22423
rect 12173 22389 12207 22423
rect 14841 22389 14875 22423
rect 21097 22389 21131 22423
rect 21833 22389 21867 22423
rect 22753 22389 22787 22423
rect 23213 22389 23247 22423
rect 23489 22389 23523 22423
rect 6272 22185 6306 22219
rect 7757 22185 7791 22219
rect 14736 22185 14770 22219
rect 21649 22185 21683 22219
rect 22109 22185 22143 22219
rect 23765 22185 23799 22219
rect 22477 22117 22511 22151
rect 6009 22049 6043 22083
rect 10333 22049 10367 22083
rect 14473 22049 14507 22083
rect 22569 22049 22603 22083
rect 23009 22049 23043 22083
rect 23305 22049 23339 22083
rect 24777 22049 24811 22083
rect 4169 21981 4203 22015
rect 4445 21981 4479 22015
rect 5365 21981 5399 22015
rect 7849 21981 7883 22015
rect 9045 21981 9079 22015
rect 9413 21981 9447 22015
rect 9689 21981 9723 22015
rect 10425 21981 10459 22015
rect 10518 21981 10552 22015
rect 10793 21981 10827 22015
rect 10931 21981 10965 22015
rect 17325 21981 17359 22015
rect 20085 21981 20119 22015
rect 20177 21981 20211 22015
rect 20269 21981 20303 22015
rect 20545 21981 20579 22015
rect 20821 21981 20855 22015
rect 21097 21981 21131 22015
rect 21281 21981 21315 22015
rect 21373 21981 21407 22015
rect 21465 21981 21499 22015
rect 21741 21981 21775 22015
rect 21925 21981 21959 22015
rect 22385 21981 22419 22015
rect 22661 21981 22695 22015
rect 22845 21981 22879 22015
rect 23213 21981 23247 22015
rect 23489 21981 23523 22015
rect 23857 21981 23891 22015
rect 23949 21981 23983 22015
rect 24133 21981 24167 22015
rect 24225 21981 24259 22015
rect 24409 21981 24443 22015
rect 24593 21981 24627 22015
rect 24869 21981 24903 22015
rect 25145 21981 25179 22015
rect 25421 21981 25455 22015
rect 25697 21981 25731 22015
rect 25973 21981 26007 22015
rect 9229 21913 9263 21947
rect 9321 21913 9355 21947
rect 10701 21913 10735 21947
rect 22937 21913 22971 21947
rect 25329 21913 25363 21947
rect 25881 21913 25915 21947
rect 4077 21845 4111 21879
rect 5917 21845 5951 21879
rect 8493 21845 8527 21879
rect 9597 21845 9631 21879
rect 11069 21845 11103 21879
rect 16221 21845 16255 21879
rect 17877 21845 17911 21879
rect 20361 21845 20395 21879
rect 20729 21845 20763 21879
rect 22201 21845 22235 21879
rect 23121 21845 23155 21879
rect 24047 21845 24081 21879
rect 24961 21845 24995 21879
rect 25513 21845 25547 21879
rect 5549 21641 5583 21675
rect 6193 21641 6227 21675
rect 18429 21641 18463 21675
rect 20177 21641 20211 21675
rect 20821 21641 20855 21675
rect 21557 21641 21591 21675
rect 23397 21641 23431 21675
rect 23673 21641 23707 21675
rect 3341 21573 3375 21607
rect 3433 21573 3467 21607
rect 8401 21573 8435 21607
rect 8493 21573 8527 21607
rect 12449 21573 12483 21607
rect 3157 21505 3191 21539
rect 3525 21505 3559 21539
rect 5641 21505 5675 21539
rect 5825 21505 5859 21539
rect 5917 21505 5951 21539
rect 6009 21505 6043 21539
rect 6377 21505 6411 21539
rect 8217 21505 8251 21539
rect 8585 21505 8619 21539
rect 9045 21505 9079 21539
rect 12081 21505 12115 21539
rect 12174 21505 12208 21539
rect 12357 21505 12391 21539
rect 12587 21505 12621 21539
rect 12909 21505 12943 21539
rect 18797 21505 18831 21539
rect 19165 21505 19199 21539
rect 19349 21505 19383 21539
rect 21097 21505 21131 21539
rect 21465 21505 21499 21539
rect 21833 21505 21867 21539
rect 22017 21505 22051 21539
rect 22109 21505 22143 21539
rect 22385 21505 22419 21539
rect 22477 21505 22511 21539
rect 22845 21505 22879 21539
rect 23857 21505 23891 21539
rect 24317 21505 24351 21539
rect 24685 21505 24719 21539
rect 24961 21505 24995 21539
rect 25329 21505 25363 21539
rect 25513 21505 25547 21539
rect 26985 21505 27019 21539
rect 27169 21505 27203 21539
rect 27537 21505 27571 21539
rect 27721 21505 27755 21539
rect 3801 21437 3835 21471
rect 4077 21437 4111 21471
rect 6653 21437 6687 21471
rect 9321 21437 9355 21471
rect 13185 21437 13219 21471
rect 16681 21437 16715 21471
rect 16957 21437 16991 21471
rect 18705 21437 18739 21471
rect 18889 21437 18923 21471
rect 18981 21437 19015 21471
rect 20545 21437 20579 21471
rect 20637 21437 20671 21471
rect 21281 21437 21315 21471
rect 21373 21437 21407 21471
rect 22201 21437 22235 21471
rect 22569 21437 22603 21471
rect 22661 21437 22695 21471
rect 22937 21437 22971 21471
rect 23489 21437 23523 21471
rect 8769 21369 8803 21403
rect 18521 21369 18555 21403
rect 20913 21369 20947 21403
rect 21833 21369 21867 21403
rect 23213 21369 23247 21403
rect 24409 21369 24443 21403
rect 27077 21369 27111 21403
rect 3709 21301 3743 21335
rect 8125 21301 8159 21335
rect 10793 21301 10827 21335
rect 12725 21301 12759 21335
rect 14657 21301 14691 21335
rect 19533 21301 19567 21335
rect 23949 21301 23983 21335
rect 25329 21301 25363 21335
rect 27629 21301 27663 21335
rect 4058 21097 4092 21131
rect 5549 21097 5583 21131
rect 14749 21097 14783 21131
rect 16497 21097 16531 21131
rect 23489 21097 23523 21131
rect 25881 21097 25915 21131
rect 27077 21097 27111 21131
rect 27813 21097 27847 21131
rect 21557 21029 21591 21063
rect 23305 21029 23339 21063
rect 3801 20961 3835 20995
rect 9597 20961 9631 20995
rect 12173 20961 12207 20995
rect 12449 20961 12483 20995
rect 18337 20961 18371 20995
rect 18521 20961 18555 20995
rect 20361 20961 20395 20995
rect 23949 20961 23983 20995
rect 25237 20961 25271 20995
rect 26709 20961 26743 20995
rect 27629 20961 27663 20995
rect 6009 20893 6043 20927
rect 6102 20893 6136 20927
rect 6515 20893 6549 20927
rect 7297 20893 7331 20927
rect 7390 20893 7424 20927
rect 7762 20893 7796 20927
rect 10425 20893 10459 20927
rect 11437 20893 11471 20927
rect 11530 20893 11564 20927
rect 11713 20893 11747 20927
rect 11902 20893 11936 20927
rect 14105 20893 14139 20927
rect 14198 20893 14232 20927
rect 14570 20893 14604 20927
rect 14841 20893 14875 20927
rect 15945 20893 15979 20927
rect 16313 20893 16347 20927
rect 16589 20893 16623 20927
rect 19441 20893 19475 20927
rect 19809 20893 19843 20927
rect 19993 20893 20027 20927
rect 20637 20893 20671 20927
rect 20913 20893 20947 20927
rect 21097 20893 21131 20927
rect 21281 20893 21315 20927
rect 21465 20893 21499 20927
rect 22201 20893 22235 20927
rect 22293 20893 22327 20927
rect 22661 20893 22695 20927
rect 23029 20893 23063 20927
rect 23673 20893 23707 20927
rect 23857 20893 23891 20927
rect 24961 20893 24995 20927
rect 26157 20893 26191 20927
rect 26801 20893 26835 20927
rect 27353 20893 27387 20927
rect 27445 20893 27479 20927
rect 27721 20893 27755 20927
rect 28457 20893 28491 20927
rect 6285 20825 6319 20859
rect 6377 20825 6411 20859
rect 7573 20825 7607 20859
rect 7665 20825 7699 20859
rect 11161 20825 11195 20859
rect 11805 20825 11839 20859
rect 14381 20825 14415 20859
rect 14473 20825 14507 20859
rect 16129 20825 16163 20859
rect 16221 20825 16255 20859
rect 16865 20825 16899 20859
rect 21189 20825 21223 20859
rect 25881 20825 25915 20859
rect 28273 20825 28307 20859
rect 6653 20757 6687 20791
rect 7941 20757 7975 20791
rect 10149 20757 10183 20791
rect 12081 20757 12115 20791
rect 13921 20757 13955 20791
rect 15485 20757 15519 20791
rect 19073 20757 19107 20791
rect 25789 20757 25823 20791
rect 26065 20757 26099 20791
rect 28181 20757 28215 20791
rect 28641 20757 28675 20791
rect 10885 20553 10919 20587
rect 14933 20553 14967 20587
rect 16957 20553 16991 20587
rect 21373 20553 21407 20587
rect 22033 20553 22067 20587
rect 22201 20553 22235 20587
rect 23121 20553 23155 20587
rect 23489 20553 23523 20587
rect 3525 20485 3559 20519
rect 3617 20485 3651 20519
rect 9965 20485 9999 20519
rect 17067 20485 17101 20519
rect 17969 20485 18003 20519
rect 21005 20485 21039 20519
rect 21833 20485 21867 20519
rect 3341 20417 3375 20451
rect 3709 20417 3743 20451
rect 4261 20417 4295 20451
rect 4445 20417 4479 20451
rect 9689 20417 9723 20451
rect 9873 20417 9907 20451
rect 10057 20417 10091 20451
rect 10333 20417 10367 20451
rect 10517 20417 10551 20451
rect 10609 20417 10643 20451
rect 10701 20417 10735 20451
rect 11805 20417 11839 20451
rect 13737 20417 13771 20451
rect 14381 20417 14415 20451
rect 14565 20417 14599 20451
rect 14657 20417 14691 20451
rect 14749 20417 14783 20451
rect 16865 20417 16899 20451
rect 17233 20417 17267 20451
rect 17325 20417 17359 20451
rect 17509 20417 17543 20451
rect 17601 20417 17635 20451
rect 17693 20417 17727 20451
rect 18153 20417 18187 20451
rect 18337 20417 18371 20451
rect 18797 20417 18831 20451
rect 19165 20417 19199 20451
rect 19441 20417 19475 20451
rect 21189 20417 21223 20451
rect 21465 20417 21499 20451
rect 21649 20417 21683 20451
rect 22753 20417 22787 20451
rect 22937 20417 22971 20451
rect 23673 20417 23707 20451
rect 23857 20417 23891 20451
rect 23949 20417 23983 20451
rect 24041 20417 24075 20451
rect 24133 20417 24167 20451
rect 26617 20417 26651 20451
rect 27077 20417 27111 20451
rect 27445 20417 27479 20451
rect 27905 20417 27939 20451
rect 27997 20417 28031 20451
rect 28181 20417 28215 20451
rect 28273 20417 28307 20451
rect 28552 20439 28586 20473
rect 28641 20417 28675 20451
rect 28825 20417 28859 20451
rect 28917 20417 28951 20451
rect 4721 20349 4755 20383
rect 6377 20349 6411 20383
rect 6653 20349 6687 20383
rect 8217 20349 8251 20383
rect 12081 20349 12115 20383
rect 13553 20349 13587 20383
rect 18429 20349 18463 20383
rect 24317 20349 24351 20383
rect 26709 20349 26743 20383
rect 10241 20281 10275 20315
rect 16681 20281 16715 20315
rect 18889 20281 18923 20315
rect 24225 20281 24259 20315
rect 3893 20213 3927 20247
rect 8125 20213 8159 20247
rect 8861 20213 8895 20247
rect 14289 20213 14323 20247
rect 17877 20213 17911 20247
rect 21557 20213 21591 20247
rect 22017 20213 22051 20247
rect 27353 20213 27387 20247
rect 27629 20213 27663 20247
rect 27721 20213 27755 20247
rect 28365 20213 28399 20247
rect 4445 20009 4479 20043
rect 6929 20009 6963 20043
rect 8769 20009 8803 20043
rect 12633 20009 12667 20043
rect 16129 20009 16163 20043
rect 27629 20009 27663 20043
rect 2145 19873 2179 19907
rect 10517 19873 10551 19907
rect 1869 19805 1903 19839
rect 3893 19805 3927 19839
rect 6377 19805 6411 19839
rect 6653 19805 6687 19839
rect 6745 19805 6779 19839
rect 7021 19805 7055 19839
rect 7169 19805 7203 19839
rect 7527 19805 7561 19839
rect 8217 19805 8251 19839
rect 8953 19805 8987 19839
rect 10241 19805 10275 19839
rect 10609 19805 10643 19839
rect 10793 19805 10827 19839
rect 10977 19805 11011 19839
rect 12081 19805 12115 19839
rect 12449 19805 12483 19839
rect 13001 19805 13035 19839
rect 15945 19805 15979 19839
rect 27261 19805 27295 19839
rect 27537 19805 27571 19839
rect 27629 19805 27663 19839
rect 27813 19805 27847 19839
rect 28089 19805 28123 19839
rect 28365 19805 28399 19839
rect 6561 19737 6595 19771
rect 7297 19737 7331 19771
rect 7389 19737 7423 19771
rect 10885 19737 10919 19771
rect 12265 19737 12299 19771
rect 12357 19737 12391 19771
rect 15761 19737 15795 19771
rect 28273 19737 28307 19771
rect 3617 19669 3651 19703
rect 7665 19669 7699 19703
rect 9597 19669 9631 19703
rect 11161 19669 11195 19703
rect 13553 19669 13587 19703
rect 27077 19669 27111 19703
rect 27445 19669 27479 19703
rect 27905 19669 27939 19703
rect 1593 19465 1627 19499
rect 12173 19465 12207 19499
rect 13369 19465 13403 19499
rect 17233 19465 17267 19499
rect 18981 19465 19015 19499
rect 19073 19465 19107 19499
rect 20545 19465 20579 19499
rect 7573 19397 7607 19431
rect 8217 19397 8251 19431
rect 15117 19397 15151 19431
rect 15209 19397 15243 19431
rect 16957 19397 16991 19431
rect 19257 19397 19291 19431
rect 19533 19397 19567 19431
rect 19625 19397 19659 19431
rect 20177 19397 20211 19431
rect 20269 19397 20303 19431
rect 1501 19329 1535 19363
rect 7297 19329 7331 19363
rect 7481 19329 7515 19363
rect 7665 19329 7699 19363
rect 7941 19329 7975 19363
rect 12817 19329 12851 19363
rect 13001 19329 13035 19363
rect 13093 19329 13127 19363
rect 13185 19329 13219 19363
rect 14933 19329 14967 19363
rect 15301 19329 15335 19363
rect 16681 19329 16715 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 18889 19329 18923 19363
rect 19349 19329 19383 19363
rect 19717 19329 19751 19363
rect 19993 19329 20027 19363
rect 20361 19329 20395 19363
rect 27537 19329 27571 19363
rect 27629 19329 27663 19363
rect 9689 19261 9723 19295
rect 11621 19261 11655 19295
rect 15853 19261 15887 19295
rect 27813 19261 27847 19295
rect 16405 19193 16439 19227
rect 18705 19193 18739 19227
rect 19901 19193 19935 19227
rect 7849 19125 7883 19159
rect 15485 19125 15519 19159
rect 8769 18921 8803 18955
rect 9597 18921 9631 18955
rect 11897 18921 11931 18955
rect 15945 18921 15979 18955
rect 19809 18921 19843 18955
rect 20269 18921 20303 18955
rect 7021 18785 7055 18819
rect 7297 18785 7331 18819
rect 10149 18785 10183 18819
rect 10425 18785 10459 18819
rect 14473 18785 14507 18819
rect 19073 18785 19107 18819
rect 4077 18717 4111 18751
rect 6193 18717 6227 18751
rect 6469 18717 6503 18751
rect 6561 18717 6595 18751
rect 8953 18717 8987 18751
rect 9046 18717 9080 18751
rect 9321 18717 9355 18751
rect 9418 18717 9452 18751
rect 12265 18717 12299 18751
rect 12449 18717 12483 18751
rect 12633 18717 12667 18751
rect 14197 18717 14231 18751
rect 16037 18717 16071 18751
rect 16589 18717 16623 18751
rect 17417 18717 17451 18751
rect 17693 18717 17727 18751
rect 17785 18717 17819 18751
rect 18521 18717 18555 18751
rect 19257 18717 19291 18751
rect 19441 18717 19475 18751
rect 19625 18717 19659 18751
rect 19901 18717 19935 18751
rect 28825 18717 28859 18751
rect 6377 18649 6411 18683
rect 9229 18649 9263 18683
rect 12541 18649 12575 18683
rect 17601 18649 17635 18683
rect 19533 18649 19567 18683
rect 20085 18649 20119 18683
rect 4721 18581 4755 18615
rect 6745 18581 6779 18615
rect 12817 18581 12851 18615
rect 16129 18581 16163 18615
rect 17969 18581 18003 18615
rect 29009 18581 29043 18615
rect 8217 18377 8251 18411
rect 11345 18377 11379 18411
rect 14013 18377 14047 18411
rect 18797 18377 18831 18411
rect 21005 18377 21039 18411
rect 5917 18309 5951 18343
rect 12173 18309 12207 18343
rect 13001 18309 13035 18343
rect 17325 18309 17359 18343
rect 20637 18309 20671 18343
rect 1869 18241 1903 18275
rect 3709 18241 3743 18275
rect 5641 18241 5675 18275
rect 5825 18241 5859 18275
rect 6009 18241 6043 18275
rect 6837 18241 6871 18275
rect 7297 18241 7331 18275
rect 9413 18241 9447 18275
rect 9597 18241 9631 18275
rect 9689 18241 9723 18275
rect 9781 18241 9815 18275
rect 10057 18241 10091 18275
rect 10241 18241 10275 18275
rect 10333 18241 10367 18275
rect 10425 18241 10459 18275
rect 12633 18241 12667 18275
rect 12781 18241 12815 18275
rect 12909 18241 12943 18275
rect 13139 18241 13173 18275
rect 14749 18241 14783 18275
rect 17049 18241 17083 18275
rect 19349 18241 19383 18275
rect 19441 18241 19475 18275
rect 19809 18241 19843 18275
rect 20361 18241 20395 18275
rect 20454 18241 20488 18275
rect 20729 18241 20763 18275
rect 20826 18241 20860 18275
rect 22937 18241 22971 18275
rect 2145 18173 2179 18207
rect 3985 18173 4019 18207
rect 7481 18173 7515 18207
rect 7665 18173 7699 18207
rect 10793 18173 10827 18207
rect 11529 18173 11563 18207
rect 13461 18173 13495 18207
rect 15025 18173 15059 18207
rect 19257 18173 19291 18207
rect 23213 18173 23247 18207
rect 24961 18173 24995 18207
rect 25053 18173 25087 18207
rect 26985 18173 27019 18207
rect 27261 18173 27295 18207
rect 29009 18173 29043 18207
rect 20269 18105 20303 18139
rect 3617 18037 3651 18071
rect 5457 18037 5491 18071
rect 6193 18037 6227 18071
rect 9965 18037 9999 18071
rect 10609 18037 10643 18071
rect 13277 18037 13311 18071
rect 16497 18037 16531 18071
rect 25697 18037 25731 18071
rect 12081 17833 12115 17867
rect 13921 17833 13955 17867
rect 15669 17833 15703 17867
rect 19809 17833 19843 17867
rect 23305 17833 23339 17867
rect 27169 17833 27203 17867
rect 11345 17765 11379 17799
rect 22385 17765 22419 17799
rect 22937 17765 22971 17799
rect 25053 17765 25087 17799
rect 25881 17765 25915 17799
rect 27997 17765 28031 17799
rect 5273 17697 5307 17731
rect 7021 17697 7055 17731
rect 9597 17697 9631 17731
rect 12173 17697 12207 17731
rect 17325 17697 17359 17731
rect 20085 17697 20119 17731
rect 20361 17697 20395 17731
rect 21833 17697 21867 17731
rect 23029 17697 23063 17731
rect 23949 17697 23983 17731
rect 25789 17697 25823 17731
rect 26065 17697 26099 17731
rect 26157 17697 26191 17731
rect 26525 17697 26559 17731
rect 4445 17629 4479 17663
rect 7297 17629 7331 17663
rect 7389 17629 7423 17663
rect 7573 17629 7607 17663
rect 7665 17629 7699 17663
rect 11437 17629 11471 17663
rect 11530 17629 11564 17663
rect 11805 17629 11839 17663
rect 11902 17629 11936 17663
rect 16129 17629 16163 17663
rect 19257 17629 19291 17663
rect 19441 17629 19475 17663
rect 19533 17629 19567 17663
rect 19625 17629 19659 17663
rect 22293 17629 22327 17663
rect 22753 17629 22787 17663
rect 23489 17629 23523 17663
rect 24409 17629 24443 17663
rect 25330 17607 25364 17641
rect 25513 17629 25547 17663
rect 25651 17629 25685 17663
rect 26617 17629 26651 17663
rect 26893 17629 26927 17663
rect 26985 17629 27019 17663
rect 27629 17629 27663 17663
rect 27905 17629 27939 17663
rect 28181 17629 28215 17663
rect 28365 17629 28399 17663
rect 5549 17561 5583 17595
rect 7113 17561 7147 17595
rect 9873 17561 9907 17595
rect 11713 17561 11747 17595
rect 12449 17561 12483 17595
rect 14197 17561 14231 17595
rect 17601 17561 17635 17595
rect 23581 17561 23615 17595
rect 23673 17561 23707 17595
rect 23811 17561 23845 17595
rect 25421 17561 25455 17595
rect 26801 17561 26835 17595
rect 27445 17561 27479 17595
rect 4997 17493 5031 17527
rect 16681 17493 16715 17527
rect 19073 17493 19107 17527
rect 22569 17493 22603 17527
rect 25145 17493 25179 17527
rect 26249 17493 26283 17527
rect 26433 17493 26467 17527
rect 27813 17493 27847 17527
rect 28273 17493 28307 17527
rect 4537 17289 4571 17323
rect 5181 17289 5215 17323
rect 13921 17289 13955 17323
rect 18797 17289 18831 17323
rect 19257 17289 19291 17323
rect 20821 17289 20855 17323
rect 21833 17289 21867 17323
rect 23397 17289 23431 17323
rect 25881 17289 25915 17323
rect 26801 17289 26835 17323
rect 3525 17221 3559 17255
rect 4261 17221 4295 17255
rect 4813 17221 4847 17255
rect 5457 17221 5491 17255
rect 12449 17221 12483 17255
rect 15209 17221 15243 17255
rect 18889 17221 18923 17255
rect 22293 17221 22327 17255
rect 23765 17221 23799 17255
rect 26249 17221 26283 17255
rect 28273 17221 28307 17255
rect 3341 17153 3375 17187
rect 3617 17153 3651 17187
rect 3709 17153 3743 17187
rect 3985 17153 4019 17187
rect 4169 17153 4203 17187
rect 4353 17153 4387 17187
rect 4629 17153 4663 17187
rect 4905 17153 4939 17187
rect 4997 17153 5031 17187
rect 5273 17153 5307 17187
rect 5545 17153 5579 17187
rect 5641 17153 5675 17187
rect 9597 17153 9631 17187
rect 12173 17153 12207 17187
rect 14013 17153 14047 17187
rect 15025 17153 15059 17187
rect 15301 17153 15335 17187
rect 15393 17153 15427 17187
rect 16957 17153 16991 17187
rect 17049 17153 17083 17187
rect 17141 17153 17175 17187
rect 17325 17153 17359 17187
rect 17601 17153 17635 17187
rect 18153 17153 18187 17187
rect 18245 17153 18279 17187
rect 18429 17153 18463 17187
rect 18521 17153 18555 17187
rect 18613 17153 18647 17187
rect 19073 17153 19107 17187
rect 21005 17153 21039 17187
rect 21281 17153 21315 17187
rect 22201 17153 22235 17187
rect 22845 17153 22879 17187
rect 25421 17153 25455 17187
rect 25605 17153 25639 17187
rect 26065 17153 26099 17187
rect 26341 17153 26375 17187
rect 26433 17153 26467 17187
rect 26617 17153 26651 17187
rect 27169 17153 27203 17187
rect 27629 17153 27663 17187
rect 27905 17153 27939 17187
rect 28457 17153 28491 17187
rect 9873 17085 9907 17119
rect 16681 17085 16715 17119
rect 21373 17085 21407 17119
rect 22477 17085 22511 17119
rect 23121 17085 23155 17119
rect 23489 17085 23523 17119
rect 27261 17085 27295 17119
rect 27353 17085 27387 17119
rect 27445 17085 27479 17119
rect 28181 17085 28215 17119
rect 11345 17017 11379 17051
rect 15577 17017 15611 17051
rect 21649 17017 21683 17051
rect 25789 17017 25823 17051
rect 26985 17017 27019 17051
rect 27721 17017 27755 17051
rect 3893 16949 3927 16983
rect 5825 16949 5859 16983
rect 14657 16949 14691 16983
rect 23121 16949 23155 16983
rect 25237 16949 25271 16983
rect 26433 16949 26467 16983
rect 28089 16949 28123 16983
rect 28641 16949 28675 16983
rect 6285 16745 6319 16779
rect 14657 16745 14691 16779
rect 22017 16745 22051 16779
rect 22385 16745 22419 16779
rect 22753 16745 22787 16779
rect 23121 16745 23155 16779
rect 23765 16745 23799 16779
rect 24409 16745 24443 16779
rect 27813 16745 27847 16779
rect 23305 16677 23339 16711
rect 23673 16677 23707 16711
rect 3157 16609 3191 16643
rect 3801 16609 3835 16643
rect 10701 16609 10735 16643
rect 22845 16609 22879 16643
rect 23857 16609 23891 16643
rect 26157 16609 26191 16643
rect 1409 16541 1443 16575
rect 4997 16541 5031 16575
rect 5181 16541 5215 16575
rect 5365 16541 5399 16575
rect 5733 16541 5767 16575
rect 9873 16541 9907 16575
rect 10241 16541 10275 16575
rect 14105 16541 14139 16575
rect 14289 16541 14323 16575
rect 14473 16541 14507 16575
rect 15117 16541 15151 16575
rect 15209 16541 15243 16575
rect 15301 16541 15335 16575
rect 15485 16541 15519 16575
rect 22201 16541 22235 16575
rect 22477 16541 22511 16575
rect 22753 16541 22787 16575
rect 23213 16541 23247 16575
rect 23489 16541 23523 16575
rect 23581 16541 23615 16575
rect 24593 16541 24627 16575
rect 24869 16541 24903 16575
rect 24961 16541 24995 16575
rect 25513 16541 25547 16575
rect 25697 16541 25731 16575
rect 26341 16541 26375 16575
rect 26525 16541 26559 16575
rect 26617 16541 26651 16575
rect 26893 16541 26927 16575
rect 27445 16541 27479 16575
rect 27629 16541 27663 16575
rect 27721 16541 27755 16575
rect 28089 16541 28123 16575
rect 28181 16541 28215 16575
rect 28373 16541 28407 16575
rect 1685 16473 1719 16507
rect 5265 16473 5299 16507
rect 10057 16473 10091 16507
rect 10149 16473 10183 16507
rect 11253 16473 11287 16507
rect 14381 16473 14415 16507
rect 25053 16473 25087 16507
rect 25605 16473 25639 16507
rect 26709 16473 26743 16507
rect 27813 16473 27847 16507
rect 28273 16473 28307 16507
rect 4445 16405 4479 16439
rect 5549 16405 5583 16439
rect 10425 16405 10459 16439
rect 14841 16405 14875 16439
rect 23213 16405 23247 16439
rect 24777 16405 24811 16439
rect 27077 16405 27111 16439
rect 27261 16405 27295 16439
rect 27997 16405 28031 16439
rect 1409 16201 1443 16235
rect 4997 16201 5031 16235
rect 6193 16201 6227 16235
rect 2789 16133 2823 16167
rect 9321 16133 9355 16167
rect 10057 16133 10091 16167
rect 10149 16133 10183 16167
rect 12173 16133 12207 16167
rect 13277 16133 13311 16167
rect 16037 16133 16071 16167
rect 23305 16133 23339 16167
rect 1593 16065 1627 16099
rect 6377 16065 6411 16099
rect 6470 16065 6504 16099
rect 6653 16065 6687 16099
rect 6745 16065 6779 16099
rect 6883 16065 6917 16099
rect 7113 16065 7147 16099
rect 7297 16065 7331 16099
rect 7389 16065 7423 16099
rect 7481 16065 7515 16099
rect 7941 16065 7975 16099
rect 8309 16065 8343 16099
rect 9873 16065 9907 16099
rect 10241 16065 10275 16099
rect 13001 16065 13035 16099
rect 13185 16065 13219 16099
rect 13369 16065 13403 16099
rect 15669 16065 15703 16099
rect 15761 16065 15795 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 23489 16065 23523 16099
rect 25697 16065 25731 16099
rect 25881 16065 25915 16099
rect 2513 15997 2547 16031
rect 4445 15997 4479 16031
rect 5641 15997 5675 16031
rect 8677 15997 8711 16031
rect 10517 15997 10551 16031
rect 11529 15997 11563 16031
rect 15117 15997 15151 16031
rect 7021 15929 7055 15963
rect 23673 15929 23707 15963
rect 4261 15861 4295 15895
rect 7665 15861 7699 15895
rect 10425 15861 10459 15895
rect 11161 15861 11195 15895
rect 13553 15861 13587 15895
rect 16313 15861 16347 15895
rect 25789 15861 25823 15895
rect 3617 15657 3651 15691
rect 6009 15657 6043 15691
rect 8401 15657 8435 15691
rect 9492 15657 9526 15691
rect 10977 15657 11011 15691
rect 16129 15657 16163 15691
rect 23581 15657 23615 15691
rect 26249 15657 26283 15691
rect 26985 15657 27019 15691
rect 18797 15589 18831 15623
rect 23213 15589 23247 15623
rect 26525 15589 26559 15623
rect 1869 15521 1903 15555
rect 2145 15521 2179 15555
rect 4537 15521 4571 15555
rect 6929 15521 6963 15555
rect 13185 15521 13219 15555
rect 14381 15521 14415 15555
rect 14657 15521 14691 15555
rect 16497 15521 16531 15555
rect 18705 15521 18739 15555
rect 23765 15521 23799 15555
rect 24041 15521 24075 15555
rect 27172 15521 27206 15555
rect 4261 15453 4295 15487
rect 6653 15453 6687 15487
rect 9229 15453 9263 15487
rect 11897 15453 11931 15487
rect 12081 15453 12115 15487
rect 12265 15453 12299 15487
rect 12633 15453 12667 15487
rect 13369 15453 13403 15487
rect 18429 15453 18463 15487
rect 19625 15453 19659 15487
rect 19717 15453 19751 15487
rect 19809 15453 19843 15487
rect 19901 15453 19935 15487
rect 19993 15453 20027 15487
rect 20177 15453 20211 15487
rect 23213 15453 23247 15487
rect 23397 15453 23431 15487
rect 23857 15453 23891 15487
rect 23949 15453 23983 15487
rect 26801 15453 26835 15487
rect 26893 15453 26927 15487
rect 27261 15453 27295 15487
rect 27445 15453 27479 15487
rect 26295 15419 26329 15453
rect 12173 15385 12207 15419
rect 16773 15385 16807 15419
rect 19257 15385 19291 15419
rect 19441 15385 19475 15419
rect 26065 15385 26099 15419
rect 26525 15385 26559 15419
rect 12449 15317 12483 15351
rect 13921 15317 13955 15351
rect 18245 15317 18279 15351
rect 20085 15317 20119 15351
rect 26433 15317 26467 15351
rect 26709 15317 26743 15351
rect 27169 15317 27203 15351
rect 27353 15317 27387 15351
rect 5825 15113 5859 15147
rect 10977 15113 11011 15147
rect 13921 15113 13955 15147
rect 19625 15113 19659 15147
rect 26249 15113 26283 15147
rect 27905 15113 27939 15147
rect 4353 15045 4387 15079
rect 8769 15045 8803 15079
rect 9505 15045 9539 15079
rect 12449 15045 12483 15079
rect 16681 15045 16715 15079
rect 17417 15045 17451 15079
rect 17693 15045 17727 15079
rect 19073 15045 19107 15079
rect 24041 15045 24075 15079
rect 24777 15045 24811 15079
rect 24869 15045 24903 15079
rect 24987 15045 25021 15079
rect 27261 15045 27295 15079
rect 27471 15045 27505 15079
rect 8401 14977 8435 15011
rect 8494 14977 8528 15011
rect 8677 14977 8711 15011
rect 8907 14977 8941 15011
rect 11529 14977 11563 15011
rect 11713 14977 11747 15011
rect 11805 14977 11839 15011
rect 11897 14977 11931 15011
rect 16313 14977 16347 15011
rect 18245 14977 18279 15011
rect 19441 14977 19475 15011
rect 19717 14977 19751 15011
rect 19901 14977 19935 15011
rect 22109 14977 22143 15011
rect 22937 14977 22971 15011
rect 23305 14977 23339 15011
rect 23765 14977 23799 15011
rect 24686 14999 24720 15033
rect 25145 14977 25179 15011
rect 26065 14977 26099 15011
rect 26157 14977 26191 15011
rect 26341 14977 26375 15011
rect 27169 14977 27203 15011
rect 27353 14977 27387 15011
rect 27721 14977 27755 15011
rect 27997 14977 28031 15011
rect 4077 14909 4111 14943
rect 6561 14909 6595 14943
rect 6837 14909 6871 14943
rect 9229 14909 9263 14943
rect 12173 14909 12207 14943
rect 14473 14909 14507 14943
rect 14749 14909 14783 14943
rect 20177 14909 20211 14943
rect 21649 14909 21683 14943
rect 22293 14909 22327 14943
rect 25421 14909 25455 14943
rect 27629 14909 27663 14943
rect 9045 14841 9079 14875
rect 17969 14841 18003 14875
rect 27721 14841 27755 14875
rect 8309 14773 8343 14807
rect 12081 14773 12115 14807
rect 16221 14773 16255 14807
rect 16405 14773 16439 14807
rect 18153 14773 18187 14807
rect 19257 14773 19291 14807
rect 24501 14773 24535 14807
rect 26985 14773 27019 14807
rect 7665 14569 7699 14603
rect 11884 14569 11918 14603
rect 13369 14569 13403 14603
rect 16037 14569 16071 14603
rect 18797 14569 18831 14603
rect 20085 14569 20119 14603
rect 20729 14569 20763 14603
rect 23121 14569 23155 14603
rect 23581 14569 23615 14603
rect 24758 14569 24792 14603
rect 22293 14501 22327 14535
rect 8125 14433 8159 14467
rect 11621 14433 11655 14467
rect 15117 14433 15151 14467
rect 20269 14433 20303 14467
rect 22753 14433 22787 14467
rect 24501 14433 24535 14467
rect 26801 14433 26835 14467
rect 27077 14433 27111 14467
rect 28825 14433 28859 14467
rect 7113 14365 7147 14399
rect 7389 14365 7423 14399
rect 7481 14365 7515 14399
rect 10425 14365 10459 14399
rect 10573 14365 10607 14399
rect 10793 14365 10827 14399
rect 10890 14365 10924 14399
rect 14197 14365 14231 14399
rect 15761 14365 15795 14399
rect 16497 14365 16531 14399
rect 16589 14365 16623 14399
rect 18521 14365 18555 14399
rect 18613 14365 18647 14399
rect 18889 14365 18923 14399
rect 19441 14365 19475 14399
rect 19625 14365 19659 14399
rect 19763 14365 19797 14399
rect 19901 14365 19935 14399
rect 20453 14365 20487 14399
rect 20913 14365 20947 14399
rect 21373 14365 21407 14399
rect 21557 14365 21591 14399
rect 21649 14365 21683 14399
rect 21742 14365 21776 14399
rect 22155 14365 22189 14399
rect 22385 14365 22419 14399
rect 22569 14365 22603 14399
rect 22661 14365 22695 14399
rect 22937 14365 22971 14399
rect 23489 14365 23523 14399
rect 7297 14297 7331 14331
rect 10701 14297 10735 14331
rect 14565 14297 14599 14331
rect 19533 14297 19567 14331
rect 19993 14297 20027 14331
rect 21465 14297 21499 14331
rect 21925 14297 21959 14331
rect 22017 14297 22051 14331
rect 26525 14297 26559 14331
rect 8677 14229 8711 14263
rect 11069 14229 11103 14263
rect 15669 14229 15703 14263
rect 16221 14229 16255 14263
rect 16773 14229 16807 14263
rect 18337 14229 18371 14263
rect 19257 14229 19291 14263
rect 20637 14229 20671 14263
rect 23949 14229 23983 14263
rect 6377 14025 6411 14059
rect 20545 14025 20579 14059
rect 21557 14025 21591 14059
rect 23673 14025 23707 14059
rect 26249 14025 26283 14059
rect 3617 13957 3651 13991
rect 15209 13957 15243 13991
rect 19717 13957 19751 13991
rect 19901 13957 19935 13991
rect 1593 13889 1627 13923
rect 6561 13889 6595 13923
rect 6745 13889 6779 13923
rect 9873 13889 9907 13923
rect 10057 13889 10091 13923
rect 10149 13889 10183 13923
rect 10241 13889 10275 13923
rect 14105 13889 14139 13923
rect 14197 13889 14231 13923
rect 14473 13889 14507 13923
rect 14933 13889 14967 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 18613 13889 18647 13923
rect 18705 13889 18739 13923
rect 18889 13889 18923 13923
rect 18981 13889 19015 13923
rect 19073 13889 19107 13923
rect 19257 13889 19291 13923
rect 19349 13889 19383 13923
rect 19533 13889 19567 13923
rect 19625 13889 19659 13923
rect 20177 13889 20211 13923
rect 22661 13889 22695 13923
rect 23489 13889 23523 13923
rect 24501 13889 24535 13923
rect 27997 13889 28031 13923
rect 1869 13821 1903 13855
rect 6653 13821 6687 13855
rect 6837 13821 6871 13855
rect 10793 13821 10827 13855
rect 11345 13821 11379 13855
rect 14381 13821 14415 13855
rect 20269 13821 20303 13855
rect 21097 13821 21131 13855
rect 24041 13821 24075 13855
rect 24133 13821 24167 13855
rect 24317 13821 24351 13855
rect 24777 13821 24811 13855
rect 28365 13821 28399 13855
rect 13921 13753 13955 13787
rect 15485 13753 15519 13787
rect 20085 13753 20119 13787
rect 21373 13753 21407 13787
rect 10425 13685 10459 13719
rect 18429 13685 18463 13719
rect 20177 13685 20211 13719
rect 2237 13481 2271 13515
rect 6285 13481 6319 13515
rect 8493 13481 8527 13515
rect 18797 13481 18831 13515
rect 19533 13481 19567 13515
rect 25789 13481 25823 13515
rect 29009 13481 29043 13515
rect 2605 13413 2639 13447
rect 12081 13413 12115 13447
rect 15301 13413 15335 13447
rect 15853 13413 15887 13447
rect 22477 13413 22511 13447
rect 3249 13345 3283 13379
rect 17325 13345 17359 13379
rect 19349 13345 19383 13379
rect 25145 13345 25179 13379
rect 2421 13277 2455 13311
rect 2973 13277 3007 13311
rect 3433 13277 3467 13311
rect 3617 13277 3651 13311
rect 6193 13277 6227 13311
rect 6561 13277 6595 13311
rect 7297 13277 7331 13311
rect 7573 13277 7607 13311
rect 8125 13277 8159 13311
rect 8401 13277 8435 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9689 13277 9723 13311
rect 10425 13277 10459 13311
rect 10518 13277 10552 13311
rect 10793 13277 10827 13311
rect 10890 13277 10924 13311
rect 11529 13277 11563 13311
rect 11897 13277 11931 13311
rect 15577 13277 15611 13311
rect 15761 13277 15795 13311
rect 16313 13277 16347 13311
rect 16957 13277 16991 13311
rect 17141 13277 17175 13311
rect 18797 13277 18831 13311
rect 18981 13277 19015 13311
rect 19257 13277 19291 13311
rect 19533 13277 19567 13311
rect 21741 13277 21775 13311
rect 21925 13277 21959 13311
rect 22845 13277 22879 13311
rect 23305 13277 23339 13311
rect 28825 13277 28859 13311
rect 7849 13209 7883 13243
rect 10701 13209 10735 13243
rect 11713 13209 11747 13243
rect 11805 13209 11839 13243
rect 16129 13209 16163 13243
rect 3065 13141 3099 13175
rect 3525 13141 3559 13175
rect 7113 13141 7147 13175
rect 9137 13141 9171 13175
rect 11069 13141 11103 13175
rect 16865 13141 16899 13175
rect 19717 13141 19751 13175
rect 21833 13141 21867 13175
rect 10977 12937 11011 12971
rect 12173 12937 12207 12971
rect 14657 12937 14691 12971
rect 16497 12937 16531 12971
rect 21189 12937 21223 12971
rect 5365 12869 5399 12903
rect 5917 12869 5951 12903
rect 7481 12869 7515 12903
rect 9505 12869 9539 12903
rect 14013 12869 14047 12903
rect 14289 12869 14323 12903
rect 16957 12869 16991 12903
rect 18337 12869 18371 12903
rect 22017 12869 22051 12903
rect 1777 12801 1811 12835
rect 3893 12801 3927 12835
rect 4077 12801 4111 12835
rect 4629 12801 4663 12835
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 6009 12801 6043 12835
rect 6929 12801 6963 12835
rect 7205 12801 7239 12835
rect 7573 12801 7607 12835
rect 12265 12801 12299 12835
rect 12449 12801 12483 12835
rect 12541 12801 12575 12835
rect 12633 12801 12667 12835
rect 13461 12801 13495 12835
rect 14105 12801 14139 12835
rect 14381 12801 14415 12835
rect 14473 12801 14507 12835
rect 16681 12801 16715 12835
rect 16865 12801 16899 12835
rect 17049 12801 17083 12835
rect 18061 12801 18095 12835
rect 21465 12801 21499 12835
rect 23029 12801 23063 12835
rect 23121 12801 23155 12835
rect 2053 12733 2087 12767
rect 3801 12733 3835 12767
rect 7849 12733 7883 12767
rect 9229 12733 9263 12767
rect 11529 12733 11563 12767
rect 14749 12733 14783 12767
rect 15025 12733 15059 12767
rect 20085 12733 20119 12767
rect 21373 12733 21407 12767
rect 21557 12733 21591 12767
rect 22753 12733 22787 12767
rect 17233 12665 17267 12699
rect 4261 12597 4295 12631
rect 6193 12597 6227 12631
rect 12817 12597 12851 12631
rect 23029 12597 23063 12631
rect 23397 12597 23431 12631
rect 2697 12393 2731 12427
rect 3525 12393 3559 12427
rect 6929 12393 6963 12427
rect 7941 12393 7975 12427
rect 10977 12393 11011 12427
rect 15393 12325 15427 12359
rect 16221 12325 16255 12359
rect 3341 12257 3375 12291
rect 4629 12257 4663 12291
rect 5181 12257 5215 12291
rect 5457 12257 5491 12291
rect 7389 12257 7423 12291
rect 9229 12257 9263 12291
rect 11805 12257 11839 12291
rect 12173 12257 12207 12291
rect 12449 12257 12483 12291
rect 16773 12257 16807 12291
rect 23029 12257 23063 12291
rect 2881 12189 2915 12223
rect 2973 12189 3007 12223
rect 3065 12189 3099 12223
rect 3203 12189 3237 12223
rect 3433 12189 3467 12223
rect 3617 12189 3651 12223
rect 4445 12189 4479 12223
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 7205 12189 7239 12223
rect 7297 12189 7331 12223
rect 7665 12189 7699 12223
rect 7757 12189 7791 12223
rect 14197 12189 14231 12223
rect 14749 12189 14783 12223
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 15209 12189 15243 12223
rect 16129 12189 16163 12223
rect 16681 12189 16715 12223
rect 19993 12189 20027 12223
rect 22477 12189 22511 12223
rect 22937 12189 22971 12223
rect 24041 12189 24075 12223
rect 9505 12121 9539 12155
rect 11069 12121 11103 12155
rect 15117 12121 15151 12155
rect 23397 12121 23431 12155
rect 4261 12053 4295 12087
rect 7021 12053 7055 12087
rect 13921 12053 13955 12087
rect 19809 12053 19843 12087
rect 23673 12053 23707 12087
rect 23857 12053 23891 12087
rect 4077 11849 4111 11883
rect 7021 11849 7055 11883
rect 13829 11849 13863 11883
rect 16497 11849 16531 11883
rect 19993 11849 20027 11883
rect 23765 11849 23799 11883
rect 24409 11849 24443 11883
rect 6469 11781 6503 11815
rect 10885 11781 10919 11815
rect 12357 11781 12391 11815
rect 13921 11781 13955 11815
rect 16221 11781 16255 11815
rect 1409 11713 1443 11747
rect 1777 11713 1811 11747
rect 2237 11713 2271 11747
rect 4261 11713 4295 11747
rect 4905 11713 4939 11747
rect 6929 11713 6963 11747
rect 7573 11713 7607 11747
rect 10471 11713 10505 11747
rect 10609 11713 10643 11747
rect 12081 11713 12115 11747
rect 14105 11713 14139 11747
rect 15945 11713 15979 11747
rect 16129 11713 16163 11747
rect 16313 11713 16347 11747
rect 18521 11713 18555 11747
rect 19533 11713 19567 11747
rect 19809 11713 19843 11747
rect 20269 11713 20303 11747
rect 20545 11713 20579 11747
rect 21833 11713 21867 11747
rect 22661 11713 22695 11747
rect 22845 11713 22879 11747
rect 23489 11713 23523 11747
rect 23949 11713 23983 11747
rect 24225 11713 24259 11747
rect 25697 11713 25731 11747
rect 2329 11645 2363 11679
rect 2605 11645 2639 11679
rect 5641 11645 5675 11679
rect 8677 11645 8711 11679
rect 9045 11645 9079 11679
rect 17049 11645 17083 11679
rect 23305 11645 23339 11679
rect 23581 11645 23615 11679
rect 25605 11645 25639 11679
rect 6469 11577 6503 11611
rect 18429 11577 18463 11611
rect 4813 11509 4847 11543
rect 7205 11509 7239 11543
rect 8217 11509 8251 11543
rect 14289 11509 14323 11543
rect 17601 11509 17635 11543
rect 24133 11509 24167 11543
rect 26065 11509 26099 11543
rect 4353 11305 4387 11339
rect 5720 11305 5754 11339
rect 7849 11305 7883 11339
rect 18061 11305 18095 11339
rect 20250 11305 20284 11339
rect 22109 11305 22143 11339
rect 26709 11305 26743 11339
rect 7205 11237 7239 11271
rect 16221 11237 16255 11271
rect 18889 11237 18923 11271
rect 22477 11237 22511 11271
rect 24685 11237 24719 11271
rect 1869 11169 1903 11203
rect 5457 11169 5491 11203
rect 16313 11169 16347 11203
rect 19993 11169 20027 11203
rect 24961 11169 24995 11203
rect 26893 11169 26927 11203
rect 29009 11169 29043 11203
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 4169 11101 4203 11135
rect 4537 11101 4571 11135
rect 7297 11101 7331 11135
rect 7665 11101 7699 11135
rect 9965 11101 9999 11135
rect 15669 11101 15703 11135
rect 16037 11101 16071 11135
rect 18521 11101 18555 11135
rect 18705 11101 18739 11135
rect 19441 11101 19475 11135
rect 22109 11101 22143 11135
rect 22293 11101 22327 11135
rect 22385 11101 22419 11135
rect 22661 11101 22695 11135
rect 23397 11101 23431 11135
rect 28733 11101 28767 11135
rect 2145 11033 2179 11067
rect 4077 11033 4111 11067
rect 7481 11033 7515 11067
rect 7573 11033 7607 11067
rect 10701 11033 10735 11067
rect 15853 11033 15887 11067
rect 15945 11033 15979 11067
rect 16589 11033 16623 11067
rect 19717 11033 19751 11067
rect 22017 11033 22051 11067
rect 23121 11033 23155 11067
rect 24041 11033 24075 11067
rect 24409 11033 24443 11067
rect 25237 11033 25271 11067
rect 3617 10965 3651 10999
rect 5089 10965 5123 10999
rect 24869 10965 24903 10999
rect 27537 10965 27571 10999
rect 5181 10761 5215 10795
rect 5917 10761 5951 10795
rect 6009 10761 6043 10795
rect 9689 10761 9723 10795
rect 14473 10761 14507 10795
rect 14565 10761 14599 10795
rect 17877 10761 17911 10795
rect 19993 10761 20027 10795
rect 20361 10761 20395 10795
rect 22753 10761 22787 10795
rect 25421 10761 25455 10795
rect 26157 10761 26191 10795
rect 3985 10693 4019 10727
rect 4813 10693 4847 10727
rect 4905 10693 4939 10727
rect 5457 10693 5491 10727
rect 6377 10693 6411 10727
rect 17141 10693 17175 10727
rect 17233 10693 17267 10727
rect 23121 10693 23155 10727
rect 24869 10693 24903 10727
rect 25973 10693 26007 10727
rect 3801 10625 3835 10659
rect 4077 10625 4111 10659
rect 4169 10625 4203 10659
rect 4629 10625 4663 10659
rect 4997 10625 5031 10659
rect 6653 10625 6687 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 10241 10625 10275 10659
rect 10333 10625 10367 10659
rect 10517 10625 10551 10659
rect 13737 10625 13771 10659
rect 13829 10625 13863 10659
rect 14381 10625 14415 10659
rect 16313 10625 16347 10659
rect 16497 10625 16531 10659
rect 16865 10625 16899 10659
rect 17013 10625 17047 10659
rect 17330 10625 17364 10659
rect 17874 10625 17908 10659
rect 18245 10625 18279 10659
rect 18613 10625 18647 10659
rect 18797 10625 18831 10659
rect 18981 10625 19015 10659
rect 19165 10625 19199 10659
rect 19257 10625 19291 10659
rect 20177 10625 20211 10659
rect 20637 10625 20671 10659
rect 20821 10625 20855 10659
rect 22109 10625 22143 10659
rect 22569 10625 22603 10659
rect 22845 10625 22879 10659
rect 25697 10625 25731 10659
rect 26341 10625 26375 10659
rect 26433 10625 26467 10659
rect 26525 10625 26559 10659
rect 26709 10625 26743 10659
rect 26801 10625 26835 10659
rect 6193 10557 6227 10591
rect 6469 10557 6503 10591
rect 13921 10557 13955 10591
rect 14013 10557 14047 10591
rect 16129 10557 16163 10591
rect 18337 10557 18371 10591
rect 19717 10557 19751 10591
rect 22385 10557 22419 10591
rect 25605 10557 25639 10591
rect 26065 10557 26099 10591
rect 5457 10489 5491 10523
rect 6837 10489 6871 10523
rect 14197 10489 14231 10523
rect 17693 10489 17727 10523
rect 4353 10421 4387 10455
rect 6561 10421 6595 10455
rect 10701 10421 10735 10455
rect 13553 10421 13587 10455
rect 14749 10421 14783 10455
rect 17509 10421 17543 10455
rect 19625 10421 19659 10455
rect 22385 10421 22419 10455
rect 4721 10217 4755 10251
rect 10609 10217 10643 10251
rect 13575 10217 13609 10251
rect 20729 10217 20763 10251
rect 22845 10217 22879 10251
rect 23305 10217 23339 10251
rect 25881 10217 25915 10251
rect 13277 10149 13311 10183
rect 20361 10149 20395 10183
rect 9597 10081 9631 10115
rect 10241 10081 10275 10115
rect 10701 10081 10735 10115
rect 11345 10081 11379 10115
rect 11989 10081 12023 10115
rect 16589 10081 16623 10115
rect 20453 10081 20487 10115
rect 23029 10081 23063 10115
rect 4077 10013 4111 10047
rect 9413 10013 9447 10047
rect 9873 10013 9907 10047
rect 10057 10013 10091 10047
rect 10149 10013 10183 10047
rect 10425 10013 10459 10047
rect 10885 10013 10919 10047
rect 11161 10013 11195 10047
rect 11259 10013 11293 10047
rect 11437 10015 11471 10049
rect 11713 10013 11747 10047
rect 12633 10013 12667 10047
rect 12817 10013 12851 10047
rect 14289 10013 14323 10047
rect 15393 10013 15427 10047
rect 15486 10013 15520 10047
rect 15669 10013 15703 10047
rect 15899 10013 15933 10047
rect 18429 10013 18463 10047
rect 19901 10013 19935 10047
rect 19993 10013 20027 10047
rect 22293 10013 22327 10047
rect 22477 10013 22511 10047
rect 23121 10013 23155 10047
rect 26065 10013 26099 10047
rect 26157 10013 26191 10047
rect 9505 9945 9539 9979
rect 13369 9945 13403 9979
rect 15761 9945 15795 9979
rect 16865 9945 16899 9979
rect 22845 9945 22879 9979
rect 25881 9945 25915 9979
rect 9045 9877 9079 9911
rect 11069 9877 11103 9911
rect 12817 9877 12851 9911
rect 13569 9877 13603 9911
rect 13737 9877 13771 9911
rect 14105 9877 14139 9911
rect 16037 9877 16071 9911
rect 18337 9877 18371 9911
rect 19073 9877 19107 9911
rect 22385 9877 22419 9911
rect 3709 9673 3743 9707
rect 9689 9673 9723 9707
rect 10609 9673 10643 9707
rect 17233 9673 17267 9707
rect 17785 9673 17819 9707
rect 18521 9673 18555 9707
rect 6469 9605 6503 9639
rect 7021 9605 7055 9639
rect 10149 9605 10183 9639
rect 10241 9605 10275 9639
rect 10379 9605 10413 9639
rect 11161 9605 11195 9639
rect 13185 9605 13219 9639
rect 13553 9605 13587 9639
rect 1961 9537 1995 9571
rect 4997 9537 5031 9571
rect 5089 9537 5123 9571
rect 5273 9537 5307 9571
rect 5365 9537 5399 9571
rect 5457 9537 5491 9571
rect 6929 9537 6963 9571
rect 8769 9537 8803 9571
rect 9321 9537 9355 9571
rect 9551 9537 9585 9571
rect 10057 9537 10091 9571
rect 10517 9537 10551 9571
rect 10609 9537 10643 9571
rect 10977 9537 11011 9571
rect 11253 9537 11287 9571
rect 11897 9537 11931 9571
rect 12541 9537 12575 9571
rect 13277 9537 13311 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 16957 9537 16991 9571
rect 17049 9537 17083 9571
rect 17782 9537 17816 9571
rect 18153 9537 18187 9571
rect 18518 9537 18552 9571
rect 26341 9537 26375 9571
rect 26433 9537 26467 9571
rect 26985 9537 27019 9571
rect 27905 9537 27939 9571
rect 27997 9537 28031 9571
rect 28181 9537 28215 9571
rect 28273 9537 28307 9571
rect 2237 9469 2271 9503
rect 4353 9469 4387 9503
rect 8677 9469 8711 9503
rect 8861 9469 8895 9503
rect 8953 9469 8987 9503
rect 9137 9469 9171 9503
rect 9413 9469 9447 9503
rect 9781 9469 9815 9503
rect 10885 9469 10919 9503
rect 15301 9469 15335 9503
rect 18245 9469 18279 9503
rect 18981 9469 19015 9503
rect 26617 9469 26651 9503
rect 6469 9401 6503 9435
rect 8493 9401 8527 9435
rect 9873 9401 9907 9435
rect 10701 9401 10735 9435
rect 10977 9401 11011 9435
rect 27629 9401 27663 9435
rect 5641 9333 5675 9367
rect 7205 9333 7239 9367
rect 17601 9333 17635 9367
rect 18337 9333 18371 9367
rect 18889 9333 18923 9367
rect 27721 9333 27755 9367
rect 2132 9129 2166 9163
rect 13093 9129 13127 9163
rect 22569 9129 22603 9163
rect 23029 9129 23063 9163
rect 27997 9129 28031 9163
rect 5365 9061 5399 9095
rect 1869 8993 1903 9027
rect 3617 8993 3651 9027
rect 5825 8993 5859 9027
rect 5917 8993 5951 9027
rect 6193 8993 6227 9027
rect 9321 8993 9355 9027
rect 11161 8993 11195 9027
rect 11370 8993 11404 9027
rect 14657 8993 14691 9027
rect 22201 8993 22235 9027
rect 22293 8993 22327 9027
rect 22661 8993 22695 9027
rect 26249 8993 26283 9027
rect 4261 8925 4295 8959
rect 6561 8925 6595 8959
rect 8953 8925 8987 8959
rect 10885 8925 10919 8959
rect 11621 8925 11655 8959
rect 11897 8925 11931 8959
rect 13001 8925 13035 8959
rect 13829 8925 13863 8959
rect 17969 8925 18003 8959
rect 18337 8925 18371 8959
rect 19349 8925 19383 8959
rect 22109 8925 22143 8959
rect 22845 8925 22879 8959
rect 25698 8925 25732 8959
rect 25999 8925 26033 8959
rect 26157 8925 26191 8959
rect 28365 8925 28399 8959
rect 5365 8857 5399 8891
rect 11253 8857 11287 8891
rect 13553 8857 13587 8891
rect 18153 8857 18187 8891
rect 18245 8857 18279 8891
rect 19901 8857 19935 8891
rect 22569 8857 22603 8891
rect 25789 8857 25823 8891
rect 25881 8857 25915 8891
rect 26525 8857 26559 8891
rect 28181 8857 28215 8891
rect 28549 8857 28583 8891
rect 4905 8789 4939 8823
rect 6101 8789 6135 8823
rect 7987 8789 8021 8823
rect 10747 8789 10781 8823
rect 11529 8789 11563 8823
rect 13651 8789 13685 8823
rect 13737 8789 13771 8823
rect 15209 8789 15243 8823
rect 18521 8789 18555 8823
rect 21741 8789 21775 8823
rect 25513 8789 25547 8823
rect 5457 8585 5491 8619
rect 5641 8585 5675 8619
rect 13369 8585 13403 8619
rect 20637 8585 20671 8619
rect 4997 8517 5031 8551
rect 7665 8517 7699 8551
rect 8309 8517 8343 8551
rect 9045 8517 9079 8551
rect 9229 8517 9263 8551
rect 13737 8517 13771 8551
rect 15485 8517 15519 8551
rect 23397 8517 23431 8551
rect 27077 8517 27111 8551
rect 2145 8449 2179 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 4261 8449 4295 8483
rect 4353 8449 4387 8483
rect 5273 8449 5307 8483
rect 6837 8449 6871 8483
rect 7297 8449 7331 8483
rect 13093 8449 13127 8483
rect 16681 8449 16715 8483
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 17141 8449 17175 8483
rect 17289 8449 17323 8483
rect 17417 8449 17451 8483
rect 17509 8449 17543 8483
rect 17647 8449 17681 8483
rect 18889 8449 18923 8483
rect 21097 8449 21131 8483
rect 22845 8449 22879 8483
rect 23029 8449 23063 8483
rect 23581 8449 23615 8483
rect 23949 8449 23983 8483
rect 24133 8449 24167 8483
rect 26065 8449 26099 8483
rect 26985 8449 27019 8483
rect 27261 8449 27295 8483
rect 27537 8449 27571 8483
rect 27813 8449 27847 8483
rect 2421 8381 2455 8415
rect 5089 8381 5123 8415
rect 5825 8381 5859 8415
rect 5917 8381 5951 8415
rect 6009 8381 6043 8415
rect 6101 8381 6135 8415
rect 6561 8381 6595 8415
rect 6653 8381 6687 8415
rect 6745 8381 6779 8415
rect 8769 8381 8803 8415
rect 8861 8381 8895 8415
rect 9965 8381 9999 8415
rect 13369 8381 13403 8415
rect 13461 8381 13495 8415
rect 19165 8381 19199 8415
rect 23765 8381 23799 8415
rect 25881 8381 25915 8415
rect 26341 8381 26375 8415
rect 26801 8381 26835 8415
rect 3893 8313 3927 8347
rect 4537 8313 4571 8347
rect 8309 8313 8343 8347
rect 13185 8313 13219 8347
rect 23673 8313 23707 8347
rect 23949 8313 23983 8347
rect 26617 8313 26651 8347
rect 5089 8245 5123 8279
rect 6377 8245 6411 8279
rect 17785 8245 17819 8279
rect 20913 8245 20947 8279
rect 23213 8245 23247 8279
rect 23857 8245 23891 8279
rect 26249 8245 26283 8279
rect 5181 8041 5215 8075
rect 5549 8041 5583 8075
rect 6101 8041 6135 8075
rect 13737 8041 13771 8075
rect 21833 8041 21867 8075
rect 25237 8041 25271 8075
rect 27537 8041 27571 8075
rect 6745 7973 6779 8007
rect 1961 7905 1995 7939
rect 5733 7905 5767 7939
rect 6285 7905 6319 7939
rect 20361 7905 20395 7939
rect 26249 7905 26283 7939
rect 27169 7905 27203 7939
rect 27537 7905 27571 7939
rect 1685 7837 1719 7871
rect 3985 7837 4019 7871
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 4997 7837 5031 7871
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 6377 7837 6411 7871
rect 7481 7837 7515 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14565 7837 14599 7871
rect 14749 7837 14783 7871
rect 16405 7837 16439 7871
rect 16589 7837 16623 7871
rect 16865 7837 16899 7871
rect 17049 7837 17083 7871
rect 17417 7837 17451 7871
rect 17693 7837 17727 7871
rect 17785 7837 17819 7871
rect 17933 7837 17967 7871
rect 18061 7837 18095 7871
rect 18250 7837 18284 7871
rect 20085 7837 20119 7871
rect 22017 7837 22051 7871
rect 22201 7837 22235 7871
rect 22293 7837 22327 7871
rect 22569 7837 22603 7871
rect 22871 7837 22905 7871
rect 23029 7837 23063 7871
rect 23121 7837 23155 7871
rect 23305 7837 23339 7871
rect 23673 7837 23707 7871
rect 23765 7837 23799 7871
rect 23857 7837 23891 7871
rect 24041 7837 24075 7871
rect 24409 7837 24443 7871
rect 24593 7837 24627 7871
rect 24869 7837 24903 7871
rect 25053 7837 25087 7871
rect 25789 7837 25823 7871
rect 26091 7837 26125 7871
rect 26525 7837 26559 7871
rect 27261 7837 27295 7871
rect 4813 7769 4847 7803
rect 4905 7769 4939 7803
rect 6101 7769 6135 7803
rect 6745 7769 6779 7803
rect 7297 7769 7331 7803
rect 13553 7769 13587 7803
rect 13769 7769 13803 7803
rect 17233 7769 17267 7803
rect 18153 7769 18187 7803
rect 22661 7769 22695 7803
rect 22753 7769 22787 7803
rect 25881 7769 25915 7803
rect 25973 7769 26007 7803
rect 3433 7701 3467 7735
rect 6561 7701 6595 7735
rect 7205 7701 7239 7735
rect 13921 7701 13955 7735
rect 14473 7701 14507 7735
rect 14657 7701 14691 7735
rect 16773 7701 16807 7735
rect 18429 7701 18463 7735
rect 22293 7701 22327 7735
rect 22385 7701 22419 7735
rect 23305 7701 23339 7735
rect 23397 7701 23431 7735
rect 24777 7701 24811 7735
rect 25605 7701 25639 7735
rect 27813 7701 27847 7735
rect 5641 7497 5675 7531
rect 16957 7497 16991 7531
rect 22569 7497 22603 7531
rect 22937 7497 22971 7531
rect 27169 7497 27203 7531
rect 11529 7429 11563 7463
rect 13001 7429 13035 7463
rect 13829 7429 13863 7463
rect 22477 7429 22511 7463
rect 23765 7429 23799 7463
rect 24133 7429 24167 7463
rect 25237 7429 25271 7463
rect 6009 7361 6043 7395
rect 10333 7361 10367 7395
rect 10609 7361 10643 7395
rect 10885 7361 10919 7395
rect 11805 7361 11839 7395
rect 12265 7361 12299 7395
rect 13185 7361 13219 7395
rect 13369 7361 13403 7395
rect 13553 7361 13587 7395
rect 16773 7361 16807 7395
rect 17049 7361 17083 7395
rect 17141 7361 17175 7395
rect 17289 7361 17323 7395
rect 17417 7361 17451 7395
rect 17509 7361 17543 7395
rect 17601 7361 17635 7395
rect 17877 7361 17911 7395
rect 18061 7361 18095 7395
rect 18245 7361 18279 7395
rect 18429 7361 18463 7395
rect 22753 7361 22787 7395
rect 23029 7361 23063 7395
rect 23857 7361 23891 7395
rect 24041 7361 24075 7395
rect 24225 7361 24259 7395
rect 24501 7361 24535 7395
rect 24685 7361 24719 7395
rect 24961 7361 24995 7395
rect 26985 7361 27019 7395
rect 27261 7361 27295 7395
rect 27445 7361 27479 7395
rect 27537 7361 27571 7395
rect 27721 7361 27755 7395
rect 28733 7361 28767 7395
rect 5825 7293 5859 7327
rect 5917 7293 5951 7327
rect 11069 7293 11103 7327
rect 13461 7293 13495 7327
rect 15577 7293 15611 7327
rect 18337 7293 18371 7327
rect 21925 7293 21959 7327
rect 23213 7293 23247 7327
rect 24593 7293 24627 7327
rect 12081 7225 12115 7259
rect 26709 7225 26743 7259
rect 27537 7225 27571 7259
rect 11897 7157 11931 7191
rect 11989 7157 12023 7191
rect 16773 7157 16807 7191
rect 17141 7157 17175 7191
rect 17877 7157 17911 7191
rect 24409 7157 24443 7191
rect 29009 7157 29043 7191
rect 11161 6953 11195 6987
rect 12173 6953 12207 6987
rect 14473 6953 14507 6987
rect 20808 6953 20842 6987
rect 22740 6953 22774 6987
rect 5089 6885 5123 6919
rect 7389 6885 7423 6919
rect 11345 6885 11379 6919
rect 22293 6885 22327 6919
rect 24225 6885 24259 6919
rect 5365 6817 5399 6851
rect 11437 6817 11471 6851
rect 13829 6817 13863 6851
rect 20545 6817 20579 6851
rect 22477 6817 22511 6851
rect 24501 6817 24535 6851
rect 4537 6749 4571 6783
rect 4905 6749 4939 6783
rect 6009 6749 6043 6783
rect 6377 6749 6411 6783
rect 6837 6749 6871 6783
rect 7113 6749 7147 6783
rect 7251 6749 7285 6783
rect 7481 6749 7515 6783
rect 7665 6749 7699 6783
rect 7895 6749 7929 6783
rect 9965 6749 9999 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 10793 6749 10827 6783
rect 12081 6749 12115 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 17049 6749 17083 6783
rect 17325 6749 17359 6783
rect 17417 6749 17451 6783
rect 17601 6749 17635 6783
rect 17877 6749 17911 6783
rect 18061 6749 18095 6783
rect 24409 6749 24443 6783
rect 24593 6749 24627 6783
rect 4721 6681 4755 6715
rect 4813 6681 4847 6715
rect 5917 6681 5951 6715
rect 6193 6681 6227 6715
rect 6285 6681 6319 6715
rect 7021 6681 7055 6715
rect 7757 6681 7791 6715
rect 10057 6681 10091 6715
rect 10517 6681 10551 6715
rect 11621 6681 11655 6715
rect 11713 6681 11747 6715
rect 11805 6681 11839 6715
rect 6561 6613 6595 6647
rect 8033 6613 8067 6647
rect 11161 6613 11195 6647
rect 11989 6613 12023 6647
rect 14105 6613 14139 6647
rect 16865 6613 16899 6647
rect 17233 6613 17267 6647
rect 17785 6613 17819 6647
rect 17969 6613 18003 6647
rect 5641 6409 5675 6443
rect 7021 6409 7055 6443
rect 8769 6409 8803 6443
rect 10885 6409 10919 6443
rect 11069 6409 11103 6443
rect 17141 6409 17175 6443
rect 20085 6409 20119 6443
rect 20637 6409 20671 6443
rect 4169 6341 4203 6375
rect 8033 6341 8067 6375
rect 10057 6341 10091 6375
rect 10517 6341 10551 6375
rect 13737 6341 13771 6375
rect 15485 6341 15519 6375
rect 16957 6341 16991 6375
rect 3893 6273 3927 6307
rect 7389 6273 7423 6307
rect 8217 6273 8251 6307
rect 9965 6273 9999 6307
rect 10241 6273 10275 6307
rect 10726 6273 10760 6307
rect 10983 6273 11017 6307
rect 11161 6273 11195 6307
rect 11529 6273 11563 6307
rect 17233 6273 17267 6307
rect 20269 6273 20303 6307
rect 20453 6273 20487 6307
rect 20545 6273 20579 6307
rect 20821 6273 20855 6307
rect 21005 6273 21039 6307
rect 21097 6273 21131 6307
rect 6377 6205 6411 6239
rect 10609 6205 10643 6239
rect 11713 6205 11747 6239
rect 13461 6205 13495 6239
rect 16957 6069 16991 6103
rect 4248 5865 4282 5899
rect 8033 5865 8067 5899
rect 10793 5865 10827 5899
rect 11069 5865 11103 5899
rect 17693 5865 17727 5899
rect 5733 5797 5767 5831
rect 17877 5797 17911 5831
rect 6285 5729 6319 5763
rect 6561 5729 6595 5763
rect 10057 5729 10091 5763
rect 10149 5729 10183 5763
rect 10885 5729 10919 5763
rect 3985 5661 4019 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 9965 5661 9999 5695
rect 10241 5661 10275 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 10977 5661 11011 5695
rect 11161 5661 11195 5695
rect 11253 5661 11287 5695
rect 11529 5661 11563 5695
rect 11621 5661 11655 5695
rect 17601 5661 17635 5695
rect 18153 5661 18187 5695
rect 18245 5661 18279 5695
rect 18429 5663 18463 5697
rect 9597 5593 9631 5627
rect 11437 5593 11471 5627
rect 17417 5593 17451 5627
rect 17877 5593 17911 5627
rect 9229 5525 9263 5559
rect 9781 5525 9815 5559
rect 11805 5525 11839 5559
rect 18061 5525 18095 5559
rect 18337 5525 18371 5559
rect 8125 5321 8159 5355
rect 16891 5321 16925 5355
rect 17325 5321 17359 5355
rect 20361 5321 20395 5355
rect 28273 5321 28307 5355
rect 10333 5253 10367 5287
rect 16681 5253 16715 5287
rect 6377 5185 6411 5219
rect 8493 5185 8527 5219
rect 11529 5185 11563 5219
rect 11897 5185 11931 5219
rect 17141 5185 17175 5219
rect 17785 5185 17819 5219
rect 18061 5185 18095 5219
rect 18245 5185 18279 5219
rect 18521 5185 18555 5219
rect 18705 5185 18739 5219
rect 18981 5185 19015 5219
rect 19165 5185 19199 5219
rect 19625 5185 19659 5219
rect 20269 5185 20303 5219
rect 28089 5185 28123 5219
rect 6653 5117 6687 5151
rect 8861 5117 8895 5151
rect 10425 5117 10459 5151
rect 13323 5117 13357 5151
rect 17509 5117 17543 5151
rect 20085 5117 20119 5151
rect 11069 5049 11103 5083
rect 17049 5049 17083 5083
rect 16865 4981 16899 5015
rect 17509 4981 17543 5015
rect 17877 4981 17911 5015
rect 18889 4981 18923 5015
rect 18981 4981 19015 5015
rect 19717 4981 19751 5015
rect 10701 4777 10735 4811
rect 11345 4777 11379 4811
rect 16037 4777 16071 4811
rect 16957 4777 16991 4811
rect 17601 4777 17635 4811
rect 17785 4777 17819 4811
rect 19993 4777 20027 4811
rect 20453 4777 20487 4811
rect 16221 4709 16255 4743
rect 18797 4709 18831 4743
rect 8953 4641 8987 4675
rect 9321 4641 9355 4675
rect 11161 4641 11195 4675
rect 13369 4641 13403 4675
rect 17693 4641 17727 4675
rect 18153 4641 18187 4675
rect 18245 4641 18279 4675
rect 18429 4641 18463 4675
rect 18889 4641 18923 4675
rect 19442 4641 19476 4675
rect 19533 4641 19567 4675
rect 19625 4641 19659 4675
rect 11069 4573 11103 4607
rect 13093 4573 13127 4607
rect 13277 4573 13311 4607
rect 15945 4573 15979 4607
rect 16129 4573 16163 4607
rect 16497 4573 16531 4607
rect 16589 4573 16623 4607
rect 17417 4573 17451 4607
rect 17969 4573 18003 4607
rect 18613 4573 18647 4607
rect 19717 4573 19751 4607
rect 19901 4573 19935 4607
rect 20177 4573 20211 4607
rect 20545 4573 20579 4607
rect 20729 4573 20763 4607
rect 16221 4505 16255 4539
rect 20637 4505 20671 4539
rect 12909 4437 12943 4471
rect 16405 4437 16439 4471
rect 16957 4437 16991 4471
rect 17141 4437 17175 4471
rect 17233 4437 17267 4471
rect 19257 4437 19291 4471
rect 13185 4233 13219 4267
rect 13921 4233 13955 4267
rect 14473 4233 14507 4267
rect 19993 4233 20027 4267
rect 24041 4165 24075 4199
rect 24225 4165 24259 4199
rect 24777 4165 24811 4199
rect 2421 4097 2455 4131
rect 13123 4097 13157 4131
rect 13645 4097 13679 4131
rect 13737 4097 13771 4131
rect 14381 4097 14415 4131
rect 14565 4097 14599 4131
rect 15577 4097 15611 4131
rect 15761 4097 15795 4131
rect 16037 4097 16071 4131
rect 16313 4097 16347 4131
rect 16681 4097 16715 4131
rect 17325 4097 17359 4131
rect 17601 4097 17635 4131
rect 18797 4097 18831 4131
rect 19257 4097 19291 4131
rect 19717 4097 19751 4131
rect 20085 4097 20119 4131
rect 24593 4097 24627 4131
rect 14105 4029 14139 4063
rect 16221 4029 16255 4063
rect 17417 4029 17451 4063
rect 19533 4029 19567 4063
rect 19993 4029 20027 4063
rect 13001 3961 13035 3995
rect 15853 3961 15887 3995
rect 2237 3893 2271 3927
rect 13553 3893 13587 3927
rect 14289 3893 14323 3927
rect 15669 3893 15703 3927
rect 19809 3893 19843 3927
rect 20177 3893 20211 3927
rect 24409 3893 24443 3927
rect 24961 3893 24995 3927
rect 12633 3689 12667 3723
rect 14565 3689 14599 3723
rect 14749 3621 14783 3655
rect 15117 3621 15151 3655
rect 15485 3621 15519 3655
rect 16405 3553 16439 3587
rect 18061 3553 18095 3587
rect 18981 3553 19015 3587
rect 1501 3485 1535 3519
rect 2421 3485 2455 3519
rect 12541 3485 12575 3519
rect 13001 3485 13035 3519
rect 13277 3485 13311 3519
rect 13461 3485 13495 3519
rect 13737 3485 13771 3519
rect 14473 3485 14507 3519
rect 14565 3485 14599 3519
rect 14841 3485 14875 3519
rect 15393 3485 15427 3519
rect 15577 3485 15611 3519
rect 16681 3485 16715 3519
rect 16773 3485 16807 3519
rect 16865 3485 16899 3519
rect 17049 3485 17083 3519
rect 18705 3485 18739 3519
rect 25421 3485 25455 3519
rect 14105 3417 14139 3451
rect 17877 3417 17911 3451
rect 1593 3349 1627 3383
rect 2237 3349 2271 3383
rect 12817 3349 12851 3383
rect 13829 3349 13863 3383
rect 15301 3349 15335 3383
rect 17509 3349 17543 3383
rect 17969 3349 18003 3383
rect 18337 3349 18371 3383
rect 18797 3349 18831 3383
rect 25237 3349 25271 3383
rect 13001 3145 13035 3179
rect 14565 3145 14599 3179
rect 17601 3145 17635 3179
rect 17969 3145 18003 3179
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 13369 3009 13403 3043
rect 13461 3009 13495 3043
rect 13645 3009 13679 3043
rect 13737 3009 13771 3043
rect 14013 3009 14047 3043
rect 14197 3009 14231 3043
rect 14289 3009 14323 3043
rect 14381 3009 14415 3043
rect 14565 3009 14599 3043
rect 16865 3009 16899 3043
rect 17049 3009 17083 3043
rect 17141 3009 17175 3043
rect 17233 3009 17267 3043
rect 17693 3009 17727 3043
rect 17785 3009 17819 3043
rect 18061 3009 18095 3043
rect 18245 3009 18279 3043
rect 28825 3009 28859 3043
rect 16957 2941 16991 2975
rect 17417 2941 17451 2975
rect 17509 2941 17543 2975
rect 17969 2941 18003 2975
rect 13829 2873 13863 2907
rect 13185 2805 13219 2839
rect 18061 2805 18095 2839
rect 29009 2805 29043 2839
rect 13461 2601 13495 2635
rect 1501 2397 1535 2431
rect 3893 2397 3927 2431
rect 13461 2397 13495 2431
rect 13645 2397 13679 2431
rect 15025 2397 15059 2431
rect 25973 2397 26007 2431
rect 28733 2397 28767 2431
rect 7297 2329 7331 2363
rect 11621 2329 11655 2363
rect 19349 2329 19383 2363
rect 22109 2329 22143 2363
rect 29101 2329 29135 2363
rect 1593 2261 1627 2295
rect 4169 2261 4203 2295
rect 7389 2261 7423 2295
rect 11713 2261 11747 2295
rect 15301 2261 15335 2295
rect 19441 2261 19475 2295
rect 22201 2261 22235 2295
rect 26249 2261 26283 2295
<< metal1 >>
rect 1104 30490 29440 30512
rect 1104 30438 5151 30490
rect 5203 30438 5215 30490
rect 5267 30438 5279 30490
rect 5331 30438 5343 30490
rect 5395 30438 5407 30490
rect 5459 30438 12234 30490
rect 12286 30438 12298 30490
rect 12350 30438 12362 30490
rect 12414 30438 12426 30490
rect 12478 30438 12490 30490
rect 12542 30438 19317 30490
rect 19369 30438 19381 30490
rect 19433 30438 19445 30490
rect 19497 30438 19509 30490
rect 19561 30438 19573 30490
rect 19625 30438 26400 30490
rect 26452 30438 26464 30490
rect 26516 30438 26528 30490
rect 26580 30438 26592 30490
rect 26644 30438 26656 30490
rect 26708 30438 29440 30490
rect 1104 30416 29440 30438
rect 6730 30336 6736 30388
rect 6788 30336 6794 30388
rect 9674 30268 9680 30320
rect 9732 30308 9738 30320
rect 10229 30311 10287 30317
rect 10229 30308 10241 30311
rect 9732 30280 10241 30308
rect 9732 30268 9738 30280
rect 10229 30277 10241 30280
rect 10275 30277 10287 30311
rect 10229 30271 10287 30277
rect 21266 30268 21272 30320
rect 21324 30308 21330 30320
rect 22281 30311 22339 30317
rect 22281 30308 22293 30311
rect 21324 30280 22293 30308
rect 21324 30268 21330 30280
rect 22281 30277 22293 30280
rect 22327 30277 22339 30311
rect 22281 30271 22339 30277
rect 25406 30268 25412 30320
rect 25464 30308 25470 30320
rect 25685 30311 25743 30317
rect 25685 30308 25697 30311
rect 25464 30280 25697 30308
rect 25464 30268 25470 30280
rect 25685 30277 25697 30280
rect 25731 30277 25743 30311
rect 28994 30308 29000 30320
rect 25685 30271 25743 30277
rect 28368 30280 29000 30308
rect 1578 30200 1584 30252
rect 1636 30200 1642 30252
rect 2777 30243 2835 30249
rect 2777 30209 2789 30243
rect 2823 30240 2835 30243
rect 3326 30240 3332 30252
rect 2823 30212 3332 30240
rect 2823 30209 2835 30212
rect 2777 30203 2835 30209
rect 3326 30200 3332 30212
rect 3384 30200 3390 30252
rect 6086 30200 6092 30252
rect 6144 30240 6150 30252
rect 6641 30243 6699 30249
rect 6641 30240 6653 30243
rect 6144 30212 6653 30240
rect 6144 30200 6150 30212
rect 6641 30209 6653 30212
rect 6687 30209 6699 30243
rect 6641 30203 6699 30209
rect 9858 30200 9864 30252
rect 9916 30200 9922 30252
rect 14182 30200 14188 30252
rect 14240 30200 14246 30252
rect 17586 30200 17592 30252
rect 17644 30200 17650 30252
rect 21910 30200 21916 30252
rect 21968 30200 21974 30252
rect 25314 30200 25320 30252
rect 25372 30200 25378 30252
rect 28368 30249 28396 30280
rect 28994 30268 29000 30280
rect 29052 30268 29058 30320
rect 28353 30243 28411 30249
rect 28353 30209 28365 30243
rect 28399 30209 28411 30243
rect 28353 30203 28411 30209
rect 28718 30200 28724 30252
rect 28776 30200 28782 30252
rect 28902 30132 28908 30184
rect 28960 30172 28966 30184
rect 28997 30175 29055 30181
rect 28997 30172 29009 30175
rect 28960 30144 29009 30172
rect 28960 30132 28966 30144
rect 28997 30141 29009 30144
rect 29043 30141 29055 30175
rect 28997 30135 29055 30141
rect 13814 30064 13820 30116
rect 13872 30104 13878 30116
rect 14369 30107 14427 30113
rect 14369 30104 14381 30107
rect 13872 30076 14381 30104
rect 13872 30064 13878 30076
rect 14369 30073 14381 30076
rect 14415 30073 14427 30107
rect 14369 30067 14427 30073
rect 17402 30064 17408 30116
rect 17460 30104 17466 30116
rect 17773 30107 17831 30113
rect 17773 30104 17785 30107
rect 17460 30076 17785 30104
rect 17460 30064 17466 30076
rect 17773 30073 17785 30076
rect 17819 30073 17831 30107
rect 17773 30067 17831 30073
rect 1397 30039 1455 30045
rect 1397 30005 1409 30039
rect 1443 30036 1455 30039
rect 1578 30036 1584 30048
rect 1443 30008 1584 30036
rect 1443 30005 1455 30008
rect 1397 29999 1455 30005
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 2866 29996 2872 30048
rect 2924 29996 2930 30048
rect 28534 29996 28540 30048
rect 28592 29996 28598 30048
rect 1104 29946 29440 29968
rect 1104 29894 4491 29946
rect 4543 29894 4555 29946
rect 4607 29894 4619 29946
rect 4671 29894 4683 29946
rect 4735 29894 4747 29946
rect 4799 29894 11574 29946
rect 11626 29894 11638 29946
rect 11690 29894 11702 29946
rect 11754 29894 11766 29946
rect 11818 29894 11830 29946
rect 11882 29894 18657 29946
rect 18709 29894 18721 29946
rect 18773 29894 18785 29946
rect 18837 29894 18849 29946
rect 18901 29894 18913 29946
rect 18965 29894 25740 29946
rect 25792 29894 25804 29946
rect 25856 29894 25868 29946
rect 25920 29894 25932 29946
rect 25984 29894 25996 29946
rect 26048 29894 29440 29946
rect 1104 29872 29440 29894
rect 21910 29792 21916 29844
rect 21968 29832 21974 29844
rect 23661 29835 23719 29841
rect 23661 29832 23673 29835
rect 21968 29804 23673 29832
rect 21968 29792 21974 29804
rect 23661 29801 23673 29804
rect 23707 29801 23719 29835
rect 23661 29795 23719 29801
rect 23934 29764 23940 29776
rect 14844 29736 23940 29764
rect 5537 29699 5595 29705
rect 5537 29696 5549 29699
rect 5000 29668 5549 29696
rect 5000 29640 5028 29668
rect 5537 29665 5549 29668
rect 5583 29665 5595 29699
rect 14090 29696 14096 29708
rect 5537 29659 5595 29665
rect 9048 29668 14096 29696
rect 9048 29640 9076 29668
rect 14090 29656 14096 29668
rect 14148 29696 14154 29708
rect 14844 29696 14872 29736
rect 23934 29724 23940 29736
rect 23992 29724 23998 29776
rect 14148 29668 14872 29696
rect 14148 29656 14154 29668
rect 4982 29588 4988 29640
rect 5040 29588 5046 29640
rect 5077 29631 5135 29637
rect 5077 29597 5089 29631
rect 5123 29597 5135 29631
rect 5077 29591 5135 29597
rect 5092 29560 5120 29591
rect 5166 29588 5172 29640
rect 5224 29628 5230 29640
rect 5445 29631 5503 29637
rect 5445 29628 5457 29631
rect 5224 29600 5457 29628
rect 5224 29588 5230 29600
rect 5445 29597 5457 29600
rect 5491 29597 5503 29631
rect 5445 29591 5503 29597
rect 5626 29588 5632 29640
rect 5684 29588 5690 29640
rect 5718 29588 5724 29640
rect 5776 29588 5782 29640
rect 8478 29628 8484 29640
rect 7300 29600 8484 29628
rect 5994 29560 6000 29572
rect 5092 29532 6000 29560
rect 5994 29520 6000 29532
rect 6052 29520 6058 29572
rect 7300 29504 7328 29600
rect 8478 29588 8484 29600
rect 8536 29588 8542 29640
rect 9030 29588 9036 29640
rect 9088 29588 9094 29640
rect 11241 29631 11299 29637
rect 11241 29597 11253 29631
rect 11287 29628 11299 29631
rect 11330 29628 11336 29640
rect 11287 29600 11336 29628
rect 11287 29597 11299 29600
rect 11241 29591 11299 29597
rect 11330 29588 11336 29600
rect 11388 29628 11394 29640
rect 13262 29628 13268 29640
rect 11388 29600 13268 29628
rect 11388 29588 11394 29600
rect 13262 29588 13268 29600
rect 13320 29588 13326 29640
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29628 14795 29631
rect 14844 29628 14872 29668
rect 16206 29656 16212 29708
rect 16264 29696 16270 29708
rect 16761 29699 16819 29705
rect 16761 29696 16773 29699
rect 16264 29668 16773 29696
rect 16264 29656 16270 29668
rect 16761 29665 16773 29668
rect 16807 29665 16819 29699
rect 19150 29696 19156 29708
rect 16761 29659 16819 29665
rect 16868 29668 19156 29696
rect 16868 29637 16896 29668
rect 19150 29656 19156 29668
rect 19208 29656 19214 29708
rect 14783 29600 14872 29628
rect 16853 29631 16911 29637
rect 14783 29597 14795 29600
rect 14737 29591 14795 29597
rect 16853 29597 16865 29631
rect 16899 29597 16911 29631
rect 16853 29591 16911 29597
rect 17497 29631 17555 29637
rect 17497 29597 17509 29631
rect 17543 29597 17555 29631
rect 17497 29591 17555 29597
rect 7377 29563 7435 29569
rect 7377 29529 7389 29563
rect 7423 29529 7435 29563
rect 7377 29523 7435 29529
rect 4890 29452 4896 29504
rect 4948 29452 4954 29504
rect 5261 29495 5319 29501
rect 5261 29461 5273 29495
rect 5307 29492 5319 29495
rect 5810 29492 5816 29504
rect 5307 29464 5816 29492
rect 5307 29461 5319 29464
rect 5261 29455 5319 29461
rect 5810 29452 5816 29464
rect 5868 29452 5874 29504
rect 5902 29452 5908 29504
rect 5960 29492 5966 29504
rect 7282 29492 7288 29504
rect 5960 29464 7288 29492
rect 5960 29452 5966 29464
rect 7282 29452 7288 29464
rect 7340 29452 7346 29504
rect 7392 29492 7420 29523
rect 7558 29520 7564 29572
rect 7616 29520 7622 29572
rect 8496 29560 8524 29588
rect 9401 29563 9459 29569
rect 9401 29560 9413 29563
rect 8496 29532 9413 29560
rect 9401 29529 9413 29532
rect 9447 29529 9459 29563
rect 9401 29523 9459 29529
rect 14274 29520 14280 29572
rect 14332 29560 14338 29572
rect 15105 29563 15163 29569
rect 15105 29560 15117 29563
rect 14332 29532 15117 29560
rect 14332 29520 14338 29532
rect 15105 29529 15117 29532
rect 15151 29529 15163 29563
rect 15105 29523 15163 29529
rect 16482 29520 16488 29572
rect 16540 29560 16546 29572
rect 17512 29560 17540 29591
rect 20806 29588 20812 29640
rect 20864 29588 20870 29640
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29628 23903 29631
rect 25222 29628 25228 29640
rect 23891 29600 25228 29628
rect 23891 29597 23903 29600
rect 23845 29591 23903 29597
rect 25222 29588 25228 29600
rect 25280 29588 25286 29640
rect 16540 29532 17540 29560
rect 16540 29520 16546 29532
rect 7466 29492 7472 29504
rect 7392 29464 7472 29492
rect 7466 29452 7472 29464
rect 7524 29452 7530 29504
rect 7742 29452 7748 29504
rect 7800 29452 7806 29504
rect 11238 29452 11244 29504
rect 11296 29492 11302 29504
rect 11793 29495 11851 29501
rect 11793 29492 11805 29495
rect 11296 29464 11805 29492
rect 11296 29452 11302 29464
rect 11793 29461 11805 29464
rect 11839 29461 11851 29495
rect 11793 29455 11851 29461
rect 17126 29452 17132 29504
rect 17184 29492 17190 29504
rect 17221 29495 17279 29501
rect 17221 29492 17233 29495
rect 17184 29464 17233 29492
rect 17184 29452 17190 29464
rect 17221 29461 17233 29464
rect 17267 29461 17279 29495
rect 17221 29455 17279 29461
rect 17310 29452 17316 29504
rect 17368 29452 17374 29504
rect 20438 29452 20444 29504
rect 20496 29492 20502 29504
rect 20625 29495 20683 29501
rect 20625 29492 20637 29495
rect 20496 29464 20637 29492
rect 20496 29452 20502 29464
rect 20625 29461 20637 29464
rect 20671 29461 20683 29495
rect 20625 29455 20683 29461
rect 1104 29402 29440 29424
rect 1104 29350 5151 29402
rect 5203 29350 5215 29402
rect 5267 29350 5279 29402
rect 5331 29350 5343 29402
rect 5395 29350 5407 29402
rect 5459 29350 12234 29402
rect 12286 29350 12298 29402
rect 12350 29350 12362 29402
rect 12414 29350 12426 29402
rect 12478 29350 12490 29402
rect 12542 29350 19317 29402
rect 19369 29350 19381 29402
rect 19433 29350 19445 29402
rect 19497 29350 19509 29402
rect 19561 29350 19573 29402
rect 19625 29350 26400 29402
rect 26452 29350 26464 29402
rect 26516 29350 26528 29402
rect 26580 29350 26592 29402
rect 26644 29350 26656 29402
rect 26708 29350 29440 29402
rect 1104 29328 29440 29350
rect 5902 29288 5908 29300
rect 3896 29260 5908 29288
rect 1578 29180 1584 29232
rect 1636 29220 1642 29232
rect 1673 29223 1731 29229
rect 1673 29220 1685 29223
rect 1636 29192 1685 29220
rect 1636 29180 1642 29192
rect 1673 29189 1685 29192
rect 1719 29189 1731 29223
rect 3050 29220 3056 29232
rect 2898 29192 3056 29220
rect 1673 29183 1731 29189
rect 3050 29180 3056 29192
rect 3108 29180 3114 29232
rect 3234 29180 3240 29232
rect 3292 29220 3298 29232
rect 3896 29220 3924 29260
rect 5902 29248 5908 29260
rect 5960 29248 5966 29300
rect 6641 29291 6699 29297
rect 6641 29257 6653 29291
rect 6687 29288 6699 29291
rect 6687 29260 7236 29288
rect 6687 29257 6699 29260
rect 6641 29251 6699 29257
rect 7098 29220 7104 29232
rect 3292 29192 4002 29220
rect 6840 29192 7104 29220
rect 3292 29180 3298 29192
rect 6840 29161 6868 29192
rect 7098 29180 7104 29192
rect 7156 29180 7162 29232
rect 7208 29229 7236 29260
rect 7466 29248 7472 29300
rect 7524 29288 7530 29300
rect 7524 29260 9076 29288
rect 7524 29248 7530 29260
rect 7193 29223 7251 29229
rect 7193 29189 7205 29223
rect 7239 29189 7251 29223
rect 7193 29183 7251 29189
rect 7282 29180 7288 29232
rect 7340 29220 7346 29232
rect 8941 29223 8999 29229
rect 8941 29220 8953 29223
rect 7340 29192 7682 29220
rect 8680 29192 8953 29220
rect 7340 29180 7346 29192
rect 6825 29155 6883 29161
rect 6825 29121 6837 29155
rect 6871 29121 6883 29155
rect 6825 29115 6883 29121
rect 1397 29087 1455 29093
rect 1397 29053 1409 29087
rect 1443 29084 1455 29087
rect 3237 29087 3295 29093
rect 3237 29084 3249 29087
rect 1443 29056 3249 29084
rect 1443 29053 1455 29056
rect 1397 29047 1455 29053
rect 3237 29053 3249 29056
rect 3283 29053 3295 29087
rect 3237 29047 3295 29053
rect 3142 28976 3148 29028
rect 3200 28976 3206 29028
rect 3252 28948 3280 29047
rect 3510 29044 3516 29096
rect 3568 29044 3574 29096
rect 5077 29087 5135 29093
rect 5077 29053 5089 29087
rect 5123 29084 5135 29087
rect 5626 29084 5632 29096
rect 5123 29056 5632 29084
rect 5123 29053 5135 29056
rect 5077 29047 5135 29053
rect 5626 29044 5632 29056
rect 5684 29084 5690 29096
rect 6178 29084 6184 29096
rect 5684 29056 6184 29084
rect 5684 29044 5690 29056
rect 6178 29044 6184 29056
rect 6236 29044 6242 29096
rect 6917 29087 6975 29093
rect 6917 29053 6929 29087
rect 6963 29053 6975 29087
rect 6917 29047 6975 29053
rect 5166 28976 5172 29028
rect 5224 29016 5230 29028
rect 5721 29019 5779 29025
rect 5721 29016 5733 29019
rect 5224 28988 5733 29016
rect 5224 28976 5230 28988
rect 5721 28985 5733 28988
rect 5767 28985 5779 29019
rect 5721 28979 5779 28985
rect 4154 28948 4160 28960
rect 3252 28920 4160 28948
rect 4154 28908 4160 28920
rect 4212 28908 4218 28960
rect 4982 28908 4988 28960
rect 5040 28908 5046 28960
rect 6932 28948 6960 29047
rect 7650 29044 7656 29096
rect 7708 29084 7714 29096
rect 8680 29093 8708 29192
rect 8941 29189 8953 29192
rect 8987 29189 8999 29223
rect 8941 29183 8999 29189
rect 9048 29161 9076 29260
rect 11238 29248 11244 29300
rect 11296 29248 11302 29300
rect 12618 29288 12624 29300
rect 11348 29260 12624 29288
rect 8761 29155 8819 29161
rect 8761 29121 8773 29155
rect 8807 29152 8819 29155
rect 9033 29155 9091 29161
rect 8807 29124 8984 29152
rect 8807 29121 8819 29124
rect 8761 29115 8819 29121
rect 8665 29087 8723 29093
rect 8665 29084 8677 29087
rect 7708 29056 8677 29084
rect 7708 29044 7714 29056
rect 8665 29053 8677 29056
rect 8711 29053 8723 29087
rect 8956 29084 8984 29124
rect 9033 29121 9045 29155
rect 9079 29121 9091 29155
rect 9033 29115 9091 29121
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29152 10747 29155
rect 11256 29152 11284 29248
rect 11348 29161 11376 29260
rect 12618 29248 12624 29260
rect 12676 29248 12682 29300
rect 13262 29248 13268 29300
rect 13320 29248 13326 29300
rect 16482 29248 16488 29300
rect 16540 29248 16546 29300
rect 17310 29288 17316 29300
rect 16960 29260 17316 29288
rect 11793 29223 11851 29229
rect 11793 29220 11805 29223
rect 11440 29192 11805 29220
rect 10735 29124 11284 29152
rect 11333 29155 11391 29161
rect 10735 29121 10747 29124
rect 10689 29115 10747 29121
rect 11333 29121 11345 29155
rect 11379 29121 11391 29155
rect 11333 29115 11391 29121
rect 9766 29084 9772 29096
rect 8956 29056 9772 29084
rect 8665 29047 8723 29053
rect 9766 29044 9772 29056
rect 9824 29044 9830 29096
rect 10781 29087 10839 29093
rect 10781 29053 10793 29087
rect 10827 29084 10839 29087
rect 11238 29084 11244 29096
rect 10827 29056 11244 29084
rect 10827 29053 10839 29056
rect 10781 29047 10839 29053
rect 11238 29044 11244 29056
rect 11296 29044 11302 29096
rect 11057 29019 11115 29025
rect 11057 28985 11069 29019
rect 11103 29016 11115 29019
rect 11440 29016 11468 29192
rect 11793 29189 11805 29192
rect 11839 29189 11851 29223
rect 11793 29183 11851 29189
rect 12250 29180 12256 29232
rect 12308 29180 12314 29232
rect 14274 29180 14280 29232
rect 14332 29180 14338 29232
rect 16666 29220 16672 29232
rect 16316 29192 16672 29220
rect 16206 29112 16212 29164
rect 16264 29112 16270 29164
rect 16316 29161 16344 29192
rect 16666 29180 16672 29192
rect 16724 29180 16730 29232
rect 16960 29229 16988 29260
rect 17310 29248 17316 29260
rect 17368 29248 17374 29300
rect 19150 29248 19156 29300
rect 19208 29248 19214 29300
rect 28534 29248 28540 29300
rect 28592 29248 28598 29300
rect 16945 29223 17003 29229
rect 16945 29189 16957 29223
rect 16991 29189 17003 29223
rect 16945 29183 17003 29189
rect 20165 29223 20223 29229
rect 20165 29189 20177 29223
rect 20211 29220 20223 29223
rect 20438 29220 20444 29232
rect 20211 29192 20444 29220
rect 20211 29189 20223 29192
rect 20165 29183 20223 29189
rect 20438 29180 20444 29192
rect 20496 29180 20502 29232
rect 24029 29223 24087 29229
rect 24029 29220 24041 29223
rect 22664 29192 24041 29220
rect 16301 29155 16359 29161
rect 16301 29121 16313 29155
rect 16347 29121 16359 29155
rect 18230 29152 18236 29164
rect 18078 29124 18236 29152
rect 16301 29115 16359 29121
rect 18230 29112 18236 29124
rect 18288 29112 18294 29164
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29121 19947 29155
rect 19889 29115 19947 29121
rect 11517 29087 11575 29093
rect 11517 29053 11529 29087
rect 11563 29084 11575 29087
rect 13446 29084 13452 29096
rect 11563 29056 13452 29084
rect 11563 29053 11575 29056
rect 11517 29047 11575 29053
rect 13446 29044 13452 29056
rect 13504 29044 13510 29096
rect 13722 29044 13728 29096
rect 13780 29044 13786 29096
rect 15289 29087 15347 29093
rect 15289 29053 15301 29087
rect 15335 29053 15347 29087
rect 15289 29047 15347 29053
rect 11103 28988 11468 29016
rect 11103 28985 11115 28988
rect 11057 28979 11115 28985
rect 7834 28948 7840 28960
rect 6932 28920 7840 28948
rect 7834 28908 7840 28920
rect 7892 28908 7898 28960
rect 8754 28908 8760 28960
rect 8812 28908 8818 28960
rect 11146 28908 11152 28960
rect 11204 28908 11210 28960
rect 15197 28951 15255 28957
rect 15197 28917 15209 28951
rect 15243 28948 15255 28951
rect 15304 28948 15332 29047
rect 16574 29044 16580 29096
rect 16632 29084 16638 29096
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 16632 29056 16681 29084
rect 16632 29044 16638 29056
rect 16669 29053 16681 29056
rect 16715 29053 16727 29087
rect 16669 29047 16727 29053
rect 18414 29044 18420 29096
rect 18472 29084 18478 29096
rect 18509 29087 18567 29093
rect 18509 29084 18521 29087
rect 18472 29056 18521 29084
rect 18472 29044 18478 29056
rect 18509 29053 18521 29056
rect 18555 29053 18567 29087
rect 18509 29047 18567 29053
rect 19904 28960 19932 29115
rect 21174 29112 21180 29164
rect 21232 29152 21238 29164
rect 22664 29161 22692 29192
rect 24029 29189 24041 29192
rect 24075 29189 24087 29223
rect 24029 29183 24087 29189
rect 22649 29155 22707 29161
rect 21232 29124 22094 29152
rect 21232 29112 21238 29124
rect 22066 29096 22094 29124
rect 22649 29121 22661 29155
rect 22695 29121 22707 29155
rect 22649 29115 22707 29121
rect 22830 29112 22836 29164
rect 22888 29152 22894 29164
rect 23109 29155 23167 29161
rect 23109 29152 23121 29155
rect 22888 29124 23121 29152
rect 22888 29112 22894 29124
rect 23109 29121 23121 29124
rect 23155 29121 23167 29155
rect 23109 29115 23167 29121
rect 23293 29155 23351 29161
rect 23293 29121 23305 29155
rect 23339 29121 23351 29155
rect 23293 29115 23351 29121
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29152 24455 29155
rect 28552 29152 28580 29248
rect 24443 29124 28580 29152
rect 24443 29121 24455 29124
rect 24397 29115 24455 29121
rect 22066 29056 22100 29096
rect 22094 29044 22100 29056
rect 22152 29044 22158 29096
rect 22186 29044 22192 29096
rect 22244 29084 22250 29096
rect 22557 29087 22615 29093
rect 22557 29084 22569 29087
rect 22244 29056 22569 29084
rect 22244 29044 22250 29056
rect 22557 29053 22569 29056
rect 22603 29084 22615 29087
rect 23308 29084 23336 29115
rect 22603 29056 23336 29084
rect 22603 29053 22615 29056
rect 22557 29047 22615 29053
rect 23382 29044 23388 29096
rect 23440 29044 23446 29096
rect 24486 29044 24492 29096
rect 24544 29084 24550 29096
rect 24673 29087 24731 29093
rect 24673 29084 24685 29087
rect 24544 29056 24685 29084
rect 24544 29044 24550 29056
rect 24673 29053 24685 29056
rect 24719 29053 24731 29087
rect 24673 29047 24731 29053
rect 21910 29016 21916 29028
rect 21652 28988 21916 29016
rect 15470 28948 15476 28960
rect 15243 28920 15476 28948
rect 15243 28917 15255 28920
rect 15197 28911 15255 28917
rect 15470 28908 15476 28920
rect 15528 28908 15534 28960
rect 15930 28908 15936 28960
rect 15988 28908 15994 28960
rect 18322 28908 18328 28960
rect 18380 28948 18386 28960
rect 18417 28951 18475 28957
rect 18417 28948 18429 28951
rect 18380 28920 18429 28948
rect 18380 28908 18386 28920
rect 18417 28917 18429 28920
rect 18463 28917 18475 28951
rect 18417 28911 18475 28917
rect 19886 28908 19892 28960
rect 19944 28948 19950 28960
rect 21266 28948 21272 28960
rect 19944 28920 21272 28948
rect 19944 28908 19950 28920
rect 21266 28908 21272 28920
rect 21324 28908 21330 28960
rect 21358 28908 21364 28960
rect 21416 28948 21422 28960
rect 21652 28957 21680 28988
rect 21910 28976 21916 28988
rect 21968 28976 21974 29028
rect 22370 29016 22376 29028
rect 22112 28988 22376 29016
rect 21637 28951 21695 28957
rect 21637 28948 21649 28951
rect 21416 28920 21649 28948
rect 21416 28908 21422 28920
rect 21637 28917 21649 28920
rect 21683 28917 21695 28951
rect 21637 28911 21695 28917
rect 21726 28908 21732 28960
rect 21784 28948 21790 28960
rect 22112 28948 22140 28988
rect 22370 28976 22376 28988
rect 22428 29016 22434 29028
rect 23400 29016 23428 29044
rect 22428 28988 23428 29016
rect 22428 28976 22434 28988
rect 21784 28920 22140 28948
rect 21784 28908 21790 28920
rect 23014 28908 23020 28960
rect 23072 28908 23078 28960
rect 23106 28908 23112 28960
rect 23164 28908 23170 28960
rect 1104 28858 29440 28880
rect 1104 28806 4491 28858
rect 4543 28806 4555 28858
rect 4607 28806 4619 28858
rect 4671 28806 4683 28858
rect 4735 28806 4747 28858
rect 4799 28806 11574 28858
rect 11626 28806 11638 28858
rect 11690 28806 11702 28858
rect 11754 28806 11766 28858
rect 11818 28806 11830 28858
rect 11882 28806 18657 28858
rect 18709 28806 18721 28858
rect 18773 28806 18785 28858
rect 18837 28806 18849 28858
rect 18901 28806 18913 28858
rect 18965 28806 25740 28858
rect 25792 28806 25804 28858
rect 25856 28806 25868 28858
rect 25920 28806 25932 28858
rect 25984 28806 25996 28858
rect 26048 28806 29440 28858
rect 1104 28784 29440 28806
rect 5166 28744 5172 28756
rect 3252 28716 5172 28744
rect 3252 28549 3280 28716
rect 5166 28704 5172 28716
rect 5224 28704 5230 28756
rect 5718 28704 5724 28756
rect 5776 28744 5782 28756
rect 6089 28747 6147 28753
rect 6089 28744 6101 28747
rect 5776 28716 6101 28744
rect 5776 28704 5782 28716
rect 6089 28713 6101 28716
rect 6135 28744 6147 28747
rect 6454 28744 6460 28756
rect 6135 28716 6460 28744
rect 6135 28713 6147 28716
rect 6089 28707 6147 28713
rect 6454 28704 6460 28716
rect 6512 28704 6518 28756
rect 7098 28704 7104 28756
rect 7156 28704 7162 28756
rect 7377 28747 7435 28753
rect 7377 28713 7389 28747
rect 7423 28744 7435 28747
rect 7742 28744 7748 28756
rect 7423 28716 7748 28744
rect 7423 28713 7435 28716
rect 7377 28707 7435 28713
rect 7742 28704 7748 28716
rect 7800 28704 7806 28756
rect 7837 28747 7895 28753
rect 7837 28713 7849 28747
rect 7883 28713 7895 28747
rect 7837 28707 7895 28713
rect 3896 28648 4384 28676
rect 3329 28611 3387 28617
rect 3329 28577 3341 28611
rect 3375 28608 3387 28611
rect 3375 28580 3832 28608
rect 3375 28577 3387 28580
rect 3329 28571 3387 28577
rect 3237 28543 3295 28549
rect 3237 28509 3249 28543
rect 3283 28509 3295 28543
rect 3237 28503 3295 28509
rect 3602 28364 3608 28416
rect 3660 28364 3666 28416
rect 3804 28404 3832 28580
rect 3896 28481 3924 28648
rect 4246 28608 4252 28620
rect 3988 28580 4252 28608
rect 3881 28475 3939 28481
rect 3881 28441 3893 28475
rect 3927 28441 3939 28475
rect 3881 28435 3939 28441
rect 3988 28404 4016 28580
rect 4246 28568 4252 28580
rect 4304 28568 4310 28620
rect 4356 28608 4384 28648
rect 6270 28636 6276 28688
rect 6328 28676 6334 28688
rect 6733 28679 6791 28685
rect 6733 28676 6745 28679
rect 6328 28648 6745 28676
rect 6328 28636 6334 28648
rect 6733 28645 6745 28648
rect 6779 28645 6791 28679
rect 7116 28676 7144 28704
rect 7561 28679 7619 28685
rect 7561 28676 7573 28679
rect 7116 28648 7573 28676
rect 6733 28639 6791 28645
rect 7561 28645 7573 28648
rect 7607 28645 7619 28679
rect 7852 28676 7880 28707
rect 9766 28704 9772 28756
rect 9824 28704 9830 28756
rect 10321 28747 10379 28753
rect 10321 28713 10333 28747
rect 10367 28744 10379 28747
rect 12437 28747 12495 28753
rect 12437 28744 12449 28747
rect 10367 28716 12449 28744
rect 10367 28713 10379 28716
rect 10321 28707 10379 28713
rect 12437 28713 12449 28716
rect 12483 28713 12495 28747
rect 12437 28707 12495 28713
rect 12618 28704 12624 28756
rect 12676 28704 12682 28756
rect 12894 28704 12900 28756
rect 12952 28744 12958 28756
rect 13449 28747 13507 28753
rect 13449 28744 13461 28747
rect 12952 28716 13461 28744
rect 12952 28704 12958 28716
rect 13449 28713 13461 28716
rect 13495 28713 13507 28747
rect 13449 28707 13507 28713
rect 13722 28704 13728 28756
rect 13780 28744 13786 28756
rect 14921 28747 14979 28753
rect 14921 28744 14933 28747
rect 13780 28716 14933 28744
rect 13780 28704 13786 28716
rect 14921 28713 14933 28716
rect 14967 28713 14979 28747
rect 14921 28707 14979 28713
rect 16117 28747 16175 28753
rect 16117 28713 16129 28747
rect 16163 28744 16175 28747
rect 16206 28744 16212 28756
rect 16163 28716 16212 28744
rect 16163 28713 16175 28716
rect 16117 28707 16175 28713
rect 16206 28704 16212 28716
rect 16264 28704 16270 28756
rect 16666 28704 16672 28756
rect 16724 28704 16730 28756
rect 20349 28747 20407 28753
rect 20349 28713 20361 28747
rect 20395 28713 20407 28747
rect 20349 28707 20407 28713
rect 20533 28747 20591 28753
rect 20533 28713 20545 28747
rect 20579 28744 20591 28747
rect 20806 28744 20812 28756
rect 20579 28716 20812 28744
rect 20579 28713 20591 28716
rect 20533 28707 20591 28713
rect 15841 28679 15899 28685
rect 15841 28676 15853 28679
rect 7852 28648 9168 28676
rect 7561 28639 7619 28645
rect 5074 28608 5080 28620
rect 4356 28580 5080 28608
rect 5074 28568 5080 28580
rect 5132 28608 5138 28620
rect 8205 28611 8263 28617
rect 5132 28580 6592 28608
rect 5132 28568 5138 28580
rect 4154 28500 4160 28552
rect 4212 28540 4218 28552
rect 4341 28543 4399 28549
rect 4341 28540 4353 28543
rect 4212 28512 4353 28540
rect 4212 28500 4218 28512
rect 4341 28509 4353 28512
rect 4387 28509 4399 28543
rect 5902 28540 5908 28552
rect 5750 28512 5908 28540
rect 4341 28503 4399 28509
rect 5902 28500 5908 28512
rect 5960 28500 5966 28552
rect 6454 28500 6460 28552
rect 6512 28500 6518 28552
rect 6564 28549 6592 28580
rect 8205 28577 8217 28611
rect 8251 28608 8263 28611
rect 8754 28608 8760 28620
rect 8251 28580 8760 28608
rect 8251 28577 8263 28580
rect 8205 28571 8263 28577
rect 8754 28568 8760 28580
rect 8812 28568 8818 28620
rect 9140 28617 9168 28648
rect 13188 28648 15853 28676
rect 9125 28611 9183 28617
rect 9125 28577 9137 28611
rect 9171 28608 9183 28611
rect 9398 28608 9404 28620
rect 9171 28580 9404 28608
rect 9171 28577 9183 28580
rect 9125 28571 9183 28577
rect 9398 28568 9404 28580
rect 9456 28568 9462 28620
rect 10689 28611 10747 28617
rect 10689 28577 10701 28611
rect 10735 28608 10747 28611
rect 11146 28608 11152 28620
rect 10735 28580 11152 28608
rect 10735 28577 10747 28580
rect 10689 28571 10747 28577
rect 11146 28568 11152 28580
rect 11204 28568 11210 28620
rect 11238 28568 11244 28620
rect 11296 28608 11302 28620
rect 11296 28580 12496 28608
rect 11296 28568 11302 28580
rect 6549 28543 6607 28549
rect 6549 28509 6561 28543
rect 6595 28509 6607 28543
rect 6549 28503 6607 28509
rect 6917 28543 6975 28549
rect 6917 28509 6929 28543
rect 6963 28540 6975 28543
rect 7006 28540 7012 28552
rect 6963 28512 7012 28540
rect 6963 28509 6975 28512
rect 6917 28503 6975 28509
rect 7006 28500 7012 28512
rect 7064 28500 7070 28552
rect 7101 28543 7159 28549
rect 7101 28509 7113 28543
rect 7147 28509 7159 28543
rect 7101 28503 7159 28509
rect 10413 28543 10471 28549
rect 10413 28509 10425 28543
rect 10459 28509 10471 28543
rect 12158 28540 12164 28552
rect 11822 28512 12164 28540
rect 10413 28503 10471 28509
rect 4065 28475 4123 28481
rect 4065 28441 4077 28475
rect 4111 28472 4123 28475
rect 4617 28475 4675 28481
rect 4111 28444 4568 28472
rect 4111 28441 4123 28444
rect 4065 28435 4123 28441
rect 3804 28376 4016 28404
rect 4249 28407 4307 28413
rect 4249 28373 4261 28407
rect 4295 28404 4307 28407
rect 4338 28404 4344 28416
rect 4295 28376 4344 28404
rect 4295 28373 4307 28376
rect 4249 28367 4307 28373
rect 4338 28364 4344 28376
rect 4396 28364 4402 28416
rect 4540 28404 4568 28444
rect 4617 28441 4629 28475
rect 4663 28472 4675 28475
rect 4890 28472 4896 28484
rect 4663 28444 4896 28472
rect 4663 28441 4675 28444
rect 4617 28435 4675 28441
rect 4890 28432 4896 28444
rect 4948 28432 4954 28484
rect 6178 28432 6184 28484
rect 6236 28472 6242 28484
rect 6822 28472 6828 28484
rect 6236 28444 6828 28472
rect 6236 28432 6242 28444
rect 6822 28432 6828 28444
rect 6880 28432 6886 28484
rect 4982 28404 4988 28416
rect 4540 28376 4988 28404
rect 4982 28364 4988 28376
rect 5040 28364 5046 28416
rect 6362 28364 6368 28416
rect 6420 28364 6426 28416
rect 7006 28364 7012 28416
rect 7064 28364 7070 28416
rect 7116 28404 7144 28503
rect 7190 28432 7196 28484
rect 7248 28432 7254 28484
rect 7409 28475 7467 28481
rect 7409 28441 7421 28475
rect 7455 28472 7467 28475
rect 7558 28472 7564 28484
rect 7455 28444 7564 28472
rect 7455 28441 7467 28444
rect 7409 28435 7467 28441
rect 7558 28432 7564 28444
rect 7616 28432 7622 28484
rect 7650 28432 7656 28484
rect 7708 28432 7714 28484
rect 7742 28432 7748 28484
rect 7800 28472 7806 28484
rect 7853 28475 7911 28481
rect 7853 28472 7865 28475
rect 7800 28444 7865 28472
rect 7800 28432 7806 28444
rect 7853 28441 7865 28444
rect 7899 28441 7911 28475
rect 7853 28435 7911 28441
rect 8754 28432 8760 28484
rect 8812 28432 8818 28484
rect 9950 28432 9956 28484
rect 10008 28432 10014 28484
rect 10137 28475 10195 28481
rect 10137 28441 10149 28475
rect 10183 28472 10195 28475
rect 10428 28472 10456 28503
rect 12158 28500 12164 28512
rect 12216 28500 12222 28552
rect 12468 28515 12496 28580
rect 13188 28549 13216 28648
rect 15841 28645 15853 28648
rect 15887 28676 15899 28679
rect 18414 28676 18420 28688
rect 15887 28648 16068 28676
rect 15887 28645 15899 28648
rect 15841 28639 15899 28645
rect 13630 28568 13636 28620
rect 13688 28568 13694 28620
rect 15381 28611 15439 28617
rect 15381 28577 15393 28611
rect 15427 28608 15439 28611
rect 15930 28608 15936 28620
rect 15427 28580 15936 28608
rect 15427 28577 15439 28580
rect 15381 28571 15439 28577
rect 15930 28568 15936 28580
rect 15988 28568 15994 28620
rect 13173 28543 13231 28549
rect 12468 28509 12541 28515
rect 10183 28444 10364 28472
rect 10428 28444 10824 28472
rect 10183 28441 10195 28444
rect 10137 28435 10195 28441
rect 10336 28416 10364 28444
rect 10796 28416 10824 28444
rect 12066 28432 12072 28484
rect 12124 28472 12130 28484
rect 12253 28475 12311 28481
rect 12468 28478 12495 28509
rect 12253 28472 12265 28475
rect 12124 28444 12265 28472
rect 12124 28432 12130 28444
rect 12253 28441 12265 28444
rect 12299 28441 12311 28475
rect 12483 28475 12495 28478
rect 12529 28475 12541 28509
rect 13173 28509 13185 28543
rect 13219 28509 13231 28543
rect 13173 28503 13231 28509
rect 13357 28543 13415 28549
rect 13357 28509 13369 28543
rect 13403 28540 13415 28543
rect 13538 28540 13544 28552
rect 13403 28512 13544 28540
rect 13403 28509 13415 28512
rect 13357 28503 13415 28509
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 13725 28543 13783 28549
rect 13725 28509 13737 28543
rect 13771 28540 13783 28543
rect 13998 28540 14004 28552
rect 13771 28512 14004 28540
rect 13771 28509 13783 28512
rect 13725 28503 13783 28509
rect 13998 28500 14004 28512
rect 14056 28500 14062 28552
rect 14185 28543 14243 28549
rect 14185 28509 14197 28543
rect 14231 28540 14243 28543
rect 14458 28540 14464 28552
rect 14231 28512 14464 28540
rect 14231 28509 14243 28512
rect 14185 28503 14243 28509
rect 14458 28500 14464 28512
rect 14516 28500 14522 28552
rect 15105 28543 15163 28549
rect 15105 28509 15117 28543
rect 15151 28509 15163 28543
rect 15105 28503 15163 28509
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28509 15347 28543
rect 15289 28503 15347 28509
rect 12483 28469 12541 28475
rect 13449 28475 13507 28481
rect 12253 28435 12311 28441
rect 13449 28441 13461 28475
rect 13495 28472 13507 28475
rect 13630 28472 13636 28484
rect 13495 28444 13636 28472
rect 13495 28441 13507 28444
rect 13449 28435 13507 28441
rect 13630 28432 13636 28444
rect 13688 28432 13694 28484
rect 15120 28472 15148 28503
rect 13832 28444 15148 28472
rect 15304 28472 15332 28503
rect 15470 28500 15476 28552
rect 15528 28500 15534 28552
rect 16040 28549 16068 28648
rect 18156 28648 18420 28676
rect 17037 28611 17095 28617
rect 17037 28577 17049 28611
rect 17083 28608 17095 28611
rect 17126 28608 17132 28620
rect 17083 28580 17132 28608
rect 17083 28577 17095 28580
rect 17037 28571 17095 28577
rect 17126 28568 17132 28580
rect 17184 28568 17190 28620
rect 17770 28568 17776 28620
rect 17828 28608 17834 28620
rect 18156 28608 18184 28648
rect 18414 28636 18420 28648
rect 18472 28676 18478 28688
rect 18509 28679 18567 28685
rect 18509 28676 18521 28679
rect 18472 28648 18521 28676
rect 18472 28636 18478 28648
rect 18509 28645 18521 28648
rect 18555 28645 18567 28679
rect 20364 28676 20392 28707
rect 20806 28704 20812 28716
rect 20864 28704 20870 28756
rect 20916 28716 21496 28744
rect 20916 28676 20944 28716
rect 20364 28648 20944 28676
rect 21468 28676 21496 28716
rect 21726 28704 21732 28756
rect 21784 28704 21790 28756
rect 22002 28704 22008 28756
rect 22060 28704 22066 28756
rect 22094 28704 22100 28756
rect 22152 28744 22158 28756
rect 22152 28716 23888 28744
rect 22152 28704 22158 28716
rect 22189 28679 22247 28685
rect 22189 28676 22201 28679
rect 21468 28648 22201 28676
rect 18509 28639 18567 28645
rect 22189 28645 22201 28648
rect 22235 28645 22247 28679
rect 22189 28639 22247 28645
rect 17828 28580 18184 28608
rect 17828 28568 17834 28580
rect 18230 28568 18236 28620
rect 18288 28568 18294 28620
rect 19521 28611 19579 28617
rect 19521 28577 19533 28611
rect 19567 28608 19579 28611
rect 19567 28580 19840 28608
rect 19567 28577 19579 28580
rect 19521 28571 19579 28577
rect 15657 28543 15715 28549
rect 15657 28509 15669 28543
rect 15703 28509 15715 28543
rect 15657 28503 15715 28509
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28509 16083 28543
rect 16025 28503 16083 28509
rect 16209 28543 16267 28549
rect 16209 28509 16221 28543
rect 16255 28540 16267 28543
rect 16482 28540 16488 28552
rect 16255 28512 16488 28540
rect 16255 28509 16267 28512
rect 16209 28503 16267 28509
rect 15672 28472 15700 28503
rect 15304 28444 15700 28472
rect 16040 28472 16068 28503
rect 16482 28500 16488 28512
rect 16540 28500 16546 28552
rect 16574 28500 16580 28552
rect 16632 28540 16638 28552
rect 16761 28543 16819 28549
rect 16761 28540 16773 28543
rect 16632 28512 16773 28540
rect 16632 28500 16638 28512
rect 16761 28509 16773 28512
rect 16807 28509 16819 28543
rect 18248 28540 18276 28568
rect 19812 28552 19840 28580
rect 21266 28568 21272 28620
rect 21324 28608 21330 28620
rect 22741 28611 22799 28617
rect 21324 28580 22508 28608
rect 21324 28568 21330 28580
rect 18170 28512 18276 28540
rect 19245 28543 19303 28549
rect 16761 28503 16819 28509
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 16298 28472 16304 28484
rect 16040 28444 16304 28472
rect 8021 28407 8079 28413
rect 8021 28404 8033 28407
rect 7116 28376 8033 28404
rect 8021 28373 8033 28376
rect 8067 28404 8079 28407
rect 8570 28404 8576 28416
rect 8067 28376 8576 28404
rect 8067 28373 8079 28376
rect 8021 28367 8079 28373
rect 8570 28364 8576 28376
rect 8628 28364 8634 28416
rect 10318 28364 10324 28416
rect 10376 28364 10382 28416
rect 10778 28364 10784 28416
rect 10836 28364 10842 28416
rect 11698 28364 11704 28416
rect 11756 28404 11762 28416
rect 12161 28407 12219 28413
rect 12161 28404 12173 28407
rect 11756 28376 12173 28404
rect 11756 28364 11762 28376
rect 12161 28373 12173 28376
rect 12207 28373 12219 28407
rect 12161 28367 12219 28373
rect 13265 28407 13323 28413
rect 13265 28373 13277 28407
rect 13311 28404 13323 28407
rect 13832 28404 13860 28444
rect 15304 28416 15332 28444
rect 16298 28432 16304 28444
rect 16356 28432 16362 28484
rect 19260 28472 19288 28503
rect 19334 28500 19340 28552
rect 19392 28500 19398 28552
rect 19794 28500 19800 28552
rect 19852 28540 19858 28552
rect 19852 28512 20208 28540
rect 19852 28500 19858 28512
rect 20180 28481 20208 28512
rect 20806 28500 20812 28552
rect 20864 28500 20870 28552
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28509 20959 28543
rect 20901 28503 20959 28509
rect 20993 28543 21051 28549
rect 20993 28509 21005 28543
rect 21039 28509 21051 28543
rect 20993 28503 21051 28509
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28540 21143 28543
rect 21358 28540 21364 28552
rect 21131 28512 21364 28540
rect 21131 28509 21143 28512
rect 21085 28503 21143 28509
rect 20165 28475 20223 28481
rect 19260 28444 19840 28472
rect 13311 28376 13860 28404
rect 13311 28373 13323 28376
rect 13265 28367 13323 28373
rect 13906 28364 13912 28416
rect 13964 28364 13970 28416
rect 14734 28364 14740 28416
rect 14792 28364 14798 28416
rect 15286 28364 15292 28416
rect 15344 28364 15350 28416
rect 16316 28404 16344 28432
rect 18046 28404 18052 28416
rect 16316 28376 18052 28404
rect 18046 28364 18052 28376
rect 18104 28364 18110 28416
rect 19521 28407 19579 28413
rect 19521 28373 19533 28407
rect 19567 28404 19579 28407
rect 19702 28404 19708 28416
rect 19567 28376 19708 28404
rect 19567 28373 19579 28376
rect 19521 28367 19579 28373
rect 19702 28364 19708 28376
rect 19760 28364 19766 28416
rect 19812 28404 19840 28444
rect 20165 28441 20177 28475
rect 20211 28441 20223 28475
rect 20165 28435 20223 28441
rect 20381 28475 20439 28481
rect 20381 28441 20393 28475
rect 20427 28472 20439 28475
rect 20427 28444 20668 28472
rect 20427 28441 20439 28444
rect 20381 28435 20439 28441
rect 20254 28404 20260 28416
rect 19812 28376 20260 28404
rect 20254 28364 20260 28376
rect 20312 28364 20318 28416
rect 20640 28413 20668 28444
rect 20625 28407 20683 28413
rect 20625 28373 20637 28407
rect 20671 28373 20683 28407
rect 20916 28404 20944 28503
rect 21008 28472 21036 28503
rect 21358 28500 21364 28512
rect 21416 28500 21422 28552
rect 21453 28543 21511 28549
rect 21453 28509 21465 28543
rect 21499 28542 21511 28543
rect 21499 28540 21588 28542
rect 21634 28540 21640 28552
rect 21499 28514 21640 28540
rect 21499 28509 21511 28514
rect 21560 28512 21640 28514
rect 21453 28503 21511 28509
rect 21634 28500 21640 28512
rect 21692 28500 21698 28552
rect 21821 28543 21879 28549
rect 21821 28542 21833 28543
rect 21744 28514 21833 28542
rect 21744 28472 21772 28514
rect 21821 28509 21833 28514
rect 21867 28509 21879 28543
rect 21821 28503 21879 28509
rect 21910 28500 21916 28552
rect 21968 28540 21974 28552
rect 22281 28543 22339 28549
rect 22281 28540 22293 28543
rect 21968 28512 22293 28540
rect 21968 28500 21974 28512
rect 22281 28509 22293 28512
rect 22327 28509 22339 28543
rect 22281 28503 22339 28509
rect 22370 28500 22376 28552
rect 22428 28500 22434 28552
rect 22480 28549 22508 28580
rect 22741 28577 22753 28611
rect 22787 28608 22799 28611
rect 23106 28608 23112 28620
rect 22787 28580 23112 28608
rect 22787 28577 22799 28580
rect 22741 28571 22799 28577
rect 23106 28568 23112 28580
rect 23164 28568 23170 28620
rect 23860 28608 23888 28716
rect 24210 28636 24216 28688
rect 24268 28676 24274 28688
rect 24268 28648 25268 28676
rect 24268 28636 24274 28648
rect 25240 28617 25268 28648
rect 24765 28611 24823 28617
rect 24765 28608 24777 28611
rect 23860 28580 24777 28608
rect 22465 28543 22523 28549
rect 22465 28509 22477 28543
rect 22511 28509 22523 28543
rect 23860 28526 23888 28580
rect 24765 28577 24777 28580
rect 24811 28577 24823 28611
rect 24765 28571 24823 28577
rect 25225 28611 25283 28617
rect 25225 28577 25237 28611
rect 25271 28577 25283 28611
rect 25225 28571 25283 28577
rect 22465 28503 22523 28509
rect 22002 28472 22008 28484
rect 21008 28444 22008 28472
rect 22002 28432 22008 28444
rect 22060 28432 22066 28484
rect 22097 28475 22155 28481
rect 22097 28441 22109 28475
rect 22143 28472 22155 28475
rect 22186 28472 22192 28484
rect 22143 28444 22192 28472
rect 22143 28441 22155 28444
rect 22097 28435 22155 28441
rect 22186 28432 22192 28444
rect 22244 28432 22250 28484
rect 22480 28472 22508 28503
rect 24302 28500 24308 28552
rect 24360 28540 24366 28552
rect 24489 28543 24547 28549
rect 24489 28540 24501 28543
rect 24360 28512 24501 28540
rect 24360 28500 24366 28512
rect 24489 28509 24501 28512
rect 24535 28509 24547 28543
rect 24489 28503 24547 28509
rect 22480 28444 22600 28472
rect 21726 28404 21732 28416
rect 20916 28376 21732 28404
rect 20625 28367 20683 28373
rect 21726 28364 21732 28376
rect 21784 28364 21790 28416
rect 22572 28404 22600 28444
rect 22738 28432 22744 28484
rect 22796 28472 22802 28484
rect 22796 28444 23152 28472
rect 22796 28432 22802 28444
rect 22922 28404 22928 28416
rect 22572 28376 22928 28404
rect 22922 28364 22928 28376
rect 22980 28364 22986 28416
rect 23124 28404 23152 28444
rect 24210 28404 24216 28416
rect 23124 28376 24216 28404
rect 24210 28364 24216 28376
rect 24268 28364 24274 28416
rect 24394 28364 24400 28416
rect 24452 28404 24458 28416
rect 25869 28407 25927 28413
rect 25869 28404 25881 28407
rect 24452 28376 25881 28404
rect 24452 28364 24458 28376
rect 25869 28373 25881 28376
rect 25915 28373 25927 28407
rect 25869 28367 25927 28373
rect 1104 28314 29440 28336
rect 1104 28262 5151 28314
rect 5203 28262 5215 28314
rect 5267 28262 5279 28314
rect 5331 28262 5343 28314
rect 5395 28262 5407 28314
rect 5459 28262 12234 28314
rect 12286 28262 12298 28314
rect 12350 28262 12362 28314
rect 12414 28262 12426 28314
rect 12478 28262 12490 28314
rect 12542 28262 19317 28314
rect 19369 28262 19381 28314
rect 19433 28262 19445 28314
rect 19497 28262 19509 28314
rect 19561 28262 19573 28314
rect 19625 28262 26400 28314
rect 26452 28262 26464 28314
rect 26516 28262 26528 28314
rect 26580 28262 26592 28314
rect 26644 28262 26656 28314
rect 26708 28262 29440 28314
rect 1104 28240 29440 28262
rect 3421 28203 3479 28209
rect 3421 28169 3433 28203
rect 3467 28200 3479 28203
rect 3510 28200 3516 28212
rect 3467 28172 3516 28200
rect 3467 28169 3479 28172
rect 3421 28163 3479 28169
rect 3510 28160 3516 28172
rect 3568 28160 3574 28212
rect 3602 28160 3608 28212
rect 3660 28200 3666 28212
rect 5445 28203 5503 28209
rect 3660 28172 4016 28200
rect 3660 28160 3666 28172
rect 3988 28141 4016 28172
rect 5445 28169 5457 28203
rect 5491 28169 5503 28203
rect 5445 28163 5503 28169
rect 3973 28135 4031 28141
rect 3973 28101 3985 28135
rect 4019 28101 4031 28135
rect 5460 28132 5488 28163
rect 5994 28160 6000 28212
rect 6052 28160 6058 28212
rect 6178 28160 6184 28212
rect 6236 28160 6242 28212
rect 7285 28203 7343 28209
rect 7285 28169 7297 28203
rect 7331 28200 7343 28203
rect 7558 28200 7564 28212
rect 7331 28172 7564 28200
rect 7331 28169 7343 28172
rect 7285 28163 7343 28169
rect 7558 28160 7564 28172
rect 7616 28160 7622 28212
rect 8570 28160 8576 28212
rect 8628 28200 8634 28212
rect 8628 28172 9260 28200
rect 8628 28160 8634 28172
rect 6196 28132 6224 28160
rect 7466 28132 7472 28144
rect 5460 28104 6224 28132
rect 6288 28104 7472 28132
rect 3973 28095 4031 28101
rect 3602 28024 3608 28076
rect 3660 28024 3666 28076
rect 5626 28064 5632 28076
rect 5106 28036 5632 28064
rect 5626 28024 5632 28036
rect 5684 28064 5690 28076
rect 5902 28064 5908 28076
rect 5684 28036 5908 28064
rect 5684 28024 5690 28036
rect 5902 28024 5908 28036
rect 5960 28024 5966 28076
rect 6288 28008 6316 28104
rect 6365 28067 6423 28073
rect 6365 28033 6377 28067
rect 6411 28033 6423 28067
rect 6365 28027 6423 28033
rect 3697 27999 3755 28005
rect 3697 27965 3709 27999
rect 3743 27965 3755 27999
rect 3697 27959 3755 27965
rect 5537 27999 5595 28005
rect 5537 27965 5549 27999
rect 5583 27996 5595 27999
rect 6270 27996 6276 28008
rect 5583 27968 6276 27996
rect 5583 27965 5595 27968
rect 5537 27959 5595 27965
rect 3712 27860 3740 27959
rect 6270 27956 6276 27968
rect 6328 27956 6334 28008
rect 5810 27888 5816 27940
rect 5868 27888 5874 27940
rect 6380 27928 6408 28027
rect 6454 28024 6460 28076
rect 6512 28064 6518 28076
rect 6641 28067 6699 28073
rect 6641 28064 6653 28067
rect 6512 28036 6653 28064
rect 6512 28024 6518 28036
rect 6641 28033 6653 28036
rect 6687 28033 6699 28067
rect 6641 28027 6699 28033
rect 6822 28024 6828 28076
rect 6880 28024 6886 28076
rect 7006 28024 7012 28076
rect 7064 28024 7070 28076
rect 7116 28073 7144 28104
rect 7466 28092 7472 28104
rect 7524 28092 7530 28144
rect 7834 28132 7840 28144
rect 7668 28104 7840 28132
rect 7101 28067 7159 28073
rect 7101 28033 7113 28067
rect 7147 28033 7159 28067
rect 7101 28027 7159 28033
rect 7190 28024 7196 28076
rect 7248 28064 7254 28076
rect 7285 28067 7343 28073
rect 7285 28064 7297 28067
rect 7248 28036 7297 28064
rect 7248 28024 7254 28036
rect 7285 28033 7297 28036
rect 7331 28064 7343 28067
rect 7558 28064 7564 28076
rect 7331 28036 7564 28064
rect 7331 28033 7343 28036
rect 7285 28027 7343 28033
rect 7558 28024 7564 28036
rect 7616 28024 7622 28076
rect 7668 28073 7696 28104
rect 7834 28092 7840 28104
rect 7892 28092 7898 28144
rect 7653 28067 7711 28073
rect 7653 28033 7665 28067
rect 7699 28033 7711 28067
rect 7653 28027 7711 28033
rect 9030 28024 9036 28076
rect 9088 28024 9094 28076
rect 9232 28064 9260 28172
rect 9398 28160 9404 28212
rect 9456 28160 9462 28212
rect 9861 28203 9919 28209
rect 9861 28169 9873 28203
rect 9907 28200 9919 28203
rect 9950 28200 9956 28212
rect 9907 28172 9956 28200
rect 9907 28169 9919 28172
rect 9861 28163 9919 28169
rect 9950 28160 9956 28172
rect 10008 28200 10014 28212
rect 10965 28203 11023 28209
rect 10008 28172 10916 28200
rect 10008 28160 10014 28172
rect 9416 28132 9444 28160
rect 9416 28104 10824 28132
rect 9306 28064 9312 28076
rect 9232 28036 9312 28064
rect 9306 28024 9312 28036
rect 9364 28064 9370 28076
rect 10796 28073 10824 28104
rect 9677 28067 9735 28073
rect 9677 28064 9689 28067
rect 9364 28036 9689 28064
rect 9364 28024 9370 28036
rect 9677 28033 9689 28036
rect 9723 28033 9735 28067
rect 10413 28067 10471 28073
rect 10413 28064 10425 28067
rect 9677 28027 9735 28033
rect 9784 28036 10425 28064
rect 7024 27996 7052 28024
rect 9784 28008 9812 28036
rect 10413 28033 10425 28036
rect 10459 28033 10471 28067
rect 10413 28027 10471 28033
rect 10781 28067 10839 28073
rect 10781 28033 10793 28067
rect 10827 28033 10839 28067
rect 10888 28064 10916 28172
rect 10965 28169 10977 28203
rect 11011 28200 11023 28203
rect 12894 28200 12900 28212
rect 11011 28172 12900 28200
rect 11011 28169 11023 28172
rect 10965 28163 11023 28169
rect 12894 28160 12900 28172
rect 12952 28160 12958 28212
rect 13357 28203 13415 28209
rect 13357 28169 13369 28203
rect 13403 28200 13415 28203
rect 15286 28200 15292 28212
rect 13403 28172 15292 28200
rect 13403 28169 13415 28172
rect 13357 28163 13415 28169
rect 15286 28160 15292 28172
rect 15344 28160 15350 28212
rect 16298 28160 16304 28212
rect 16356 28200 16362 28212
rect 17037 28203 17095 28209
rect 17037 28200 17049 28203
rect 16356 28172 17049 28200
rect 16356 28160 16362 28172
rect 17037 28169 17049 28172
rect 17083 28169 17095 28203
rect 17770 28200 17776 28212
rect 17037 28163 17095 28169
rect 17604 28172 17776 28200
rect 11330 28092 11336 28144
rect 11388 28132 11394 28144
rect 11517 28135 11575 28141
rect 11517 28132 11529 28135
rect 11388 28104 11529 28132
rect 11388 28092 11394 28104
rect 11517 28101 11529 28104
rect 11563 28101 11575 28135
rect 11517 28095 11575 28101
rect 11698 28092 11704 28144
rect 11756 28092 11762 28144
rect 11793 28135 11851 28141
rect 11793 28101 11805 28135
rect 11839 28132 11851 28135
rect 12989 28135 13047 28141
rect 11839 28104 12296 28132
rect 11839 28101 11851 28104
rect 11793 28095 11851 28101
rect 11057 28067 11115 28073
rect 11057 28064 11069 28067
rect 10888 28036 11069 28064
rect 10781 28027 10839 28033
rect 11057 28033 11069 28036
rect 11103 28033 11115 28067
rect 11057 28027 11115 28033
rect 11241 28067 11299 28073
rect 11241 28033 11253 28067
rect 11287 28064 11299 28067
rect 11422 28064 11428 28076
rect 11287 28036 11428 28064
rect 11287 28033 11299 28036
rect 11241 28027 11299 28033
rect 7929 27999 7987 28005
rect 7929 27996 7941 27999
rect 7024 27968 7941 27996
rect 7929 27965 7941 27968
rect 7975 27965 7987 27999
rect 7929 27959 7987 27965
rect 9493 27999 9551 28005
rect 9493 27965 9505 27999
rect 9539 27996 9551 27999
rect 9766 27996 9772 28008
rect 9539 27968 9772 27996
rect 9539 27965 9551 27968
rect 9493 27959 9551 27965
rect 9766 27956 9772 27968
rect 9824 27956 9830 28008
rect 10318 27956 10324 28008
rect 10376 27956 10382 28008
rect 11072 27996 11100 28027
rect 11422 28024 11428 28036
rect 11480 28064 11486 28076
rect 11716 28064 11744 28092
rect 12268 28076 12296 28104
rect 12989 28101 13001 28135
rect 13035 28132 13047 28135
rect 13078 28132 13084 28144
rect 13035 28104 13084 28132
rect 13035 28101 13047 28104
rect 12989 28095 13047 28101
rect 13078 28092 13084 28104
rect 13136 28092 13142 28144
rect 13189 28135 13247 28141
rect 13189 28132 13201 28135
rect 13188 28101 13201 28132
rect 13235 28101 13247 28135
rect 13188 28095 13247 28101
rect 11480 28036 11744 28064
rect 11885 28067 11943 28073
rect 11480 28024 11486 28036
rect 11885 28033 11897 28067
rect 11931 28033 11943 28067
rect 11885 28027 11943 28033
rect 11900 27996 11928 28027
rect 12250 28024 12256 28076
rect 12308 28024 12314 28076
rect 12710 28024 12716 28076
rect 12768 28064 12774 28076
rect 13188 28064 13216 28095
rect 14274 28092 14280 28144
rect 14332 28092 14338 28144
rect 15304 28132 15332 28160
rect 16669 28135 16727 28141
rect 15304 28104 16252 28132
rect 12768 28036 13216 28064
rect 12768 28024 12774 28036
rect 13446 28024 13452 28076
rect 13504 28024 13510 28076
rect 16224 28073 16252 28104
rect 16669 28101 16681 28135
rect 16715 28132 16727 28135
rect 17604 28132 17632 28172
rect 17770 28160 17776 28172
rect 17828 28160 17834 28212
rect 17862 28160 17868 28212
rect 17920 28200 17926 28212
rect 20717 28203 20775 28209
rect 20717 28200 20729 28203
rect 17920 28172 20729 28200
rect 17920 28160 17926 28172
rect 20717 28169 20729 28172
rect 20763 28169 20775 28203
rect 20717 28163 20775 28169
rect 16715 28104 17632 28132
rect 16715 28101 16727 28104
rect 16669 28095 16727 28101
rect 20732 28076 20760 28163
rect 22094 28160 22100 28212
rect 22152 28200 22158 28212
rect 22738 28200 22744 28212
rect 22152 28172 22744 28200
rect 22152 28160 22158 28172
rect 22738 28160 22744 28172
rect 22796 28160 22802 28212
rect 23014 28160 23020 28212
rect 23072 28160 23078 28212
rect 23382 28160 23388 28212
rect 23440 28200 23446 28212
rect 24673 28203 24731 28209
rect 24673 28200 24685 28203
rect 23440 28172 24685 28200
rect 23440 28160 23446 28172
rect 24673 28169 24685 28172
rect 24719 28169 24731 28203
rect 24673 28163 24731 28169
rect 23032 28132 23060 28160
rect 23201 28135 23259 28141
rect 23201 28132 23213 28135
rect 23032 28104 23213 28132
rect 23201 28101 23213 28104
rect 23247 28101 23259 28135
rect 23201 28095 23259 28101
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28064 15991 28067
rect 16025 28067 16083 28073
rect 16025 28064 16037 28067
rect 15979 28036 16037 28064
rect 15979 28033 15991 28036
rect 15933 28027 15991 28033
rect 16025 28033 16037 28036
rect 16071 28033 16083 28067
rect 16025 28027 16083 28033
rect 16209 28067 16267 28073
rect 16209 28033 16221 28067
rect 16255 28033 16267 28067
rect 16209 28027 16267 28033
rect 16482 28024 16488 28076
rect 16540 28064 16546 28076
rect 16853 28067 16911 28073
rect 16853 28064 16865 28067
rect 16540 28036 16865 28064
rect 16540 28024 16546 28036
rect 16853 28033 16865 28036
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 16945 28067 17003 28073
rect 16945 28033 16957 28067
rect 16991 28033 17003 28067
rect 16945 28027 17003 28033
rect 17313 28067 17371 28073
rect 17313 28033 17325 28067
rect 17359 28064 17371 28067
rect 17678 28064 17684 28076
rect 17359 28036 17684 28064
rect 17359 28033 17371 28036
rect 17313 28027 17371 28033
rect 11072 27968 11928 27996
rect 13725 27999 13783 28005
rect 13725 27965 13737 27999
rect 13771 27996 13783 27999
rect 13771 27968 14964 27996
rect 13771 27965 13783 27968
rect 13725 27959 13783 27965
rect 7190 27928 7196 27940
rect 6380 27900 7196 27928
rect 7190 27888 7196 27900
rect 7248 27888 7254 27940
rect 10336 27928 10364 27956
rect 11422 27928 11428 27940
rect 10336 27900 11428 27928
rect 11422 27888 11428 27900
rect 11480 27888 11486 27940
rect 14936 27928 14964 27968
rect 15286 27956 15292 28008
rect 15344 27956 15350 28008
rect 16025 27931 16083 27937
rect 16025 27928 16037 27931
rect 13188 27900 13584 27928
rect 14936 27900 16037 27928
rect 4154 27860 4160 27872
rect 3712 27832 4160 27860
rect 4154 27820 4160 27832
rect 4212 27820 4218 27872
rect 6362 27820 6368 27872
rect 6420 27860 6426 27872
rect 6457 27863 6515 27869
rect 6457 27860 6469 27863
rect 6420 27832 6469 27860
rect 6420 27820 6426 27832
rect 6457 27829 6469 27832
rect 6503 27829 6515 27863
rect 6457 27823 6515 27829
rect 6546 27820 6552 27872
rect 6604 27860 6610 27872
rect 7009 27863 7067 27869
rect 7009 27860 7021 27863
rect 6604 27832 7021 27860
rect 6604 27820 6610 27832
rect 7009 27829 7021 27832
rect 7055 27829 7067 27863
rect 7009 27823 7067 27829
rect 10781 27863 10839 27869
rect 10781 27829 10793 27863
rect 10827 27860 10839 27863
rect 11054 27860 11060 27872
rect 10827 27832 11060 27860
rect 10827 27829 10839 27832
rect 10781 27823 10839 27829
rect 11054 27820 11060 27832
rect 11112 27820 11118 27872
rect 11149 27863 11207 27869
rect 11149 27829 11161 27863
rect 11195 27860 11207 27863
rect 11238 27860 11244 27872
rect 11195 27832 11244 27860
rect 11195 27829 11207 27832
rect 11149 27823 11207 27829
rect 11238 27820 11244 27832
rect 11296 27820 11302 27872
rect 12066 27820 12072 27872
rect 12124 27820 12130 27872
rect 13188 27869 13216 27900
rect 13173 27863 13231 27869
rect 13173 27829 13185 27863
rect 13219 27829 13231 27863
rect 13556 27860 13584 27900
rect 16025 27897 16037 27900
rect 16071 27897 16083 27931
rect 16868 27928 16896 28027
rect 16960 27996 16988 28027
rect 17678 28024 17684 28036
rect 17736 28024 17742 28076
rect 17770 28024 17776 28076
rect 17828 28024 17834 28076
rect 18138 28064 18144 28076
rect 17880 28036 18144 28064
rect 17589 27999 17647 28005
rect 17589 27996 17601 27999
rect 16960 27968 17601 27996
rect 17589 27965 17601 27968
rect 17635 27996 17647 27999
rect 17880 27996 17908 28036
rect 18138 28024 18144 28036
rect 18196 28064 18202 28076
rect 18509 28067 18567 28073
rect 18509 28064 18521 28067
rect 18196 28036 18521 28064
rect 18196 28024 18202 28036
rect 18509 28033 18521 28036
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 17635 27968 17908 27996
rect 17635 27965 17647 27968
rect 17589 27959 17647 27965
rect 18046 27956 18052 28008
rect 18104 27996 18110 28008
rect 18233 27999 18291 28005
rect 18233 27996 18245 27999
rect 18104 27968 18245 27996
rect 18104 27956 18110 27968
rect 18233 27965 18245 27968
rect 18279 27965 18291 27999
rect 18233 27959 18291 27965
rect 18322 27956 18328 28008
rect 18380 27956 18386 28008
rect 18414 27956 18420 28008
rect 18472 27956 18478 28008
rect 18969 27999 19027 28005
rect 18969 27965 18981 27999
rect 19015 27965 19027 27999
rect 18969 27959 19027 27965
rect 19245 27999 19303 28005
rect 19245 27965 19257 27999
rect 19291 27996 19303 27999
rect 19334 27996 19340 28008
rect 19291 27968 19340 27996
rect 19291 27965 19303 27968
rect 19245 27959 19303 27965
rect 18340 27928 18368 27956
rect 16868 27900 18368 27928
rect 16025 27891 16083 27897
rect 14458 27860 14464 27872
rect 13556 27832 14464 27860
rect 13173 27823 13231 27829
rect 14458 27820 14464 27832
rect 14516 27860 14522 27872
rect 15197 27863 15255 27869
rect 15197 27860 15209 27863
rect 14516 27832 15209 27860
rect 14516 27820 14522 27832
rect 15197 27829 15209 27832
rect 15243 27829 15255 27863
rect 15197 27823 15255 27829
rect 17126 27820 17132 27872
rect 17184 27860 17190 27872
rect 17788 27869 17816 27900
rect 17221 27863 17279 27869
rect 17221 27860 17233 27863
rect 17184 27832 17233 27860
rect 17184 27820 17190 27832
rect 17221 27829 17233 27832
rect 17267 27829 17279 27863
rect 17221 27823 17279 27829
rect 17773 27863 17831 27869
rect 17773 27829 17785 27863
rect 17819 27829 17831 27863
rect 17773 27823 17831 27829
rect 17954 27820 17960 27872
rect 18012 27820 18018 27872
rect 18046 27820 18052 27872
rect 18104 27820 18110 27872
rect 18984 27860 19012 27959
rect 19334 27956 19340 27968
rect 19392 27956 19398 28008
rect 20364 27996 20392 28050
rect 20714 28024 20720 28076
rect 20772 28064 20778 28076
rect 20809 28067 20867 28073
rect 20809 28064 20821 28067
rect 20772 28036 20821 28064
rect 20772 28024 20778 28036
rect 20809 28033 20821 28036
rect 20855 28033 20867 28067
rect 20809 28027 20867 28033
rect 21174 28024 21180 28076
rect 21232 28024 21238 28076
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22557 28067 22615 28073
rect 22557 28064 22569 28067
rect 22336 28036 22569 28064
rect 22336 28024 22342 28036
rect 22557 28033 22569 28036
rect 22603 28033 22615 28067
rect 22557 28027 22615 28033
rect 22922 28024 22928 28076
rect 22980 28024 22986 28076
rect 24302 28024 24308 28076
rect 24360 28024 24366 28076
rect 21192 27996 21220 28024
rect 20364 27968 21220 27996
rect 21634 27956 21640 28008
rect 21692 27996 21698 28008
rect 21821 27999 21879 28005
rect 21821 27996 21833 27999
rect 21692 27968 21833 27996
rect 21692 27956 21698 27968
rect 21821 27965 21833 27968
rect 21867 27965 21879 27999
rect 21821 27959 21879 27965
rect 21910 27956 21916 28008
rect 21968 27996 21974 28008
rect 22833 27999 22891 28005
rect 22833 27996 22845 27999
rect 21968 27968 22845 27996
rect 21968 27956 21974 27968
rect 22833 27965 22845 27968
rect 22879 27965 22891 27999
rect 22833 27959 22891 27965
rect 20254 27888 20260 27940
rect 20312 27928 20318 27940
rect 21453 27931 21511 27937
rect 21453 27928 21465 27931
rect 20312 27900 21465 27928
rect 20312 27888 20318 27900
rect 21453 27897 21465 27900
rect 21499 27897 21511 27931
rect 21453 27891 21511 27897
rect 22646 27888 22652 27940
rect 22704 27888 22710 27940
rect 19886 27860 19892 27872
rect 18984 27832 19892 27860
rect 19886 27820 19892 27832
rect 19944 27820 19950 27872
rect 22462 27820 22468 27872
rect 22520 27820 22526 27872
rect 22554 27820 22560 27872
rect 22612 27820 22618 27872
rect 1104 27770 29440 27792
rect 1104 27718 4491 27770
rect 4543 27718 4555 27770
rect 4607 27718 4619 27770
rect 4671 27718 4683 27770
rect 4735 27718 4747 27770
rect 4799 27718 11574 27770
rect 11626 27718 11638 27770
rect 11690 27718 11702 27770
rect 11754 27718 11766 27770
rect 11818 27718 11830 27770
rect 11882 27718 18657 27770
rect 18709 27718 18721 27770
rect 18773 27718 18785 27770
rect 18837 27718 18849 27770
rect 18901 27718 18913 27770
rect 18965 27718 25740 27770
rect 25792 27718 25804 27770
rect 25856 27718 25868 27770
rect 25920 27718 25932 27770
rect 25984 27718 25996 27770
rect 26048 27718 29440 27770
rect 1104 27696 29440 27718
rect 3602 27616 3608 27668
rect 3660 27656 3666 27668
rect 4982 27656 4988 27668
rect 3660 27628 4660 27656
rect 3660 27616 3666 27628
rect 4632 27597 4660 27628
rect 4908 27628 4988 27656
rect 4617 27591 4675 27597
rect 4617 27557 4629 27591
rect 4663 27557 4675 27591
rect 4617 27551 4675 27557
rect 2685 27523 2743 27529
rect 2685 27489 2697 27523
rect 2731 27520 2743 27523
rect 3142 27520 3148 27532
rect 2731 27492 3148 27520
rect 2731 27489 2743 27492
rect 2685 27483 2743 27489
rect 3142 27480 3148 27492
rect 3200 27480 3206 27532
rect 4246 27480 4252 27532
rect 4304 27520 4310 27532
rect 4801 27523 4859 27529
rect 4801 27520 4813 27523
rect 4304 27492 4813 27520
rect 4304 27480 4310 27492
rect 4801 27489 4813 27492
rect 4847 27489 4859 27523
rect 4801 27483 4859 27489
rect 4338 27412 4344 27464
rect 4396 27452 4402 27464
rect 4908 27461 4936 27628
rect 4982 27616 4988 27628
rect 5040 27656 5046 27668
rect 6362 27656 6368 27668
rect 5040 27628 6368 27656
rect 5040 27616 5046 27628
rect 6362 27616 6368 27628
rect 6420 27616 6426 27668
rect 11054 27616 11060 27668
rect 11112 27656 11118 27668
rect 11330 27656 11336 27668
rect 11112 27628 11336 27656
rect 11112 27616 11118 27628
rect 11330 27616 11336 27628
rect 11388 27616 11394 27668
rect 11882 27616 11888 27668
rect 11940 27656 11946 27668
rect 12066 27656 12072 27668
rect 11940 27628 12072 27656
rect 11940 27616 11946 27628
rect 12066 27616 12072 27628
rect 12124 27616 12130 27668
rect 13998 27616 14004 27668
rect 14056 27616 14062 27668
rect 14458 27616 14464 27668
rect 14516 27656 14522 27668
rect 14553 27659 14611 27665
rect 14553 27656 14565 27659
rect 14516 27628 14565 27656
rect 14516 27616 14522 27628
rect 14553 27625 14565 27628
rect 14599 27625 14611 27659
rect 14553 27619 14611 27625
rect 18138 27616 18144 27668
rect 18196 27656 18202 27668
rect 18233 27659 18291 27665
rect 18233 27656 18245 27659
rect 18196 27628 18245 27656
rect 18196 27616 18202 27628
rect 18233 27625 18245 27628
rect 18279 27625 18291 27659
rect 18233 27619 18291 27625
rect 19245 27659 19303 27665
rect 19245 27625 19257 27659
rect 19291 27656 19303 27659
rect 19334 27656 19340 27668
rect 19291 27628 19340 27656
rect 19291 27625 19303 27628
rect 19245 27619 19303 27625
rect 19334 27616 19340 27628
rect 19392 27616 19398 27668
rect 20152 27659 20210 27665
rect 20152 27625 20164 27659
rect 20198 27656 20210 27659
rect 22554 27656 22560 27668
rect 20198 27628 22560 27656
rect 20198 27625 20210 27628
rect 20152 27619 20210 27625
rect 22554 27616 22560 27628
rect 22612 27616 22618 27668
rect 7374 27548 7380 27600
rect 7432 27588 7438 27600
rect 8113 27591 8171 27597
rect 8113 27588 8125 27591
rect 7432 27560 8125 27588
rect 7432 27548 7438 27560
rect 8113 27557 8125 27560
rect 8159 27588 8171 27591
rect 11146 27588 11152 27600
rect 8159 27560 11152 27588
rect 8159 27557 8171 27560
rect 8113 27551 8171 27557
rect 8496 27461 8524 27560
rect 11146 27548 11152 27560
rect 11204 27548 11210 27600
rect 11348 27588 11376 27616
rect 12161 27591 12219 27597
rect 11348 27560 11744 27588
rect 9306 27480 9312 27532
rect 9364 27480 9370 27532
rect 11716 27529 11744 27560
rect 12161 27557 12173 27591
rect 12207 27588 12219 27591
rect 13909 27591 13967 27597
rect 13909 27588 13921 27591
rect 12207 27560 12434 27588
rect 12207 27557 12219 27560
rect 12161 27551 12219 27557
rect 9401 27523 9459 27529
rect 9401 27489 9413 27523
rect 9447 27520 9459 27523
rect 10229 27523 10287 27529
rect 10229 27520 10241 27523
rect 9447 27492 10241 27520
rect 9447 27489 9459 27492
rect 9401 27483 9459 27489
rect 10229 27489 10241 27492
rect 10275 27489 10287 27523
rect 11517 27523 11575 27529
rect 11517 27520 11529 27523
rect 10229 27483 10287 27489
rect 10336 27492 11529 27520
rect 4433 27455 4491 27461
rect 4433 27452 4445 27455
rect 4396 27424 4445 27452
rect 4396 27412 4402 27424
rect 4433 27421 4445 27424
rect 4479 27421 4491 27455
rect 4433 27415 4491 27421
rect 4709 27455 4767 27461
rect 4709 27421 4721 27455
rect 4755 27421 4767 27455
rect 4709 27415 4767 27421
rect 4893 27455 4951 27461
rect 4893 27421 4905 27455
rect 4939 27421 4951 27455
rect 4893 27415 4951 27421
rect 8481 27455 8539 27461
rect 8481 27421 8493 27455
rect 8527 27421 8539 27455
rect 8481 27415 8539 27421
rect 9125 27455 9183 27461
rect 9125 27421 9137 27455
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 9677 27455 9735 27461
rect 9677 27421 9689 27455
rect 9723 27452 9735 27455
rect 9766 27452 9772 27464
rect 9723 27424 9772 27452
rect 9723 27421 9735 27424
rect 9677 27415 9735 27421
rect 1486 27344 1492 27396
rect 1544 27344 1550 27396
rect 4724 27384 4752 27415
rect 5074 27384 5080 27396
rect 4724 27356 5080 27384
rect 5074 27344 5080 27356
rect 5132 27344 5138 27396
rect 7745 27387 7803 27393
rect 7745 27353 7757 27387
rect 7791 27353 7803 27387
rect 7745 27347 7803 27353
rect 934 27276 940 27328
rect 992 27316 998 27328
rect 1581 27319 1639 27325
rect 1581 27316 1593 27319
rect 992 27288 1593 27316
rect 992 27276 998 27288
rect 1581 27285 1593 27288
rect 1627 27285 1639 27319
rect 1581 27279 1639 27285
rect 3050 27276 3056 27328
rect 3108 27316 3114 27328
rect 3329 27319 3387 27325
rect 3329 27316 3341 27319
rect 3108 27288 3341 27316
rect 3108 27276 3114 27288
rect 3329 27285 3341 27288
rect 3375 27285 3387 27319
rect 7760 27316 7788 27347
rect 7926 27344 7932 27396
rect 7984 27344 7990 27396
rect 9030 27384 9036 27396
rect 8496 27356 9036 27384
rect 8496 27316 8524 27356
rect 9030 27344 9036 27356
rect 9088 27344 9094 27396
rect 9140 27384 9168 27415
rect 9766 27412 9772 27424
rect 9824 27412 9830 27464
rect 9950 27412 9956 27464
rect 10008 27452 10014 27464
rect 10336 27461 10364 27492
rect 11517 27489 11529 27492
rect 11563 27489 11575 27523
rect 11517 27483 11575 27489
rect 11701 27523 11759 27529
rect 11701 27489 11713 27523
rect 11747 27489 11759 27523
rect 11701 27483 11759 27489
rect 11793 27523 11851 27529
rect 11793 27489 11805 27523
rect 11839 27520 11851 27523
rect 11839 27492 12296 27520
rect 11839 27489 11851 27492
rect 11793 27483 11851 27489
rect 12268 27464 12296 27492
rect 10321 27455 10379 27461
rect 10321 27452 10333 27455
rect 10008 27424 10333 27452
rect 10008 27412 10014 27424
rect 10321 27421 10333 27424
rect 10367 27421 10379 27455
rect 10321 27415 10379 27421
rect 10505 27455 10563 27461
rect 10505 27421 10517 27455
rect 10551 27421 10563 27455
rect 10505 27415 10563 27421
rect 10413 27387 10471 27393
rect 10413 27384 10425 27387
rect 9140 27356 10425 27384
rect 10413 27353 10425 27356
rect 10459 27353 10471 27387
rect 10520 27384 10548 27415
rect 11422 27412 11428 27464
rect 11480 27452 11486 27464
rect 11609 27455 11667 27461
rect 11609 27452 11621 27455
rect 11480 27424 11621 27452
rect 11480 27412 11486 27424
rect 11609 27421 11621 27424
rect 11655 27421 11667 27455
rect 11609 27415 11667 27421
rect 11882 27412 11888 27464
rect 11940 27452 11946 27464
rect 11977 27455 12035 27461
rect 11977 27452 11989 27455
rect 11940 27424 11989 27452
rect 11940 27412 11946 27424
rect 11977 27421 11989 27424
rect 12023 27421 12035 27455
rect 11977 27415 12035 27421
rect 12250 27412 12256 27464
rect 12308 27412 12314 27464
rect 12406 27452 12434 27560
rect 12636 27560 13921 27588
rect 12636 27461 12664 27560
rect 13909 27557 13921 27560
rect 13955 27557 13967 27591
rect 14016 27588 14044 27616
rect 14829 27591 14887 27597
rect 14829 27588 14841 27591
rect 14016 27560 14841 27588
rect 13909 27551 13967 27557
rect 14829 27557 14841 27560
rect 14875 27557 14887 27591
rect 14829 27551 14887 27557
rect 21729 27591 21787 27597
rect 21729 27557 21741 27591
rect 21775 27588 21787 27591
rect 22646 27588 22652 27600
rect 21775 27560 22652 27588
rect 21775 27557 21787 27560
rect 21729 27551 21787 27557
rect 22646 27548 22652 27560
rect 22704 27548 22710 27600
rect 22830 27588 22836 27600
rect 22756 27560 22836 27588
rect 12710 27480 12716 27532
rect 12768 27480 12774 27532
rect 12989 27523 13047 27529
rect 12989 27489 13001 27523
rect 13035 27489 13047 27523
rect 12989 27483 13047 27489
rect 12621 27455 12679 27461
rect 12406 27424 12572 27452
rect 12544 27384 12572 27424
rect 12621 27421 12633 27455
rect 12667 27421 12679 27455
rect 12621 27415 12679 27421
rect 12728 27384 12756 27480
rect 13004 27396 13032 27483
rect 13078 27480 13084 27532
rect 13136 27520 13142 27532
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 13136 27492 13277 27520
rect 13136 27480 13142 27492
rect 13265 27489 13277 27492
rect 13311 27520 13323 27523
rect 13998 27520 14004 27532
rect 13311 27492 14004 27520
rect 13311 27489 13323 27492
rect 13265 27483 13323 27489
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 14185 27523 14243 27529
rect 14185 27489 14197 27523
rect 14231 27520 14243 27523
rect 15470 27520 15476 27532
rect 14231 27492 15476 27520
rect 14231 27489 14243 27492
rect 14185 27483 14243 27489
rect 15470 27480 15476 27492
rect 15528 27480 15534 27532
rect 17126 27480 17132 27532
rect 17184 27520 17190 27532
rect 19426 27520 19432 27532
rect 17184 27492 19432 27520
rect 17184 27480 17190 27492
rect 19426 27480 19432 27492
rect 19484 27520 19490 27532
rect 19794 27520 19800 27532
rect 19484 27492 19800 27520
rect 19484 27480 19490 27492
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13372 27424 14289 27452
rect 10520 27356 12020 27384
rect 12544 27356 12756 27384
rect 10413 27347 10471 27353
rect 11992 27328 12020 27356
rect 12986 27344 12992 27396
rect 13044 27344 13050 27396
rect 7760 27288 8524 27316
rect 3329 27279 3387 27285
rect 8570 27276 8576 27328
rect 8628 27276 8634 27328
rect 8938 27276 8944 27328
rect 8996 27276 9002 27328
rect 11333 27319 11391 27325
rect 11333 27285 11345 27319
rect 11379 27316 11391 27319
rect 11882 27316 11888 27328
rect 11379 27288 11888 27316
rect 11379 27285 11391 27288
rect 11333 27279 11391 27285
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 11974 27276 11980 27328
rect 12032 27276 12038 27328
rect 12250 27276 12256 27328
rect 12308 27316 12314 27328
rect 13372 27316 13400 27424
rect 14277 27421 14289 27424
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 12308 27288 13400 27316
rect 12308 27276 12314 27288
rect 13998 27276 14004 27328
rect 14056 27316 14062 27328
rect 14550 27316 14556 27328
rect 14056 27288 14556 27316
rect 14056 27276 14062 27288
rect 14550 27276 14556 27288
rect 14608 27316 14614 27328
rect 14660 27316 14688 27415
rect 16390 27412 16396 27464
rect 16448 27412 16454 27464
rect 16482 27412 16488 27464
rect 16540 27412 16546 27464
rect 17770 27412 17776 27464
rect 17828 27452 17834 27464
rect 18230 27452 18236 27464
rect 17828 27424 18236 27452
rect 17828 27412 17834 27424
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 19536 27461 19564 27492
rect 19794 27480 19800 27492
rect 19852 27480 19858 27532
rect 19886 27480 19892 27532
rect 19944 27480 19950 27532
rect 20714 27480 20720 27532
rect 20772 27520 20778 27532
rect 20772 27492 21956 27520
rect 20772 27480 20778 27492
rect 19521 27455 19579 27461
rect 19521 27421 19533 27455
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 19702 27412 19708 27464
rect 19760 27412 19766 27464
rect 21928 27461 21956 27492
rect 22094 27480 22100 27532
rect 22152 27520 22158 27532
rect 22756 27529 22784 27560
rect 22830 27548 22836 27560
rect 22888 27548 22894 27600
rect 22189 27523 22247 27529
rect 22189 27520 22201 27523
rect 22152 27492 22201 27520
rect 22152 27480 22158 27492
rect 22189 27489 22201 27492
rect 22235 27489 22247 27523
rect 22189 27483 22247 27489
rect 22741 27523 22799 27529
rect 22741 27489 22753 27523
rect 22787 27489 22799 27523
rect 22741 27483 22799 27489
rect 21913 27455 21971 27461
rect 21913 27421 21925 27455
rect 21959 27421 21971 27455
rect 21913 27415 21971 27421
rect 22002 27412 22008 27464
rect 22060 27412 22066 27464
rect 22278 27412 22284 27464
rect 22336 27452 22342 27464
rect 22373 27455 22431 27461
rect 22373 27452 22385 27455
rect 22336 27424 22385 27452
rect 22336 27412 22342 27424
rect 22373 27421 22385 27424
rect 22419 27452 22431 27455
rect 22649 27455 22707 27461
rect 22649 27452 22661 27455
rect 22419 27424 22661 27452
rect 22419 27421 22431 27424
rect 22373 27415 22431 27421
rect 22649 27421 22661 27424
rect 22695 27421 22707 27455
rect 22649 27415 22707 27421
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 24394 27452 24400 27464
rect 22879 27424 24400 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 24394 27412 24400 27424
rect 24452 27412 24458 27464
rect 16761 27387 16819 27393
rect 16761 27353 16773 27387
rect 16807 27353 16819 27387
rect 16761 27347 16819 27353
rect 19245 27387 19303 27393
rect 19245 27353 19257 27387
rect 19291 27384 19303 27387
rect 19720 27384 19748 27412
rect 19291 27356 19748 27384
rect 19291 27353 19303 27356
rect 19245 27347 19303 27353
rect 14608 27288 14688 27316
rect 16209 27319 16267 27325
rect 14608 27276 14614 27288
rect 16209 27285 16221 27319
rect 16255 27316 16267 27319
rect 16776 27316 16804 27347
rect 20254 27344 20260 27396
rect 20312 27344 20318 27396
rect 21174 27344 21180 27396
rect 21232 27344 21238 27396
rect 21729 27387 21787 27393
rect 21729 27353 21741 27387
rect 21775 27384 21787 27387
rect 22462 27384 22468 27396
rect 21775 27356 22468 27384
rect 21775 27353 21787 27356
rect 21729 27347 21787 27353
rect 22462 27344 22468 27356
rect 22520 27344 22526 27396
rect 16255 27288 16804 27316
rect 19429 27319 19487 27325
rect 16255 27285 16267 27288
rect 16209 27279 16267 27285
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 20272 27316 20300 27344
rect 19475 27288 20300 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 20990 27276 20996 27328
rect 21048 27316 21054 27328
rect 21634 27316 21640 27328
rect 21048 27288 21640 27316
rect 21048 27276 21054 27288
rect 21634 27276 21640 27288
rect 21692 27276 21698 27328
rect 22186 27276 22192 27328
rect 22244 27316 22250 27328
rect 22557 27319 22615 27325
rect 22557 27316 22569 27319
rect 22244 27288 22569 27316
rect 22244 27276 22250 27288
rect 22557 27285 22569 27288
rect 22603 27285 22615 27319
rect 22557 27279 22615 27285
rect 1104 27226 29440 27248
rect 1104 27174 5151 27226
rect 5203 27174 5215 27226
rect 5267 27174 5279 27226
rect 5331 27174 5343 27226
rect 5395 27174 5407 27226
rect 5459 27174 12234 27226
rect 12286 27174 12298 27226
rect 12350 27174 12362 27226
rect 12414 27174 12426 27226
rect 12478 27174 12490 27226
rect 12542 27174 19317 27226
rect 19369 27174 19381 27226
rect 19433 27174 19445 27226
rect 19497 27174 19509 27226
rect 19561 27174 19573 27226
rect 19625 27174 26400 27226
rect 26452 27174 26464 27226
rect 26516 27174 26528 27226
rect 26580 27174 26592 27226
rect 26644 27174 26656 27226
rect 26708 27174 29440 27226
rect 1104 27152 29440 27174
rect 8938 27112 8944 27124
rect 8220 27084 8944 27112
rect 8220 27053 8248 27084
rect 8938 27072 8944 27084
rect 8996 27072 9002 27124
rect 9030 27072 9036 27124
rect 9088 27112 9094 27124
rect 9677 27115 9735 27121
rect 9088 27084 9628 27112
rect 9088 27072 9094 27084
rect 8205 27047 8263 27053
rect 8205 27013 8217 27047
rect 8251 27013 8263 27047
rect 9600 27044 9628 27084
rect 9677 27081 9689 27115
rect 9723 27112 9735 27115
rect 9766 27112 9772 27124
rect 9723 27084 9772 27112
rect 9723 27081 9735 27084
rect 9677 27075 9735 27081
rect 9766 27072 9772 27084
rect 9824 27072 9830 27124
rect 13630 27112 13636 27124
rect 10060 27084 13636 27112
rect 10060 27044 10088 27084
rect 13630 27072 13636 27084
rect 13688 27072 13694 27124
rect 14550 27072 14556 27124
rect 14608 27072 14614 27124
rect 16390 27072 16396 27124
rect 16448 27112 16454 27124
rect 17589 27115 17647 27121
rect 17589 27112 17601 27115
rect 16448 27084 17601 27112
rect 16448 27072 16454 27084
rect 17589 27081 17601 27084
rect 17635 27081 17647 27115
rect 17589 27075 17647 27081
rect 19794 27072 19800 27124
rect 19852 27072 19858 27124
rect 20898 27072 20904 27124
rect 20956 27112 20962 27124
rect 21177 27115 21235 27121
rect 21177 27112 21189 27115
rect 20956 27084 21189 27112
rect 20956 27072 20962 27084
rect 21177 27081 21189 27084
rect 21223 27112 21235 27115
rect 22278 27112 22284 27124
rect 21223 27084 22284 27112
rect 21223 27081 21235 27084
rect 21177 27075 21235 27081
rect 22278 27072 22284 27084
rect 22336 27072 22342 27124
rect 9600 27016 10088 27044
rect 8205 27007 8263 27013
rect 11330 27004 11336 27056
rect 11388 27044 11394 27056
rect 12066 27044 12072 27056
rect 11388 27016 12072 27044
rect 11388 27004 11394 27016
rect 12066 27004 12072 27016
rect 12124 27044 12130 27056
rect 12894 27044 12900 27056
rect 12124 27016 12900 27044
rect 12124 27004 12130 27016
rect 12894 27004 12900 27016
rect 12952 27004 12958 27056
rect 14369 27047 14427 27053
rect 14369 27013 14381 27047
rect 14415 27044 14427 27047
rect 14734 27044 14740 27056
rect 14415 27016 14740 27044
rect 14415 27013 14427 27016
rect 14369 27007 14427 27013
rect 14734 27004 14740 27016
rect 14792 27004 14798 27056
rect 17126 27004 17132 27056
rect 17184 27004 17190 27056
rect 9582 26976 9588 26988
rect 9338 26948 9588 26976
rect 9582 26936 9588 26948
rect 9640 26936 9646 26988
rect 11793 26979 11851 26985
rect 11793 26976 11805 26979
rect 11624 26948 11805 26976
rect 7834 26868 7840 26920
rect 7892 26908 7898 26920
rect 7929 26911 7987 26917
rect 7929 26908 7941 26911
rect 7892 26880 7941 26908
rect 7892 26868 7898 26880
rect 7929 26877 7941 26880
rect 7975 26877 7987 26911
rect 7929 26871 7987 26877
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 11624 26908 11652 26948
rect 11793 26945 11805 26948
rect 11839 26945 11851 26979
rect 11793 26939 11851 26945
rect 11882 26936 11888 26988
rect 11940 26936 11946 26988
rect 12250 26936 12256 26988
rect 12308 26976 12314 26988
rect 12518 26979 12576 26985
rect 12518 26976 12530 26979
rect 12308 26948 12530 26976
rect 12308 26936 12314 26948
rect 12518 26945 12530 26948
rect 12564 26945 12576 26979
rect 12518 26939 12576 26945
rect 13906 26936 13912 26988
rect 13964 26976 13970 26988
rect 14274 26976 14280 26988
rect 13964 26948 14280 26976
rect 13964 26936 13970 26948
rect 14274 26936 14280 26948
rect 14332 26936 14338 26988
rect 14645 26979 14703 26985
rect 14645 26945 14657 26979
rect 14691 26945 14703 26979
rect 19812 26976 19840 27072
rect 20714 27004 20720 27056
rect 20772 27044 20778 27056
rect 20809 27047 20867 27053
rect 20809 27044 20821 27047
rect 20772 27016 20821 27044
rect 20772 27004 20778 27016
rect 20809 27013 20821 27016
rect 20855 27013 20867 27047
rect 21009 27047 21067 27053
rect 21009 27044 21021 27047
rect 20809 27007 20867 27013
rect 20916 27016 21021 27044
rect 20916 26976 20944 27016
rect 21009 27013 21021 27016
rect 21055 27044 21067 27047
rect 22002 27044 22008 27056
rect 21055 27016 22008 27044
rect 21055 27013 21067 27016
rect 21009 27007 21067 27013
rect 22002 27004 22008 27016
rect 22060 27004 22066 27056
rect 19812 26948 20944 26976
rect 14645 26939 14703 26945
rect 8628 26880 11652 26908
rect 8628 26868 8634 26880
rect 11624 26840 11652 26880
rect 11701 26911 11759 26917
rect 11701 26877 11713 26911
rect 11747 26908 11759 26911
rect 12802 26908 12808 26920
rect 11747 26880 12480 26908
rect 11747 26877 11759 26880
rect 11701 26871 11759 26877
rect 11974 26840 11980 26852
rect 11624 26812 11980 26840
rect 11974 26800 11980 26812
rect 12032 26800 12038 26852
rect 12452 26840 12480 26880
rect 12636 26880 12808 26908
rect 12636 26840 12664 26880
rect 12802 26868 12808 26880
rect 12860 26908 12866 26920
rect 14660 26908 14688 26939
rect 28258 26936 28264 26988
rect 28316 26976 28322 26988
rect 28813 26979 28871 26985
rect 28813 26976 28825 26979
rect 28316 26948 28825 26976
rect 28316 26936 28322 26948
rect 28813 26945 28825 26948
rect 28859 26945 28871 26979
rect 28813 26939 28871 26945
rect 12860 26880 14688 26908
rect 12860 26868 12866 26880
rect 15286 26868 15292 26920
rect 15344 26868 15350 26920
rect 12452 26812 12664 26840
rect 13906 26800 13912 26852
rect 13964 26800 13970 26852
rect 13998 26800 14004 26852
rect 14056 26840 14062 26852
rect 14277 26843 14335 26849
rect 14277 26840 14289 26843
rect 14056 26812 14289 26840
rect 14056 26800 14062 26812
rect 14277 26809 14289 26812
rect 14323 26809 14335 26843
rect 14277 26803 14335 26809
rect 14369 26843 14427 26849
rect 14369 26809 14381 26843
rect 14415 26840 14427 26843
rect 15304 26840 15332 26868
rect 14415 26812 15332 26840
rect 17497 26843 17555 26849
rect 14415 26809 14427 26812
rect 14369 26803 14427 26809
rect 17497 26809 17509 26843
rect 17543 26840 17555 26843
rect 18046 26840 18052 26852
rect 17543 26812 18052 26840
rect 17543 26809 17555 26812
rect 17497 26803 17555 26809
rect 18046 26800 18052 26812
rect 18104 26800 18110 26852
rect 11238 26732 11244 26784
rect 11296 26772 11302 26784
rect 12802 26781 12808 26784
rect 11517 26775 11575 26781
rect 11517 26772 11529 26775
rect 11296 26744 11529 26772
rect 11296 26732 11302 26744
rect 11517 26741 11529 26744
rect 11563 26741 11575 26775
rect 11517 26735 11575 26741
rect 12792 26775 12808 26781
rect 12792 26741 12804 26775
rect 12792 26735 12808 26741
rect 12802 26732 12808 26735
rect 12860 26732 12866 26784
rect 12894 26732 12900 26784
rect 12952 26772 12958 26784
rect 13924 26772 13952 26800
rect 12952 26744 13952 26772
rect 12952 26732 12958 26744
rect 20990 26732 20996 26784
rect 21048 26732 21054 26784
rect 28994 26732 29000 26784
rect 29052 26732 29058 26784
rect 1104 26682 29440 26704
rect 1104 26630 4491 26682
rect 4543 26630 4555 26682
rect 4607 26630 4619 26682
rect 4671 26630 4683 26682
rect 4735 26630 4747 26682
rect 4799 26630 11574 26682
rect 11626 26630 11638 26682
rect 11690 26630 11702 26682
rect 11754 26630 11766 26682
rect 11818 26630 11830 26682
rect 11882 26630 18657 26682
rect 18709 26630 18721 26682
rect 18773 26630 18785 26682
rect 18837 26630 18849 26682
rect 18901 26630 18913 26682
rect 18965 26630 25740 26682
rect 25792 26630 25804 26682
rect 25856 26630 25868 26682
rect 25920 26630 25932 26682
rect 25984 26630 25996 26682
rect 26048 26630 29440 26682
rect 1104 26608 29440 26630
rect 1486 26528 1492 26580
rect 1544 26568 1550 26580
rect 2225 26571 2283 26577
rect 2225 26568 2237 26571
rect 1544 26540 2237 26568
rect 1544 26528 1550 26540
rect 2225 26537 2237 26540
rect 2271 26537 2283 26571
rect 2225 26531 2283 26537
rect 11044 26571 11102 26577
rect 11044 26537 11056 26571
rect 11090 26568 11102 26571
rect 11238 26568 11244 26580
rect 11090 26540 11244 26568
rect 11090 26537 11102 26540
rect 11044 26531 11102 26537
rect 11238 26528 11244 26540
rect 11296 26528 11302 26580
rect 12158 26528 12164 26580
rect 12216 26568 12222 26580
rect 12529 26571 12587 26577
rect 12529 26568 12541 26571
rect 12216 26540 12541 26568
rect 12216 26528 12222 26540
rect 12529 26537 12541 26540
rect 12575 26537 12587 26571
rect 12529 26531 12587 26537
rect 6825 26435 6883 26441
rect 6825 26432 6837 26435
rect 5920 26404 6837 26432
rect 2406 26324 2412 26376
rect 2464 26324 2470 26376
rect 5920 26373 5948 26404
rect 6825 26401 6837 26404
rect 6871 26401 6883 26435
rect 6825 26395 6883 26401
rect 10778 26392 10784 26444
rect 10836 26432 10842 26444
rect 11422 26432 11428 26444
rect 10836 26404 11428 26432
rect 10836 26392 10842 26404
rect 11422 26392 11428 26404
rect 11480 26432 11486 26444
rect 12250 26432 12256 26444
rect 11480 26404 12256 26432
rect 11480 26392 11486 26404
rect 12250 26392 12256 26404
rect 12308 26392 12314 26444
rect 5721 26367 5779 26373
rect 5721 26333 5733 26367
rect 5767 26333 5779 26367
rect 5721 26327 5779 26333
rect 5905 26367 5963 26373
rect 5905 26333 5917 26367
rect 5951 26333 5963 26367
rect 5905 26327 5963 26333
rect 6273 26367 6331 26373
rect 6273 26333 6285 26367
rect 6319 26364 6331 26367
rect 6454 26364 6460 26376
rect 6319 26336 6460 26364
rect 6319 26333 6331 26336
rect 6273 26327 6331 26333
rect 5736 26296 5764 26327
rect 6454 26324 6460 26336
rect 6512 26324 6518 26376
rect 9582 26324 9588 26376
rect 9640 26324 9646 26376
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 19613 26367 19671 26373
rect 19613 26364 19625 26367
rect 18012 26336 19625 26364
rect 18012 26324 18018 26336
rect 19613 26333 19625 26336
rect 19659 26333 19671 26367
rect 19613 26327 19671 26333
rect 19720 26336 20024 26364
rect 7006 26296 7012 26308
rect 5736 26268 7012 26296
rect 7006 26256 7012 26268
rect 7064 26256 7070 26308
rect 9600 26296 9628 26324
rect 11330 26296 11336 26308
rect 9600 26268 11336 26296
rect 11330 26256 11336 26268
rect 11388 26296 11394 26308
rect 19245 26299 19303 26305
rect 11388 26268 11546 26296
rect 11388 26256 11394 26268
rect 19245 26265 19257 26299
rect 19291 26296 19303 26299
rect 19429 26299 19487 26305
rect 19291 26268 19380 26296
rect 19291 26265 19303 26268
rect 19245 26259 19303 26265
rect 5810 26188 5816 26240
rect 5868 26188 5874 26240
rect 19352 26228 19380 26268
rect 19429 26265 19441 26299
rect 19475 26296 19487 26299
rect 19720 26296 19748 26336
rect 19996 26308 20024 26336
rect 19475 26268 19748 26296
rect 19475 26265 19487 26268
rect 19429 26259 19487 26265
rect 19794 26256 19800 26308
rect 19852 26256 19858 26308
rect 19978 26256 19984 26308
rect 20036 26256 20042 26308
rect 19812 26228 19840 26256
rect 19352 26200 19840 26228
rect 1104 26138 29440 26160
rect 1104 26086 5151 26138
rect 5203 26086 5215 26138
rect 5267 26086 5279 26138
rect 5331 26086 5343 26138
rect 5395 26086 5407 26138
rect 5459 26086 12234 26138
rect 12286 26086 12298 26138
rect 12350 26086 12362 26138
rect 12414 26086 12426 26138
rect 12478 26086 12490 26138
rect 12542 26086 19317 26138
rect 19369 26086 19381 26138
rect 19433 26086 19445 26138
rect 19497 26086 19509 26138
rect 19561 26086 19573 26138
rect 19625 26086 26400 26138
rect 26452 26086 26464 26138
rect 26516 26086 26528 26138
rect 26580 26086 26592 26138
rect 26644 26086 26656 26138
rect 26708 26086 29440 26138
rect 1104 26064 29440 26086
rect 5810 25984 5816 26036
rect 5868 25984 5874 26036
rect 6181 26027 6239 26033
rect 6181 25993 6193 26027
rect 6227 26024 6239 26027
rect 7926 26024 7932 26036
rect 6227 25996 7932 26024
rect 6227 25993 6239 25996
rect 6181 25987 6239 25993
rect 7926 25984 7932 25996
rect 7984 25984 7990 26036
rect 5828 25956 5856 25984
rect 6454 25956 6460 25968
rect 5000 25928 5856 25956
rect 6012 25928 6460 25956
rect 5000 25897 5028 25928
rect 4985 25891 5043 25897
rect 4985 25857 4997 25891
rect 5031 25857 5043 25891
rect 4985 25851 5043 25857
rect 5074 25848 5080 25900
rect 5132 25888 5138 25900
rect 5169 25891 5227 25897
rect 5169 25888 5181 25891
rect 5132 25860 5181 25888
rect 5132 25848 5138 25860
rect 5169 25857 5181 25860
rect 5215 25857 5227 25891
rect 5169 25851 5227 25857
rect 5261 25891 5319 25897
rect 5261 25857 5273 25891
rect 5307 25857 5319 25891
rect 5261 25851 5319 25857
rect 4338 25712 4344 25764
rect 4396 25752 4402 25764
rect 5276 25752 5304 25851
rect 5442 25848 5448 25900
rect 5500 25848 5506 25900
rect 5626 25848 5632 25900
rect 5684 25888 5690 25900
rect 6012 25897 6040 25928
rect 6454 25916 6460 25928
rect 6512 25916 6518 25968
rect 8128 25928 8432 25956
rect 5721 25891 5779 25897
rect 5721 25888 5733 25891
rect 5684 25860 5733 25888
rect 5684 25848 5690 25860
rect 5721 25857 5733 25860
rect 5767 25857 5779 25891
rect 5721 25851 5779 25857
rect 5997 25891 6055 25897
rect 5997 25857 6009 25891
rect 6043 25857 6055 25891
rect 6546 25888 6552 25900
rect 5997 25851 6055 25857
rect 6380 25860 6552 25888
rect 5905 25823 5963 25829
rect 5905 25789 5917 25823
rect 5951 25820 5963 25823
rect 6380 25820 6408 25860
rect 6546 25848 6552 25860
rect 6604 25848 6610 25900
rect 6914 25848 6920 25900
rect 6972 25888 6978 25900
rect 7101 25891 7159 25897
rect 7101 25888 7113 25891
rect 6972 25860 7113 25888
rect 6972 25848 6978 25860
rect 7101 25857 7113 25860
rect 7147 25857 7159 25891
rect 7101 25851 7159 25857
rect 7190 25848 7196 25900
rect 7248 25888 7254 25900
rect 8128 25897 8156 25928
rect 8404 25897 8432 25928
rect 18230 25916 18236 25968
rect 18288 25956 18294 25968
rect 19061 25959 19119 25965
rect 19061 25956 19073 25959
rect 18288 25928 19073 25956
rect 18288 25916 18294 25928
rect 19061 25925 19073 25928
rect 19107 25925 19119 25959
rect 19061 25919 19119 25925
rect 7285 25891 7343 25897
rect 7285 25888 7297 25891
rect 7248 25860 7297 25888
rect 7248 25848 7254 25860
rect 7285 25857 7297 25860
rect 7331 25857 7343 25891
rect 7285 25851 7343 25857
rect 7377 25891 7435 25897
rect 7377 25857 7389 25891
rect 7423 25888 7435 25891
rect 8113 25891 8171 25897
rect 8113 25888 8125 25891
rect 7423 25860 8125 25888
rect 7423 25857 7435 25860
rect 7377 25851 7435 25857
rect 8113 25857 8125 25860
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 8205 25891 8263 25897
rect 8205 25857 8217 25891
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 8389 25891 8447 25897
rect 8389 25857 8401 25891
rect 8435 25857 8447 25891
rect 8389 25851 8447 25857
rect 5951 25792 6408 25820
rect 6457 25823 6515 25829
rect 5951 25789 5963 25792
rect 5905 25783 5963 25789
rect 6457 25789 6469 25823
rect 6503 25789 6515 25823
rect 6457 25783 6515 25789
rect 6472 25752 6500 25783
rect 6822 25780 6828 25832
rect 6880 25820 6886 25832
rect 7561 25823 7619 25829
rect 7561 25820 7573 25823
rect 6880 25792 7573 25820
rect 6880 25780 6886 25792
rect 7561 25789 7573 25792
rect 7607 25789 7619 25823
rect 8220 25820 8248 25851
rect 20070 25848 20076 25900
rect 20128 25888 20134 25900
rect 20128 25860 20194 25888
rect 20128 25848 20134 25860
rect 8570 25820 8576 25832
rect 8220 25792 8576 25820
rect 7561 25783 7619 25789
rect 7101 25755 7159 25761
rect 7101 25752 7113 25755
rect 4396 25724 5856 25752
rect 6472 25724 7113 25752
rect 4396 25712 4402 25724
rect 4982 25644 4988 25696
rect 5040 25644 5046 25696
rect 5626 25644 5632 25696
rect 5684 25644 5690 25696
rect 5718 25644 5724 25696
rect 5776 25644 5782 25696
rect 5828 25684 5856 25724
rect 7101 25721 7113 25724
rect 7147 25721 7159 25755
rect 7101 25715 7159 25721
rect 7576 25696 7604 25783
rect 8570 25780 8576 25792
rect 8628 25780 8634 25832
rect 17862 25780 17868 25832
rect 17920 25820 17926 25832
rect 18785 25823 18843 25829
rect 18785 25820 18797 25823
rect 17920 25792 18797 25820
rect 17920 25780 17926 25792
rect 18785 25789 18797 25792
rect 18831 25789 18843 25823
rect 18785 25783 18843 25789
rect 7742 25712 7748 25764
rect 7800 25752 7806 25764
rect 8205 25755 8263 25761
rect 8205 25752 8217 25755
rect 7800 25724 8217 25752
rect 7800 25712 7806 25724
rect 8205 25721 8217 25724
rect 8251 25721 8263 25755
rect 8205 25715 8263 25721
rect 6822 25684 6828 25696
rect 5828 25656 6828 25684
rect 6822 25644 6828 25656
rect 6880 25644 6886 25696
rect 7009 25687 7067 25693
rect 7009 25653 7021 25687
rect 7055 25684 7067 25687
rect 7282 25684 7288 25696
rect 7055 25656 7288 25684
rect 7055 25653 7067 25656
rect 7009 25647 7067 25653
rect 7282 25644 7288 25656
rect 7340 25644 7346 25696
rect 7558 25644 7564 25696
rect 7616 25684 7622 25696
rect 8754 25684 8760 25696
rect 7616 25656 8760 25684
rect 7616 25644 7622 25656
rect 8754 25644 8760 25656
rect 8812 25644 8818 25696
rect 20533 25687 20591 25693
rect 20533 25653 20545 25687
rect 20579 25684 20591 25687
rect 20714 25684 20720 25696
rect 20579 25656 20720 25684
rect 20579 25653 20591 25656
rect 20533 25647 20591 25653
rect 20714 25644 20720 25656
rect 20772 25644 20778 25696
rect 1104 25594 29440 25616
rect 1104 25542 4491 25594
rect 4543 25542 4555 25594
rect 4607 25542 4619 25594
rect 4671 25542 4683 25594
rect 4735 25542 4747 25594
rect 4799 25542 11574 25594
rect 11626 25542 11638 25594
rect 11690 25542 11702 25594
rect 11754 25542 11766 25594
rect 11818 25542 11830 25594
rect 11882 25542 18657 25594
rect 18709 25542 18721 25594
rect 18773 25542 18785 25594
rect 18837 25542 18849 25594
rect 18901 25542 18913 25594
rect 18965 25542 25740 25594
rect 25792 25542 25804 25594
rect 25856 25542 25868 25594
rect 25920 25542 25932 25594
rect 25984 25542 25996 25594
rect 26048 25542 29440 25594
rect 1104 25520 29440 25542
rect 3605 25483 3663 25489
rect 3605 25449 3617 25483
rect 3651 25480 3663 25483
rect 6362 25480 6368 25492
rect 3651 25452 6368 25480
rect 3651 25449 3663 25452
rect 3605 25443 3663 25449
rect 6362 25440 6368 25452
rect 6420 25440 6426 25492
rect 6733 25483 6791 25489
rect 6733 25449 6745 25483
rect 6779 25480 6791 25483
rect 6822 25480 6828 25492
rect 6779 25452 6828 25480
rect 6779 25449 6791 25452
rect 6733 25443 6791 25449
rect 6822 25440 6828 25452
rect 6880 25440 6886 25492
rect 6917 25483 6975 25489
rect 6917 25449 6929 25483
rect 6963 25480 6975 25483
rect 7006 25480 7012 25492
rect 6963 25452 7012 25480
rect 6963 25449 6975 25452
rect 6917 25443 6975 25449
rect 7006 25440 7012 25452
rect 7064 25440 7070 25492
rect 7272 25483 7330 25489
rect 7272 25449 7284 25483
rect 7318 25480 7330 25483
rect 7742 25480 7748 25492
rect 7318 25452 7748 25480
rect 7318 25449 7330 25452
rect 7272 25443 7330 25449
rect 7742 25440 7748 25452
rect 7800 25440 7806 25492
rect 8754 25440 8760 25492
rect 8812 25440 8818 25492
rect 18874 25480 18880 25492
rect 18156 25452 18880 25480
rect 18156 25424 18184 25452
rect 18874 25440 18880 25452
rect 18932 25440 18938 25492
rect 18138 25372 18144 25424
rect 18196 25372 18202 25424
rect 18616 25384 19748 25412
rect 1857 25347 1915 25353
rect 1857 25313 1869 25347
rect 1903 25344 1915 25347
rect 4154 25344 4160 25356
rect 1903 25316 4160 25344
rect 1903 25313 1915 25316
rect 1857 25307 1915 25313
rect 4154 25304 4160 25316
rect 4212 25344 4218 25356
rect 4212 25316 4752 25344
rect 4212 25304 4218 25316
rect 4338 25236 4344 25288
rect 4396 25276 4402 25288
rect 4433 25279 4491 25285
rect 4433 25276 4445 25279
rect 4396 25248 4445 25276
rect 4396 25236 4402 25248
rect 4433 25245 4445 25248
rect 4479 25245 4491 25279
rect 4433 25239 4491 25245
rect 4614 25236 4620 25288
rect 4672 25236 4678 25288
rect 4724 25285 4752 25316
rect 4982 25304 4988 25356
rect 5040 25304 5046 25356
rect 5442 25304 5448 25356
rect 5500 25344 5506 25356
rect 7009 25347 7067 25353
rect 5500 25316 6592 25344
rect 5500 25304 5506 25316
rect 4709 25279 4767 25285
rect 4709 25245 4721 25279
rect 4755 25245 4767 25279
rect 4709 25239 4767 25245
rect 6564 25276 6592 25316
rect 7009 25313 7021 25347
rect 7055 25344 7067 25347
rect 7055 25316 9168 25344
rect 7055 25313 7067 25316
rect 7009 25307 7067 25313
rect 9140 25288 9168 25316
rect 13446 25304 13452 25356
rect 13504 25344 13510 25356
rect 15010 25344 15016 25356
rect 13504 25316 15016 25344
rect 13504 25304 13510 25316
rect 15010 25304 15016 25316
rect 15068 25304 15074 25356
rect 17770 25344 17776 25356
rect 16408 25316 17776 25344
rect 6564 25248 6868 25276
rect 2133 25211 2191 25217
rect 2133 25177 2145 25211
rect 2179 25177 2191 25211
rect 4724 25208 4752 25239
rect 4890 25208 4896 25220
rect 3358 25180 4568 25208
rect 4724 25180 4896 25208
rect 2133 25171 2191 25177
rect 2148 25140 2176 25171
rect 4540 25152 4568 25180
rect 4890 25168 4896 25180
rect 4948 25168 4954 25220
rect 5534 25168 5540 25220
rect 5592 25168 5598 25220
rect 6564 25217 6592 25248
rect 6549 25211 6607 25217
rect 6549 25177 6561 25211
rect 6595 25177 6607 25211
rect 6840 25208 6868 25248
rect 8386 25236 8392 25288
rect 8444 25236 8450 25288
rect 9122 25236 9128 25288
rect 9180 25236 9186 25288
rect 12069 25279 12127 25285
rect 12069 25245 12081 25279
rect 12115 25276 12127 25279
rect 12986 25276 12992 25288
rect 12115 25248 12992 25276
rect 12115 25245 12127 25248
rect 12069 25239 12127 25245
rect 12986 25236 12992 25248
rect 13044 25236 13050 25288
rect 16408 25262 16436 25316
rect 17770 25304 17776 25316
rect 17828 25304 17834 25356
rect 17862 25276 17868 25288
rect 16592 25248 17868 25276
rect 16592 25220 16620 25248
rect 17862 25236 17868 25248
rect 17920 25276 17926 25288
rect 18616 25285 18644 25384
rect 19720 25356 19748 25384
rect 19242 25344 19248 25356
rect 18708 25316 19248 25344
rect 18708 25285 18736 25316
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 19352 25316 19656 25344
rect 18141 25279 18199 25285
rect 18141 25276 18153 25279
rect 17920 25248 18153 25276
rect 17920 25236 17926 25248
rect 18141 25245 18153 25248
rect 18187 25245 18199 25279
rect 18141 25239 18199 25245
rect 18601 25279 18659 25285
rect 18601 25245 18613 25279
rect 18647 25245 18659 25279
rect 18601 25239 18659 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25245 18751 25279
rect 18693 25239 18751 25245
rect 18782 25236 18788 25288
rect 18840 25236 18846 25288
rect 18874 25236 18880 25288
rect 18932 25285 18938 25288
rect 18932 25279 18961 25285
rect 18949 25245 18961 25279
rect 18932 25239 18961 25245
rect 18932 25236 18938 25239
rect 19058 25236 19064 25288
rect 19116 25236 19122 25288
rect 19352 25285 19380 25316
rect 19337 25279 19395 25285
rect 19337 25245 19349 25279
rect 19383 25245 19395 25279
rect 19337 25239 19395 25245
rect 19518 25236 19524 25288
rect 19576 25236 19582 25288
rect 19628 25276 19656 25316
rect 19702 25304 19708 25356
rect 19760 25304 19766 25356
rect 19886 25304 19892 25356
rect 19944 25344 19950 25356
rect 20349 25347 20407 25353
rect 20349 25344 20361 25347
rect 19944 25316 20361 25344
rect 19944 25304 19950 25316
rect 20349 25313 20361 25316
rect 20395 25344 20407 25347
rect 20625 25347 20683 25353
rect 20625 25344 20637 25347
rect 20395 25316 20637 25344
rect 20395 25313 20407 25316
rect 20349 25307 20407 25313
rect 20625 25313 20637 25316
rect 20671 25313 20683 25347
rect 20625 25307 20683 25313
rect 20901 25347 20959 25353
rect 20901 25313 20913 25347
rect 20947 25344 20959 25347
rect 21910 25344 21916 25356
rect 20947 25316 21916 25344
rect 20947 25313 20959 25316
rect 20901 25307 20959 25313
rect 21910 25304 21916 25316
rect 21968 25304 21974 25356
rect 19794 25276 19800 25288
rect 19628 25248 19800 25276
rect 19794 25236 19800 25248
rect 19852 25276 19858 25288
rect 19852 25248 20208 25276
rect 19852 25236 19858 25248
rect 7190 25208 7196 25220
rect 6840 25180 7196 25208
rect 6549 25171 6607 25177
rect 7190 25168 7196 25180
rect 7248 25168 7254 25220
rect 14918 25168 14924 25220
rect 14976 25208 14982 25220
rect 15289 25211 15347 25217
rect 15289 25208 15301 25211
rect 14976 25180 15301 25208
rect 14976 25168 14982 25180
rect 15289 25177 15301 25180
rect 15335 25177 15347 25211
rect 15289 25171 15347 25177
rect 16574 25168 16580 25220
rect 16632 25168 16638 25220
rect 16945 25211 17003 25217
rect 16945 25208 16957 25211
rect 16776 25180 16957 25208
rect 3050 25140 3056 25152
rect 2148 25112 3056 25140
rect 3050 25100 3056 25112
rect 3108 25100 3114 25152
rect 4522 25100 4528 25152
rect 4580 25100 4586 25152
rect 4617 25143 4675 25149
rect 4617 25109 4629 25143
rect 4663 25140 4675 25143
rect 4798 25140 4804 25152
rect 4663 25112 4804 25140
rect 4663 25109 4675 25112
rect 4617 25103 4675 25109
rect 4798 25100 4804 25112
rect 4856 25100 4862 25152
rect 5074 25100 5080 25152
rect 5132 25140 5138 25152
rect 5350 25140 5356 25152
rect 5132 25112 5356 25140
rect 5132 25100 5138 25112
rect 5350 25100 5356 25112
rect 5408 25100 5414 25152
rect 6454 25100 6460 25152
rect 6512 25100 6518 25152
rect 6759 25143 6817 25149
rect 6759 25109 6771 25143
rect 6805 25140 6817 25143
rect 7374 25140 7380 25152
rect 6805 25112 7380 25140
rect 6805 25109 6817 25112
rect 6759 25103 6817 25109
rect 7374 25100 7380 25112
rect 7432 25100 7438 25152
rect 11882 25100 11888 25152
rect 11940 25100 11946 25152
rect 16776 25149 16804 25180
rect 16945 25177 16957 25180
rect 16991 25177 17003 25211
rect 16945 25171 17003 25177
rect 17402 25168 17408 25220
rect 17460 25208 17466 25220
rect 19613 25211 19671 25217
rect 19613 25208 19625 25211
rect 17460 25180 18552 25208
rect 17460 25168 17466 25180
rect 16761 25143 16819 25149
rect 16761 25109 16773 25143
rect 16807 25109 16819 25143
rect 16761 25103 16819 25109
rect 17034 25100 17040 25152
rect 17092 25100 17098 25152
rect 18414 25100 18420 25152
rect 18472 25100 18478 25152
rect 18524 25140 18552 25180
rect 18892 25180 19625 25208
rect 18892 25140 18920 25180
rect 19613 25177 19625 25180
rect 19659 25177 19671 25211
rect 19613 25171 19671 25177
rect 20180 25152 20208 25248
rect 20254 25236 20260 25288
rect 20312 25236 20318 25288
rect 20272 25208 20300 25236
rect 21174 25208 21180 25220
rect 20272 25180 21180 25208
rect 21174 25168 21180 25180
rect 21232 25208 21238 25220
rect 21232 25180 21390 25208
rect 21232 25168 21238 25180
rect 22278 25168 22284 25220
rect 22336 25208 22342 25220
rect 22649 25211 22707 25217
rect 22649 25208 22661 25211
rect 22336 25180 22661 25208
rect 22336 25168 22342 25180
rect 22649 25177 22661 25180
rect 22695 25177 22707 25211
rect 22649 25171 22707 25177
rect 18524 25112 18920 25140
rect 19150 25100 19156 25152
rect 19208 25140 19214 25152
rect 19429 25143 19487 25149
rect 19429 25140 19441 25143
rect 19208 25112 19441 25140
rect 19208 25100 19214 25112
rect 19429 25109 19441 25112
rect 19475 25109 19487 25143
rect 19429 25103 19487 25109
rect 19518 25100 19524 25152
rect 19576 25140 19582 25152
rect 19978 25140 19984 25152
rect 19576 25112 19984 25140
rect 19576 25100 19582 25112
rect 19978 25100 19984 25112
rect 20036 25100 20042 25152
rect 20162 25100 20168 25152
rect 20220 25100 20226 25152
rect 1104 25050 29440 25072
rect 1104 24998 5151 25050
rect 5203 24998 5215 25050
rect 5267 24998 5279 25050
rect 5331 24998 5343 25050
rect 5395 24998 5407 25050
rect 5459 24998 12234 25050
rect 12286 24998 12298 25050
rect 12350 24998 12362 25050
rect 12414 24998 12426 25050
rect 12478 24998 12490 25050
rect 12542 24998 19317 25050
rect 19369 24998 19381 25050
rect 19433 24998 19445 25050
rect 19497 24998 19509 25050
rect 19561 24998 19573 25050
rect 19625 24998 26400 25050
rect 26452 24998 26464 25050
rect 26516 24998 26528 25050
rect 26580 24998 26592 25050
rect 26644 24998 26656 25050
rect 26708 24998 29440 25050
rect 1104 24976 29440 24998
rect 4890 24936 4896 24948
rect 3160 24908 4896 24936
rect 3160 24809 3188 24908
rect 4890 24896 4896 24908
rect 4948 24896 4954 24948
rect 5718 24896 5724 24948
rect 5776 24896 5782 24948
rect 6454 24896 6460 24948
rect 6512 24936 6518 24948
rect 7377 24939 7435 24945
rect 7377 24936 7389 24939
rect 6512 24908 7389 24936
rect 6512 24896 6518 24908
rect 7377 24905 7389 24908
rect 7423 24905 7435 24939
rect 7377 24899 7435 24905
rect 7558 24896 7564 24948
rect 7616 24896 7622 24948
rect 14918 24896 14924 24948
rect 14976 24896 14982 24948
rect 15286 24896 15292 24948
rect 15344 24936 15350 24948
rect 16114 24936 16120 24948
rect 15344 24908 16120 24936
rect 15344 24896 15350 24908
rect 16114 24896 16120 24908
rect 16172 24896 16178 24948
rect 19058 24936 19064 24948
rect 17972 24908 19064 24936
rect 4798 24828 4804 24880
rect 4856 24868 4862 24880
rect 4856 24840 5212 24868
rect 4856 24828 4862 24840
rect 3145 24803 3203 24809
rect 3145 24769 3157 24803
rect 3191 24769 3203 24803
rect 3145 24763 3203 24769
rect 4522 24760 4528 24812
rect 4580 24760 4586 24812
rect 5074 24800 5080 24812
rect 4908 24772 5080 24800
rect 3418 24692 3424 24744
rect 3476 24692 3482 24744
rect 4540 24664 4568 24760
rect 4614 24692 4620 24744
rect 4672 24732 4678 24744
rect 4908 24741 4936 24772
rect 5074 24760 5080 24772
rect 5132 24760 5138 24812
rect 5184 24809 5212 24840
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24769 5227 24803
rect 5626 24800 5632 24812
rect 5169 24763 5227 24769
rect 5460 24772 5632 24800
rect 4893 24735 4951 24741
rect 4893 24732 4905 24735
rect 4672 24704 4905 24732
rect 4672 24692 4678 24704
rect 4893 24701 4905 24704
rect 4939 24701 4951 24735
rect 4893 24695 4951 24701
rect 4985 24735 5043 24741
rect 4985 24701 4997 24735
rect 5031 24732 5043 24735
rect 5460 24732 5488 24772
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 5031 24704 5488 24732
rect 5537 24735 5595 24741
rect 5031 24701 5043 24704
rect 4985 24695 5043 24701
rect 5537 24701 5549 24735
rect 5583 24732 5595 24735
rect 5736 24732 5764 24896
rect 7101 24871 7159 24877
rect 7101 24837 7113 24871
rect 7147 24868 7159 24871
rect 7190 24868 7196 24880
rect 7147 24840 7196 24868
rect 7147 24837 7159 24840
rect 7101 24831 7159 24837
rect 7190 24828 7196 24840
rect 7248 24828 7254 24880
rect 7285 24871 7343 24877
rect 7285 24837 7297 24871
rect 7331 24868 7343 24871
rect 7576 24868 7604 24896
rect 9582 24868 9588 24880
rect 7331 24840 7604 24868
rect 9338 24840 9588 24868
rect 7331 24837 7343 24840
rect 7285 24831 7343 24837
rect 9582 24828 9588 24840
rect 9640 24828 9646 24880
rect 11793 24871 11851 24877
rect 11793 24837 11805 24871
rect 11839 24868 11851 24871
rect 11882 24868 11888 24880
rect 11839 24840 11888 24868
rect 11839 24837 11851 24840
rect 11793 24831 11851 24837
rect 11882 24828 11888 24840
rect 11940 24828 11946 24880
rect 14090 24868 14096 24880
rect 13018 24854 14096 24868
rect 13004 24840 14096 24854
rect 6362 24760 6368 24812
rect 6420 24760 6426 24812
rect 7374 24760 7380 24812
rect 7432 24800 7438 24812
rect 7469 24803 7527 24809
rect 7469 24800 7481 24803
rect 7432 24772 7481 24800
rect 7432 24760 7438 24772
rect 7469 24769 7481 24772
rect 7515 24769 7527 24803
rect 7469 24763 7527 24769
rect 7650 24760 7656 24812
rect 7708 24760 7714 24812
rect 9677 24803 9735 24809
rect 9677 24800 9689 24803
rect 9324 24772 9689 24800
rect 6638 24732 6644 24744
rect 5583 24704 6644 24732
rect 5583 24701 5595 24704
rect 5537 24695 5595 24701
rect 6638 24692 6644 24704
rect 6696 24692 6702 24744
rect 7009 24735 7067 24741
rect 7009 24701 7021 24735
rect 7055 24732 7067 24735
rect 7055 24704 7788 24732
rect 7055 24701 7067 24704
rect 7009 24695 7067 24701
rect 5074 24664 5080 24676
rect 4540 24636 5080 24664
rect 5074 24624 5080 24636
rect 5132 24664 5138 24676
rect 6181 24667 6239 24673
rect 5132 24636 5580 24664
rect 5132 24624 5138 24636
rect 5552 24608 5580 24636
rect 6181 24633 6193 24667
rect 6227 24664 6239 24667
rect 6914 24664 6920 24676
rect 6227 24636 6920 24664
rect 6227 24633 6239 24636
rect 6181 24627 6239 24633
rect 6914 24624 6920 24636
rect 6972 24624 6978 24676
rect 7760 24664 7788 24704
rect 7834 24692 7840 24744
rect 7892 24692 7898 24744
rect 8113 24735 8171 24741
rect 8113 24732 8125 24735
rect 7944 24704 8125 24732
rect 7944 24664 7972 24704
rect 8113 24701 8125 24704
rect 8159 24701 8171 24735
rect 8113 24695 8171 24701
rect 7760 24636 7972 24664
rect 5166 24556 5172 24608
rect 5224 24596 5230 24608
rect 5353 24599 5411 24605
rect 5353 24596 5365 24599
rect 5224 24568 5365 24596
rect 5224 24556 5230 24568
rect 5353 24565 5365 24568
rect 5399 24565 5411 24599
rect 5353 24559 5411 24565
rect 5534 24556 5540 24608
rect 5592 24556 5598 24608
rect 6362 24556 6368 24608
rect 6420 24596 6426 24608
rect 9324 24596 9352 24772
rect 9677 24769 9689 24772
rect 9723 24769 9735 24803
rect 9677 24763 9735 24769
rect 11422 24760 11428 24812
rect 11480 24800 11486 24812
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 11480 24772 11529 24800
rect 11480 24760 11486 24772
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 10594 24692 10600 24744
rect 10652 24732 10658 24744
rect 13004 24732 13032 24840
rect 14090 24828 14096 24840
rect 14148 24828 14154 24880
rect 14185 24871 14243 24877
rect 14185 24837 14197 24871
rect 14231 24868 14243 24871
rect 15562 24868 15568 24880
rect 14231 24840 15568 24868
rect 14231 24837 14243 24840
rect 14185 24831 14243 24837
rect 15562 24828 15568 24840
rect 15620 24828 15626 24880
rect 17034 24868 17040 24880
rect 16040 24840 16252 24868
rect 14108 24800 14136 24828
rect 16040 24812 16068 24840
rect 14274 24800 14280 24812
rect 14108 24772 14280 24800
rect 14274 24760 14280 24772
rect 14332 24760 14338 24812
rect 15105 24803 15163 24809
rect 15105 24769 15117 24803
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 15197 24803 15255 24809
rect 15197 24769 15209 24803
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 10652 24704 13032 24732
rect 13541 24735 13599 24741
rect 10652 24692 10658 24704
rect 13541 24701 13553 24735
rect 13587 24732 13599 24735
rect 13722 24732 13728 24744
rect 13587 24704 13728 24732
rect 13587 24701 13599 24704
rect 13541 24695 13599 24701
rect 13722 24692 13728 24704
rect 13780 24692 13786 24744
rect 14369 24735 14427 24741
rect 14369 24701 14381 24735
rect 14415 24701 14427 24735
rect 14369 24695 14427 24701
rect 6420 24568 9352 24596
rect 9585 24599 9643 24605
rect 6420 24556 6426 24568
rect 9585 24565 9597 24599
rect 9631 24596 9643 24599
rect 9769 24599 9827 24605
rect 9769 24596 9781 24599
rect 9631 24568 9781 24596
rect 9631 24565 9643 24568
rect 9585 24559 9643 24565
rect 9769 24565 9781 24568
rect 9815 24565 9827 24599
rect 9769 24559 9827 24565
rect 10137 24599 10195 24605
rect 10137 24565 10149 24599
rect 10183 24596 10195 24599
rect 10410 24596 10416 24608
rect 10183 24568 10416 24596
rect 10183 24565 10195 24568
rect 10137 24559 10195 24565
rect 10410 24556 10416 24568
rect 10468 24556 10474 24608
rect 14384 24596 14412 24695
rect 14458 24692 14464 24744
rect 14516 24692 14522 24744
rect 14550 24692 14556 24744
rect 14608 24692 14614 24744
rect 14918 24624 14924 24676
rect 14976 24664 14982 24676
rect 15120 24664 15148 24763
rect 15212 24732 15240 24763
rect 15286 24760 15292 24812
rect 15344 24760 15350 24812
rect 15378 24760 15384 24812
rect 15436 24809 15442 24812
rect 15436 24803 15465 24809
rect 15453 24769 15465 24803
rect 15436 24763 15465 24769
rect 15436 24760 15442 24763
rect 15654 24760 15660 24812
rect 15712 24760 15718 24812
rect 15841 24803 15899 24809
rect 15841 24769 15853 24803
rect 15887 24800 15899 24803
rect 16022 24800 16028 24812
rect 15887 24772 16028 24800
rect 15887 24769 15899 24772
rect 15841 24763 15899 24769
rect 15565 24735 15623 24741
rect 15212 24704 15332 24732
rect 15304 24664 15332 24704
rect 15565 24701 15577 24735
rect 15611 24732 15623 24735
rect 15856 24732 15884 24763
rect 16022 24760 16028 24772
rect 16080 24760 16086 24812
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24769 16175 24803
rect 16224 24800 16252 24840
rect 16776 24840 17040 24868
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 16224 24772 16313 24800
rect 16117 24763 16175 24769
rect 16301 24769 16313 24772
rect 16347 24800 16359 24803
rect 16776 24800 16804 24840
rect 17034 24828 17040 24840
rect 17092 24828 17098 24880
rect 17972 24868 18000 24908
rect 19058 24896 19064 24908
rect 19116 24896 19122 24948
rect 17880 24840 18000 24868
rect 18049 24871 18107 24877
rect 17880 24809 17908 24840
rect 18049 24837 18061 24871
rect 18095 24868 18107 24871
rect 18322 24868 18328 24880
rect 18095 24840 18328 24868
rect 18095 24837 18107 24840
rect 18049 24831 18107 24837
rect 18322 24828 18328 24840
rect 18380 24828 18386 24880
rect 18414 24828 18420 24880
rect 18472 24868 18478 24880
rect 18693 24871 18751 24877
rect 18693 24868 18705 24871
rect 18472 24840 18705 24868
rect 18472 24828 18478 24840
rect 18693 24837 18705 24840
rect 18739 24837 18751 24871
rect 18693 24831 18751 24837
rect 20162 24828 20168 24880
rect 20220 24868 20226 24880
rect 22278 24868 22284 24880
rect 20220 24840 22284 24868
rect 20220 24828 20226 24840
rect 22278 24828 22284 24840
rect 22336 24828 22342 24880
rect 16347 24772 16804 24800
rect 16861 24803 16919 24809
rect 16347 24769 16359 24772
rect 16301 24763 16359 24769
rect 16861 24769 16873 24803
rect 16907 24800 16919 24803
rect 17865 24803 17923 24809
rect 16907 24772 16988 24800
rect 16907 24769 16919 24772
rect 16861 24763 16919 24769
rect 15611 24704 15884 24732
rect 15611 24701 15623 24704
rect 15565 24695 15623 24701
rect 15930 24692 15936 24744
rect 15988 24732 15994 24744
rect 16132 24732 16160 24763
rect 16960 24744 16988 24772
rect 17865 24769 17877 24803
rect 17911 24769 17923 24803
rect 17865 24763 17923 24769
rect 17954 24760 17960 24812
rect 18012 24760 18018 24812
rect 18138 24760 18144 24812
rect 18196 24809 18202 24812
rect 18196 24803 18225 24809
rect 18213 24769 18225 24803
rect 18196 24763 18225 24769
rect 18196 24760 18202 24763
rect 19794 24760 19800 24812
rect 19852 24800 19858 24812
rect 20070 24800 20076 24812
rect 19852 24772 20076 24800
rect 19852 24760 19858 24772
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20349 24803 20407 24809
rect 20349 24800 20361 24803
rect 20180 24772 20361 24800
rect 16942 24732 16948 24744
rect 15988 24704 16948 24732
rect 15988 24692 15994 24704
rect 16942 24692 16948 24704
rect 17000 24692 17006 24744
rect 18325 24735 18383 24741
rect 18325 24732 18337 24735
rect 17604 24704 18337 24732
rect 16025 24667 16083 24673
rect 16025 24664 16037 24667
rect 14976 24636 15240 24664
rect 15304 24636 16037 24664
rect 14976 24624 14982 24636
rect 15102 24596 15108 24608
rect 14384 24568 15108 24596
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 15212 24596 15240 24636
rect 16025 24633 16037 24636
rect 16071 24633 16083 24667
rect 16025 24627 16083 24633
rect 17604 24608 17632 24704
rect 18325 24701 18337 24704
rect 18371 24701 18383 24735
rect 18325 24695 18383 24701
rect 18417 24735 18475 24741
rect 18417 24701 18429 24735
rect 18463 24732 18475 24735
rect 19886 24732 19892 24744
rect 18463 24704 19892 24732
rect 18463 24701 18475 24704
rect 18417 24695 18475 24701
rect 19886 24692 19892 24704
rect 19944 24692 19950 24744
rect 19978 24692 19984 24744
rect 20036 24692 20042 24744
rect 20180 24741 20208 24772
rect 20349 24769 20361 24772
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 20714 24760 20720 24812
rect 20772 24800 20778 24812
rect 20809 24803 20867 24809
rect 20809 24800 20821 24803
rect 20772 24772 20821 24800
rect 20772 24760 20778 24772
rect 20809 24769 20821 24772
rect 20855 24769 20867 24803
rect 20809 24763 20867 24769
rect 20165 24735 20223 24741
rect 20165 24701 20177 24735
rect 20211 24701 20223 24735
rect 20165 24695 20223 24701
rect 20993 24735 21051 24741
rect 20993 24701 21005 24735
rect 21039 24701 21051 24735
rect 20993 24695 21051 24701
rect 17681 24667 17739 24673
rect 17681 24633 17693 24667
rect 17727 24664 17739 24667
rect 18230 24664 18236 24676
rect 17727 24636 18236 24664
rect 17727 24633 17739 24636
rect 17681 24627 17739 24633
rect 18230 24624 18236 24636
rect 18288 24624 18294 24676
rect 19996 24664 20024 24692
rect 21008 24664 21036 24695
rect 19996 24636 21036 24664
rect 16209 24599 16267 24605
rect 16209 24596 16221 24599
rect 15212 24568 16221 24596
rect 16209 24565 16221 24568
rect 16255 24565 16267 24599
rect 16209 24559 16267 24565
rect 16298 24556 16304 24608
rect 16356 24596 16362 24608
rect 16945 24599 17003 24605
rect 16945 24596 16957 24599
rect 16356 24568 16957 24596
rect 16356 24556 16362 24568
rect 16945 24565 16957 24568
rect 16991 24565 17003 24599
rect 16945 24559 17003 24565
rect 17586 24556 17592 24608
rect 17644 24556 17650 24608
rect 20070 24556 20076 24608
rect 20128 24596 20134 24608
rect 20441 24599 20499 24605
rect 20441 24596 20453 24599
rect 20128 24568 20453 24596
rect 20128 24556 20134 24568
rect 20441 24565 20453 24568
rect 20487 24565 20499 24599
rect 20441 24559 20499 24565
rect 1104 24506 29440 24528
rect 1104 24454 4491 24506
rect 4543 24454 4555 24506
rect 4607 24454 4619 24506
rect 4671 24454 4683 24506
rect 4735 24454 4747 24506
rect 4799 24454 11574 24506
rect 11626 24454 11638 24506
rect 11690 24454 11702 24506
rect 11754 24454 11766 24506
rect 11818 24454 11830 24506
rect 11882 24454 18657 24506
rect 18709 24454 18721 24506
rect 18773 24454 18785 24506
rect 18837 24454 18849 24506
rect 18901 24454 18913 24506
rect 18965 24454 25740 24506
rect 25792 24454 25804 24506
rect 25856 24454 25868 24506
rect 25920 24454 25932 24506
rect 25984 24454 25996 24506
rect 26048 24454 29440 24506
rect 1104 24432 29440 24454
rect 3418 24352 3424 24404
rect 3476 24392 3482 24404
rect 4065 24395 4123 24401
rect 4065 24392 4077 24395
rect 3476 24364 4077 24392
rect 3476 24352 3482 24364
rect 4065 24361 4077 24364
rect 4111 24361 4123 24395
rect 4065 24355 4123 24361
rect 4982 24352 4988 24404
rect 5040 24392 5046 24404
rect 5040 24364 6592 24392
rect 5040 24352 5046 24364
rect 5166 24324 5172 24336
rect 4264 24296 5172 24324
rect 4264 24197 4292 24296
rect 5166 24284 5172 24296
rect 5224 24284 5230 24336
rect 6564 24324 6592 24364
rect 6638 24352 6644 24404
rect 6696 24392 6702 24404
rect 7009 24395 7067 24401
rect 7009 24392 7021 24395
rect 6696 24364 7021 24392
rect 6696 24352 6702 24364
rect 7009 24361 7021 24364
rect 7055 24392 7067 24395
rect 7374 24392 7380 24404
rect 7055 24364 7380 24392
rect 7055 24361 7067 24364
rect 7009 24355 7067 24361
rect 7374 24352 7380 24364
rect 7432 24352 7438 24404
rect 7650 24352 7656 24404
rect 7708 24352 7714 24404
rect 14458 24392 14464 24404
rect 13188 24364 14464 24392
rect 7668 24324 7696 24352
rect 13188 24336 13216 24364
rect 14458 24352 14464 24364
rect 14516 24352 14522 24404
rect 15286 24352 15292 24404
rect 15344 24392 15350 24404
rect 15654 24392 15660 24404
rect 15344 24364 15660 24392
rect 15344 24352 15350 24364
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 15838 24352 15844 24404
rect 15896 24392 15902 24404
rect 16650 24395 16708 24401
rect 16650 24392 16662 24395
rect 15896 24364 16662 24392
rect 15896 24352 15902 24364
rect 16650 24361 16662 24364
rect 16696 24361 16708 24395
rect 16650 24355 16708 24361
rect 19242 24352 19248 24404
rect 19300 24352 19306 24404
rect 19702 24352 19708 24404
rect 19760 24392 19766 24404
rect 19889 24395 19947 24401
rect 19889 24392 19901 24395
rect 19760 24364 19901 24392
rect 19760 24352 19766 24364
rect 19889 24361 19901 24364
rect 19935 24361 19947 24395
rect 19889 24355 19947 24361
rect 6564 24296 7696 24324
rect 13170 24284 13176 24336
rect 13228 24284 13234 24336
rect 16206 24284 16212 24336
rect 16264 24284 16270 24336
rect 16316 24296 16528 24324
rect 4890 24216 4896 24268
rect 4948 24256 4954 24268
rect 5261 24259 5319 24265
rect 5261 24256 5273 24259
rect 4948 24228 5273 24256
rect 4948 24216 4954 24228
rect 5261 24225 5273 24228
rect 5307 24256 5319 24259
rect 7834 24256 7840 24268
rect 5307 24228 7840 24256
rect 5307 24225 5319 24228
rect 5261 24219 5319 24225
rect 6564 24200 6592 24228
rect 7834 24216 7840 24228
rect 7892 24216 7898 24268
rect 11609 24259 11667 24265
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 15010 24256 15016 24268
rect 11655 24228 15016 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 15010 24216 15016 24228
rect 15068 24256 15074 24268
rect 15289 24259 15347 24265
rect 15289 24256 15301 24259
rect 15068 24228 15301 24256
rect 15068 24216 15074 24228
rect 15289 24225 15301 24228
rect 15335 24225 15347 24259
rect 16224 24256 16252 24284
rect 16316 24265 16344 24296
rect 15289 24219 15347 24225
rect 15764 24228 16252 24256
rect 16301 24259 16359 24265
rect 4249 24191 4307 24197
rect 4249 24157 4261 24191
rect 4295 24157 4307 24191
rect 4249 24151 4307 24157
rect 6546 24148 6552 24200
rect 6604 24148 6610 24200
rect 7006 24148 7012 24200
rect 7064 24188 7070 24200
rect 7101 24191 7159 24197
rect 7101 24188 7113 24191
rect 7064 24160 7113 24188
rect 7064 24148 7070 24160
rect 7101 24157 7113 24160
rect 7147 24157 7159 24191
rect 7101 24151 7159 24157
rect 7282 24148 7288 24200
rect 7340 24148 7346 24200
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24188 10103 24191
rect 10778 24188 10784 24200
rect 10091 24160 10784 24188
rect 10091 24157 10103 24160
rect 10045 24151 10103 24157
rect 10778 24148 10784 24160
rect 10836 24148 10842 24200
rect 13906 24188 13912 24200
rect 13556 24160 13912 24188
rect 13556 24132 13584 24160
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 15764 24188 15792 24228
rect 16301 24225 16313 24259
rect 16347 24225 16359 24259
rect 16301 24219 16359 24225
rect 16390 24216 16396 24268
rect 16448 24216 16454 24268
rect 16500 24256 16528 24296
rect 17218 24256 17224 24268
rect 16500 24228 17224 24256
rect 17218 24216 17224 24228
rect 17276 24216 17282 24268
rect 19812 24228 20208 24256
rect 16206 24197 16212 24200
rect 15841 24191 15899 24197
rect 15841 24188 15853 24191
rect 15764 24160 15853 24188
rect 15841 24157 15853 24160
rect 15887 24157 15899 24191
rect 15841 24151 15899 24157
rect 16163 24191 16212 24197
rect 16163 24157 16175 24191
rect 16209 24157 16212 24191
rect 16163 24151 16212 24157
rect 16206 24148 16212 24151
rect 16264 24148 16270 24200
rect 17770 24148 17776 24200
rect 17828 24148 17834 24200
rect 19058 24148 19064 24200
rect 19116 24188 19122 24200
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 19116 24160 19441 24188
rect 19116 24148 19122 24160
rect 19429 24157 19441 24160
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 5537 24123 5595 24129
rect 5537 24089 5549 24123
rect 5583 24089 5595 24123
rect 5537 24083 5595 24089
rect 5552 24052 5580 24083
rect 5626 24080 5632 24132
rect 5684 24120 5690 24132
rect 7193 24123 7251 24129
rect 7193 24120 7205 24123
rect 5684 24092 6026 24120
rect 6840 24092 7205 24120
rect 5684 24080 5690 24092
rect 6840 24052 6868 24092
rect 7193 24089 7205 24092
rect 7239 24089 7251 24123
rect 7193 24083 7251 24089
rect 11790 24080 11796 24132
rect 11848 24080 11854 24132
rect 11882 24080 11888 24132
rect 11940 24080 11946 24132
rect 13538 24120 13544 24132
rect 13110 24092 13544 24120
rect 13538 24080 13544 24092
rect 13596 24080 13602 24132
rect 13633 24123 13691 24129
rect 13633 24089 13645 24123
rect 13679 24089 13691 24123
rect 13633 24083 13691 24089
rect 14553 24123 14611 24129
rect 14553 24089 14565 24123
rect 14599 24120 14611 24123
rect 15102 24120 15108 24132
rect 14599 24092 15108 24120
rect 14599 24089 14611 24092
rect 14553 24083 14611 24089
rect 5552 24024 6868 24052
rect 9674 24012 9680 24064
rect 9732 24052 9738 24064
rect 10597 24055 10655 24061
rect 10597 24052 10609 24055
rect 9732 24024 10609 24052
rect 9732 24012 9738 24024
rect 10597 24021 10609 24024
rect 10643 24021 10655 24055
rect 11808 24052 11836 24080
rect 13648 24052 13676 24083
rect 15102 24080 15108 24092
rect 15160 24080 15166 24132
rect 15933 24123 15991 24129
rect 15933 24089 15945 24123
rect 15979 24089 15991 24123
rect 15933 24083 15991 24089
rect 14274 24052 14280 24064
rect 11808 24024 14280 24052
rect 10597 24015 10655 24021
rect 14274 24012 14280 24024
rect 14332 24012 14338 24064
rect 15657 24055 15715 24061
rect 15657 24021 15669 24055
rect 15703 24052 15715 24055
rect 15838 24052 15844 24064
rect 15703 24024 15844 24052
rect 15703 24021 15715 24024
rect 15657 24015 15715 24021
rect 15838 24012 15844 24024
rect 15896 24012 15902 24064
rect 15948 24052 15976 24083
rect 16022 24080 16028 24132
rect 16080 24080 16086 24132
rect 18046 24080 18052 24132
rect 18104 24120 18110 24132
rect 18417 24123 18475 24129
rect 18417 24120 18429 24123
rect 18104 24092 18429 24120
rect 18104 24080 18110 24092
rect 18417 24089 18429 24092
rect 18463 24089 18475 24123
rect 19444 24120 19472 24151
rect 19702 24148 19708 24200
rect 19760 24188 19766 24200
rect 19812 24197 19840 24228
rect 20180 24200 20208 24228
rect 19797 24191 19855 24197
rect 19797 24188 19809 24191
rect 19760 24160 19809 24188
rect 19760 24148 19766 24160
rect 19797 24157 19809 24160
rect 19843 24157 19855 24191
rect 20073 24191 20131 24197
rect 20073 24188 20085 24191
rect 19797 24151 19855 24157
rect 19904 24160 20085 24188
rect 19904 24120 19932 24160
rect 20073 24157 20085 24160
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 19444 24092 19932 24120
rect 18417 24083 18475 24089
rect 19978 24080 19984 24132
rect 20036 24080 20042 24132
rect 16758 24052 16764 24064
rect 15948 24024 16764 24052
rect 16758 24012 16764 24024
rect 16816 24012 16822 24064
rect 17586 24012 17592 24064
rect 17644 24052 17650 24064
rect 19613 24055 19671 24061
rect 19613 24052 19625 24055
rect 17644 24024 19625 24052
rect 17644 24012 17650 24024
rect 19613 24021 19625 24024
rect 19659 24052 19671 24055
rect 19996 24052 20024 24080
rect 20088 24064 20116 24151
rect 20162 24148 20168 24200
rect 20220 24148 20226 24200
rect 19659 24024 20024 24052
rect 19659 24021 19671 24024
rect 19613 24015 19671 24021
rect 20070 24012 20076 24064
rect 20128 24012 20134 24064
rect 1104 23962 29440 23984
rect 1104 23910 5151 23962
rect 5203 23910 5215 23962
rect 5267 23910 5279 23962
rect 5331 23910 5343 23962
rect 5395 23910 5407 23962
rect 5459 23910 12234 23962
rect 12286 23910 12298 23962
rect 12350 23910 12362 23962
rect 12414 23910 12426 23962
rect 12478 23910 12490 23962
rect 12542 23910 19317 23962
rect 19369 23910 19381 23962
rect 19433 23910 19445 23962
rect 19497 23910 19509 23962
rect 19561 23910 19573 23962
rect 19625 23910 26400 23962
rect 26452 23910 26464 23962
rect 26516 23910 26528 23962
rect 26580 23910 26592 23962
rect 26644 23910 26656 23962
rect 26708 23910 29440 23962
rect 1104 23888 29440 23910
rect 5810 23808 5816 23860
rect 5868 23848 5874 23860
rect 11790 23848 11796 23860
rect 5868 23820 11796 23848
rect 5868 23808 5874 23820
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 11882 23808 11888 23860
rect 11940 23848 11946 23860
rect 11940 23820 12434 23848
rect 11940 23808 11946 23820
rect 12406 23780 12434 23820
rect 12986 23808 12992 23860
rect 13044 23808 13050 23860
rect 14737 23851 14795 23857
rect 14737 23848 14749 23851
rect 13280 23820 14749 23848
rect 13280 23780 13308 23820
rect 14737 23817 14749 23820
rect 14783 23817 14795 23851
rect 14737 23811 14795 23817
rect 15562 23808 15568 23860
rect 15620 23848 15626 23860
rect 15620 23820 15700 23848
rect 15620 23808 15626 23820
rect 15672 23789 15700 23820
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 17589 23851 17647 23857
rect 17589 23848 17601 23851
rect 16816 23820 17601 23848
rect 16816 23808 16822 23820
rect 17589 23817 17601 23820
rect 17635 23817 17647 23851
rect 17589 23811 17647 23817
rect 12406 23752 13308 23780
rect 13357 23783 13415 23789
rect 13357 23749 13369 23783
rect 13403 23749 13415 23783
rect 15657 23783 15715 23789
rect 13357 23743 13415 23749
rect 14844 23752 15608 23780
rect 1486 23672 1492 23724
rect 1544 23672 1550 23724
rect 10594 23672 10600 23724
rect 10652 23672 10658 23724
rect 12802 23712 12808 23724
rect 10980 23684 12808 23712
rect 9122 23604 9128 23656
rect 9180 23644 9186 23656
rect 9217 23647 9275 23653
rect 9217 23644 9229 23647
rect 9180 23616 9229 23644
rect 9180 23604 9186 23616
rect 9217 23613 9229 23616
rect 9263 23613 9275 23647
rect 9217 23607 9275 23613
rect 9493 23647 9551 23653
rect 9493 23613 9505 23647
rect 9539 23644 9551 23647
rect 10980 23644 11008 23684
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 9539 23616 11008 23644
rect 11517 23647 11575 23653
rect 9539 23613 9551 23616
rect 9493 23607 9551 23613
rect 11517 23613 11529 23647
rect 11563 23613 11575 23647
rect 11517 23607 11575 23613
rect 11532 23576 11560 23607
rect 10980 23548 11560 23576
rect 10980 23520 11008 23548
rect 1578 23468 1584 23520
rect 1636 23468 1642 23520
rect 10962 23468 10968 23520
rect 11020 23468 11026 23520
rect 12158 23468 12164 23520
rect 12216 23468 12222 23520
rect 13372 23508 13400 23743
rect 14844 23721 14872 23752
rect 15580 23724 15608 23752
rect 15657 23749 15669 23783
rect 15703 23749 15715 23783
rect 15657 23743 15715 23749
rect 16298 23740 16304 23792
rect 16356 23740 16362 23792
rect 16942 23740 16948 23792
rect 17000 23780 17006 23792
rect 17497 23783 17555 23789
rect 17497 23780 17509 23783
rect 17000 23752 17509 23780
rect 17000 23740 17006 23752
rect 17497 23749 17509 23752
rect 17543 23749 17555 23783
rect 17497 23743 17555 23749
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 14553 23715 14611 23721
rect 14553 23712 14565 23715
rect 13495 23684 14565 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 14553 23681 14565 23684
rect 14599 23681 14611 23715
rect 14553 23675 14611 23681
rect 14829 23715 14887 23721
rect 14829 23681 14841 23715
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 13633 23647 13691 23653
rect 13633 23613 13645 23647
rect 13679 23644 13691 23647
rect 13722 23644 13728 23656
rect 13679 23616 13728 23644
rect 13679 23613 13691 23616
rect 13633 23607 13691 23613
rect 13722 23604 13728 23616
rect 13780 23604 13786 23656
rect 14093 23647 14151 23653
rect 14093 23613 14105 23647
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 14108 23576 14136 23607
rect 14274 23604 14280 23656
rect 14332 23644 14338 23656
rect 14458 23644 14464 23656
rect 14332 23616 14464 23644
rect 14332 23604 14338 23616
rect 14458 23604 14464 23616
rect 14516 23604 14522 23656
rect 14568 23644 14596 23675
rect 15010 23672 15016 23724
rect 15068 23672 15074 23724
rect 15289 23715 15347 23721
rect 15289 23681 15301 23715
rect 15335 23712 15347 23715
rect 15378 23712 15384 23724
rect 15335 23684 15384 23712
rect 15335 23681 15347 23684
rect 15289 23675 15347 23681
rect 15378 23672 15384 23684
rect 15436 23672 15442 23724
rect 15473 23715 15531 23721
rect 15473 23681 15485 23715
rect 15519 23681 15531 23715
rect 15473 23675 15531 23681
rect 15105 23647 15163 23653
rect 15105 23644 15117 23647
rect 14568 23616 15117 23644
rect 15105 23613 15117 23616
rect 15151 23613 15163 23647
rect 15105 23607 15163 23613
rect 15194 23576 15200 23588
rect 14108 23548 15200 23576
rect 15194 23536 15200 23548
rect 15252 23536 15258 23588
rect 14829 23511 14887 23517
rect 14829 23508 14841 23511
rect 13372 23480 14841 23508
rect 14829 23477 14841 23480
rect 14875 23477 14887 23511
rect 15396 23508 15424 23672
rect 15488 23644 15516 23675
rect 15562 23672 15568 23724
rect 15620 23672 15626 23724
rect 16316 23712 16344 23740
rect 17129 23715 17187 23721
rect 17129 23712 17141 23715
rect 16316 23684 17141 23712
rect 17129 23681 17141 23684
rect 17175 23681 17187 23715
rect 17129 23675 17187 23681
rect 16022 23644 16028 23656
rect 15488 23616 16028 23644
rect 16022 23604 16028 23616
rect 16080 23604 16086 23656
rect 17144 23644 17172 23675
rect 17218 23672 17224 23724
rect 17276 23672 17282 23724
rect 17313 23715 17371 23721
rect 17313 23681 17325 23715
rect 17359 23712 17371 23715
rect 17773 23715 17831 23721
rect 17773 23712 17785 23715
rect 17359 23684 17785 23712
rect 17359 23681 17371 23684
rect 17313 23675 17371 23681
rect 17773 23681 17785 23684
rect 17819 23712 17831 23715
rect 19702 23712 19708 23724
rect 17819 23684 19708 23712
rect 17819 23681 17831 23684
rect 17773 23675 17831 23681
rect 19702 23672 19708 23684
rect 19760 23672 19766 23724
rect 17586 23644 17592 23656
rect 17144 23616 17592 23644
rect 17586 23604 17592 23616
rect 17644 23644 17650 23656
rect 17865 23647 17923 23653
rect 17865 23644 17877 23647
rect 17644 23616 17877 23644
rect 17644 23604 17650 23616
rect 17865 23613 17877 23616
rect 17911 23613 17923 23647
rect 17865 23607 17923 23613
rect 17957 23647 18015 23653
rect 17957 23613 17969 23647
rect 18003 23613 18015 23647
rect 17957 23607 18015 23613
rect 15838 23536 15844 23588
rect 15896 23576 15902 23588
rect 15933 23579 15991 23585
rect 15933 23576 15945 23579
rect 15896 23548 15945 23576
rect 15896 23536 15902 23548
rect 15933 23545 15945 23548
rect 15979 23545 15991 23579
rect 15933 23539 15991 23545
rect 16206 23536 16212 23588
rect 16264 23576 16270 23588
rect 16945 23579 17003 23585
rect 16945 23576 16957 23579
rect 16264 23548 16957 23576
rect 16264 23536 16270 23548
rect 16945 23545 16957 23548
rect 16991 23576 17003 23579
rect 17972 23576 18000 23607
rect 18046 23604 18052 23656
rect 18104 23604 18110 23656
rect 19058 23604 19064 23656
rect 19116 23604 19122 23656
rect 19076 23576 19104 23604
rect 16991 23548 19104 23576
rect 16991 23545 17003 23548
rect 16945 23539 17003 23545
rect 19702 23536 19708 23588
rect 19760 23576 19766 23588
rect 19978 23576 19984 23588
rect 19760 23548 19984 23576
rect 19760 23536 19766 23548
rect 19978 23536 19984 23548
rect 20036 23536 20042 23588
rect 16114 23508 16120 23520
rect 15396 23480 16120 23508
rect 14829 23471 14887 23477
rect 16114 23468 16120 23480
rect 16172 23468 16178 23520
rect 1104 23418 29440 23440
rect 1104 23366 4491 23418
rect 4543 23366 4555 23418
rect 4607 23366 4619 23418
rect 4671 23366 4683 23418
rect 4735 23366 4747 23418
rect 4799 23366 11574 23418
rect 11626 23366 11638 23418
rect 11690 23366 11702 23418
rect 11754 23366 11766 23418
rect 11818 23366 11830 23418
rect 11882 23366 18657 23418
rect 18709 23366 18721 23418
rect 18773 23366 18785 23418
rect 18837 23366 18849 23418
rect 18901 23366 18913 23418
rect 18965 23366 25740 23418
rect 25792 23366 25804 23418
rect 25856 23366 25868 23418
rect 25920 23366 25932 23418
rect 25984 23366 25996 23418
rect 26048 23366 29440 23418
rect 1104 23344 29440 23366
rect 9122 23304 9128 23316
rect 9048 23276 9128 23304
rect 6546 23128 6552 23180
rect 6604 23168 6610 23180
rect 9048 23177 9076 23276
rect 9122 23264 9128 23276
rect 9180 23304 9186 23316
rect 11422 23304 11428 23316
rect 9180 23276 11428 23304
rect 9180 23264 9186 23276
rect 11422 23264 11428 23276
rect 11480 23264 11486 23316
rect 14550 23264 14556 23316
rect 14608 23304 14614 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14608 23276 14657 23304
rect 14608 23264 14614 23276
rect 14645 23273 14657 23276
rect 14691 23273 14703 23307
rect 14645 23267 14703 23273
rect 15010 23264 15016 23316
rect 15068 23264 15074 23316
rect 15102 23264 15108 23316
rect 15160 23304 15166 23316
rect 15378 23304 15384 23316
rect 15160 23276 15384 23304
rect 15160 23264 15166 23276
rect 15378 23264 15384 23276
rect 15436 23304 15442 23316
rect 17402 23304 17408 23316
rect 15436 23276 17408 23304
rect 15436 23264 15442 23276
rect 17402 23264 17408 23276
rect 17460 23264 17466 23316
rect 25222 23264 25228 23316
rect 25280 23264 25286 23316
rect 10594 23196 10600 23248
rect 10652 23196 10658 23248
rect 10778 23196 10784 23248
rect 10836 23196 10842 23248
rect 15120 23236 15148 23264
rect 10888 23208 15148 23236
rect 6733 23171 6791 23177
rect 6733 23168 6745 23171
rect 6604 23140 6745 23168
rect 6604 23128 6610 23140
rect 6733 23137 6745 23140
rect 6779 23137 6791 23171
rect 6733 23131 6791 23137
rect 9033 23171 9091 23177
rect 9033 23137 9045 23171
rect 9079 23137 9091 23171
rect 9033 23131 9091 23137
rect 4525 23103 4583 23109
rect 4525 23069 4537 23103
rect 4571 23100 4583 23103
rect 6178 23100 6184 23112
rect 4571 23072 6184 23100
rect 4571 23069 4583 23072
rect 4525 23063 4583 23069
rect 6178 23060 6184 23072
rect 6236 23060 6242 23112
rect 10612 23100 10640 23196
rect 10442 23072 10640 23100
rect 10888 23044 10916 23208
rect 15194 23196 15200 23248
rect 15252 23196 15258 23248
rect 15562 23196 15568 23248
rect 15620 23196 15626 23248
rect 15838 23196 15844 23248
rect 15896 23236 15902 23248
rect 17589 23239 17647 23245
rect 17589 23236 17601 23239
rect 15896 23208 17601 23236
rect 15896 23196 15902 23208
rect 17589 23205 17601 23208
rect 17635 23236 17647 23239
rect 18138 23236 18144 23248
rect 17635 23208 18144 23236
rect 17635 23205 17647 23208
rect 17589 23199 17647 23205
rect 18138 23196 18144 23208
rect 18196 23196 18202 23248
rect 11422 23128 11428 23180
rect 11480 23168 11486 23180
rect 11609 23171 11667 23177
rect 11609 23168 11621 23171
rect 11480 23140 11621 23168
rect 11480 23128 11486 23140
rect 11609 23137 11621 23140
rect 11655 23137 11667 23171
rect 11609 23131 11667 23137
rect 14550 23128 14556 23180
rect 14608 23168 14614 23180
rect 14829 23171 14887 23177
rect 14829 23168 14841 23171
rect 14608 23140 14841 23168
rect 14608 23128 14614 23140
rect 14829 23137 14841 23140
rect 14875 23168 14887 23171
rect 14875 23140 15884 23168
rect 14875 23137 14887 23140
rect 14829 23131 14887 23137
rect 14093 23103 14151 23109
rect 14093 23069 14105 23103
rect 14139 23100 14151 23103
rect 14274 23100 14280 23112
rect 14139 23072 14280 23100
rect 14139 23069 14151 23072
rect 14093 23063 14151 23069
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 14458 23060 14464 23112
rect 14516 23060 14522 23112
rect 14737 23103 14795 23109
rect 14737 23069 14749 23103
rect 14783 23100 14795 23103
rect 14918 23100 14924 23112
rect 14783 23072 14924 23100
rect 14783 23069 14795 23072
rect 14737 23063 14795 23069
rect 14918 23060 14924 23072
rect 14976 23060 14982 23112
rect 15013 23103 15071 23109
rect 15013 23069 15025 23103
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 5997 23035 6055 23041
rect 5997 23001 6009 23035
rect 6043 23001 6055 23035
rect 5997 22995 6055 23001
rect 5074 22924 5080 22976
rect 5132 22924 5138 22976
rect 5902 22924 5908 22976
rect 5960 22964 5966 22976
rect 6012 22964 6040 22995
rect 9306 22992 9312 23044
rect 9364 22992 9370 23044
rect 10870 23032 10876 23044
rect 10612 23004 10876 23032
rect 10612 22964 10640 23004
rect 10870 22992 10876 23004
rect 10928 22992 10934 23044
rect 14369 23035 14427 23041
rect 14369 23032 14381 23035
rect 13740 23004 14381 23032
rect 13740 22976 13768 23004
rect 14369 23001 14381 23004
rect 14415 23001 14427 23035
rect 14476 23032 14504 23060
rect 15028 23032 15056 23063
rect 15286 23060 15292 23112
rect 15344 23060 15350 23112
rect 15856 23109 15884 23140
rect 16022 23128 16028 23180
rect 16080 23168 16086 23180
rect 20993 23171 21051 23177
rect 16080 23140 18368 23168
rect 16080 23128 16086 23140
rect 15749 23103 15807 23109
rect 15563 23081 15621 23087
rect 15563 23047 15575 23081
rect 15609 23047 15621 23081
rect 15749 23069 15761 23103
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 15841 23103 15899 23109
rect 15841 23069 15853 23103
rect 15887 23069 15899 23103
rect 15841 23063 15899 23069
rect 15563 23044 15621 23047
rect 15194 23032 15200 23044
rect 14476 23004 15200 23032
rect 14369 22995 14427 23001
rect 15194 22992 15200 23004
rect 15252 23032 15258 23044
rect 15473 23035 15531 23041
rect 15473 23032 15485 23035
rect 15252 23004 15485 23032
rect 15252 22992 15258 23004
rect 15473 23001 15485 23004
rect 15519 23001 15531 23035
rect 15473 22995 15531 23001
rect 15562 22992 15568 23044
rect 15620 22992 15626 23044
rect 15764 23032 15792 23063
rect 16114 23060 16120 23112
rect 16172 23060 16178 23112
rect 17604 23109 17632 23140
rect 18340 23112 18368 23140
rect 20993 23137 21005 23171
rect 21039 23168 21051 23171
rect 21634 23168 21640 23180
rect 21039 23140 21640 23168
rect 21039 23137 21051 23140
rect 20993 23131 21051 23137
rect 21634 23128 21640 23140
rect 21692 23128 21698 23180
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 17773 23103 17831 23109
rect 17773 23069 17785 23103
rect 17819 23069 17831 23103
rect 17773 23063 17831 23069
rect 16132 23032 16160 23060
rect 15764 23004 16160 23032
rect 5960 22936 10640 22964
rect 5960 22924 5966 22936
rect 13722 22924 13728 22976
rect 13780 22924 13786 22976
rect 14277 22967 14335 22973
rect 14277 22933 14289 22967
rect 14323 22964 14335 22967
rect 14642 22964 14648 22976
rect 14323 22936 14648 22964
rect 14323 22933 14335 22936
rect 14277 22927 14335 22933
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 15010 22924 15016 22976
rect 15068 22964 15074 22976
rect 15764 22964 15792 23004
rect 17310 22992 17316 23044
rect 17368 23032 17374 23044
rect 17788 23032 17816 23063
rect 18322 23060 18328 23112
rect 18380 23060 18386 23112
rect 20714 23060 20720 23112
rect 20772 23060 20778 23112
rect 20806 23060 20812 23112
rect 20864 23060 20870 23112
rect 21082 23060 21088 23112
rect 21140 23060 21146 23112
rect 23750 23060 23756 23112
rect 23808 23100 23814 23112
rect 24486 23100 24492 23112
rect 23808 23072 24492 23100
rect 23808 23060 23814 23072
rect 24486 23060 24492 23072
rect 24544 23060 24550 23112
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23100 24639 23103
rect 24670 23100 24676 23112
rect 24627 23072 24676 23100
rect 24627 23069 24639 23072
rect 24581 23063 24639 23069
rect 17368 23004 17816 23032
rect 17368 22992 17374 23004
rect 21174 22992 21180 23044
rect 21232 22992 21238 23044
rect 22554 22992 22560 23044
rect 22612 23032 22618 23044
rect 24596 23032 24624 23063
rect 24670 23060 24676 23072
rect 24728 23060 24734 23112
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23100 24823 23103
rect 24857 23103 24915 23109
rect 24857 23100 24869 23103
rect 24811 23072 24869 23100
rect 24811 23069 24823 23072
rect 24765 23063 24823 23069
rect 24857 23069 24869 23072
rect 24903 23100 24915 23103
rect 24903 23072 25544 23100
rect 24903 23069 24915 23072
rect 24857 23063 24915 23069
rect 25516 23044 25544 23072
rect 22612 23004 24624 23032
rect 25041 23035 25099 23041
rect 22612 22992 22618 23004
rect 25041 23001 25053 23035
rect 25087 23001 25099 23035
rect 25041 22995 25099 23001
rect 15068 22936 15792 22964
rect 15068 22924 15074 22936
rect 17218 22924 17224 22976
rect 17276 22964 17282 22976
rect 17586 22964 17592 22976
rect 17276 22936 17592 22964
rect 17276 22924 17282 22936
rect 17586 22924 17592 22936
rect 17644 22964 17650 22976
rect 18046 22964 18052 22976
rect 17644 22936 18052 22964
rect 17644 22924 17650 22936
rect 18046 22924 18052 22936
rect 18104 22924 18110 22976
rect 20990 22924 20996 22976
rect 21048 22924 21054 22976
rect 23842 22924 23848 22976
rect 23900 22964 23906 22976
rect 24394 22964 24400 22976
rect 23900 22936 24400 22964
rect 23900 22924 23906 22936
rect 24394 22924 24400 22936
rect 24452 22924 24458 22976
rect 24762 22924 24768 22976
rect 24820 22964 24826 22976
rect 25056 22964 25084 22995
rect 25498 22992 25504 23044
rect 25556 22992 25562 23044
rect 25406 22964 25412 22976
rect 24820 22936 25412 22964
rect 24820 22924 24826 22936
rect 25406 22924 25412 22936
rect 25464 22924 25470 22976
rect 1104 22874 29440 22896
rect 1104 22822 5151 22874
rect 5203 22822 5215 22874
rect 5267 22822 5279 22874
rect 5331 22822 5343 22874
rect 5395 22822 5407 22874
rect 5459 22822 12234 22874
rect 12286 22822 12298 22874
rect 12350 22822 12362 22874
rect 12414 22822 12426 22874
rect 12478 22822 12490 22874
rect 12542 22822 19317 22874
rect 19369 22822 19381 22874
rect 19433 22822 19445 22874
rect 19497 22822 19509 22874
rect 19561 22822 19573 22874
rect 19625 22822 26400 22874
rect 26452 22822 26464 22874
rect 26516 22822 26528 22874
rect 26580 22822 26592 22874
rect 26644 22822 26656 22874
rect 26708 22822 29440 22874
rect 1104 22800 29440 22822
rect 9217 22763 9275 22769
rect 9217 22729 9229 22763
rect 9263 22760 9275 22763
rect 9306 22760 9312 22772
rect 9263 22732 9312 22760
rect 9263 22729 9275 22732
rect 9217 22723 9275 22729
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 9548 22732 12480 22760
rect 9548 22720 9554 22732
rect 5261 22695 5319 22701
rect 5261 22661 5273 22695
rect 5307 22692 5319 22695
rect 5902 22692 5908 22704
rect 5307 22664 5908 22692
rect 5307 22661 5319 22664
rect 5261 22655 5319 22661
rect 5902 22652 5908 22664
rect 5960 22652 5966 22704
rect 8205 22695 8263 22701
rect 8205 22692 8217 22695
rect 6748 22664 8217 22692
rect 6748 22633 6776 22664
rect 8205 22661 8217 22664
rect 8251 22661 8263 22695
rect 8205 22655 8263 22661
rect 8941 22695 8999 22701
rect 8941 22661 8953 22695
rect 8987 22692 8999 22695
rect 9674 22692 9680 22704
rect 8987 22664 9680 22692
rect 8987 22661 8999 22664
rect 8941 22655 8999 22661
rect 9674 22652 9680 22664
rect 9732 22652 9738 22704
rect 10962 22692 10968 22704
rect 10810 22664 10968 22692
rect 10962 22652 10968 22664
rect 11020 22652 11026 22704
rect 12452 22701 12480 22732
rect 12802 22720 12808 22772
rect 12860 22720 12866 22772
rect 15838 22760 15844 22772
rect 15120 22732 15844 22760
rect 12437 22695 12495 22701
rect 12437 22661 12449 22695
rect 12483 22661 12495 22695
rect 12437 22655 12495 22661
rect 12529 22695 12587 22701
rect 12529 22661 12541 22695
rect 12575 22692 12587 22695
rect 12575 22664 13216 22692
rect 12575 22661 12587 22664
rect 12529 22655 12587 22661
rect 6733 22627 6791 22633
rect 6733 22593 6745 22627
rect 6779 22593 6791 22627
rect 6733 22587 6791 22593
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 7009 22627 7067 22633
rect 7009 22593 7021 22627
rect 7055 22593 7067 22627
rect 7009 22587 7067 22593
rect 4525 22559 4583 22565
rect 4525 22525 4537 22559
rect 4571 22556 4583 22559
rect 5718 22556 5724 22568
rect 4571 22528 5724 22556
rect 4571 22525 4583 22528
rect 4525 22519 4583 22525
rect 5718 22516 5724 22528
rect 5776 22516 5782 22568
rect 5994 22516 6000 22568
rect 6052 22516 6058 22568
rect 6932 22488 6960 22587
rect 7024 22556 7052 22587
rect 7098 22584 7104 22636
rect 7156 22584 7162 22636
rect 8110 22624 8116 22636
rect 7208 22596 8116 22624
rect 7208 22556 7236 22596
rect 8110 22584 8116 22596
rect 8168 22584 8174 22636
rect 8662 22584 8668 22636
rect 8720 22584 8726 22636
rect 8846 22584 8852 22636
rect 8904 22584 8910 22636
rect 9033 22627 9091 22633
rect 9033 22593 9045 22627
rect 9079 22593 9091 22627
rect 9033 22587 9091 22593
rect 7024 22528 7236 22556
rect 7650 22516 7656 22568
rect 7708 22516 7714 22568
rect 9048 22556 9076 22587
rect 9122 22584 9128 22636
rect 9180 22624 9186 22636
rect 9309 22627 9367 22633
rect 9309 22624 9321 22627
rect 9180 22596 9321 22624
rect 9180 22584 9186 22596
rect 9309 22593 9321 22596
rect 9355 22593 9367 22627
rect 11330 22624 11336 22636
rect 9309 22587 9367 22593
rect 10796 22596 11336 22624
rect 10796 22568 10824 22596
rect 11330 22584 11336 22596
rect 11388 22584 11394 22636
rect 12158 22584 12164 22636
rect 12216 22624 12222 22636
rect 12253 22627 12311 22633
rect 12253 22624 12265 22627
rect 12216 22596 12265 22624
rect 12216 22584 12222 22596
rect 12253 22593 12265 22596
rect 12299 22593 12311 22627
rect 12253 22587 12311 22593
rect 8588 22528 9076 22556
rect 9585 22559 9643 22565
rect 8588 22500 8616 22528
rect 9585 22525 9597 22559
rect 9631 22556 9643 22559
rect 10134 22556 10140 22568
rect 9631 22528 10140 22556
rect 9631 22525 9643 22528
rect 9585 22519 9643 22525
rect 10134 22516 10140 22528
rect 10192 22516 10198 22568
rect 10778 22516 10784 22568
rect 10836 22516 10842 22568
rect 11057 22559 11115 22565
rect 11057 22525 11069 22559
rect 11103 22556 11115 22559
rect 11422 22556 11428 22568
rect 11103 22528 11428 22556
rect 11103 22525 11115 22528
rect 11057 22519 11115 22525
rect 11422 22516 11428 22528
rect 11480 22556 11486 22568
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 11480 22528 11529 22556
rect 11480 22516 11486 22528
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 11517 22519 11575 22525
rect 6932 22460 7420 22488
rect 7392 22432 7420 22460
rect 8570 22448 8576 22500
rect 8628 22448 8634 22500
rect 11238 22448 11244 22500
rect 11296 22488 11302 22500
rect 12544 22488 12572 22655
rect 13188 22636 13216 22664
rect 12618 22584 12624 22636
rect 12676 22584 12682 22636
rect 13170 22584 13176 22636
rect 13228 22584 13234 22636
rect 14274 22584 14280 22636
rect 14332 22584 14338 22636
rect 15013 22627 15071 22633
rect 15013 22593 15025 22627
rect 15059 22624 15071 22627
rect 15120 22624 15148 22732
rect 15838 22720 15844 22732
rect 15896 22720 15902 22772
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 20901 22763 20959 22769
rect 20901 22760 20913 22763
rect 20772 22732 20913 22760
rect 20772 22720 20778 22732
rect 20901 22729 20913 22732
rect 20947 22729 20959 22763
rect 20901 22723 20959 22729
rect 15378 22652 15384 22704
rect 15436 22692 15442 22704
rect 15930 22692 15936 22704
rect 15436 22664 15936 22692
rect 15436 22652 15442 22664
rect 15930 22652 15936 22664
rect 15988 22652 15994 22704
rect 15059 22596 15148 22624
rect 15289 22627 15347 22633
rect 15059 22593 15071 22596
rect 15013 22587 15071 22593
rect 15289 22593 15301 22627
rect 15335 22624 15347 22627
rect 17313 22627 17371 22633
rect 17313 22624 17325 22627
rect 15335 22596 17325 22624
rect 15335 22593 15347 22596
rect 15289 22587 15347 22593
rect 17313 22593 17325 22596
rect 17359 22593 17371 22627
rect 17313 22587 17371 22593
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22593 20775 22627
rect 20717 22587 20775 22593
rect 14292 22556 14320 22584
rect 15197 22559 15255 22565
rect 14292 22528 15148 22556
rect 11296 22460 12572 22488
rect 11296 22448 11302 22460
rect 13722 22448 13728 22500
rect 13780 22488 13786 22500
rect 15120 22488 15148 22528
rect 15197 22525 15209 22559
rect 15243 22556 15255 22559
rect 15470 22556 15476 22568
rect 15243 22528 15476 22556
rect 15243 22525 15255 22528
rect 15197 22519 15255 22525
rect 15470 22516 15476 22528
rect 15528 22516 15534 22568
rect 16209 22559 16267 22565
rect 16209 22525 16221 22559
rect 16255 22556 16267 22559
rect 16482 22556 16488 22568
rect 16255 22528 16488 22556
rect 16255 22525 16267 22528
rect 16209 22519 16267 22525
rect 16482 22516 16488 22528
rect 16540 22516 16546 22568
rect 16666 22516 16672 22568
rect 16724 22516 16730 22568
rect 20530 22516 20536 22568
rect 20588 22516 20594 22568
rect 15562 22488 15568 22500
rect 13780 22460 14964 22488
rect 15120 22460 15568 22488
rect 13780 22448 13786 22460
rect 4154 22380 4160 22432
rect 4212 22420 4218 22432
rect 5077 22423 5135 22429
rect 5077 22420 5089 22423
rect 4212 22392 5089 22420
rect 4212 22380 4218 22392
rect 5077 22389 5089 22392
rect 5123 22389 5135 22423
rect 5077 22383 5135 22389
rect 7282 22380 7288 22432
rect 7340 22380 7346 22432
rect 7374 22380 7380 22432
rect 7432 22420 7438 22432
rect 9398 22420 9404 22432
rect 7432 22392 9404 22420
rect 7432 22380 7438 22392
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 10226 22380 10232 22432
rect 10284 22420 10290 22432
rect 12161 22423 12219 22429
rect 12161 22420 12173 22423
rect 10284 22392 12173 22420
rect 10284 22380 10290 22392
rect 12161 22389 12173 22392
rect 12207 22389 12219 22423
rect 12161 22383 12219 22389
rect 14826 22380 14832 22432
rect 14884 22380 14890 22432
rect 14936 22420 14964 22460
rect 15562 22448 15568 22460
rect 15620 22448 15626 22500
rect 16390 22448 16396 22500
rect 16448 22448 16454 22500
rect 20732 22488 20760 22587
rect 20806 22584 20812 22636
rect 20864 22584 20870 22636
rect 20916 22624 20944 22723
rect 22830 22720 22836 22772
rect 22888 22760 22894 22772
rect 24397 22763 24455 22769
rect 22888 22732 24348 22760
rect 22888 22720 22894 22732
rect 21082 22652 21088 22704
rect 21140 22692 21146 22704
rect 21726 22692 21732 22704
rect 21140 22664 21732 22692
rect 21140 22652 21146 22664
rect 21560 22633 21588 22664
rect 21726 22652 21732 22664
rect 21784 22652 21790 22704
rect 22020 22664 22968 22692
rect 21269 22627 21327 22633
rect 21269 22624 21281 22627
rect 20916 22596 21281 22624
rect 21269 22593 21281 22596
rect 21315 22593 21327 22627
rect 21269 22587 21327 22593
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 21545 22627 21603 22633
rect 21545 22593 21557 22627
rect 21591 22593 21603 22627
rect 21545 22587 21603 22593
rect 20824 22556 20852 22584
rect 21174 22556 21180 22568
rect 20824 22528 21180 22556
rect 21174 22516 21180 22528
rect 21232 22556 21238 22568
rect 21361 22559 21419 22565
rect 21361 22556 21373 22559
rect 21232 22528 21373 22556
rect 21232 22516 21238 22528
rect 21361 22525 21373 22528
rect 21407 22525 21419 22559
rect 21468 22556 21496 22587
rect 21634 22584 21640 22636
rect 21692 22624 21698 22636
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21692 22596 21833 22624
rect 21692 22584 21698 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 22020 22633 22048 22664
rect 22940 22633 22968 22664
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21968 22596 22017 22624
rect 21968 22584 21974 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22741 22627 22799 22633
rect 22741 22593 22753 22627
rect 22787 22593 22799 22627
rect 22741 22587 22799 22593
rect 22925 22627 22983 22633
rect 22925 22593 22937 22627
rect 22971 22624 22983 22627
rect 23014 22624 23020 22636
rect 22971 22596 23020 22624
rect 22971 22593 22983 22596
rect 22925 22587 22983 22593
rect 22646 22556 22652 22568
rect 21468 22528 22652 22556
rect 21361 22519 21419 22525
rect 22646 22516 22652 22528
rect 22704 22516 22710 22568
rect 22756 22556 22784 22587
rect 23014 22584 23020 22596
rect 23072 22584 23078 22636
rect 23106 22584 23112 22636
rect 23164 22584 23170 22636
rect 23198 22584 23204 22636
rect 23256 22584 23262 22636
rect 23290 22584 23296 22636
rect 23348 22584 23354 22636
rect 23768 22633 23796 22732
rect 24320 22692 24348 22732
rect 24397 22729 24409 22763
rect 24443 22760 24455 22763
rect 25314 22760 25320 22772
rect 24443 22732 25320 22760
rect 24443 22729 24455 22732
rect 24397 22723 24455 22729
rect 25314 22720 25320 22732
rect 25372 22720 25378 22772
rect 25406 22720 25412 22772
rect 25464 22720 25470 22772
rect 24320 22664 25084 22692
rect 23661 22627 23719 22633
rect 23661 22624 23673 22627
rect 23400 22596 23673 22624
rect 23216 22556 23244 22584
rect 22756 22528 23244 22556
rect 20732 22460 20852 22488
rect 16408 22420 16436 22448
rect 20824 22432 20852 22460
rect 21634 22448 21640 22500
rect 21692 22488 21698 22500
rect 23400 22488 23428 22596
rect 23661 22593 23673 22596
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 23753 22627 23811 22633
rect 23753 22593 23765 22627
rect 23799 22593 23811 22627
rect 23753 22587 23811 22593
rect 23842 22584 23848 22636
rect 23900 22633 23906 22636
rect 23900 22627 23954 22633
rect 23900 22593 23908 22627
rect 23942 22593 23954 22627
rect 23900 22587 23954 22593
rect 23900 22584 23906 22587
rect 24026 22584 24032 22636
rect 24084 22584 24090 22636
rect 24320 22633 24348 22664
rect 25056 22636 25084 22664
rect 24121 22627 24179 22633
rect 24121 22593 24133 22627
rect 24167 22593 24179 22627
rect 24121 22587 24179 22593
rect 24305 22627 24363 22633
rect 24305 22593 24317 22627
rect 24351 22593 24363 22627
rect 24305 22587 24363 22593
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 24136 22556 24164 22587
rect 24394 22584 24400 22636
rect 24452 22584 24458 22636
rect 24568 22627 24626 22633
rect 24568 22624 24580 22627
rect 24504 22596 24580 22624
rect 23532 22528 24164 22556
rect 24213 22559 24271 22565
rect 23532 22516 23538 22528
rect 24213 22525 24225 22559
rect 24259 22556 24271 22559
rect 24412 22556 24440 22584
rect 24259 22528 24440 22556
rect 24259 22525 24271 22528
rect 24213 22519 24271 22525
rect 21692 22460 23428 22488
rect 21692 22448 21698 22460
rect 24026 22448 24032 22500
rect 24084 22448 24090 22500
rect 24394 22448 24400 22500
rect 24452 22488 24458 22500
rect 24504 22488 24532 22596
rect 24568 22593 24580 22596
rect 24614 22593 24626 22627
rect 24568 22587 24626 22593
rect 24673 22627 24731 22633
rect 24673 22593 24685 22627
rect 24719 22593 24731 22627
rect 24673 22587 24731 22593
rect 24688 22556 24716 22587
rect 24762 22584 24768 22636
rect 24820 22584 24826 22636
rect 24857 22630 24915 22633
rect 24857 22627 24992 22630
rect 24857 22593 24869 22627
rect 24903 22602 24992 22627
rect 24903 22593 24915 22602
rect 24857 22587 24915 22593
rect 24964 22568 24992 22602
rect 25038 22584 25044 22636
rect 25096 22584 25102 22636
rect 25222 22584 25228 22636
rect 25280 22584 25286 22636
rect 28810 22584 28816 22636
rect 28868 22584 28874 22636
rect 24596 22528 24716 22556
rect 24596 22500 24624 22528
rect 24946 22516 24952 22568
rect 25004 22516 25010 22568
rect 24452 22460 24532 22488
rect 24452 22448 24458 22460
rect 24578 22448 24584 22500
rect 24636 22448 24642 22500
rect 28994 22448 29000 22500
rect 29052 22448 29058 22500
rect 14936 22392 16436 22420
rect 20806 22380 20812 22432
rect 20864 22380 20870 22432
rect 21082 22380 21088 22432
rect 21140 22380 21146 22432
rect 21821 22423 21879 22429
rect 21821 22389 21833 22423
rect 21867 22420 21879 22423
rect 22094 22420 22100 22432
rect 21867 22392 22100 22420
rect 21867 22389 21879 22392
rect 21821 22383 21879 22389
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 22738 22380 22744 22432
rect 22796 22380 22802 22432
rect 23198 22380 23204 22432
rect 23256 22380 23262 22432
rect 23382 22380 23388 22432
rect 23440 22420 23446 22432
rect 23477 22423 23535 22429
rect 23477 22420 23489 22423
rect 23440 22392 23489 22420
rect 23440 22380 23446 22392
rect 23477 22389 23489 22392
rect 23523 22389 23535 22423
rect 24044 22420 24072 22448
rect 24946 22420 24952 22432
rect 24044 22392 24952 22420
rect 23477 22383 23535 22389
rect 24946 22380 24952 22392
rect 25004 22380 25010 22432
rect 1104 22330 29440 22352
rect 1104 22278 4491 22330
rect 4543 22278 4555 22330
rect 4607 22278 4619 22330
rect 4671 22278 4683 22330
rect 4735 22278 4747 22330
rect 4799 22278 11574 22330
rect 11626 22278 11638 22330
rect 11690 22278 11702 22330
rect 11754 22278 11766 22330
rect 11818 22278 11830 22330
rect 11882 22278 18657 22330
rect 18709 22278 18721 22330
rect 18773 22278 18785 22330
rect 18837 22278 18849 22330
rect 18901 22278 18913 22330
rect 18965 22278 25740 22330
rect 25792 22278 25804 22330
rect 25856 22278 25868 22330
rect 25920 22278 25932 22330
rect 25984 22278 25996 22330
rect 26048 22278 29440 22330
rect 1104 22256 29440 22278
rect 6260 22219 6318 22225
rect 6260 22185 6272 22219
rect 6306 22216 6318 22219
rect 7282 22216 7288 22228
rect 6306 22188 7288 22216
rect 6306 22185 6318 22188
rect 6260 22179 6318 22185
rect 7282 22176 7288 22188
rect 7340 22176 7346 22228
rect 7650 22176 7656 22228
rect 7708 22216 7714 22228
rect 7745 22219 7803 22225
rect 7745 22216 7757 22219
rect 7708 22188 7757 22216
rect 7708 22176 7714 22188
rect 7745 22185 7757 22188
rect 7791 22185 7803 22219
rect 7745 22179 7803 22185
rect 8662 22176 8668 22228
rect 8720 22216 8726 22228
rect 11238 22216 11244 22228
rect 8720 22188 11244 22216
rect 8720 22176 8726 22188
rect 11238 22176 11244 22188
rect 11296 22176 11302 22228
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 12618 22216 12624 22228
rect 11388 22188 12624 22216
rect 11388 22176 11394 22188
rect 12618 22176 12624 22188
rect 12676 22176 12682 22228
rect 13722 22176 13728 22228
rect 13780 22176 13786 22228
rect 14724 22219 14782 22225
rect 14724 22185 14736 22219
rect 14770 22216 14782 22219
rect 14826 22216 14832 22228
rect 14770 22188 14832 22216
rect 14770 22185 14782 22188
rect 14724 22179 14782 22185
rect 14826 22176 14832 22188
rect 14884 22176 14890 22228
rect 21634 22176 21640 22228
rect 21692 22176 21698 22228
rect 21726 22176 21732 22228
rect 21784 22216 21790 22228
rect 22097 22219 22155 22225
rect 21784 22188 22064 22216
rect 21784 22176 21790 22188
rect 8110 22108 8116 22160
rect 8168 22148 8174 22160
rect 9950 22148 9956 22160
rect 8168 22120 9956 22148
rect 8168 22108 8174 22120
rect 9950 22108 9956 22120
rect 10008 22148 10014 22160
rect 13740 22148 13768 22176
rect 10008 22120 13768 22148
rect 10008 22108 10014 22120
rect 21266 22108 21272 22160
rect 21324 22148 21330 22160
rect 21542 22148 21548 22160
rect 21324 22120 21548 22148
rect 21324 22108 21330 22120
rect 3694 22040 3700 22092
rect 3752 22080 3758 22092
rect 5442 22080 5448 22092
rect 3752 22052 5448 22080
rect 3752 22040 3758 22052
rect 4264 22024 4292 22052
rect 5442 22040 5448 22052
rect 5500 22040 5506 22092
rect 5994 22040 6000 22092
rect 6052 22080 6058 22092
rect 6362 22080 6368 22092
rect 6052 22052 6368 22080
rect 6052 22040 6058 22052
rect 6362 22040 6368 22052
rect 6420 22040 6426 22092
rect 10042 22080 10048 22092
rect 8588 22052 9168 22080
rect 8588 22024 8616 22052
rect 4157 22015 4215 22021
rect 4157 21981 4169 22015
rect 4203 21981 4215 22015
rect 4157 21975 4215 21981
rect 4172 21944 4200 21975
rect 4246 21972 4252 22024
rect 4304 22012 4310 22024
rect 4433 22015 4491 22021
rect 4433 22012 4445 22015
rect 4304 21984 4445 22012
rect 4304 21972 4310 21984
rect 4433 21981 4445 21984
rect 4479 21981 4491 22015
rect 4982 22012 4988 22024
rect 4433 21975 4491 21981
rect 4540 21984 4988 22012
rect 4540 21944 4568 21984
rect 4982 21972 4988 21984
rect 5040 21972 5046 22024
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 22012 5411 22015
rect 5534 22012 5540 22024
rect 5399 21984 5540 22012
rect 5399 21981 5411 21984
rect 5353 21975 5411 21981
rect 5534 21972 5540 21984
rect 5592 21972 5598 22024
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 4172 21916 4568 21944
rect 4890 21904 4896 21956
rect 4948 21944 4954 21956
rect 4948 21916 6762 21944
rect 4948 21904 4954 21916
rect 3234 21836 3240 21888
rect 3292 21876 3298 21888
rect 4065 21879 4123 21885
rect 4065 21876 4077 21879
rect 3292 21848 4077 21876
rect 3292 21836 3298 21848
rect 4065 21845 4077 21848
rect 4111 21876 4123 21879
rect 4706 21876 4712 21888
rect 4111 21848 4712 21876
rect 4111 21845 4123 21848
rect 4065 21839 4123 21845
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 5902 21836 5908 21888
rect 5960 21836 5966 21888
rect 6656 21876 6684 21916
rect 7852 21888 7880 21975
rect 8570 21972 8576 22024
rect 8628 21972 8634 22024
rect 9033 22015 9091 22021
rect 9033 21981 9045 22015
rect 9079 21981 9091 22015
rect 9140 22012 9168 22052
rect 9508 22052 10048 22080
rect 9401 22015 9459 22021
rect 9401 22012 9413 22015
rect 9140 21984 9413 22012
rect 9033 21975 9091 21981
rect 9401 21981 9413 21984
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 7098 21876 7104 21888
rect 6656 21848 7104 21876
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 7834 21836 7840 21888
rect 7892 21836 7898 21888
rect 8478 21836 8484 21888
rect 8536 21836 8542 21888
rect 9048 21876 9076 21975
rect 9122 21904 9128 21956
rect 9180 21944 9186 21956
rect 9217 21947 9275 21953
rect 9217 21944 9229 21947
rect 9180 21916 9229 21944
rect 9180 21904 9186 21916
rect 9217 21913 9229 21916
rect 9263 21913 9275 21947
rect 9217 21907 9275 21913
rect 9309 21947 9367 21953
rect 9309 21913 9321 21947
rect 9355 21944 9367 21947
rect 9508 21944 9536 22052
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 10134 22040 10140 22092
rect 10192 22080 10198 22092
rect 10321 22083 10379 22089
rect 10321 22080 10333 22083
rect 10192 22052 10333 22080
rect 10192 22040 10198 22052
rect 10321 22049 10333 22052
rect 10367 22049 10379 22083
rect 10321 22043 10379 22049
rect 10594 22040 10600 22092
rect 10652 22080 10658 22092
rect 12894 22080 12900 22092
rect 10652 22052 12900 22080
rect 10652 22040 10658 22052
rect 12894 22040 12900 22052
rect 12952 22040 12958 22092
rect 14458 22040 14464 22092
rect 14516 22080 14522 22092
rect 16482 22080 16488 22092
rect 14516 22052 16488 22080
rect 14516 22040 14522 22052
rect 16482 22040 16488 22052
rect 16540 22040 16546 22092
rect 20088 22052 20849 22080
rect 9677 22015 9735 22021
rect 9677 22012 9689 22015
rect 9355 21916 9536 21944
rect 9600 21984 9689 22012
rect 9355 21913 9367 21916
rect 9309 21907 9367 21913
rect 9490 21876 9496 21888
rect 9048 21848 9496 21876
rect 9490 21836 9496 21848
rect 9548 21836 9554 21888
rect 9600 21885 9628 21984
rect 9677 21981 9689 21984
rect 9723 21981 9735 22015
rect 9677 21975 9735 21981
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 9585 21879 9643 21885
rect 9585 21845 9597 21879
rect 9631 21845 9643 21879
rect 9585 21839 9643 21845
rect 10226 21836 10232 21888
rect 10284 21876 10290 21888
rect 10428 21876 10456 21975
rect 10502 21972 10508 22024
rect 10560 21972 10566 22024
rect 10778 21972 10784 22024
rect 10836 21972 10842 22024
rect 10919 22015 10977 22021
rect 10919 21981 10931 22015
rect 10965 22012 10977 22015
rect 17313 22015 17371 22021
rect 10965 21984 12020 22012
rect 10965 21981 10977 21984
rect 10919 21975 10977 21981
rect 11992 21956 12020 21984
rect 17313 21981 17325 22015
rect 17359 22012 17371 22015
rect 18414 22012 18420 22024
rect 17359 21984 18420 22012
rect 17359 21981 17371 21984
rect 17313 21975 17371 21981
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 20088 22021 20116 22052
rect 20821 22024 20849 22052
rect 21008 22052 21312 22080
rect 21008 22024 21036 22052
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 21981 20131 22015
rect 20073 21975 20131 21981
rect 20165 22015 20223 22021
rect 20165 21981 20177 22015
rect 20211 21981 20223 22015
rect 20165 21975 20223 21981
rect 20257 22015 20315 22021
rect 20257 21981 20269 22015
rect 20303 22012 20315 22015
rect 20438 22012 20444 22024
rect 20303 21984 20444 22012
rect 20303 21981 20315 21984
rect 20257 21975 20315 21981
rect 10689 21947 10747 21953
rect 10689 21944 10701 21947
rect 10520 21916 10701 21944
rect 10520 21888 10548 21916
rect 10689 21913 10701 21916
rect 10735 21913 10747 21947
rect 10689 21907 10747 21913
rect 11974 21904 11980 21956
rect 12032 21904 12038 21956
rect 12618 21904 12624 21956
rect 12676 21944 12682 21956
rect 13446 21944 13452 21956
rect 12676 21916 13452 21944
rect 12676 21904 12682 21916
rect 13446 21904 13452 21916
rect 13504 21904 13510 21956
rect 17770 21944 17776 21956
rect 15962 21916 17776 21944
rect 17770 21904 17776 21916
rect 17828 21944 17834 21956
rect 19794 21944 19800 21956
rect 17828 21916 19800 21944
rect 17828 21904 17834 21916
rect 19794 21904 19800 21916
rect 19852 21904 19858 21956
rect 20180 21944 20208 21975
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 22012 20591 22015
rect 20714 22012 20720 22024
rect 20579 21984 20720 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 20806 21972 20812 22024
rect 20864 21972 20870 22024
rect 20990 21972 20996 22024
rect 21048 21972 21054 22024
rect 21082 21972 21088 22024
rect 21140 21972 21146 22024
rect 21284 22021 21312 22052
rect 21376 22021 21404 22120
rect 21542 22108 21548 22120
rect 21600 22148 21606 22160
rect 22036 22148 22064 22188
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22554 22216 22560 22228
rect 22143 22188 22560 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22554 22176 22560 22188
rect 22612 22176 22618 22228
rect 23753 22219 23811 22225
rect 23753 22185 23765 22219
rect 23799 22216 23811 22219
rect 24578 22216 24584 22228
rect 23799 22188 24584 22216
rect 23799 22185 23811 22188
rect 23753 22179 23811 22185
rect 22465 22151 22523 22157
rect 22465 22148 22477 22151
rect 21600 22120 21956 22148
rect 22036 22120 22477 22148
rect 21600 22108 21606 22120
rect 21269 22015 21327 22021
rect 21269 21981 21281 22015
rect 21315 21981 21327 22015
rect 21269 21975 21327 21981
rect 21361 22015 21419 22021
rect 21361 21981 21373 22015
rect 21407 21981 21419 22015
rect 21361 21975 21419 21981
rect 21450 21972 21456 22024
rect 21508 21972 21514 22024
rect 21542 21972 21548 22024
rect 21600 22012 21606 22024
rect 21729 22015 21787 22021
rect 21729 22012 21741 22015
rect 21600 21984 21741 22012
rect 21600 21972 21606 21984
rect 21729 21981 21741 21984
rect 21775 22012 21787 22015
rect 21818 22012 21824 22024
rect 21775 21984 21824 22012
rect 21775 21981 21787 21984
rect 21729 21975 21787 21981
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 21928 22021 21956 22120
rect 22465 22117 22477 22120
rect 22511 22148 22523 22151
rect 23934 22148 23940 22160
rect 22511 22120 23940 22148
rect 22511 22117 22523 22120
rect 22465 22111 22523 22117
rect 23934 22108 23940 22120
rect 23992 22108 23998 22160
rect 22554 22040 22560 22092
rect 22612 22040 22618 22092
rect 22997 22083 23055 22089
rect 22997 22080 23009 22083
rect 22664 22052 23009 22080
rect 21913 22015 21971 22021
rect 21913 21981 21925 22015
rect 21959 21981 21971 22015
rect 21913 21975 21971 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22664 22021 22692 22052
rect 22997 22049 23009 22052
rect 23043 22049 23055 22083
rect 23293 22083 23351 22089
rect 23293 22080 23305 22083
rect 22997 22043 23055 22049
rect 23124 22052 23305 22080
rect 23124 22024 23152 22052
rect 23293 22049 23305 22052
rect 23339 22049 23351 22083
rect 23293 22043 23351 22049
rect 23952 22024 23980 22108
rect 24136 22024 24164 22188
rect 24578 22176 24584 22188
rect 24636 22216 24642 22228
rect 24636 22188 26096 22216
rect 24636 22176 24642 22188
rect 24320 22120 25820 22148
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22152 21984 22385 22012
rect 22152 21972 22158 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22649 22015 22707 22021
rect 22649 21981 22661 22015
rect 22695 21981 22707 22015
rect 22649 21975 22707 21981
rect 22738 21972 22744 22024
rect 22796 21972 22802 22024
rect 22830 21972 22836 22024
rect 22888 21972 22894 22024
rect 23106 21972 23112 22024
rect 23164 21972 23170 22024
rect 23198 21972 23204 22024
rect 23256 22012 23262 22024
rect 23477 22015 23535 22021
rect 23477 22012 23489 22015
rect 23256 21984 23489 22012
rect 23256 21972 23262 21984
rect 23477 21981 23489 21984
rect 23523 21981 23535 22015
rect 23477 21975 23535 21981
rect 23750 21972 23756 22024
rect 23808 22012 23814 22024
rect 23845 22015 23903 22021
rect 23845 22012 23857 22015
rect 23808 21984 23857 22012
rect 23808 21972 23814 21984
rect 23845 21981 23857 21984
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 23934 21972 23940 22024
rect 23992 21972 23998 22024
rect 24118 21972 24124 22024
rect 24176 21972 24182 22024
rect 24213 22015 24271 22021
rect 24213 21981 24225 22015
rect 24259 22012 24271 22015
rect 24320 22012 24348 22120
rect 24765 22083 24823 22089
rect 24765 22049 24777 22083
rect 24811 22049 24823 22083
rect 24765 22043 24823 22049
rect 24964 22052 25176 22080
rect 24259 21984 24348 22012
rect 24259 21981 24271 21984
rect 24213 21975 24271 21981
rect 24394 21972 24400 22024
rect 24452 21972 24458 22024
rect 24486 21972 24492 22024
rect 24544 22006 24550 22024
rect 24581 22015 24639 22021
rect 24581 22006 24593 22015
rect 24544 21981 24593 22006
rect 24627 21981 24639 22015
rect 24544 21978 24639 21981
rect 24544 21972 24550 21978
rect 24581 21975 24639 21978
rect 21174 21944 21180 21956
rect 20180 21916 21180 21944
rect 21174 21904 21180 21916
rect 21232 21904 21238 21956
rect 22756 21944 22784 21972
rect 22925 21947 22983 21953
rect 22925 21944 22937 21947
rect 21284 21916 22600 21944
rect 22756 21916 22937 21944
rect 10284 21848 10456 21876
rect 10284 21836 10290 21848
rect 10502 21836 10508 21888
rect 10560 21836 10566 21888
rect 11057 21879 11115 21885
rect 11057 21845 11069 21879
rect 11103 21876 11115 21879
rect 12066 21876 12072 21888
rect 11103 21848 12072 21876
rect 11103 21845 11115 21848
rect 11057 21839 11115 21845
rect 12066 21836 12072 21848
rect 12124 21836 12130 21888
rect 12710 21836 12716 21888
rect 12768 21876 12774 21888
rect 13538 21876 13544 21888
rect 12768 21848 13544 21876
rect 12768 21836 12774 21848
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 16209 21879 16267 21885
rect 16209 21845 16221 21879
rect 16255 21876 16267 21879
rect 16482 21876 16488 21888
rect 16255 21848 16488 21876
rect 16255 21845 16267 21848
rect 16209 21839 16267 21845
rect 16482 21836 16488 21848
rect 16540 21876 16546 21888
rect 16666 21876 16672 21888
rect 16540 21848 16672 21876
rect 16540 21836 16546 21848
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 17862 21836 17868 21888
rect 17920 21836 17926 21888
rect 20346 21836 20352 21888
rect 20404 21836 20410 21888
rect 20438 21836 20444 21888
rect 20496 21876 20502 21888
rect 20717 21879 20775 21885
rect 20717 21876 20729 21879
rect 20496 21848 20729 21876
rect 20496 21836 20502 21848
rect 20717 21845 20729 21848
rect 20763 21876 20775 21879
rect 20990 21876 20996 21888
rect 20763 21848 20996 21876
rect 20763 21845 20775 21848
rect 20717 21839 20775 21845
rect 20990 21836 20996 21848
rect 21048 21876 21054 21888
rect 21284 21876 21312 21916
rect 21048 21848 21312 21876
rect 22189 21879 22247 21885
rect 21048 21836 21054 21848
rect 22189 21845 22201 21879
rect 22235 21876 22247 21879
rect 22462 21876 22468 21888
rect 22235 21848 22468 21876
rect 22235 21845 22247 21848
rect 22189 21839 22247 21845
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 22572 21876 22600 21916
rect 22925 21913 22937 21916
rect 22971 21913 22983 21947
rect 24781 21944 24809 22043
rect 24964 22024 24992 22052
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 22925 21907 22983 21913
rect 23492 21916 24809 21944
rect 23492 21888 23520 21916
rect 23109 21879 23167 21885
rect 23109 21876 23121 21879
rect 22572 21848 23121 21876
rect 23109 21845 23121 21848
rect 23155 21845 23167 21879
rect 23109 21839 23167 21845
rect 23474 21836 23480 21888
rect 23532 21836 23538 21888
rect 24035 21879 24093 21885
rect 24035 21845 24047 21879
rect 24081 21876 24093 21879
rect 24578 21876 24584 21888
rect 24081 21848 24584 21876
rect 24081 21845 24093 21848
rect 24035 21839 24093 21845
rect 24578 21836 24584 21848
rect 24636 21836 24642 21888
rect 24762 21836 24768 21888
rect 24820 21876 24826 21888
rect 24872 21876 24900 21975
rect 24946 21972 24952 22024
rect 25004 21972 25010 22024
rect 25038 21972 25044 22024
rect 25096 21972 25102 22024
rect 25148 22021 25176 22052
rect 25133 22015 25191 22021
rect 25133 21981 25145 22015
rect 25179 21981 25191 22015
rect 25133 21975 25191 21981
rect 25222 21972 25228 22024
rect 25280 22012 25286 22024
rect 25409 22015 25467 22021
rect 25409 22012 25421 22015
rect 25280 21984 25421 22012
rect 25280 21972 25286 21984
rect 25409 21981 25421 21984
rect 25455 21981 25467 22015
rect 25409 21975 25467 21981
rect 25498 21972 25504 22024
rect 25556 22012 25562 22024
rect 25685 22015 25743 22021
rect 25685 22012 25697 22015
rect 25556 21984 25697 22012
rect 25556 21972 25562 21984
rect 25685 21981 25697 21984
rect 25731 21981 25743 22015
rect 25685 21975 25743 21981
rect 25792 22012 25820 22120
rect 25961 22015 26019 22021
rect 25961 22012 25973 22015
rect 25792 21984 25973 22012
rect 25056 21944 25084 21972
rect 25317 21947 25375 21953
rect 25317 21944 25329 21947
rect 25056 21916 25329 21944
rect 25317 21913 25329 21916
rect 25363 21913 25375 21947
rect 25792 21944 25820 21984
rect 25961 21981 25973 21984
rect 26007 21981 26019 22015
rect 25961 21975 26019 21981
rect 25317 21907 25375 21913
rect 25424 21916 25820 21944
rect 25869 21947 25927 21953
rect 24820 21848 24900 21876
rect 24949 21879 25007 21885
rect 24820 21836 24826 21848
rect 24949 21845 24961 21879
rect 24995 21876 25007 21879
rect 25424 21876 25452 21916
rect 25869 21913 25881 21947
rect 25915 21944 25927 21947
rect 26068 21944 26096 22188
rect 28810 21972 28816 22024
rect 28868 21972 28874 22024
rect 28828 21944 28856 21972
rect 25915 21916 28856 21944
rect 25915 21913 25927 21916
rect 25869 21907 25927 21913
rect 24995 21848 25452 21876
rect 25501 21879 25559 21885
rect 24995 21845 25007 21848
rect 24949 21839 25007 21845
rect 25501 21845 25513 21879
rect 25547 21876 25559 21879
rect 25590 21876 25596 21888
rect 25547 21848 25596 21876
rect 25547 21845 25559 21848
rect 25501 21839 25559 21845
rect 25590 21836 25596 21848
rect 25648 21836 25654 21888
rect 1104 21786 29440 21808
rect 1104 21734 5151 21786
rect 5203 21734 5215 21786
rect 5267 21734 5279 21786
rect 5331 21734 5343 21786
rect 5395 21734 5407 21786
rect 5459 21734 12234 21786
rect 12286 21734 12298 21786
rect 12350 21734 12362 21786
rect 12414 21734 12426 21786
rect 12478 21734 12490 21786
rect 12542 21734 19317 21786
rect 19369 21734 19381 21786
rect 19433 21734 19445 21786
rect 19497 21734 19509 21786
rect 19561 21734 19573 21786
rect 19625 21734 26400 21786
rect 26452 21734 26464 21786
rect 26516 21734 26528 21786
rect 26580 21734 26592 21786
rect 26644 21734 26656 21786
rect 26708 21734 29440 21786
rect 1104 21712 29440 21734
rect 4154 21672 4160 21684
rect 3160 21644 4160 21672
rect 3160 21545 3188 21644
rect 4154 21632 4160 21644
rect 4212 21632 4218 21684
rect 4890 21672 4896 21684
rect 4448 21644 4896 21672
rect 3329 21607 3387 21613
rect 3329 21604 3341 21607
rect 3252 21576 3341 21604
rect 3252 21548 3280 21576
rect 3329 21573 3341 21576
rect 3375 21573 3387 21607
rect 3329 21567 3387 21573
rect 3421 21607 3479 21613
rect 3421 21573 3433 21607
rect 3467 21604 3479 21607
rect 4062 21604 4068 21616
rect 3467 21576 4068 21604
rect 3467 21573 3479 21576
rect 3421 21567 3479 21573
rect 4062 21564 4068 21576
rect 4120 21564 4126 21616
rect 4338 21564 4344 21616
rect 4396 21604 4402 21616
rect 4448 21604 4476 21644
rect 4890 21632 4896 21644
rect 4948 21632 4954 21684
rect 5534 21632 5540 21684
rect 5592 21632 5598 21684
rect 5626 21632 5632 21684
rect 5684 21672 5690 21684
rect 5684 21644 5764 21672
rect 5684 21632 5690 21644
rect 4396 21576 4554 21604
rect 4396 21564 4402 21576
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21505 3203 21539
rect 3145 21499 3203 21505
rect 3234 21496 3240 21548
rect 3292 21496 3298 21548
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21536 3571 21539
rect 3694 21536 3700 21548
rect 3559 21508 3700 21536
rect 3559 21505 3571 21508
rect 3513 21499 3571 21505
rect 3694 21496 3700 21508
rect 3752 21496 3758 21548
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21505 5687 21539
rect 5736 21536 5764 21644
rect 5902 21632 5908 21684
rect 5960 21632 5966 21684
rect 6178 21632 6184 21684
rect 6236 21632 6242 21684
rect 7926 21672 7932 21684
rect 6380 21644 7932 21672
rect 5920 21545 5948 21632
rect 5813 21539 5871 21545
rect 5813 21536 5825 21539
rect 5736 21508 5825 21536
rect 5629 21499 5687 21505
rect 5813 21505 5825 21508
rect 5859 21505 5871 21539
rect 5813 21499 5871 21505
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 3789 21471 3847 21477
rect 3789 21437 3801 21471
rect 3835 21437 3847 21471
rect 3789 21431 3847 21437
rect 4065 21471 4123 21477
rect 4065 21437 4077 21471
rect 4111 21468 4123 21471
rect 5074 21468 5080 21480
rect 4111 21440 5080 21468
rect 4111 21437 4123 21440
rect 4065 21431 4123 21437
rect 3804 21344 3832 21431
rect 5074 21428 5080 21440
rect 5132 21428 5138 21480
rect 5644 21468 5672 21499
rect 5994 21496 6000 21548
rect 6052 21496 6058 21548
rect 6380 21545 6408 21644
rect 7926 21632 7932 21644
rect 7984 21672 7990 21684
rect 9950 21672 9956 21684
rect 7984 21644 9956 21672
rect 7984 21632 7990 21644
rect 7098 21564 7104 21616
rect 7156 21564 7162 21616
rect 8386 21564 8392 21616
rect 8444 21564 8450 21616
rect 8478 21564 8484 21616
rect 8536 21564 8542 21616
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 8110 21496 8116 21548
rect 8168 21536 8174 21548
rect 8205 21539 8263 21545
rect 8205 21536 8217 21539
rect 8168 21508 8217 21536
rect 8168 21496 8174 21508
rect 8205 21505 8217 21508
rect 8251 21505 8263 21539
rect 8404 21536 8432 21564
rect 8404 21508 8524 21536
rect 8205 21499 8263 21505
rect 6641 21471 6699 21477
rect 5644 21440 6500 21468
rect 5828 21412 5856 21440
rect 5810 21360 5816 21412
rect 5868 21360 5874 21412
rect 3694 21292 3700 21344
rect 3752 21292 3758 21344
rect 3786 21292 3792 21344
rect 3844 21292 3850 21344
rect 4062 21292 4068 21344
rect 4120 21332 4126 21344
rect 5828 21332 5856 21360
rect 6472 21344 6500 21440
rect 6641 21437 6653 21471
rect 6687 21468 6699 21471
rect 8496 21468 8524 21508
rect 8570 21496 8576 21548
rect 8628 21496 8634 21548
rect 9048 21545 9076 21644
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 10778 21632 10784 21684
rect 10836 21672 10842 21684
rect 11054 21672 11060 21684
rect 10836 21644 11060 21672
rect 10836 21632 10842 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 14458 21672 14464 21684
rect 12912 21644 14464 21672
rect 10594 21604 10600 21616
rect 10534 21576 10600 21604
rect 10594 21564 10600 21576
rect 10652 21604 10658 21616
rect 10962 21604 10968 21616
rect 10652 21576 10968 21604
rect 10652 21564 10658 21576
rect 10962 21564 10968 21576
rect 11020 21564 11026 21616
rect 12437 21607 12495 21613
rect 12437 21573 12449 21607
rect 12483 21604 12495 21607
rect 12483 21576 12848 21604
rect 12483 21573 12495 21576
rect 12437 21567 12495 21573
rect 9033 21539 9091 21545
rect 9033 21505 9045 21539
rect 9079 21505 9091 21539
rect 9033 21499 9091 21505
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 12158 21496 12164 21548
rect 12216 21496 12222 21548
rect 12618 21545 12624 21548
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 12575 21539 12624 21545
rect 12575 21505 12587 21539
rect 12621 21505 12624 21539
rect 12575 21499 12624 21505
rect 9309 21471 9367 21477
rect 6687 21440 8248 21468
rect 8496 21440 9168 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 4120 21304 5856 21332
rect 4120 21292 4126 21304
rect 6454 21292 6460 21344
rect 6512 21292 6518 21344
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 7834 21332 7840 21344
rect 7432 21304 7840 21332
rect 7432 21292 7438 21304
rect 7834 21292 7840 21304
rect 7892 21332 7898 21344
rect 8113 21335 8171 21341
rect 8113 21332 8125 21335
rect 7892 21304 8125 21332
rect 7892 21292 7898 21304
rect 8113 21301 8125 21304
rect 8159 21301 8171 21335
rect 8220 21332 8248 21440
rect 8757 21403 8815 21409
rect 8757 21369 8769 21403
rect 8803 21369 8815 21403
rect 8757 21363 8815 21369
rect 8772 21332 8800 21363
rect 9140 21344 9168 21440
rect 9309 21437 9321 21471
rect 9355 21468 9367 21471
rect 10042 21468 10048 21480
rect 9355 21440 10048 21468
rect 9355 21437 9367 21440
rect 9309 21431 9367 21437
rect 10042 21428 10048 21440
rect 10100 21428 10106 21480
rect 12360 21468 12388 21499
rect 12618 21496 12624 21499
rect 12676 21496 12682 21548
rect 12710 21468 12716 21480
rect 12360 21440 12716 21468
rect 12710 21428 12716 21440
rect 12768 21428 12774 21480
rect 8220 21304 8800 21332
rect 8113 21295 8171 21301
rect 9122 21292 9128 21344
rect 9180 21292 9186 21344
rect 9490 21292 9496 21344
rect 9548 21332 9554 21344
rect 10594 21332 10600 21344
rect 9548 21304 10600 21332
rect 9548 21292 9554 21304
rect 10594 21292 10600 21304
rect 10652 21292 10658 21344
rect 10778 21292 10784 21344
rect 10836 21292 10842 21344
rect 12710 21292 12716 21344
rect 12768 21292 12774 21344
rect 12820 21332 12848 21576
rect 12912 21545 12940 21644
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 17770 21632 17776 21684
rect 17828 21672 17834 21684
rect 17828 21644 18092 21672
rect 17828 21632 17834 21644
rect 13078 21564 13084 21616
rect 13136 21604 13142 21616
rect 13630 21604 13636 21616
rect 13136 21576 13636 21604
rect 13136 21564 13142 21576
rect 13630 21564 13636 21576
rect 13688 21564 13694 21616
rect 12897 21539 12955 21545
rect 12897 21505 12909 21539
rect 12943 21505 12955 21539
rect 18064 21522 18092 21644
rect 18414 21632 18420 21684
rect 18472 21632 18478 21684
rect 20165 21675 20223 21681
rect 20165 21641 20177 21675
rect 20211 21672 20223 21675
rect 20211 21644 20760 21672
rect 20211 21641 20223 21644
rect 20165 21635 20223 21641
rect 19242 21564 19248 21616
rect 19300 21604 19306 21616
rect 20732 21604 20760 21644
rect 20806 21632 20812 21684
rect 20864 21632 20870 21684
rect 20990 21632 20996 21684
rect 21048 21672 21054 21684
rect 21545 21675 21603 21681
rect 21545 21672 21557 21675
rect 21048 21644 21557 21672
rect 21048 21632 21054 21644
rect 21545 21641 21557 21644
rect 21591 21641 21603 21675
rect 21545 21635 21603 21641
rect 22646 21632 22652 21684
rect 22704 21672 22710 21684
rect 23385 21675 23443 21681
rect 23385 21672 23397 21675
rect 22704 21644 23397 21672
rect 22704 21632 22710 21644
rect 23385 21641 23397 21644
rect 23431 21672 23443 21675
rect 23474 21672 23480 21684
rect 23431 21644 23480 21672
rect 23431 21641 23443 21644
rect 23385 21635 23443 21641
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 23566 21632 23572 21684
rect 23624 21632 23630 21684
rect 23661 21675 23719 21681
rect 23661 21641 23673 21675
rect 23707 21672 23719 21675
rect 24486 21672 24492 21684
rect 23707 21644 24492 21672
rect 23707 21641 23719 21644
rect 23661 21635 23719 21641
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 21174 21604 21180 21616
rect 19300 21576 20392 21604
rect 20732 21576 21180 21604
rect 19300 21564 19306 21576
rect 18506 21536 18512 21548
rect 12897 21499 12955 21505
rect 18156 21508 18512 21536
rect 13173 21471 13231 21477
rect 13173 21437 13185 21471
rect 13219 21468 13231 21471
rect 13262 21468 13268 21480
rect 13219 21440 13268 21468
rect 13219 21437 13231 21440
rect 13173 21431 13231 21437
rect 13262 21428 13268 21440
rect 13320 21428 13326 21480
rect 16574 21428 16580 21480
rect 16632 21468 16638 21480
rect 16669 21471 16727 21477
rect 16669 21468 16681 21471
rect 16632 21440 16681 21468
rect 16632 21428 16638 21440
rect 16669 21437 16681 21440
rect 16715 21437 16727 21471
rect 16669 21431 16727 21437
rect 16942 21428 16948 21480
rect 17000 21428 17006 21480
rect 18156 21468 18184 21508
rect 18506 21496 18512 21508
rect 18564 21536 18570 21548
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 18564 21508 18797 21536
rect 18564 21496 18570 21508
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 19150 21496 19156 21548
rect 19208 21496 19214 21548
rect 19334 21496 19340 21548
rect 19392 21496 19398 21548
rect 20364 21536 20392 21576
rect 21174 21564 21180 21576
rect 21232 21564 21238 21616
rect 21358 21564 21364 21616
rect 21416 21604 21422 21616
rect 23106 21604 23112 21616
rect 21416 21576 22140 21604
rect 21416 21564 21422 21576
rect 20364 21508 20760 21536
rect 17972 21440 18184 21468
rect 18693 21471 18751 21477
rect 12986 21332 12992 21344
rect 12820 21304 12992 21332
rect 12986 21292 12992 21304
rect 13044 21332 13050 21344
rect 14645 21335 14703 21341
rect 14645 21332 14657 21335
rect 13044 21304 14657 21332
rect 13044 21292 13050 21304
rect 14645 21301 14657 21304
rect 14691 21301 14703 21335
rect 14645 21295 14703 21301
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 17972 21332 18000 21440
rect 18693 21437 18705 21471
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 18509 21403 18567 21409
rect 18509 21369 18521 21403
rect 18555 21369 18567 21403
rect 18708 21400 18736 21431
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 18969 21471 19027 21477
rect 18969 21437 18981 21471
rect 19015 21468 19027 21471
rect 20346 21468 20352 21480
rect 19015 21440 20352 21468
rect 19015 21437 19027 21440
rect 18969 21431 19027 21437
rect 20346 21428 20352 21440
rect 20404 21428 20410 21480
rect 20530 21428 20536 21480
rect 20588 21428 20594 21480
rect 20625 21471 20683 21477
rect 20625 21437 20637 21471
rect 20671 21437 20683 21471
rect 20732 21468 20760 21508
rect 21082 21496 21088 21548
rect 21140 21536 21146 21548
rect 21453 21539 21511 21545
rect 21453 21536 21465 21539
rect 21140 21508 21465 21536
rect 21140 21496 21146 21508
rect 21453 21505 21465 21508
rect 21499 21505 21511 21539
rect 21453 21499 21511 21505
rect 21821 21539 21879 21545
rect 21821 21505 21833 21539
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 21266 21468 21272 21480
rect 20732 21440 21272 21468
rect 20625 21431 20683 21437
rect 18708 21372 19564 21400
rect 18509 21363 18567 21369
rect 14792 21304 18000 21332
rect 18524 21332 18552 21363
rect 19536 21344 19564 21372
rect 19242 21332 19248 21344
rect 18524 21304 19248 21332
rect 14792 21292 14798 21304
rect 19242 21292 19248 21304
rect 19300 21292 19306 21344
rect 19518 21292 19524 21344
rect 19576 21292 19582 21344
rect 20640 21332 20668 21431
rect 21266 21428 21272 21440
rect 21324 21428 21330 21480
rect 21358 21428 21364 21480
rect 21416 21428 21422 21480
rect 21468 21468 21496 21499
rect 21836 21468 21864 21499
rect 21910 21496 21916 21548
rect 21968 21536 21974 21548
rect 22112 21545 22140 21576
rect 22388 21576 23112 21604
rect 22388 21545 22416 21576
rect 23106 21564 23112 21576
rect 23164 21604 23170 21616
rect 23584 21604 23612 21632
rect 23164 21576 23612 21604
rect 23164 21564 23170 21576
rect 23750 21564 23756 21616
rect 23808 21604 23814 21616
rect 23808 21576 25360 21604
rect 23808 21564 23814 21576
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21968 21508 22017 21536
rect 21968 21496 21974 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 22097 21539 22155 21545
rect 22097 21505 22109 21539
rect 22143 21505 22155 21539
rect 22097 21499 22155 21505
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22462 21496 22468 21548
rect 22520 21496 22526 21548
rect 22738 21496 22744 21548
rect 22796 21536 22802 21548
rect 22833 21539 22891 21545
rect 22833 21536 22845 21539
rect 22796 21508 22845 21536
rect 22796 21496 22802 21508
rect 22833 21505 22845 21508
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 23382 21496 23388 21548
rect 23440 21496 23446 21548
rect 23566 21496 23572 21548
rect 23624 21536 23630 21548
rect 23845 21539 23903 21545
rect 23845 21536 23857 21539
rect 23624 21508 23857 21536
rect 23624 21496 23630 21508
rect 23845 21505 23857 21508
rect 23891 21536 23903 21539
rect 24026 21536 24032 21548
rect 23891 21508 24032 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 24026 21496 24032 21508
rect 24084 21496 24090 21548
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 24394 21536 24400 21548
rect 24351 21508 24400 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 24670 21496 24676 21548
rect 24728 21496 24734 21548
rect 24946 21496 24952 21548
rect 25004 21496 25010 21548
rect 25332 21545 25360 21576
rect 25317 21539 25375 21545
rect 25317 21505 25329 21539
rect 25363 21505 25375 21539
rect 25317 21499 25375 21505
rect 25498 21496 25504 21548
rect 25556 21496 25562 21548
rect 26970 21496 26976 21548
rect 27028 21496 27034 21548
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21536 27215 21539
rect 27522 21536 27528 21548
rect 27203 21508 27528 21536
rect 27203 21505 27215 21508
rect 27157 21499 27215 21505
rect 22189 21471 22247 21477
rect 22189 21468 22201 21471
rect 21468 21440 21588 21468
rect 21836 21440 22201 21468
rect 20714 21360 20720 21412
rect 20772 21400 20778 21412
rect 20901 21403 20959 21409
rect 20901 21400 20913 21403
rect 20772 21372 20913 21400
rect 20772 21360 20778 21372
rect 20901 21369 20913 21372
rect 20947 21400 20959 21403
rect 20947 21372 21496 21400
rect 20947 21369 20959 21372
rect 20901 21363 20959 21369
rect 21468 21344 21496 21372
rect 20990 21332 20996 21344
rect 20640 21304 20996 21332
rect 20990 21292 20996 21304
rect 21048 21292 21054 21344
rect 21450 21292 21456 21344
rect 21508 21292 21514 21344
rect 21560 21332 21588 21440
rect 22189 21437 22201 21440
rect 22235 21437 22247 21471
rect 22189 21431 22247 21437
rect 22554 21428 22560 21480
rect 22612 21428 22618 21480
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 22695 21440 22876 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 21818 21360 21824 21412
rect 21876 21360 21882 21412
rect 22646 21332 22652 21344
rect 21560 21304 22652 21332
rect 22646 21292 22652 21304
rect 22704 21292 22710 21344
rect 22848 21332 22876 21440
rect 22922 21428 22928 21480
rect 22980 21428 22986 21480
rect 23198 21360 23204 21412
rect 23256 21360 23262 21412
rect 23400 21400 23428 21496
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21468 23535 21471
rect 25590 21468 25596 21480
rect 23523 21440 25596 21468
rect 23523 21437 23535 21440
rect 23477 21431 23535 21437
rect 25590 21428 25596 21440
rect 25648 21428 25654 21480
rect 27172 21468 27200 21499
rect 27522 21496 27528 21508
rect 27580 21496 27586 21548
rect 27709 21539 27767 21545
rect 27709 21505 27721 21539
rect 27755 21536 27767 21539
rect 27798 21536 27804 21548
rect 27755 21508 27804 21536
rect 27755 21505 27767 21508
rect 27709 21499 27767 21505
rect 27798 21496 27804 21508
rect 27856 21496 27862 21548
rect 26252 21440 27200 21468
rect 26252 21412 26280 21440
rect 24397 21403 24455 21409
rect 23400 21372 24348 21400
rect 23658 21332 23664 21344
rect 22848 21304 23664 21332
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 23934 21292 23940 21344
rect 23992 21292 23998 21344
rect 24320 21332 24348 21372
rect 24397 21369 24409 21403
rect 24443 21400 24455 21403
rect 26234 21400 26240 21412
rect 24443 21372 26240 21400
rect 24443 21369 24455 21372
rect 24397 21363 24455 21369
rect 26234 21360 26240 21372
rect 26292 21360 26298 21412
rect 27062 21360 27068 21412
rect 27120 21360 27126 21412
rect 24946 21332 24952 21344
rect 24320 21304 24952 21332
rect 24946 21292 24952 21304
rect 25004 21292 25010 21344
rect 25317 21335 25375 21341
rect 25317 21301 25329 21335
rect 25363 21332 25375 21335
rect 27246 21332 27252 21344
rect 25363 21304 27252 21332
rect 25363 21301 25375 21304
rect 25317 21295 25375 21301
rect 27246 21292 27252 21304
rect 27304 21292 27310 21344
rect 27614 21292 27620 21344
rect 27672 21292 27678 21344
rect 1104 21242 29440 21264
rect 1104 21190 4491 21242
rect 4543 21190 4555 21242
rect 4607 21190 4619 21242
rect 4671 21190 4683 21242
rect 4735 21190 4747 21242
rect 4799 21190 11574 21242
rect 11626 21190 11638 21242
rect 11690 21190 11702 21242
rect 11754 21190 11766 21242
rect 11818 21190 11830 21242
rect 11882 21190 18657 21242
rect 18709 21190 18721 21242
rect 18773 21190 18785 21242
rect 18837 21190 18849 21242
rect 18901 21190 18913 21242
rect 18965 21190 25740 21242
rect 25792 21190 25804 21242
rect 25856 21190 25868 21242
rect 25920 21190 25932 21242
rect 25984 21190 25996 21242
rect 26048 21190 29440 21242
rect 1104 21168 29440 21190
rect 3694 21088 3700 21140
rect 3752 21128 3758 21140
rect 4046 21131 4104 21137
rect 4046 21128 4058 21131
rect 3752 21100 4058 21128
rect 3752 21088 3758 21100
rect 4046 21097 4058 21100
rect 4092 21097 4104 21131
rect 4046 21091 4104 21097
rect 5537 21131 5595 21137
rect 5537 21097 5549 21131
rect 5583 21128 5595 21131
rect 5718 21128 5724 21140
rect 5583 21100 5724 21128
rect 5583 21097 5595 21100
rect 5537 21091 5595 21097
rect 5718 21088 5724 21100
rect 5776 21088 5782 21140
rect 6362 21128 6368 21140
rect 5828 21100 6368 21128
rect 3786 20952 3792 21004
rect 3844 20992 3850 21004
rect 5828 20992 5856 21100
rect 6362 21088 6368 21100
rect 6420 21088 6426 21140
rect 7466 21088 7472 21140
rect 7524 21128 7530 21140
rect 10502 21128 10508 21140
rect 7524 21100 10508 21128
rect 7524 21088 7530 21100
rect 10502 21088 10508 21100
rect 10560 21128 10566 21140
rect 10560 21100 11652 21128
rect 10560 21088 10566 21100
rect 5902 21020 5908 21072
rect 5960 21060 5966 21072
rect 8570 21060 8576 21072
rect 5960 21032 8576 21060
rect 5960 21020 5966 21032
rect 8570 21020 8576 21032
rect 8628 21020 8634 21072
rect 10226 21020 10232 21072
rect 10284 21060 10290 21072
rect 10284 21032 11468 21060
rect 10284 21020 10290 21032
rect 9585 20995 9643 21001
rect 3844 20964 5856 20992
rect 6012 20964 7512 20992
rect 3844 20952 3850 20964
rect 1854 20884 1860 20936
rect 1912 20924 1918 20936
rect 3804 20924 3832 20952
rect 1912 20896 3832 20924
rect 1912 20884 1918 20896
rect 5534 20884 5540 20936
rect 5592 20884 5598 20936
rect 5902 20884 5908 20936
rect 5960 20924 5966 20936
rect 6012 20933 6040 20964
rect 5997 20927 6055 20933
rect 5997 20924 6009 20927
rect 5960 20896 6009 20924
rect 5960 20884 5966 20896
rect 5997 20893 6009 20896
rect 6043 20893 6055 20927
rect 5997 20887 6055 20893
rect 6090 20927 6148 20933
rect 6090 20893 6102 20927
rect 6136 20893 6148 20927
rect 6090 20887 6148 20893
rect 6503 20927 6561 20933
rect 6503 20893 6515 20927
rect 6549 20924 6561 20927
rect 6730 20924 6736 20936
rect 6549 20896 6736 20924
rect 6549 20893 6561 20896
rect 6503 20887 6561 20893
rect 5552 20856 5580 20884
rect 6104 20856 6132 20887
rect 6730 20884 6736 20896
rect 6788 20924 6794 20936
rect 7300 20933 7328 20964
rect 7285 20927 7343 20933
rect 6788 20896 7236 20924
rect 6788 20884 6794 20896
rect 4448 20828 4554 20856
rect 5552 20828 6132 20856
rect 3418 20748 3424 20800
rect 3476 20788 3482 20800
rect 4338 20788 4344 20800
rect 3476 20760 4344 20788
rect 3476 20748 3482 20760
rect 4338 20748 4344 20760
rect 4396 20788 4402 20800
rect 4448 20788 4476 20828
rect 6178 20816 6184 20868
rect 6236 20856 6242 20868
rect 6273 20859 6331 20865
rect 6273 20856 6285 20859
rect 6236 20828 6285 20856
rect 6236 20816 6242 20828
rect 6273 20825 6285 20828
rect 6319 20825 6331 20859
rect 6273 20819 6331 20825
rect 6365 20859 6423 20865
rect 6365 20825 6377 20859
rect 6411 20825 6423 20859
rect 6365 20819 6423 20825
rect 4396 20760 4476 20788
rect 4396 20748 4402 20760
rect 5718 20748 5724 20800
rect 5776 20788 5782 20800
rect 6380 20788 6408 20819
rect 5776 20760 6408 20788
rect 6641 20791 6699 20797
rect 5776 20748 5782 20760
rect 6641 20757 6653 20791
rect 6687 20788 6699 20791
rect 6914 20788 6920 20800
rect 6687 20760 6920 20788
rect 6687 20757 6699 20760
rect 6641 20751 6699 20757
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 7208 20788 7236 20896
rect 7285 20893 7297 20927
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 7374 20884 7380 20936
rect 7432 20884 7438 20936
rect 7484 20924 7512 20964
rect 7668 20964 7880 20992
rect 7668 20924 7696 20964
rect 7484 20896 7696 20924
rect 7750 20927 7808 20933
rect 7750 20893 7762 20927
rect 7796 20893 7808 20927
rect 7852 20924 7880 20964
rect 9585 20961 9597 20995
rect 9631 20992 9643 20995
rect 10778 20992 10784 21004
rect 9631 20964 10784 20992
rect 9631 20961 9643 20964
rect 9585 20955 9643 20961
rect 10778 20952 10784 20964
rect 10836 20952 10842 21004
rect 11440 20936 11468 21032
rect 10226 20924 10232 20936
rect 7852 20896 10232 20924
rect 7750 20887 7808 20893
rect 7466 20816 7472 20868
rect 7524 20856 7530 20868
rect 7561 20859 7619 20865
rect 7561 20856 7573 20859
rect 7524 20828 7573 20856
rect 7524 20816 7530 20828
rect 7561 20825 7573 20828
rect 7607 20825 7619 20859
rect 7561 20819 7619 20825
rect 7650 20816 7656 20868
rect 7708 20816 7714 20868
rect 7760 20788 7788 20887
rect 10226 20884 10232 20896
rect 10284 20884 10290 20936
rect 10413 20927 10471 20933
rect 10413 20893 10425 20927
rect 10459 20924 10471 20927
rect 10870 20924 10876 20936
rect 10459 20896 10876 20924
rect 10459 20893 10471 20896
rect 10413 20887 10471 20893
rect 10870 20884 10876 20896
rect 10928 20884 10934 20936
rect 11422 20884 11428 20936
rect 11480 20884 11486 20936
rect 11514 20884 11520 20936
rect 11572 20884 11578 20936
rect 11624 20924 11652 21100
rect 14734 21088 14740 21140
rect 14792 21088 14798 21140
rect 16485 21131 16543 21137
rect 16485 21097 16497 21131
rect 16531 21128 16543 21131
rect 16942 21128 16948 21140
rect 16531 21100 16948 21128
rect 16531 21097 16543 21100
rect 16485 21091 16543 21097
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17862 21088 17868 21140
rect 17920 21088 17926 21140
rect 19058 21128 19064 21140
rect 18064 21100 19064 21128
rect 13446 21020 13452 21072
rect 13504 21060 13510 21072
rect 13504 21032 14320 21060
rect 13504 21020 13510 21032
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 12161 20995 12219 21001
rect 12161 20992 12173 20995
rect 11848 20964 12173 20992
rect 11848 20952 11854 20964
rect 12161 20961 12173 20964
rect 12207 20961 12219 20995
rect 12161 20955 12219 20961
rect 12437 20995 12495 21001
rect 12437 20961 12449 20995
rect 12483 20992 12495 20995
rect 13906 20992 13912 21004
rect 12483 20964 13912 20992
rect 12483 20961 12495 20964
rect 12437 20955 12495 20961
rect 13906 20952 13912 20964
rect 13964 20952 13970 21004
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 11624 20896 11713 20924
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 11890 20927 11948 20933
rect 11890 20893 11902 20927
rect 11936 20924 11948 20927
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 11936 20896 12020 20924
rect 11936 20893 11948 20896
rect 11890 20887 11948 20893
rect 9950 20816 9956 20868
rect 10008 20856 10014 20868
rect 11146 20856 11152 20868
rect 10008 20828 11152 20856
rect 10008 20816 10014 20828
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 11793 20859 11851 20865
rect 11793 20825 11805 20859
rect 11839 20825 11851 20859
rect 11793 20819 11851 20825
rect 7208 20760 7788 20788
rect 7929 20791 7987 20797
rect 7929 20757 7941 20791
rect 7975 20788 7987 20791
rect 8570 20788 8576 20800
rect 7975 20760 8576 20788
rect 7975 20757 7987 20760
rect 7929 20751 7987 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 10134 20748 10140 20800
rect 10192 20748 10198 20800
rect 10778 20748 10784 20800
rect 10836 20788 10842 20800
rect 11808 20788 11836 20819
rect 11992 20800 12020 20896
rect 13740 20896 14105 20924
rect 12894 20816 12900 20868
rect 12952 20816 12958 20868
rect 10836 20760 11836 20788
rect 10836 20748 10842 20760
rect 11974 20748 11980 20800
rect 12032 20748 12038 20800
rect 12069 20791 12127 20797
rect 12069 20757 12081 20791
rect 12115 20788 12127 20791
rect 13740 20788 13768 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 14182 20884 14188 20936
rect 14240 20884 14246 20936
rect 14292 20924 14320 21032
rect 17880 20992 17908 21088
rect 18064 21004 18092 21100
rect 19058 21088 19064 21100
rect 19116 21128 19122 21140
rect 19116 21100 19334 21128
rect 19116 21088 19122 21100
rect 19306 21060 19334 21100
rect 20990 21088 20996 21140
rect 21048 21128 21054 21140
rect 22186 21128 22192 21140
rect 21048 21100 22192 21128
rect 21048 21088 21054 21100
rect 19306 21032 20024 21060
rect 15948 20964 17908 20992
rect 15948 20933 15976 20964
rect 18046 20952 18052 21004
rect 18104 20952 18110 21004
rect 18325 20995 18383 21001
rect 18325 20961 18337 20995
rect 18371 20992 18383 20995
rect 18509 20995 18567 21001
rect 18509 20992 18521 20995
rect 18371 20964 18521 20992
rect 18371 20961 18383 20964
rect 18325 20955 18383 20961
rect 18509 20961 18521 20964
rect 18555 20992 18567 20995
rect 19150 20992 19156 21004
rect 18555 20964 19156 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 19150 20952 19156 20964
rect 19208 20952 19214 21004
rect 19518 20992 19524 21004
rect 19444 20964 19524 20992
rect 14558 20927 14616 20933
rect 14558 20924 14570 20927
rect 14292 20896 14570 20924
rect 14558 20893 14570 20896
rect 14604 20893 14616 20927
rect 14558 20887 14616 20893
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20893 14887 20927
rect 14829 20887 14887 20893
rect 15933 20927 15991 20933
rect 15933 20893 15945 20927
rect 15979 20893 15991 20927
rect 15933 20887 15991 20893
rect 14369 20859 14427 20865
rect 14369 20856 14381 20859
rect 13832 20828 14381 20856
rect 13832 20800 13860 20828
rect 14369 20825 14381 20828
rect 14415 20825 14427 20859
rect 14369 20819 14427 20825
rect 14461 20859 14519 20865
rect 14461 20825 14473 20859
rect 14507 20856 14519 20859
rect 14844 20856 14872 20887
rect 16022 20884 16028 20936
rect 16080 20924 16086 20936
rect 16301 20927 16359 20933
rect 16301 20924 16313 20927
rect 16080 20896 16313 20924
rect 16080 20884 16086 20896
rect 16301 20893 16313 20896
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 16574 20884 16580 20936
rect 16632 20884 16638 20936
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 19444 20933 19472 20964
rect 19518 20952 19524 20964
rect 19576 20952 19582 21004
rect 19996 20933 20024 21032
rect 20346 20952 20352 21004
rect 20404 20952 20410 21004
rect 21192 20992 21220 21100
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 23477 21131 23535 21137
rect 23477 21097 23489 21131
rect 23523 21128 23535 21131
rect 23566 21128 23572 21140
rect 23523 21100 23572 21128
rect 23523 21097 23535 21100
rect 23477 21091 23535 21097
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 25590 21088 25596 21140
rect 25648 21088 25654 21140
rect 25869 21131 25927 21137
rect 25869 21097 25881 21131
rect 25915 21128 25927 21131
rect 26142 21128 26148 21140
rect 25915 21100 26148 21128
rect 25915 21097 25927 21100
rect 25869 21091 25927 21097
rect 26142 21088 26148 21100
rect 26200 21088 26206 21140
rect 26970 21088 26976 21140
rect 27028 21128 27034 21140
rect 27065 21131 27123 21137
rect 27065 21128 27077 21131
rect 27028 21100 27077 21128
rect 27028 21088 27034 21100
rect 27065 21097 27077 21100
rect 27111 21128 27123 21131
rect 27801 21131 27859 21137
rect 27801 21128 27813 21131
rect 27111 21100 27813 21128
rect 27111 21097 27123 21100
rect 27065 21091 27123 21097
rect 27801 21097 27813 21100
rect 27847 21097 27859 21131
rect 27801 21091 27859 21097
rect 21545 21063 21603 21069
rect 21545 21029 21557 21063
rect 21591 21060 21603 21063
rect 21726 21060 21732 21072
rect 21591 21032 21732 21060
rect 21591 21029 21603 21032
rect 21545 21023 21603 21029
rect 21726 21020 21732 21032
rect 21784 21020 21790 21072
rect 22830 21020 22836 21072
rect 22888 21060 22894 21072
rect 23293 21063 23351 21069
rect 23293 21060 23305 21063
rect 22888 21032 23305 21060
rect 22888 21020 22894 21032
rect 23293 21029 23305 21032
rect 23339 21029 23351 21063
rect 23293 21023 23351 21029
rect 23937 20995 23995 21001
rect 23937 20992 23949 20995
rect 20456 20964 21220 20992
rect 19429 20927 19487 20933
rect 17920 20896 18552 20924
rect 17920 20884 17926 20896
rect 18524 20868 18552 20896
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20893 20039 20927
rect 19981 20887 20039 20893
rect 14507 20828 14872 20856
rect 14507 20825 14519 20828
rect 14461 20819 14519 20825
rect 12115 20760 13768 20788
rect 12115 20757 12127 20760
rect 12069 20751 12127 20757
rect 13814 20748 13820 20800
rect 13872 20748 13878 20800
rect 13909 20791 13967 20797
rect 13909 20757 13921 20791
rect 13955 20788 13967 20791
rect 14476 20788 14504 20819
rect 15746 20816 15752 20868
rect 15804 20856 15810 20868
rect 16117 20859 16175 20865
rect 16117 20856 16129 20859
rect 15804 20828 16129 20856
rect 15804 20816 15810 20828
rect 16117 20825 16129 20828
rect 16163 20825 16175 20859
rect 16117 20819 16175 20825
rect 16206 20816 16212 20868
rect 16264 20816 16270 20868
rect 16853 20859 16911 20865
rect 16853 20825 16865 20859
rect 16899 20856 16911 20859
rect 16942 20856 16948 20868
rect 16899 20828 16948 20856
rect 16899 20825 16911 20828
rect 16853 20819 16911 20825
rect 16942 20816 16948 20828
rect 17000 20816 17006 20868
rect 18506 20816 18512 20868
rect 18564 20816 18570 20868
rect 18598 20816 18604 20868
rect 18656 20856 18662 20868
rect 19812 20856 19840 20887
rect 18656 20828 19840 20856
rect 18656 20816 18662 20828
rect 13955 20760 14504 20788
rect 13955 20757 13967 20760
rect 13909 20751 13967 20757
rect 14550 20748 14556 20800
rect 14608 20788 14614 20800
rect 15473 20791 15531 20797
rect 15473 20788 15485 20791
rect 14608 20760 15485 20788
rect 14608 20748 14614 20760
rect 15473 20757 15485 20760
rect 15519 20757 15531 20791
rect 15473 20751 15531 20757
rect 17494 20748 17500 20800
rect 17552 20788 17558 20800
rect 19061 20791 19119 20797
rect 19061 20788 19073 20791
rect 17552 20760 19073 20788
rect 17552 20748 17558 20760
rect 19061 20757 19073 20760
rect 19107 20757 19119 20791
rect 19061 20751 19119 20757
rect 19150 20748 19156 20800
rect 19208 20788 19214 20800
rect 20456 20788 20484 20964
rect 20530 20884 20536 20936
rect 20588 20924 20594 20936
rect 20625 20927 20683 20933
rect 20625 20924 20637 20927
rect 20588 20896 20637 20924
rect 20588 20884 20594 20896
rect 20625 20893 20637 20896
rect 20671 20924 20683 20927
rect 20901 20927 20959 20933
rect 20901 20924 20913 20927
rect 20671 20896 20913 20924
rect 20671 20893 20683 20896
rect 20625 20887 20683 20893
rect 20901 20893 20913 20896
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 21085 20927 21143 20933
rect 21085 20893 21097 20927
rect 21131 20924 21143 20927
rect 21192 20924 21220 20964
rect 21376 20964 22324 20992
rect 21376 20936 21404 20964
rect 21131 20896 21220 20924
rect 21131 20893 21143 20896
rect 21085 20887 21143 20893
rect 20916 20856 20944 20887
rect 21266 20884 21272 20936
rect 21324 20884 21330 20936
rect 21358 20884 21364 20936
rect 21416 20884 21422 20936
rect 21450 20884 21456 20936
rect 21508 20884 21514 20936
rect 22186 20924 22192 20936
rect 21652 20896 22192 20924
rect 21177 20859 21235 20865
rect 20916 20828 21036 20856
rect 19208 20760 20484 20788
rect 21008 20788 21036 20828
rect 21177 20825 21189 20859
rect 21223 20856 21235 20859
rect 21542 20856 21548 20868
rect 21223 20828 21548 20856
rect 21223 20825 21235 20828
rect 21177 20819 21235 20825
rect 21542 20816 21548 20828
rect 21600 20856 21606 20868
rect 21652 20856 21680 20896
rect 22186 20884 22192 20896
rect 22244 20884 22250 20936
rect 22296 20933 22324 20964
rect 22664 20964 23949 20992
rect 22664 20936 22692 20964
rect 23937 20961 23949 20964
rect 23983 20961 23995 20995
rect 23937 20955 23995 20961
rect 25225 20995 25283 21001
rect 25225 20961 25237 20995
rect 25271 20992 25283 20995
rect 25608 20992 25636 21088
rect 27982 21060 27988 21072
rect 27448 21032 27988 21060
rect 26697 20995 26755 21001
rect 26697 20992 26709 20995
rect 25271 20964 25636 20992
rect 26068 20964 26709 20992
rect 25271 20961 25283 20964
rect 25225 20955 25283 20961
rect 22281 20927 22339 20933
rect 22281 20893 22293 20927
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 21600 20828 21680 20856
rect 22296 20856 22324 20887
rect 22646 20884 22652 20936
rect 22704 20884 22710 20936
rect 22738 20884 22744 20936
rect 22796 20924 22802 20936
rect 23017 20927 23075 20933
rect 23017 20924 23029 20927
rect 22796 20896 23029 20924
rect 22796 20884 22802 20896
rect 23017 20893 23029 20896
rect 23063 20924 23075 20927
rect 23661 20927 23719 20933
rect 23661 20924 23673 20927
rect 23063 20896 23673 20924
rect 23063 20893 23075 20896
rect 23017 20887 23075 20893
rect 23661 20893 23673 20896
rect 23707 20893 23719 20927
rect 23661 20887 23719 20893
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20893 23903 20927
rect 23845 20887 23903 20893
rect 23860 20856 23888 20887
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 24949 20927 25007 20933
rect 24949 20924 24961 20927
rect 24912 20896 24961 20924
rect 24912 20884 24918 20896
rect 24949 20893 24961 20896
rect 24995 20893 25007 20927
rect 24949 20887 25007 20893
rect 24210 20856 24216 20868
rect 22296 20828 24216 20856
rect 21600 20816 21606 20828
rect 24210 20816 24216 20828
rect 24268 20816 24274 20868
rect 25314 20816 25320 20868
rect 25372 20856 25378 20868
rect 25866 20856 25872 20868
rect 25372 20828 25872 20856
rect 25372 20816 25378 20828
rect 25866 20816 25872 20828
rect 25924 20816 25930 20868
rect 23290 20788 23296 20800
rect 21008 20760 23296 20788
rect 19208 20748 19214 20760
rect 23290 20748 23296 20760
rect 23348 20788 23354 20800
rect 23842 20788 23848 20800
rect 23348 20760 23848 20788
rect 23348 20748 23354 20760
rect 23842 20748 23848 20760
rect 23900 20748 23906 20800
rect 26068 20797 26096 20964
rect 26697 20961 26709 20964
rect 26743 20992 26755 20995
rect 27062 20992 27068 21004
rect 26743 20964 27068 20992
rect 26743 20961 26755 20964
rect 26697 20955 26755 20961
rect 27062 20952 27068 20964
rect 27120 20992 27126 21004
rect 27448 20992 27476 21032
rect 27982 21020 27988 21032
rect 28040 21020 28046 21072
rect 27120 20964 27476 20992
rect 27120 20952 27126 20964
rect 26145 20927 26203 20933
rect 26145 20893 26157 20927
rect 26191 20924 26203 20927
rect 26234 20924 26240 20936
rect 26191 20896 26240 20924
rect 26191 20893 26203 20896
rect 26145 20887 26203 20893
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 26786 20884 26792 20936
rect 26844 20884 26850 20936
rect 27448 20933 27476 20964
rect 27522 20952 27528 21004
rect 27580 20952 27586 21004
rect 27617 20995 27675 21001
rect 27617 20961 27629 20995
rect 27663 20992 27675 20995
rect 27798 20992 27804 21004
rect 27663 20964 27804 20992
rect 27663 20961 27675 20964
rect 27617 20955 27675 20961
rect 27798 20952 27804 20964
rect 27856 20992 27862 21004
rect 28902 20992 28908 21004
rect 27856 20964 28908 20992
rect 27856 20952 27862 20964
rect 28902 20952 28908 20964
rect 28960 20952 28966 21004
rect 27341 20927 27399 20933
rect 27341 20893 27353 20927
rect 27387 20893 27399 20927
rect 27341 20887 27399 20893
rect 27433 20927 27491 20933
rect 27433 20893 27445 20927
rect 27479 20893 27491 20927
rect 27540 20924 27568 20952
rect 27709 20927 27767 20933
rect 27709 20924 27721 20927
rect 27540 20896 27721 20924
rect 27433 20887 27491 20893
rect 27709 20893 27721 20896
rect 27755 20893 27767 20927
rect 28445 20927 28503 20933
rect 28445 20924 28457 20927
rect 27709 20887 27767 20893
rect 27816 20896 28457 20924
rect 27356 20856 27384 20887
rect 27816 20856 27844 20896
rect 28445 20893 28457 20896
rect 28491 20893 28503 20927
rect 28445 20887 28503 20893
rect 27356 20828 27844 20856
rect 27448 20800 27476 20828
rect 27982 20816 27988 20868
rect 28040 20856 28046 20868
rect 28261 20859 28319 20865
rect 28261 20856 28273 20859
rect 28040 20828 28273 20856
rect 28040 20816 28046 20828
rect 28261 20825 28273 20828
rect 28307 20825 28319 20859
rect 28261 20819 28319 20825
rect 25777 20791 25835 20797
rect 25777 20757 25789 20791
rect 25823 20788 25835 20791
rect 26053 20791 26111 20797
rect 26053 20788 26065 20791
rect 25823 20760 26065 20788
rect 25823 20757 25835 20760
rect 25777 20751 25835 20757
rect 26053 20757 26065 20760
rect 26099 20757 26111 20791
rect 26053 20751 26111 20757
rect 27430 20748 27436 20800
rect 27488 20748 27494 20800
rect 28166 20748 28172 20800
rect 28224 20748 28230 20800
rect 28534 20748 28540 20800
rect 28592 20788 28598 20800
rect 28629 20791 28687 20797
rect 28629 20788 28641 20791
rect 28592 20760 28641 20788
rect 28592 20748 28598 20760
rect 28629 20757 28641 20760
rect 28675 20757 28687 20791
rect 28629 20751 28687 20757
rect 1104 20698 29440 20720
rect 1104 20646 5151 20698
rect 5203 20646 5215 20698
rect 5267 20646 5279 20698
rect 5331 20646 5343 20698
rect 5395 20646 5407 20698
rect 5459 20646 12234 20698
rect 12286 20646 12298 20698
rect 12350 20646 12362 20698
rect 12414 20646 12426 20698
rect 12478 20646 12490 20698
rect 12542 20646 19317 20698
rect 19369 20646 19381 20698
rect 19433 20646 19445 20698
rect 19497 20646 19509 20698
rect 19561 20646 19573 20698
rect 19625 20646 26400 20698
rect 26452 20646 26464 20698
rect 26516 20646 26528 20698
rect 26580 20646 26592 20698
rect 26644 20646 26656 20698
rect 26708 20646 29440 20698
rect 1104 20624 29440 20646
rect 3528 20556 4752 20584
rect 3528 20525 3556 20556
rect 3513 20519 3571 20525
rect 3513 20485 3525 20519
rect 3559 20485 3571 20519
rect 3513 20479 3571 20485
rect 3605 20519 3663 20525
rect 3605 20485 3617 20519
rect 3651 20516 3663 20519
rect 4062 20516 4068 20528
rect 3651 20488 4068 20516
rect 3651 20485 3663 20488
rect 3605 20479 3663 20485
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 4338 20516 4344 20528
rect 4172 20488 4344 20516
rect 3329 20451 3387 20457
rect 3329 20417 3341 20451
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 3697 20451 3755 20457
rect 3697 20417 3709 20451
rect 3743 20448 3755 20451
rect 4172 20448 4200 20488
rect 4338 20476 4344 20488
rect 4396 20516 4402 20528
rect 4396 20488 4476 20516
rect 4396 20476 4402 20488
rect 4448 20457 4476 20488
rect 3743 20420 4200 20448
rect 4249 20451 4307 20457
rect 3743 20417 3755 20420
rect 3697 20411 3755 20417
rect 4249 20417 4261 20451
rect 4295 20417 4307 20451
rect 4249 20411 4307 20417
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20417 4491 20451
rect 4433 20411 4491 20417
rect 3344 20380 3372 20411
rect 3344 20352 4016 20380
rect 3988 20256 4016 20352
rect 3878 20204 3884 20256
rect 3936 20204 3942 20256
rect 3970 20204 3976 20256
rect 4028 20204 4034 20256
rect 4264 20244 4292 20411
rect 4724 20389 4752 20556
rect 6178 20544 6184 20596
rect 6236 20584 6242 20596
rect 7466 20584 7472 20596
rect 6236 20556 7472 20584
rect 6236 20544 6242 20556
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 9858 20544 9864 20596
rect 9916 20584 9922 20596
rect 9916 20556 9996 20584
rect 9916 20544 9922 20556
rect 7098 20476 7104 20528
rect 7156 20476 7162 20528
rect 9692 20516 9720 20544
rect 9968 20525 9996 20556
rect 10042 20544 10048 20596
rect 10100 20584 10106 20596
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 10100 20556 10885 20584
rect 10100 20544 10106 20556
rect 10873 20553 10885 20556
rect 10919 20553 10931 20587
rect 10873 20547 10931 20553
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13136 20556 13860 20584
rect 13136 20544 13142 20556
rect 9953 20519 10011 20525
rect 9692 20488 9812 20516
rect 9674 20408 9680 20460
rect 9732 20408 9738 20460
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 4890 20380 4896 20392
rect 4755 20352 4896 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 6362 20340 6368 20392
rect 6420 20340 6426 20392
rect 6638 20340 6644 20392
rect 6696 20340 6702 20392
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 8128 20352 8217 20380
rect 4982 20244 4988 20256
rect 4264 20216 4988 20244
rect 4982 20204 4988 20216
rect 5040 20244 5046 20256
rect 7006 20244 7012 20256
rect 5040 20216 7012 20244
rect 5040 20204 5046 20216
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 8128 20253 8156 20352
rect 8205 20349 8217 20352
rect 8251 20349 8263 20383
rect 9784 20380 9812 20488
rect 9953 20485 9965 20519
rect 9999 20485 10011 20519
rect 9953 20479 10011 20485
rect 10060 20488 11008 20516
rect 9858 20408 9864 20460
rect 9916 20408 9922 20460
rect 10060 20457 10088 20488
rect 10980 20460 11008 20488
rect 12802 20476 12808 20528
rect 12860 20476 12866 20528
rect 13832 20516 13860 20556
rect 13906 20544 13912 20596
rect 13964 20584 13970 20596
rect 14921 20587 14979 20593
rect 14921 20584 14933 20587
rect 13964 20556 14933 20584
rect 13964 20544 13970 20556
rect 14921 20553 14933 20556
rect 14967 20553 14979 20587
rect 14921 20547 14979 20553
rect 15010 20544 15016 20596
rect 15068 20584 15074 20596
rect 16945 20587 17003 20593
rect 16945 20584 16957 20587
rect 15068 20556 16957 20584
rect 15068 20544 15074 20556
rect 16945 20553 16957 20556
rect 16991 20553 17003 20587
rect 21361 20587 21419 20593
rect 16945 20547 17003 20553
rect 17236 20556 17908 20584
rect 16206 20516 16212 20528
rect 13832 20488 16212 20516
rect 16206 20476 16212 20488
rect 16264 20476 16270 20528
rect 17055 20519 17113 20525
rect 17055 20485 17067 20519
rect 17101 20516 17113 20519
rect 17236 20516 17264 20556
rect 17101 20488 17264 20516
rect 17101 20485 17113 20488
rect 17055 20479 17113 20485
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 10134 20408 10140 20460
rect 10192 20448 10198 20460
rect 10321 20451 10379 20457
rect 10321 20448 10333 20451
rect 10192 20420 10333 20448
rect 10192 20408 10198 20420
rect 10321 20417 10333 20420
rect 10367 20417 10379 20451
rect 10321 20411 10379 20417
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 10520 20380 10548 20411
rect 10594 20408 10600 20460
rect 10652 20408 10658 20460
rect 10686 20408 10692 20460
rect 10744 20408 10750 20460
rect 10962 20408 10968 20460
rect 11020 20408 11026 20460
rect 11146 20408 11152 20460
rect 11204 20448 11210 20460
rect 11790 20448 11796 20460
rect 11204 20420 11796 20448
rect 11204 20408 11210 20420
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20448 13783 20451
rect 14182 20448 14188 20460
rect 13771 20420 14188 20448
rect 13771 20417 13783 20420
rect 13725 20411 13783 20417
rect 9784 20352 10548 20380
rect 8205 20343 8263 20349
rect 8478 20272 8484 20324
rect 8536 20312 8542 20324
rect 10229 20315 10287 20321
rect 10229 20312 10241 20315
rect 8536 20284 10241 20312
rect 8536 20272 8542 20284
rect 10229 20281 10241 20284
rect 10275 20281 10287 20315
rect 10229 20275 10287 20281
rect 8113 20247 8171 20253
rect 8113 20244 8125 20247
rect 7248 20216 8125 20244
rect 7248 20204 7254 20216
rect 8113 20213 8125 20216
rect 8159 20213 8171 20247
rect 8113 20207 8171 20213
rect 8202 20204 8208 20256
rect 8260 20244 8266 20256
rect 8849 20247 8907 20253
rect 8849 20244 8861 20247
rect 8260 20216 8861 20244
rect 8260 20204 8266 20216
rect 8849 20213 8861 20216
rect 8895 20213 8907 20247
rect 8849 20207 8907 20213
rect 10134 20204 10140 20256
rect 10192 20244 10198 20256
rect 10336 20244 10364 20352
rect 10192 20216 10364 20244
rect 10612 20244 10640 20408
rect 12066 20340 12072 20392
rect 12124 20340 12130 20392
rect 13541 20383 13599 20389
rect 13541 20349 13553 20383
rect 13587 20380 13599 20383
rect 13740 20380 13768 20411
rect 14182 20408 14188 20420
rect 14240 20408 14246 20460
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20448 14427 20451
rect 14458 20448 14464 20460
rect 14415 20420 14464 20448
rect 14415 20417 14427 20420
rect 14369 20411 14427 20417
rect 14458 20408 14464 20420
rect 14516 20408 14522 20460
rect 14550 20408 14556 20460
rect 14608 20408 14614 20460
rect 14645 20451 14703 20457
rect 14645 20417 14657 20451
rect 14691 20417 14703 20451
rect 14645 20411 14703 20417
rect 13587 20352 13768 20380
rect 13587 20349 13599 20352
rect 13541 20343 13599 20349
rect 14660 20324 14688 20411
rect 14734 20408 14740 20460
rect 14792 20408 14798 20460
rect 16850 20408 16856 20460
rect 16908 20408 16914 20460
rect 17218 20408 17224 20460
rect 17276 20408 17282 20460
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20448 17371 20451
rect 17402 20448 17408 20460
rect 17359 20420 17408 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 17494 20408 17500 20460
rect 17552 20408 17558 20460
rect 17586 20408 17592 20460
rect 17644 20408 17650 20460
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20448 17739 20451
rect 17770 20448 17776 20460
rect 17727 20420 17776 20448
rect 17727 20417 17739 20420
rect 17681 20411 17739 20417
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 17880 20448 17908 20556
rect 21361 20553 21373 20587
rect 21407 20584 21419 20587
rect 22021 20587 22079 20593
rect 22021 20584 22033 20587
rect 21407 20556 22033 20584
rect 21407 20553 21419 20556
rect 21361 20547 21419 20553
rect 22021 20553 22033 20556
rect 22067 20553 22079 20587
rect 22021 20547 22079 20553
rect 22189 20587 22247 20593
rect 22189 20553 22201 20587
rect 22235 20584 22247 20587
rect 22554 20584 22560 20596
rect 22235 20556 22560 20584
rect 22235 20553 22247 20556
rect 22189 20547 22247 20553
rect 22554 20544 22560 20556
rect 22612 20544 22618 20596
rect 22646 20544 22652 20596
rect 22704 20544 22710 20596
rect 23106 20544 23112 20596
rect 23164 20544 23170 20596
rect 23477 20587 23535 20593
rect 23477 20553 23489 20587
rect 23523 20584 23535 20587
rect 24670 20584 24676 20596
rect 23523 20556 24676 20584
rect 23523 20553 23535 20556
rect 23477 20547 23535 20553
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 27062 20544 27068 20596
rect 27120 20544 27126 20596
rect 27540 20556 28764 20584
rect 17957 20519 18015 20525
rect 17957 20485 17969 20519
rect 18003 20516 18015 20519
rect 20993 20519 21051 20525
rect 18003 20488 19472 20516
rect 18003 20485 18015 20488
rect 17957 20479 18015 20485
rect 18046 20448 18052 20460
rect 17880 20420 18052 20448
rect 18046 20408 18052 20420
rect 18104 20448 18110 20460
rect 18141 20451 18199 20457
rect 18141 20448 18153 20451
rect 18104 20420 18153 20448
rect 18104 20408 18110 20420
rect 18141 20417 18153 20420
rect 18187 20417 18199 20451
rect 18141 20411 18199 20417
rect 18322 20408 18328 20460
rect 18380 20408 18386 20460
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 17604 20380 17632 20408
rect 15578 20352 17632 20380
rect 14642 20272 14648 20324
rect 14700 20312 14706 20324
rect 15578 20312 15606 20352
rect 18230 20340 18236 20392
rect 18288 20380 18294 20392
rect 18417 20383 18475 20389
rect 18417 20380 18429 20383
rect 18288 20352 18429 20380
rect 18288 20340 18294 20352
rect 18417 20349 18429 20352
rect 18463 20349 18475 20383
rect 18800 20380 18828 20411
rect 19058 20408 19064 20460
rect 19116 20448 19122 20460
rect 19444 20457 19472 20488
rect 20993 20485 21005 20519
rect 21039 20516 21051 20519
rect 21542 20516 21548 20528
rect 21039 20488 21548 20516
rect 21039 20485 21051 20488
rect 20993 20479 21051 20485
rect 21542 20476 21548 20488
rect 21600 20476 21606 20528
rect 21821 20519 21879 20525
rect 21821 20516 21833 20519
rect 21744 20488 21833 20516
rect 19153 20451 19211 20457
rect 19153 20448 19165 20451
rect 19116 20420 19165 20448
rect 19116 20408 19122 20420
rect 19153 20417 19165 20420
rect 19199 20417 19211 20451
rect 19153 20411 19211 20417
rect 19429 20451 19487 20457
rect 19429 20417 19441 20451
rect 19475 20417 19487 20451
rect 19429 20411 19487 20417
rect 20898 20408 20904 20460
rect 20956 20448 20962 20460
rect 21174 20448 21180 20460
rect 20956 20420 21180 20448
rect 20956 20408 20962 20420
rect 21174 20408 21180 20420
rect 21232 20408 21238 20460
rect 21453 20451 21511 20457
rect 21453 20417 21465 20451
rect 21499 20448 21511 20451
rect 21560 20448 21588 20476
rect 21499 20420 21588 20448
rect 21637 20451 21695 20457
rect 21499 20417 21511 20420
rect 21453 20411 21511 20417
rect 21637 20417 21649 20451
rect 21683 20417 21695 20451
rect 21637 20411 21695 20417
rect 21744 20448 21772 20488
rect 21821 20485 21833 20488
rect 21867 20485 21879 20519
rect 22664 20516 22692 20544
rect 22664 20488 24072 20516
rect 21821 20479 21879 20485
rect 21910 20448 21916 20460
rect 21744 20420 21916 20448
rect 20530 20380 20536 20392
rect 18800 20352 20536 20380
rect 18417 20343 18475 20349
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 21192 20380 21220 20408
rect 21652 20380 21680 20411
rect 21744 20392 21772 20420
rect 21910 20408 21916 20420
rect 21968 20448 21974 20460
rect 22738 20448 22744 20460
rect 21968 20420 22744 20448
rect 21968 20408 21974 20420
rect 22738 20408 22744 20420
rect 22796 20408 22802 20460
rect 22940 20457 22968 20488
rect 22925 20451 22983 20457
rect 22925 20417 22937 20451
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 23658 20408 23664 20460
rect 23716 20408 23722 20460
rect 23842 20408 23848 20460
rect 23900 20408 23906 20460
rect 23934 20408 23940 20460
rect 23992 20408 23998 20460
rect 24044 20457 24072 20488
rect 25866 20476 25872 20528
rect 25924 20516 25930 20528
rect 26786 20516 26792 20528
rect 25924 20488 26792 20516
rect 25924 20476 25930 20488
rect 24029 20451 24087 20457
rect 24029 20417 24041 20451
rect 24075 20417 24087 20451
rect 24029 20411 24087 20417
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 24210 20448 24216 20460
rect 24167 20420 24216 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 26620 20457 26648 20488
rect 26786 20476 26792 20488
rect 26844 20476 26850 20528
rect 27080 20457 27108 20544
rect 27540 20516 27568 20556
rect 28534 20516 28540 20528
rect 27356 20488 27568 20516
rect 27356 20460 27384 20488
rect 26605 20451 26663 20457
rect 26605 20417 26617 20451
rect 26651 20417 26663 20451
rect 26605 20411 26663 20417
rect 27065 20451 27123 20457
rect 27065 20417 27077 20451
rect 27111 20417 27123 20451
rect 27065 20411 27123 20417
rect 27338 20408 27344 20460
rect 27396 20408 27402 20460
rect 27430 20408 27436 20460
rect 27488 20408 27494 20460
rect 21192 20352 21680 20380
rect 21726 20340 21732 20392
rect 21784 20340 21790 20392
rect 22756 20380 22784 20408
rect 24305 20383 24363 20389
rect 24305 20380 24317 20383
rect 22756 20352 24317 20380
rect 24305 20349 24317 20352
rect 24351 20349 24363 20383
rect 24305 20343 24363 20349
rect 26697 20383 26755 20389
rect 26697 20349 26709 20383
rect 26743 20380 26755 20383
rect 27448 20380 27476 20408
rect 26743 20352 27476 20380
rect 27540 20380 27568 20488
rect 27908 20488 28540 20516
rect 27908 20457 27936 20488
rect 28534 20476 28540 20488
rect 28592 20476 28598 20528
rect 28540 20473 28598 20476
rect 27893 20451 27951 20457
rect 27893 20417 27905 20451
rect 27939 20417 27951 20451
rect 27893 20411 27951 20417
rect 27985 20451 28043 20457
rect 27985 20417 27997 20451
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 28000 20380 28028 20411
rect 28074 20408 28080 20460
rect 28132 20448 28138 20460
rect 28169 20451 28227 20457
rect 28169 20448 28181 20451
rect 28132 20420 28181 20448
rect 28132 20408 28138 20420
rect 28169 20417 28181 20420
rect 28215 20417 28227 20451
rect 28169 20411 28227 20417
rect 28261 20451 28319 20457
rect 28261 20417 28273 20451
rect 28307 20417 28319 20451
rect 28540 20439 28552 20473
rect 28586 20439 28598 20473
rect 28540 20433 28598 20439
rect 28629 20451 28687 20457
rect 28261 20411 28319 20417
rect 28629 20417 28641 20451
rect 28675 20448 28687 20451
rect 28736 20448 28764 20556
rect 28675 20420 28764 20448
rect 28813 20451 28871 20457
rect 28675 20417 28687 20420
rect 28629 20411 28687 20417
rect 28813 20417 28825 20451
rect 28859 20417 28871 20451
rect 28813 20411 28871 20417
rect 27540 20352 28028 20380
rect 28276 20380 28304 20411
rect 28828 20380 28856 20411
rect 28902 20408 28908 20460
rect 28960 20408 28966 20460
rect 28276 20352 28856 20380
rect 26743 20349 26755 20352
rect 26697 20343 26755 20349
rect 14700 20284 15606 20312
rect 16669 20315 16727 20321
rect 14700 20272 14706 20284
rect 16669 20281 16681 20315
rect 16715 20312 16727 20315
rect 17034 20312 17040 20324
rect 16715 20284 17040 20312
rect 16715 20281 16727 20284
rect 16669 20275 16727 20281
rect 17034 20272 17040 20284
rect 17092 20272 17098 20324
rect 18877 20315 18935 20321
rect 18877 20281 18889 20315
rect 18923 20312 18935 20315
rect 19150 20312 19156 20324
rect 18923 20284 19156 20312
rect 18923 20281 18935 20284
rect 18877 20275 18935 20281
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 23658 20272 23664 20324
rect 23716 20312 23722 20324
rect 24213 20315 24271 20321
rect 24213 20312 24225 20315
rect 23716 20284 24225 20312
rect 23716 20272 23722 20284
rect 24213 20281 24225 20284
rect 24259 20281 24271 20315
rect 24213 20275 24271 20281
rect 27246 20272 27252 20324
rect 27304 20312 27310 20324
rect 28276 20312 28304 20352
rect 27304 20284 28304 20312
rect 27304 20272 27310 20284
rect 12526 20244 12532 20256
rect 10612 20216 12532 20244
rect 10192 20204 10198 20216
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 14274 20204 14280 20256
rect 14332 20204 14338 20256
rect 17862 20204 17868 20256
rect 17920 20204 17926 20256
rect 21545 20247 21603 20253
rect 21545 20213 21557 20247
rect 21591 20244 21603 20247
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 21591 20216 22017 20244
rect 21591 20213 21603 20216
rect 21545 20207 21603 20213
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 22005 20207 22063 20213
rect 24118 20204 24124 20256
rect 24176 20244 24182 20256
rect 24486 20244 24492 20256
rect 24176 20216 24492 20244
rect 24176 20204 24182 20216
rect 24486 20204 24492 20216
rect 24544 20204 24550 20256
rect 27338 20204 27344 20256
rect 27396 20204 27402 20256
rect 27522 20204 27528 20256
rect 27580 20244 27586 20256
rect 27617 20247 27675 20253
rect 27617 20244 27629 20247
rect 27580 20216 27629 20244
rect 27580 20204 27586 20216
rect 27617 20213 27629 20216
rect 27663 20213 27675 20247
rect 27617 20207 27675 20213
rect 27706 20204 27712 20256
rect 27764 20204 27770 20256
rect 28350 20204 28356 20256
rect 28408 20204 28414 20256
rect 1104 20154 29440 20176
rect 1104 20102 4491 20154
rect 4543 20102 4555 20154
rect 4607 20102 4619 20154
rect 4671 20102 4683 20154
rect 4735 20102 4747 20154
rect 4799 20102 11574 20154
rect 11626 20102 11638 20154
rect 11690 20102 11702 20154
rect 11754 20102 11766 20154
rect 11818 20102 11830 20154
rect 11882 20102 18657 20154
rect 18709 20102 18721 20154
rect 18773 20102 18785 20154
rect 18837 20102 18849 20154
rect 18901 20102 18913 20154
rect 18965 20102 25740 20154
rect 25792 20102 25804 20154
rect 25856 20102 25868 20154
rect 25920 20102 25932 20154
rect 25984 20102 25996 20154
rect 26048 20102 29440 20154
rect 1104 20080 29440 20102
rect 3878 20000 3884 20052
rect 3936 20000 3942 20052
rect 3970 20000 3976 20052
rect 4028 20040 4034 20052
rect 4433 20043 4491 20049
rect 4433 20040 4445 20043
rect 4028 20012 4445 20040
rect 4028 20000 4034 20012
rect 4433 20009 4445 20012
rect 4479 20009 4491 20043
rect 4433 20003 4491 20009
rect 6638 20000 6644 20052
rect 6696 20040 6702 20052
rect 6917 20043 6975 20049
rect 6917 20040 6929 20043
rect 6696 20012 6929 20040
rect 6696 20000 6702 20012
rect 6917 20009 6929 20012
rect 6963 20009 6975 20043
rect 8202 20040 8208 20052
rect 6917 20003 6975 20009
rect 7024 20012 8208 20040
rect 2133 19907 2191 19913
rect 2133 19873 2145 19907
rect 2179 19904 2191 19907
rect 3896 19904 3924 20000
rect 7024 19904 7052 20012
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 8757 20043 8815 20049
rect 8757 20009 8769 20043
rect 8803 20040 8815 20043
rect 9674 20040 9680 20052
rect 8803 20012 9680 20040
rect 8803 20009 8815 20012
rect 8757 20003 8815 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 12621 20043 12679 20049
rect 12621 20040 12633 20043
rect 12124 20012 12633 20040
rect 12124 20000 12130 20012
rect 12621 20009 12633 20012
rect 12667 20009 12679 20043
rect 12621 20003 12679 20009
rect 14274 20000 14280 20052
rect 14332 20000 14338 20052
rect 16117 20043 16175 20049
rect 16117 20009 16129 20043
rect 16163 20040 16175 20043
rect 16850 20040 16856 20052
rect 16163 20012 16856 20040
rect 16163 20009 16175 20012
rect 16117 20003 16175 20009
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 16942 20000 16948 20052
rect 17000 20000 17006 20052
rect 17034 20000 17040 20052
rect 17092 20040 17098 20052
rect 21082 20040 21088 20052
rect 17092 20012 21088 20040
rect 17092 20000 17098 20012
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 27617 20043 27675 20049
rect 27617 20009 27629 20043
rect 27663 20040 27675 20043
rect 28074 20040 28080 20052
rect 27663 20012 28080 20040
rect 27663 20009 27675 20012
rect 27617 20003 27675 20009
rect 28074 20000 28080 20012
rect 28132 20000 28138 20052
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 7616 19944 10824 19972
rect 7616 19932 7622 19944
rect 9398 19904 9404 19916
rect 2179 19876 3924 19904
rect 6380 19876 7052 19904
rect 8128 19876 9404 19904
rect 2179 19873 2191 19876
rect 2133 19867 2191 19873
rect 1854 19796 1860 19848
rect 1912 19796 1918 19848
rect 6380 19845 6408 19876
rect 3881 19839 3939 19845
rect 3881 19805 3893 19839
rect 3927 19805 3939 19839
rect 3881 19799 3939 19805
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 3418 19768 3424 19780
rect 3358 19740 3424 19768
rect 3418 19728 3424 19740
rect 3476 19728 3482 19780
rect 3605 19703 3663 19709
rect 3605 19669 3617 19703
rect 3651 19700 3663 19703
rect 3896 19700 3924 19799
rect 6454 19796 6460 19848
rect 6512 19836 6518 19848
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 6512 19808 6653 19836
rect 6512 19796 6518 19808
rect 6641 19805 6653 19808
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 6822 19836 6828 19848
rect 6779 19808 6828 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 6914 19796 6920 19848
rect 6972 19836 6978 19848
rect 7190 19845 7196 19848
rect 7009 19839 7067 19845
rect 7009 19836 7021 19839
rect 6972 19808 7021 19836
rect 6972 19796 6978 19808
rect 7009 19805 7021 19808
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7157 19839 7196 19845
rect 7157 19805 7169 19839
rect 7157 19799 7196 19805
rect 7190 19796 7196 19799
rect 7248 19796 7254 19848
rect 7515 19839 7573 19845
rect 7515 19805 7527 19839
rect 7561 19836 7573 19839
rect 8128 19836 8156 19876
rect 9398 19864 9404 19876
rect 9456 19864 9462 19916
rect 10502 19864 10508 19916
rect 10560 19864 10566 19916
rect 10796 19904 10824 19944
rect 11330 19904 11336 19916
rect 10796 19876 11336 19904
rect 7561 19808 8156 19836
rect 8205 19839 8263 19845
rect 7561 19805 7573 19808
rect 7515 19799 7573 19805
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 8846 19836 8852 19848
rect 8251 19808 8852 19836
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 8846 19796 8852 19808
rect 8904 19796 8910 19848
rect 8938 19796 8944 19848
rect 8996 19796 9002 19848
rect 10226 19796 10232 19848
rect 10284 19796 10290 19848
rect 10796 19845 10824 19876
rect 11330 19864 11336 19876
rect 11388 19864 11394 19916
rect 14292 19904 14320 20000
rect 16960 19972 16988 20000
rect 17862 19972 17868 19984
rect 16960 19944 17868 19972
rect 17862 19932 17868 19944
rect 17920 19932 17926 19984
rect 27264 19944 28028 19972
rect 18230 19904 18236 19916
rect 12084 19876 14320 19904
rect 15948 19876 18236 19904
rect 12084 19845 12112 19876
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 10965 19839 11023 19845
rect 10965 19805 10977 19839
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19805 12127 19839
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 12069 19799 12127 19805
rect 12176 19808 12449 19836
rect 6546 19728 6552 19780
rect 6604 19728 6610 19780
rect 7282 19728 7288 19780
rect 7340 19728 7346 19780
rect 7377 19771 7435 19777
rect 7377 19737 7389 19771
rect 7423 19737 7435 19771
rect 10318 19768 10324 19780
rect 7377 19731 7435 19737
rect 7668 19740 10324 19768
rect 7392 19700 7420 19731
rect 7668 19709 7696 19740
rect 10318 19728 10324 19740
rect 10376 19728 10382 19780
rect 3651 19672 7420 19700
rect 7653 19703 7711 19709
rect 3651 19669 3663 19672
rect 3605 19663 3663 19669
rect 7653 19669 7665 19703
rect 7699 19669 7711 19703
rect 7653 19663 7711 19669
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 10612 19700 10640 19799
rect 10870 19728 10876 19780
rect 10928 19728 10934 19780
rect 10980 19768 11008 19799
rect 12176 19768 12204 19808
rect 12437 19805 12449 19808
rect 12483 19836 12495 19839
rect 12710 19836 12716 19848
rect 12483 19808 12716 19836
rect 12483 19805 12495 19808
rect 12437 19799 12495 19805
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 12986 19796 12992 19848
rect 13044 19796 13050 19848
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 14734 19836 14740 19848
rect 13228 19808 14740 19836
rect 13228 19796 13234 19808
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 15102 19796 15108 19848
rect 15160 19836 15166 19848
rect 15948 19845 15976 19876
rect 18230 19864 18236 19876
rect 18288 19864 18294 19916
rect 27264 19848 27292 19944
rect 28000 19904 28028 19944
rect 27356 19876 27660 19904
rect 28000 19876 28120 19904
rect 27356 19848 27384 19876
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15160 19808 15945 19836
rect 15160 19796 15166 19808
rect 15933 19805 15945 19808
rect 15979 19805 15991 19839
rect 15933 19799 15991 19805
rect 16850 19796 16856 19848
rect 16908 19836 16914 19848
rect 19702 19836 19708 19848
rect 16908 19808 19708 19836
rect 16908 19796 16914 19808
rect 19702 19796 19708 19808
rect 19760 19836 19766 19848
rect 20162 19836 20168 19848
rect 19760 19808 20168 19836
rect 19760 19796 19766 19808
rect 20162 19796 20168 19808
rect 20220 19796 20226 19848
rect 27246 19796 27252 19848
rect 27304 19796 27310 19848
rect 27338 19796 27344 19848
rect 27396 19796 27402 19848
rect 27522 19846 27528 19848
rect 27448 19818 27528 19846
rect 10980 19740 12204 19768
rect 12253 19771 12311 19777
rect 12253 19737 12265 19771
rect 12299 19737 12311 19771
rect 12253 19731 12311 19737
rect 12345 19771 12403 19777
rect 12345 19737 12357 19771
rect 12391 19768 12403 19771
rect 12526 19768 12532 19780
rect 12391 19740 12532 19768
rect 12391 19737 12403 19740
rect 12345 19731 12403 19737
rect 11054 19700 11060 19712
rect 10612 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11146 19660 11152 19712
rect 11204 19660 11210 19712
rect 11330 19660 11336 19712
rect 11388 19700 11394 19712
rect 12268 19700 12296 19731
rect 12526 19728 12532 19740
rect 12584 19768 12590 19780
rect 14642 19768 14648 19780
rect 12584 19740 14648 19768
rect 12584 19728 12590 19740
rect 14642 19728 14648 19740
rect 14700 19728 14706 19780
rect 15749 19771 15807 19777
rect 15749 19737 15761 19771
rect 15795 19768 15807 19771
rect 15838 19768 15844 19780
rect 15795 19740 15844 19768
rect 15795 19737 15807 19740
rect 15749 19731 15807 19737
rect 15838 19728 15844 19740
rect 15896 19728 15902 19780
rect 17586 19728 17592 19780
rect 17644 19768 17650 19780
rect 19242 19768 19248 19780
rect 17644 19740 19248 19768
rect 17644 19728 17650 19740
rect 19242 19728 19248 19740
rect 19300 19728 19306 19780
rect 25038 19768 25044 19780
rect 19904 19740 25044 19768
rect 19904 19712 19932 19740
rect 25038 19728 25044 19740
rect 25096 19728 25102 19780
rect 27448 19768 27476 19818
rect 27522 19796 27528 19818
rect 27580 19796 27586 19848
rect 27632 19845 27660 19876
rect 27617 19839 27675 19845
rect 27617 19805 27629 19839
rect 27663 19805 27675 19839
rect 27617 19799 27675 19805
rect 27801 19839 27859 19845
rect 27801 19805 27813 19839
rect 27847 19836 27859 19839
rect 27982 19836 27988 19848
rect 27847 19808 27988 19836
rect 27847 19805 27859 19808
rect 27801 19799 27859 19805
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 28092 19845 28120 19876
rect 28077 19839 28135 19845
rect 28077 19805 28089 19839
rect 28123 19805 28135 19839
rect 28077 19799 28135 19805
rect 28166 19796 28172 19848
rect 28224 19836 28230 19848
rect 28353 19839 28411 19845
rect 28353 19836 28365 19839
rect 28224 19808 28365 19836
rect 28224 19796 28230 19808
rect 28353 19805 28365 19808
rect 28399 19805 28411 19839
rect 28353 19799 28411 19805
rect 28261 19771 28319 19777
rect 28261 19768 28273 19771
rect 27448 19740 28273 19768
rect 28261 19737 28273 19740
rect 28307 19737 28319 19771
rect 28261 19731 28319 19737
rect 12618 19700 12624 19712
rect 11388 19672 12624 19700
rect 11388 19660 11394 19672
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 13541 19703 13599 19709
rect 13541 19700 13553 19703
rect 12952 19672 13553 19700
rect 12952 19660 12958 19672
rect 13541 19669 13553 19672
rect 13587 19669 13599 19703
rect 13541 19663 13599 19669
rect 19886 19660 19892 19712
rect 19944 19660 19950 19712
rect 19978 19660 19984 19712
rect 20036 19700 20042 19712
rect 26326 19700 26332 19712
rect 20036 19672 26332 19700
rect 20036 19660 20042 19672
rect 26326 19660 26332 19672
rect 26384 19660 26390 19712
rect 27062 19660 27068 19712
rect 27120 19660 27126 19712
rect 27433 19703 27491 19709
rect 27433 19669 27445 19703
rect 27479 19700 27491 19703
rect 27614 19700 27620 19712
rect 27479 19672 27620 19700
rect 27479 19669 27491 19672
rect 27433 19663 27491 19669
rect 27614 19660 27620 19672
rect 27672 19660 27678 19712
rect 27893 19703 27951 19709
rect 27893 19669 27905 19703
rect 27939 19700 27951 19703
rect 28718 19700 28724 19712
rect 27939 19672 28724 19700
rect 27939 19669 27951 19672
rect 27893 19663 27951 19669
rect 28718 19660 28724 19672
rect 28776 19660 28782 19712
rect 1104 19610 29440 19632
rect 1104 19558 5151 19610
rect 5203 19558 5215 19610
rect 5267 19558 5279 19610
rect 5331 19558 5343 19610
rect 5395 19558 5407 19610
rect 5459 19558 12234 19610
rect 12286 19558 12298 19610
rect 12350 19558 12362 19610
rect 12414 19558 12426 19610
rect 12478 19558 12490 19610
rect 12542 19558 19317 19610
rect 19369 19558 19381 19610
rect 19433 19558 19445 19610
rect 19497 19558 19509 19610
rect 19561 19558 19573 19610
rect 19625 19558 26400 19610
rect 26452 19558 26464 19610
rect 26516 19558 26528 19610
rect 26580 19558 26592 19610
rect 26644 19558 26656 19610
rect 26708 19558 29440 19610
rect 1104 19536 29440 19558
rect 1578 19456 1584 19508
rect 1636 19456 1642 19508
rect 9582 19496 9588 19508
rect 7300 19468 9588 19496
rect 1486 19320 1492 19372
rect 1544 19320 1550 19372
rect 7300 19369 7328 19468
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 11054 19456 11060 19508
rect 11112 19496 11118 19508
rect 12161 19499 12219 19505
rect 12161 19496 12173 19499
rect 11112 19468 12173 19496
rect 11112 19456 11118 19468
rect 12161 19465 12173 19468
rect 12207 19465 12219 19499
rect 13078 19496 13084 19508
rect 12161 19459 12219 19465
rect 12728 19468 13084 19496
rect 7561 19431 7619 19437
rect 7561 19397 7573 19431
rect 7607 19428 7619 19431
rect 8110 19428 8116 19440
rect 7607 19400 8116 19428
rect 7607 19397 7619 19400
rect 7561 19391 7619 19397
rect 8110 19388 8116 19400
rect 8168 19388 8174 19440
rect 8205 19431 8263 19437
rect 8205 19397 8217 19431
rect 8251 19428 8263 19431
rect 8478 19428 8484 19440
rect 8251 19400 8484 19428
rect 8251 19397 8263 19400
rect 8205 19391 8263 19397
rect 8478 19388 8484 19400
rect 8536 19388 8542 19440
rect 9766 19428 9772 19440
rect 9430 19400 9772 19428
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 10870 19388 10876 19440
rect 10928 19428 10934 19440
rect 12728 19428 12756 19468
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13357 19499 13415 19505
rect 13357 19496 13369 19499
rect 13320 19468 13369 19496
rect 13320 19456 13326 19468
rect 13357 19465 13369 19468
rect 13403 19465 13415 19499
rect 13357 19459 13415 19465
rect 14550 19456 14556 19508
rect 14608 19456 14614 19508
rect 14918 19456 14924 19508
rect 14976 19496 14982 19508
rect 14976 19468 15240 19496
rect 14976 19456 14982 19468
rect 10928 19400 12756 19428
rect 10928 19388 10934 19400
rect 7285 19363 7343 19369
rect 7285 19329 7297 19363
rect 7331 19329 7343 19363
rect 7285 19323 7343 19329
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 6546 19252 6552 19304
rect 6604 19292 6610 19304
rect 7484 19292 7512 19323
rect 7650 19320 7656 19372
rect 7708 19320 7714 19372
rect 7926 19320 7932 19372
rect 7984 19320 7990 19372
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 12805 19363 12863 19369
rect 9916 19332 12756 19360
rect 9916 19320 9922 19332
rect 7558 19292 7564 19304
rect 6604 19264 7564 19292
rect 6604 19252 6610 19264
rect 7558 19252 7564 19264
rect 7616 19252 7622 19304
rect 8846 19252 8852 19304
rect 8904 19292 8910 19304
rect 9214 19292 9220 19304
rect 8904 19264 9220 19292
rect 8904 19252 8910 19264
rect 9214 19252 9220 19264
rect 9272 19292 9278 19304
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9272 19264 9689 19292
rect 9272 19252 9278 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 9677 19255 9735 19261
rect 11609 19295 11667 19301
rect 11609 19261 11621 19295
rect 11655 19292 11667 19295
rect 12158 19292 12164 19304
rect 11655 19264 12164 19292
rect 11655 19261 11667 19264
rect 11609 19255 11667 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12728 19292 12756 19332
rect 12805 19329 12817 19363
rect 12851 19360 12863 19363
rect 12894 19360 12900 19372
rect 12851 19332 12900 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 13096 19369 13124 19456
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 13004 19292 13032 19323
rect 13170 19320 13176 19372
rect 13228 19320 13234 19372
rect 14568 19360 14596 19456
rect 15102 19388 15108 19440
rect 15160 19388 15166 19440
rect 15212 19437 15240 19468
rect 15470 19456 15476 19508
rect 15528 19496 15534 19508
rect 15528 19468 16712 19496
rect 15528 19456 15534 19468
rect 15197 19431 15255 19437
rect 15197 19397 15209 19431
rect 15243 19397 15255 19431
rect 15197 19391 15255 19397
rect 15304 19400 15606 19428
rect 15304 19369 15332 19400
rect 13280 19332 14596 19360
rect 14921 19363 14979 19369
rect 13280 19292 13308 19332
rect 14921 19329 14933 19363
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15289 19363 15347 19369
rect 15289 19329 15301 19363
rect 15335 19329 15347 19363
rect 15578 19360 15606 19400
rect 16022 19360 16028 19372
rect 15578 19332 16028 19360
rect 15289 19323 15347 19329
rect 12728 19264 13308 19292
rect 4982 19184 4988 19236
rect 5040 19224 5046 19236
rect 6454 19224 6460 19236
rect 5040 19196 6460 19224
rect 5040 19184 5046 19196
rect 6454 19184 6460 19196
rect 6512 19224 6518 19236
rect 6512 19196 7972 19224
rect 6512 19184 6518 19196
rect 7834 19116 7840 19168
rect 7892 19116 7898 19168
rect 7944 19156 7972 19196
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 13814 19224 13820 19236
rect 9640 19196 13820 19224
rect 9640 19184 9646 19196
rect 13814 19184 13820 19196
rect 13872 19184 13878 19236
rect 14936 19224 14964 19323
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 16684 19369 16712 19468
rect 16850 19456 16856 19508
rect 16908 19456 16914 19508
rect 17218 19456 17224 19508
rect 17276 19456 17282 19508
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 18012 19468 18981 19496
rect 18012 19456 18018 19468
rect 18969 19465 18981 19468
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 19058 19456 19064 19508
rect 19116 19456 19122 19508
rect 19978 19496 19984 19508
rect 19168 19468 19984 19496
rect 16868 19369 16896 19456
rect 16945 19431 17003 19437
rect 16945 19397 16957 19431
rect 16991 19428 17003 19431
rect 19168 19428 19196 19468
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20530 19456 20536 19508
rect 20588 19456 20594 19508
rect 28074 19456 28080 19508
rect 28132 19456 28138 19508
rect 16991 19400 19196 19428
rect 19245 19431 19303 19437
rect 16991 19397 17003 19400
rect 16945 19391 17003 19397
rect 19245 19397 19257 19431
rect 19291 19428 19303 19431
rect 19426 19428 19432 19440
rect 19291 19400 19432 19428
rect 19291 19397 19303 19400
rect 19245 19391 19303 19397
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 19518 19388 19524 19440
rect 19576 19388 19582 19440
rect 19613 19431 19671 19437
rect 19613 19397 19625 19431
rect 19659 19428 19671 19431
rect 19886 19428 19892 19440
rect 19659 19400 19892 19428
rect 19659 19397 19671 19400
rect 19613 19391 19671 19397
rect 19886 19388 19892 19400
rect 19944 19388 19950 19440
rect 20070 19428 20076 19440
rect 19996 19400 20076 19428
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19360 17095 19363
rect 17083 19332 17954 19360
rect 17083 19329 17095 19332
rect 17037 19323 17095 19329
rect 15838 19252 15844 19304
rect 15896 19252 15902 19304
rect 17926 19292 17954 19332
rect 18874 19320 18880 19372
rect 18932 19320 18938 19372
rect 19334 19320 19340 19372
rect 19392 19320 19398 19372
rect 19996 19369 20024 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 20162 19388 20168 19440
rect 20220 19388 20226 19440
rect 20257 19431 20315 19437
rect 20257 19397 20269 19431
rect 20303 19428 20315 19431
rect 22646 19428 22652 19440
rect 20303 19400 22652 19428
rect 20303 19397 20315 19400
rect 20257 19391 20315 19397
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 28092 19428 28120 19456
rect 27540 19400 28120 19428
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19360 19763 19363
rect 19981 19363 20039 19369
rect 19751 19332 19932 19360
rect 19751 19329 19763 19332
rect 19705 19323 19763 19329
rect 17926 19264 19472 19292
rect 16393 19227 16451 19233
rect 16393 19224 16405 19227
rect 14936 19196 16405 19224
rect 16393 19193 16405 19196
rect 16439 19193 16451 19227
rect 16393 19187 16451 19193
rect 18693 19227 18751 19233
rect 18693 19193 18705 19227
rect 18739 19193 18751 19227
rect 19444 19224 19472 19264
rect 19610 19224 19616 19236
rect 19444 19196 19616 19224
rect 18693 19187 18751 19193
rect 14182 19156 14188 19168
rect 7944 19128 14188 19156
rect 14182 19116 14188 19128
rect 14240 19156 14246 19168
rect 15378 19156 15384 19168
rect 14240 19128 15384 19156
rect 14240 19116 14246 19128
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 15470 19116 15476 19168
rect 15528 19116 15534 19168
rect 18708 19156 18736 19187
rect 19610 19184 19616 19196
rect 19668 19224 19674 19236
rect 19720 19224 19748 19323
rect 19904 19292 19932 19332
rect 19981 19329 19993 19363
rect 20027 19329 20039 19363
rect 19981 19323 20039 19329
rect 20349 19363 20407 19369
rect 20349 19329 20361 19363
rect 20395 19329 20407 19363
rect 20349 19323 20407 19329
rect 20364 19292 20392 19323
rect 27430 19320 27436 19372
rect 27488 19320 27494 19372
rect 27540 19369 27568 19400
rect 27525 19363 27583 19369
rect 27525 19329 27537 19363
rect 27571 19329 27583 19363
rect 27525 19323 27583 19329
rect 27617 19363 27675 19369
rect 27617 19329 27629 19363
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 20806 19292 20812 19304
rect 19904 19264 20812 19292
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 27448 19292 27476 19320
rect 27632 19292 27660 19323
rect 27448 19264 27660 19292
rect 27798 19252 27804 19304
rect 27856 19252 27862 19304
rect 19668 19196 19748 19224
rect 19889 19227 19947 19233
rect 19668 19184 19674 19196
rect 19889 19193 19901 19227
rect 19935 19224 19947 19227
rect 20346 19224 20352 19236
rect 19935 19196 20352 19224
rect 19935 19193 19947 19196
rect 19889 19187 19947 19193
rect 20346 19184 20352 19196
rect 20404 19184 20410 19236
rect 19334 19156 19340 19168
rect 18708 19128 19340 19156
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 1104 19066 29440 19088
rect 1104 19014 4491 19066
rect 4543 19014 4555 19066
rect 4607 19014 4619 19066
rect 4671 19014 4683 19066
rect 4735 19014 4747 19066
rect 4799 19014 11574 19066
rect 11626 19014 11638 19066
rect 11690 19014 11702 19066
rect 11754 19014 11766 19066
rect 11818 19014 11830 19066
rect 11882 19014 18657 19066
rect 18709 19014 18721 19066
rect 18773 19014 18785 19066
rect 18837 19014 18849 19066
rect 18901 19014 18913 19066
rect 18965 19014 25740 19066
rect 25792 19014 25804 19066
rect 25856 19014 25868 19066
rect 25920 19014 25932 19066
rect 25984 19014 25996 19066
rect 26048 19014 29440 19066
rect 1104 18992 29440 19014
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 8757 18955 8815 18961
rect 7064 18924 8340 18952
rect 7064 18912 7070 18924
rect 6546 18884 6552 18896
rect 6288 18856 6552 18884
rect 3602 18708 3608 18760
rect 3660 18748 3666 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3660 18720 4077 18748
rect 3660 18708 3666 18720
rect 4065 18717 4077 18720
rect 4111 18748 4123 18751
rect 6181 18751 6239 18757
rect 4111 18720 5580 18748
rect 4111 18717 4123 18720
rect 4065 18711 4123 18717
rect 5552 18624 5580 18720
rect 6181 18717 6193 18751
rect 6227 18717 6239 18751
rect 6288 18748 6316 18856
rect 6546 18844 6552 18856
rect 6604 18844 6610 18896
rect 8312 18884 8340 18924
rect 8757 18921 8769 18955
rect 8803 18952 8815 18955
rect 8938 18952 8944 18964
rect 8803 18924 8944 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 9582 18912 9588 18964
rect 9640 18912 9646 18964
rect 11885 18955 11943 18961
rect 11885 18921 11897 18955
rect 11931 18952 11943 18955
rect 12158 18952 12164 18964
rect 11931 18924 12164 18952
rect 11931 18921 11943 18924
rect 11885 18915 11943 18921
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 15470 18912 15476 18964
rect 15528 18912 15534 18964
rect 15838 18912 15844 18964
rect 15896 18952 15902 18964
rect 15933 18955 15991 18961
rect 15933 18952 15945 18955
rect 15896 18924 15945 18952
rect 15896 18912 15902 18924
rect 15933 18921 15945 18924
rect 15979 18921 15991 18955
rect 15933 18915 15991 18921
rect 16022 18912 16028 18964
rect 16080 18952 16086 18964
rect 17770 18952 17776 18964
rect 16080 18924 17776 18952
rect 16080 18912 16086 18924
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19484 18924 19809 18952
rect 19484 18912 19490 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 20254 18912 20260 18964
rect 20312 18912 20318 18964
rect 21266 18912 21272 18964
rect 21324 18912 21330 18964
rect 12802 18884 12808 18896
rect 8312 18856 9628 18884
rect 6362 18776 6368 18828
rect 6420 18816 6426 18828
rect 7009 18819 7067 18825
rect 7009 18816 7021 18819
rect 6420 18788 7021 18816
rect 6420 18776 6426 18788
rect 7009 18785 7021 18788
rect 7055 18785 7067 18819
rect 7009 18779 7067 18785
rect 7285 18819 7343 18825
rect 7285 18785 7297 18819
rect 7331 18816 7343 18819
rect 7834 18816 7840 18828
rect 7331 18788 7840 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 9214 18776 9220 18828
rect 9272 18776 9278 18828
rect 6288 18720 6408 18748
rect 6181 18711 6239 18717
rect 6196 18680 6224 18711
rect 6270 18680 6276 18692
rect 6196 18652 6276 18680
rect 6270 18640 6276 18652
rect 6328 18640 6334 18692
rect 6380 18689 6408 18720
rect 6454 18708 6460 18760
rect 6512 18708 6518 18760
rect 6549 18751 6607 18757
rect 6549 18717 6561 18751
rect 6595 18748 6607 18751
rect 6914 18748 6920 18760
rect 6595 18720 6920 18748
rect 6595 18717 6607 18720
rect 6549 18711 6607 18717
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8628 18720 8953 18748
rect 8628 18708 8634 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9030 18708 9036 18760
rect 9088 18748 9094 18760
rect 9232 18748 9260 18776
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 9088 18720 9133 18748
rect 9232 18720 9321 18748
rect 9088 18708 9094 18720
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9398 18708 9404 18760
rect 9456 18757 9462 18760
rect 9456 18748 9464 18757
rect 9456 18720 9501 18748
rect 9456 18711 9464 18720
rect 9456 18708 9462 18711
rect 6365 18683 6423 18689
rect 6365 18649 6377 18683
rect 6411 18649 6423 18683
rect 6365 18643 6423 18649
rect 7374 18640 7380 18692
rect 7432 18680 7438 18692
rect 9217 18683 9275 18689
rect 7432 18652 7774 18680
rect 7432 18640 7438 18652
rect 9217 18649 9229 18683
rect 9263 18649 9275 18683
rect 9217 18643 9275 18649
rect 3970 18572 3976 18624
rect 4028 18612 4034 18624
rect 4709 18615 4767 18621
rect 4709 18612 4721 18615
rect 4028 18584 4721 18612
rect 4028 18572 4034 18584
rect 4709 18581 4721 18584
rect 4755 18581 4767 18615
rect 4709 18575 4767 18581
rect 5534 18572 5540 18624
rect 5592 18572 5598 18624
rect 5810 18572 5816 18624
rect 5868 18612 5874 18624
rect 6733 18615 6791 18621
rect 6733 18612 6745 18615
rect 5868 18584 6745 18612
rect 5868 18572 5874 18584
rect 6733 18581 6745 18584
rect 6779 18581 6791 18615
rect 6733 18575 6791 18581
rect 7282 18572 7288 18624
rect 7340 18612 7346 18624
rect 8202 18612 8208 18624
rect 7340 18584 8208 18612
rect 7340 18572 7346 18584
rect 8202 18572 8208 18584
rect 8260 18612 8266 18624
rect 9232 18612 9260 18643
rect 8260 18584 9260 18612
rect 9600 18612 9628 18856
rect 11532 18856 12808 18884
rect 9950 18776 9956 18828
rect 10008 18816 10014 18828
rect 10137 18819 10195 18825
rect 10137 18816 10149 18819
rect 10008 18788 10149 18816
rect 10008 18776 10014 18788
rect 10137 18785 10149 18788
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 10413 18819 10471 18825
rect 10413 18785 10425 18819
rect 10459 18816 10471 18819
rect 11146 18816 11152 18828
rect 10459 18788 11152 18816
rect 10459 18785 10471 18788
rect 10413 18779 10471 18785
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 11532 18734 11560 18856
rect 12802 18844 12808 18856
rect 12860 18884 12866 18896
rect 13078 18884 13084 18896
rect 12860 18856 13084 18884
rect 12860 18844 12866 18856
rect 13078 18844 13084 18856
rect 13136 18844 13142 18896
rect 11606 18776 11612 18828
rect 11664 18816 11670 18828
rect 11664 18788 12388 18816
rect 11664 18776 11670 18788
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18717 12311 18751
rect 12253 18711 12311 18717
rect 10410 18640 10416 18692
rect 10468 18680 10474 18692
rect 10686 18680 10692 18692
rect 10468 18652 10692 18680
rect 10468 18640 10474 18652
rect 10686 18640 10692 18652
rect 10744 18640 10750 18692
rect 11146 18612 11152 18624
rect 9600 18584 11152 18612
rect 8260 18572 8266 18584
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 12268 18612 12296 18711
rect 12360 18680 12388 18788
rect 12526 18776 12532 18828
rect 12584 18776 12590 18828
rect 12894 18776 12900 18828
rect 12952 18816 12958 18828
rect 13722 18816 13728 18828
rect 12952 18788 13728 18816
rect 12952 18776 12958 18788
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 14461 18819 14519 18825
rect 14461 18785 14473 18819
rect 14507 18816 14519 18819
rect 15488 18816 15516 18912
rect 15562 18844 15568 18896
rect 15620 18884 15626 18896
rect 18414 18884 18420 18896
rect 15620 18856 18420 18884
rect 15620 18844 15626 18856
rect 18414 18844 18420 18856
rect 18472 18844 18478 18896
rect 19334 18844 19340 18896
rect 19392 18884 19398 18896
rect 21284 18884 21312 18912
rect 19392 18856 21312 18884
rect 19392 18844 19398 18856
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 14507 18788 15516 18816
rect 15764 18788 16620 18816
rect 14507 18785 14519 18788
rect 14461 18779 14519 18785
rect 12437 18751 12495 18757
rect 12437 18717 12449 18751
rect 12483 18748 12495 18751
rect 12544 18748 12572 18776
rect 12483 18720 12572 18748
rect 12621 18751 12679 18757
rect 12483 18717 12495 18720
rect 12437 18711 12495 18717
rect 12621 18717 12633 18751
rect 12667 18748 12679 18751
rect 12710 18748 12716 18760
rect 12667 18720 12716 18748
rect 12667 18717 12679 18720
rect 12621 18711 12679 18717
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 14185 18751 14243 18757
rect 14185 18717 14197 18751
rect 14231 18717 14243 18751
rect 14185 18711 14243 18717
rect 12529 18683 12587 18689
rect 12529 18680 12541 18683
rect 12360 18652 12541 18680
rect 12529 18649 12541 18652
rect 12575 18680 12587 18683
rect 14090 18680 14096 18692
rect 12575 18652 14096 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 14090 18640 14096 18652
rect 14148 18640 14154 18692
rect 14200 18680 14228 18711
rect 14366 18680 14372 18692
rect 14200 18652 14372 18680
rect 14366 18640 14372 18652
rect 14424 18640 14430 18692
rect 15470 18640 15476 18692
rect 15528 18640 15534 18692
rect 12710 18612 12716 18624
rect 12268 18584 12716 18612
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 12802 18572 12808 18624
rect 12860 18572 12866 18624
rect 14642 18572 14648 18624
rect 14700 18612 14706 18624
rect 15764 18612 15792 18788
rect 16022 18708 16028 18760
rect 16080 18708 16086 18760
rect 16390 18708 16396 18760
rect 16448 18708 16454 18760
rect 16592 18757 16620 18788
rect 17420 18788 19073 18816
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 17310 18748 17316 18760
rect 16623 18720 17316 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 17310 18708 17316 18720
rect 17368 18708 17374 18760
rect 17420 18757 17448 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 19168 18788 19932 18816
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17681 18751 17739 18757
rect 17681 18748 17693 18751
rect 17405 18711 17463 18717
rect 17512 18720 17693 18748
rect 16408 18680 16436 18708
rect 17512 18680 17540 18720
rect 17681 18717 17693 18720
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 16408 18652 17540 18680
rect 17589 18683 17647 18689
rect 17589 18649 17601 18683
rect 17635 18649 17647 18683
rect 17696 18680 17724 18711
rect 17770 18708 17776 18760
rect 17828 18708 17834 18760
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 18782 18748 18788 18760
rect 18555 18720 18788 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18782 18708 18788 18720
rect 18840 18748 18846 18760
rect 19168 18748 19196 18788
rect 18840 18720 19196 18748
rect 19245 18751 19303 18757
rect 18840 18708 18846 18720
rect 19245 18717 19257 18751
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19260 18680 19288 18711
rect 19426 18708 19432 18760
rect 19484 18708 19490 18760
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 19904 18757 19932 18788
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18717 19947 18751
rect 23290 18748 23296 18760
rect 19889 18711 19947 18717
rect 20001 18720 23296 18748
rect 17696 18652 19288 18680
rect 17589 18643 17647 18649
rect 14700 18584 15792 18612
rect 14700 18572 14706 18584
rect 15838 18572 15844 18624
rect 15896 18612 15902 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 15896 18584 16129 18612
rect 15896 18572 15902 18584
rect 16117 18581 16129 18584
rect 16163 18612 16175 18615
rect 17494 18612 17500 18624
rect 16163 18584 17500 18612
rect 16163 18581 16175 18584
rect 16117 18575 16175 18581
rect 17494 18572 17500 18584
rect 17552 18612 17558 18624
rect 17604 18612 17632 18643
rect 17552 18584 17632 18612
rect 17552 18572 17558 18584
rect 17954 18572 17960 18624
rect 18012 18572 18018 18624
rect 19444 18612 19472 18708
rect 19521 18683 19579 18689
rect 19521 18649 19533 18683
rect 19567 18680 19579 18683
rect 20001 18680 20029 18720
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 27706 18708 27712 18760
rect 27764 18748 27770 18760
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 27764 18720 28825 18748
rect 27764 18708 27770 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 19567 18652 20029 18680
rect 19567 18649 19579 18652
rect 19521 18643 19579 18649
rect 20070 18640 20076 18692
rect 20128 18640 20134 18692
rect 19886 18612 19892 18624
rect 19444 18584 19892 18612
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 28994 18572 29000 18624
rect 29052 18572 29058 18624
rect 1104 18522 29440 18544
rect 1104 18470 5151 18522
rect 5203 18470 5215 18522
rect 5267 18470 5279 18522
rect 5331 18470 5343 18522
rect 5395 18470 5407 18522
rect 5459 18470 12234 18522
rect 12286 18470 12298 18522
rect 12350 18470 12362 18522
rect 12414 18470 12426 18522
rect 12478 18470 12490 18522
rect 12542 18470 19317 18522
rect 19369 18470 19381 18522
rect 19433 18470 19445 18522
rect 19497 18470 19509 18522
rect 19561 18470 19573 18522
rect 19625 18470 26400 18522
rect 26452 18470 26464 18522
rect 26516 18470 26528 18522
rect 26580 18470 26592 18522
rect 26644 18470 26656 18522
rect 26708 18470 29440 18522
rect 1104 18448 29440 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 3694 18408 3700 18420
rect 1912 18380 3700 18408
rect 1912 18368 1918 18380
rect 3694 18368 3700 18380
rect 3752 18368 3758 18420
rect 4356 18380 6040 18408
rect 1872 18281 1900 18368
rect 3418 18340 3424 18352
rect 3358 18312 3424 18340
rect 3418 18300 3424 18312
rect 3476 18340 3482 18352
rect 4356 18340 4384 18380
rect 5276 18340 5304 18380
rect 3476 18312 4384 18340
rect 5198 18312 5304 18340
rect 3476 18300 3482 18312
rect 5534 18300 5540 18352
rect 5592 18340 5598 18352
rect 5905 18343 5963 18349
rect 5905 18340 5917 18343
rect 5592 18312 5917 18340
rect 5592 18300 5598 18312
rect 5905 18309 5917 18312
rect 5951 18309 5963 18343
rect 6012 18340 6040 18380
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 6328 18380 8217 18408
rect 6328 18368 6334 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 8205 18371 8263 18377
rect 9858 18368 9864 18420
rect 9916 18408 9922 18420
rect 11333 18411 11391 18417
rect 11333 18408 11345 18411
rect 9916 18380 11345 18408
rect 9916 18368 9922 18380
rect 11333 18377 11345 18380
rect 11379 18377 11391 18411
rect 11333 18371 11391 18377
rect 12066 18368 12072 18420
rect 12124 18408 12130 18420
rect 12618 18408 12624 18420
rect 12124 18380 12624 18408
rect 12124 18368 12130 18380
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 14001 18411 14059 18417
rect 14001 18408 14013 18411
rect 12768 18380 14013 18408
rect 12768 18368 12774 18380
rect 14001 18377 14013 18380
rect 14047 18377 14059 18411
rect 14001 18371 14059 18377
rect 14366 18368 14372 18420
rect 14424 18408 14430 18420
rect 16574 18408 16580 18420
rect 14424 18380 16580 18408
rect 14424 18368 14430 18380
rect 7374 18340 7380 18352
rect 6012 18312 7380 18340
rect 5905 18303 5963 18309
rect 7374 18300 7380 18312
rect 7432 18300 7438 18352
rect 12161 18343 12219 18349
rect 12161 18340 12173 18343
rect 9416 18312 9996 18340
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 3602 18232 3608 18284
rect 3660 18232 3666 18284
rect 3694 18232 3700 18284
rect 3752 18232 3758 18284
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5460 18244 5641 18272
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18204 2191 18207
rect 3418 18204 3424 18216
rect 2179 18176 3424 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 3620 18077 3648 18232
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18204 4031 18207
rect 4019 18176 5120 18204
rect 4019 18173 4031 18176
rect 3973 18167 4031 18173
rect 5092 18148 5120 18176
rect 5074 18096 5080 18148
rect 5132 18096 5138 18148
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18037 3663 18071
rect 3605 18031 3663 18037
rect 5166 18028 5172 18080
rect 5224 18068 5230 18080
rect 5460 18077 5488 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18241 5871 18275
rect 5813 18235 5871 18241
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6546 18272 6552 18284
rect 6043 18244 6552 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 5828 18204 5856 18235
rect 6546 18232 6552 18244
rect 6604 18232 6610 18284
rect 6638 18232 6644 18284
rect 6696 18232 6702 18284
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 6178 18204 6184 18216
rect 5828 18176 6184 18204
rect 6178 18164 6184 18176
rect 6236 18204 6242 18216
rect 6656 18204 6684 18232
rect 6236 18176 6684 18204
rect 6840 18204 6868 18235
rect 6914 18232 6920 18284
rect 6972 18272 6978 18284
rect 7285 18275 7343 18281
rect 7285 18272 7297 18275
rect 6972 18244 7297 18272
rect 6972 18232 6978 18244
rect 7285 18241 7297 18244
rect 7331 18272 7343 18275
rect 7834 18272 7840 18284
rect 7331 18244 7840 18272
rect 7331 18241 7343 18244
rect 7285 18235 7343 18241
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 9416 18281 9444 18312
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18241 9459 18275
rect 9401 18235 9459 18241
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 7006 18204 7012 18216
rect 6840 18176 7012 18204
rect 6236 18164 6242 18176
rect 7006 18164 7012 18176
rect 7064 18164 7070 18216
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7558 18204 7564 18216
rect 7515 18176 7564 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7558 18164 7564 18176
rect 7616 18164 7622 18216
rect 7653 18207 7711 18213
rect 7653 18173 7665 18207
rect 7699 18204 7711 18207
rect 7926 18204 7932 18216
rect 7699 18176 7932 18204
rect 7699 18173 7711 18176
rect 7653 18167 7711 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 5994 18096 6000 18148
rect 6052 18136 6058 18148
rect 9122 18136 9128 18148
rect 6052 18108 9128 18136
rect 6052 18096 6058 18108
rect 9122 18096 9128 18108
rect 9180 18136 9186 18148
rect 9600 18136 9628 18235
rect 9692 18204 9720 18235
rect 9766 18232 9772 18284
rect 9824 18232 9830 18284
rect 9858 18232 9864 18284
rect 9916 18232 9922 18284
rect 9876 18204 9904 18232
rect 9692 18176 9904 18204
rect 9968 18204 9996 18312
rect 10060 18312 12173 18340
rect 10060 18281 10088 18312
rect 12161 18309 12173 18312
rect 12207 18309 12219 18343
rect 12161 18303 12219 18309
rect 12989 18343 13047 18349
rect 12989 18309 13001 18343
rect 13035 18340 13047 18343
rect 13906 18340 13912 18352
rect 13035 18312 13912 18340
rect 13035 18309 13047 18312
rect 12989 18303 13047 18309
rect 13906 18300 13912 18312
rect 13964 18300 13970 18352
rect 14642 18300 14648 18352
rect 14700 18300 14706 18352
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 10134 18232 10140 18284
rect 10192 18272 10198 18284
rect 10229 18275 10287 18281
rect 10229 18272 10241 18275
rect 10192 18244 10241 18272
rect 10192 18232 10198 18244
rect 10229 18241 10241 18244
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 10336 18204 10364 18235
rect 10410 18232 10416 18284
rect 10468 18232 10474 18284
rect 11606 18272 11612 18284
rect 10520 18244 11612 18272
rect 10520 18204 10548 18244
rect 11606 18232 11612 18244
rect 11664 18232 11670 18284
rect 12618 18232 12624 18284
rect 12676 18232 12682 18284
rect 12769 18275 12827 18281
rect 12769 18241 12781 18275
rect 12815 18272 12827 18275
rect 12815 18241 12848 18272
rect 12769 18235 12848 18241
rect 9968 18176 10548 18204
rect 10781 18207 10839 18213
rect 10781 18173 10793 18207
rect 10827 18204 10839 18207
rect 11238 18204 11244 18216
rect 10827 18176 11244 18204
rect 10827 18173 10839 18176
rect 10781 18167 10839 18173
rect 11238 18164 11244 18176
rect 11296 18164 11302 18216
rect 11330 18164 11336 18216
rect 11388 18204 11394 18216
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 11388 18176 11529 18204
rect 11388 18164 11394 18176
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 12820 18204 12848 18235
rect 12894 18232 12900 18284
rect 12952 18232 12958 18284
rect 13127 18275 13185 18281
rect 13127 18241 13139 18275
rect 13173 18272 13185 18275
rect 13354 18272 13360 18284
rect 13173 18244 13360 18272
rect 13173 18241 13185 18244
rect 13127 18235 13185 18241
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 13449 18207 13507 18213
rect 13449 18204 13461 18207
rect 12820 18176 13461 18204
rect 11517 18167 11575 18173
rect 13449 18173 13461 18176
rect 13495 18204 13507 18207
rect 13814 18204 13820 18216
rect 13495 18176 13820 18204
rect 13495 18173 13507 18176
rect 13449 18167 13507 18173
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 10318 18136 10324 18148
rect 9180 18108 10324 18136
rect 9180 18096 9186 18108
rect 10318 18096 10324 18108
rect 10376 18096 10382 18148
rect 14660 18136 14688 18300
rect 14752 18281 14780 18380
rect 16574 18368 16580 18380
rect 16632 18408 16638 18420
rect 17954 18408 17960 18420
rect 16632 18380 17080 18408
rect 16632 18368 16638 18380
rect 15470 18300 15476 18352
rect 15528 18300 15534 18352
rect 17052 18281 17080 18380
rect 17328 18380 17960 18408
rect 17328 18349 17356 18380
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 18046 18368 18052 18420
rect 18104 18408 18110 18420
rect 18104 18380 18644 18408
rect 18104 18368 18110 18380
rect 17313 18343 17371 18349
rect 17313 18309 17325 18343
rect 17359 18309 17371 18343
rect 17313 18303 17371 18309
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18241 17095 18275
rect 18616 18272 18644 18380
rect 18782 18368 18788 18420
rect 18840 18368 18846 18420
rect 19610 18368 19616 18420
rect 19668 18408 19674 18420
rect 19794 18408 19800 18420
rect 19668 18380 19800 18408
rect 19668 18368 19674 18380
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 19886 18368 19892 18420
rect 19944 18408 19950 18420
rect 20993 18411 21051 18417
rect 19944 18380 20668 18408
rect 19944 18368 19950 18380
rect 19812 18340 19840 18368
rect 20640 18349 20668 18380
rect 20993 18377 21005 18411
rect 21039 18408 21051 18411
rect 25314 18408 25320 18420
rect 21039 18380 25320 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 25314 18368 25320 18380
rect 25372 18368 25378 18420
rect 20625 18343 20683 18349
rect 19812 18312 20485 18340
rect 19058 18272 19064 18284
rect 17037 18235 17095 18241
rect 15013 18207 15071 18213
rect 15013 18173 15025 18207
rect 15059 18204 15071 18207
rect 15470 18204 15476 18216
rect 15059 18176 15476 18204
rect 15059 18173 15071 18176
rect 15013 18167 15071 18173
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 18046 18204 18052 18216
rect 15620 18176 18052 18204
rect 15620 18164 15626 18176
rect 18046 18164 18052 18176
rect 18104 18204 18110 18216
rect 18432 18204 18460 18258
rect 18616 18244 19064 18272
rect 19058 18232 19064 18244
rect 19116 18272 19122 18284
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 19116 18244 19349 18272
rect 19116 18232 19122 18244
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 19337 18235 19395 18241
rect 19426 18232 19432 18284
rect 19484 18232 19490 18284
rect 19794 18232 19800 18284
rect 19852 18232 19858 18284
rect 20457 18281 20485 18312
rect 20625 18309 20637 18343
rect 20671 18309 20683 18343
rect 23474 18340 23480 18352
rect 20625 18303 20683 18309
rect 22940 18312 23480 18340
rect 20349 18275 20407 18281
rect 20349 18241 20361 18275
rect 20395 18241 20407 18275
rect 20349 18235 20407 18241
rect 20442 18275 20500 18281
rect 20442 18241 20454 18275
rect 20488 18241 20500 18275
rect 20442 18235 20500 18241
rect 18506 18204 18512 18216
rect 18104 18176 18512 18204
rect 18104 18164 18110 18176
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 19242 18164 19248 18216
rect 19300 18164 19306 18216
rect 20364 18204 20392 18235
rect 20714 18232 20720 18284
rect 20772 18232 20778 18284
rect 20806 18232 20812 18284
rect 20864 18281 20870 18284
rect 20864 18272 20872 18281
rect 21266 18272 21272 18284
rect 20864 18244 21272 18272
rect 20864 18235 20872 18244
rect 20864 18232 20870 18235
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 22940 18281 22968 18312
rect 23474 18300 23480 18312
rect 23532 18300 23538 18352
rect 24486 18340 24492 18352
rect 24426 18312 24492 18340
rect 24486 18300 24492 18312
rect 24544 18340 24550 18352
rect 24946 18340 24952 18352
rect 24544 18312 24952 18340
rect 24544 18300 24550 18312
rect 24946 18300 24952 18312
rect 25004 18300 25010 18352
rect 27982 18300 27988 18352
rect 28040 18300 28046 18352
rect 22925 18275 22983 18281
rect 22925 18241 22937 18275
rect 22971 18241 22983 18275
rect 22925 18235 22983 18241
rect 19352 18176 20392 18204
rect 16758 18136 16764 18148
rect 12406 18108 14688 18136
rect 16040 18108 16764 18136
rect 5445 18071 5503 18077
rect 5445 18068 5457 18071
rect 5224 18040 5457 18068
rect 5224 18028 5230 18040
rect 5445 18037 5457 18040
rect 5491 18037 5503 18071
rect 5445 18031 5503 18037
rect 6181 18071 6239 18077
rect 6181 18037 6193 18071
rect 6227 18068 6239 18071
rect 7650 18068 7656 18080
rect 6227 18040 7656 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 9953 18071 10011 18077
rect 9953 18068 9965 18071
rect 9916 18040 9965 18068
rect 9916 18028 9922 18040
rect 9953 18037 9965 18040
rect 9999 18037 10011 18071
rect 9953 18031 10011 18037
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10192 18040 10609 18068
rect 10192 18028 10198 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 10597 18031 10655 18037
rect 11146 18028 11152 18080
rect 11204 18068 11210 18080
rect 12406 18068 12434 18108
rect 11204 18040 12434 18068
rect 13265 18071 13323 18077
rect 11204 18028 11210 18040
rect 13265 18037 13277 18071
rect 13311 18068 13323 18071
rect 16040 18068 16068 18108
rect 16758 18096 16764 18108
rect 16816 18096 16822 18148
rect 18322 18096 18328 18148
rect 18380 18136 18386 18148
rect 19352 18136 19380 18176
rect 23198 18164 23204 18216
rect 23256 18164 23262 18216
rect 24949 18207 25007 18213
rect 24949 18204 24961 18207
rect 24320 18176 24961 18204
rect 18380 18108 19380 18136
rect 20257 18139 20315 18145
rect 18380 18096 18386 18108
rect 20257 18105 20269 18139
rect 20303 18136 20315 18139
rect 20898 18136 20904 18148
rect 20303 18108 20904 18136
rect 20303 18105 20315 18108
rect 20257 18099 20315 18105
rect 20898 18096 20904 18108
rect 20956 18096 20962 18148
rect 13311 18040 16068 18068
rect 13311 18037 13323 18040
rect 13265 18031 13323 18037
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16485 18071 16543 18077
rect 16485 18068 16497 18071
rect 16172 18040 16497 18068
rect 16172 18028 16178 18040
rect 16485 18037 16497 18040
rect 16531 18037 16543 18071
rect 16485 18031 16543 18037
rect 22646 18028 22652 18080
rect 22704 18068 22710 18080
rect 24320 18068 24348 18176
rect 24949 18173 24961 18176
rect 24995 18204 25007 18207
rect 25041 18207 25099 18213
rect 25041 18204 25053 18207
rect 24995 18176 25053 18204
rect 24995 18173 25007 18176
rect 24949 18167 25007 18173
rect 25041 18173 25053 18176
rect 25087 18204 25099 18207
rect 25498 18204 25504 18216
rect 25087 18176 25504 18204
rect 25087 18173 25099 18176
rect 25041 18167 25099 18173
rect 25498 18164 25504 18176
rect 25556 18204 25562 18216
rect 26142 18204 26148 18216
rect 25556 18176 26148 18204
rect 25556 18164 25562 18176
rect 26142 18164 26148 18176
rect 26200 18164 26206 18216
rect 26878 18164 26884 18216
rect 26936 18204 26942 18216
rect 26973 18207 27031 18213
rect 26973 18204 26985 18207
rect 26936 18176 26985 18204
rect 26936 18164 26942 18176
rect 26973 18173 26985 18176
rect 27019 18173 27031 18207
rect 26973 18167 27031 18173
rect 27246 18164 27252 18216
rect 27304 18164 27310 18216
rect 28442 18164 28448 18216
rect 28500 18204 28506 18216
rect 28997 18207 29055 18213
rect 28997 18204 29009 18207
rect 28500 18176 29009 18204
rect 28500 18164 28506 18176
rect 28997 18173 29009 18176
rect 29043 18173 29055 18207
rect 28997 18167 29055 18173
rect 22704 18040 24348 18068
rect 22704 18028 22710 18040
rect 24854 18028 24860 18080
rect 24912 18068 24918 18080
rect 25685 18071 25743 18077
rect 25685 18068 25697 18071
rect 24912 18040 25697 18068
rect 24912 18028 24918 18040
rect 25685 18037 25697 18040
rect 25731 18037 25743 18071
rect 25685 18031 25743 18037
rect 26602 18028 26608 18080
rect 26660 18068 26666 18080
rect 26970 18068 26976 18080
rect 26660 18040 26976 18068
rect 26660 18028 26666 18040
rect 26970 18028 26976 18040
rect 27028 18028 27034 18080
rect 1104 17978 29440 18000
rect 1104 17926 4491 17978
rect 4543 17926 4555 17978
rect 4607 17926 4619 17978
rect 4671 17926 4683 17978
rect 4735 17926 4747 17978
rect 4799 17926 11574 17978
rect 11626 17926 11638 17978
rect 11690 17926 11702 17978
rect 11754 17926 11766 17978
rect 11818 17926 11830 17978
rect 11882 17926 18657 17978
rect 18709 17926 18721 17978
rect 18773 17926 18785 17978
rect 18837 17926 18849 17978
rect 18901 17926 18913 17978
rect 18965 17926 25740 17978
rect 25792 17926 25804 17978
rect 25856 17926 25868 17978
rect 25920 17926 25932 17978
rect 25984 17926 25996 17978
rect 26048 17926 29440 17978
rect 1104 17904 29440 17926
rect 7374 17824 7380 17876
rect 7432 17824 7438 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 11974 17864 11980 17876
rect 10652 17836 11980 17864
rect 10652 17824 10658 17836
rect 7392 17796 7420 17824
rect 6656 17768 7420 17796
rect 3694 17688 3700 17740
rect 3752 17728 3758 17740
rect 5261 17731 5319 17737
rect 5261 17728 5273 17731
rect 3752 17700 5273 17728
rect 3752 17688 3758 17700
rect 5261 17697 5273 17700
rect 5307 17697 5319 17731
rect 5261 17691 5319 17697
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 5166 17660 5172 17672
rect 4479 17632 5172 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6656 17646 6684 17768
rect 11330 17756 11336 17808
rect 11388 17796 11394 17808
rect 11388 17768 11836 17796
rect 11388 17756 11394 17768
rect 7009 17731 7067 17737
rect 7009 17697 7021 17731
rect 7055 17728 7067 17731
rect 9585 17731 9643 17737
rect 7055 17700 7972 17728
rect 7055 17697 7067 17700
rect 7009 17691 7067 17697
rect 7282 17620 7288 17672
rect 7340 17620 7346 17672
rect 7392 17669 7420 17700
rect 7944 17672 7972 17700
rect 9585 17697 9597 17731
rect 9631 17728 9643 17731
rect 9950 17728 9956 17740
rect 9631 17700 9956 17728
rect 9631 17697 9643 17700
rect 9585 17691 9643 17697
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10888 17700 11192 17728
rect 10888 17672 10916 17700
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 7561 17663 7619 17669
rect 7561 17629 7573 17663
rect 7607 17629 7619 17663
rect 7561 17623 7619 17629
rect 3418 17552 3424 17604
rect 3476 17592 3482 17604
rect 4522 17592 4528 17604
rect 3476 17564 4528 17592
rect 3476 17552 3482 17564
rect 4522 17552 4528 17564
rect 4580 17552 4586 17604
rect 5537 17595 5595 17601
rect 5537 17561 5549 17595
rect 5583 17592 5595 17595
rect 5810 17592 5816 17604
rect 5583 17564 5816 17592
rect 5583 17561 5595 17564
rect 5537 17555 5595 17561
rect 5810 17552 5816 17564
rect 5868 17552 5874 17604
rect 7098 17552 7104 17604
rect 7156 17552 7162 17604
rect 4798 17484 4804 17536
rect 4856 17524 4862 17536
rect 4985 17527 5043 17533
rect 4985 17524 4997 17527
rect 4856 17496 4997 17524
rect 4856 17484 4862 17496
rect 4985 17493 4997 17496
rect 5031 17493 5043 17527
rect 4985 17487 5043 17493
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 7576 17524 7604 17623
rect 7650 17620 7656 17672
rect 7708 17620 7714 17672
rect 7926 17620 7932 17672
rect 7984 17620 7990 17672
rect 10870 17620 10876 17672
rect 10928 17620 10934 17672
rect 9861 17595 9919 17601
rect 9861 17561 9873 17595
rect 9907 17592 9919 17595
rect 10134 17592 10140 17604
rect 9907 17564 10140 17592
rect 9907 17561 9919 17564
rect 9861 17555 9919 17561
rect 10134 17552 10140 17564
rect 10192 17552 10198 17604
rect 6420 17496 7604 17524
rect 6420 17484 6426 17496
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 10980 17524 11008 17646
rect 10928 17496 11008 17524
rect 11164 17524 11192 17700
rect 11238 17620 11244 17672
rect 11296 17620 11302 17672
rect 11422 17620 11428 17672
rect 11480 17620 11486 17672
rect 11808 17669 11836 17768
rect 11900 17669 11928 17836
rect 11974 17824 11980 17836
rect 12032 17824 12038 17876
rect 12069 17867 12127 17873
rect 12069 17833 12081 17867
rect 12115 17864 12127 17867
rect 12618 17864 12624 17876
rect 12115 17836 12624 17864
rect 12115 17833 12127 17836
rect 12069 17827 12127 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 13906 17824 13912 17876
rect 13964 17824 13970 17876
rect 15657 17867 15715 17873
rect 15657 17833 15669 17867
rect 15703 17864 15715 17867
rect 15930 17864 15936 17876
rect 15703 17836 15936 17864
rect 15703 17833 15715 17836
rect 15657 17827 15715 17833
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 19610 17864 19616 17876
rect 16040 17836 19616 17864
rect 15102 17756 15108 17808
rect 15160 17796 15166 17808
rect 16040 17796 16068 17836
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 19794 17824 19800 17876
rect 19852 17824 19858 17876
rect 23198 17824 23204 17876
rect 23256 17864 23262 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 23256 17836 23305 17864
rect 23256 17824 23262 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 25056 17836 25820 17864
rect 22373 17799 22431 17805
rect 15160 17768 16068 17796
rect 19306 17768 20116 17796
rect 15160 17756 15166 17768
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17728 12219 17731
rect 17313 17731 17371 17737
rect 17313 17728 17325 17731
rect 12207 17700 17325 17728
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 17313 17697 17325 17700
rect 17359 17728 17371 17731
rect 19306 17728 19334 17768
rect 20088 17740 20116 17768
rect 22373 17765 22385 17799
rect 22419 17796 22431 17799
rect 22738 17796 22744 17808
rect 22419 17768 22744 17796
rect 22419 17765 22431 17768
rect 22373 17759 22431 17765
rect 22738 17756 22744 17768
rect 22796 17796 22802 17808
rect 25056 17805 25084 17836
rect 22925 17799 22983 17805
rect 22925 17796 22937 17799
rect 22796 17768 22937 17796
rect 22796 17756 22802 17768
rect 22925 17765 22937 17768
rect 22971 17765 22983 17799
rect 25041 17799 25099 17805
rect 22925 17759 22983 17765
rect 23308 17768 23888 17796
rect 17359 17700 19334 17728
rect 19444 17700 19840 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 11518 17663 11576 17669
rect 11518 17629 11530 17663
rect 11564 17629 11576 17663
rect 11518 17623 11576 17629
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 11890 17663 11948 17669
rect 11890 17629 11902 17663
rect 11936 17629 11948 17663
rect 11890 17623 11948 17629
rect 11256 17592 11284 17620
rect 11532 17592 11560 17623
rect 16114 17620 16120 17672
rect 16172 17620 16178 17672
rect 19444 17669 19472 17700
rect 19812 17672 19840 17700
rect 20070 17688 20076 17740
rect 20128 17688 20134 17740
rect 20346 17688 20352 17740
rect 20404 17688 20410 17740
rect 20714 17688 20720 17740
rect 20772 17728 20778 17740
rect 21821 17731 21879 17737
rect 21821 17728 21833 17731
rect 20772 17700 21833 17728
rect 20772 17688 20778 17700
rect 21821 17697 21833 17700
rect 21867 17728 21879 17731
rect 22002 17728 22008 17740
rect 21867 17700 22008 17728
rect 21867 17697 21879 17700
rect 21821 17691 21879 17697
rect 22002 17688 22008 17700
rect 22060 17728 22066 17740
rect 23017 17731 23075 17737
rect 23017 17728 23029 17731
rect 22060 17700 23029 17728
rect 22060 17688 22066 17700
rect 23017 17697 23029 17700
rect 23063 17697 23075 17731
rect 23017 17691 23075 17697
rect 23308 17672 23336 17768
rect 23750 17728 23756 17740
rect 23492 17700 23756 17728
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18892 17632 19257 17660
rect 11256 17564 11560 17592
rect 11701 17595 11759 17601
rect 11701 17561 11713 17595
rect 11747 17561 11759 17595
rect 11701 17555 11759 17561
rect 12437 17595 12495 17601
rect 12437 17561 12449 17595
rect 12483 17561 12495 17595
rect 12437 17555 12495 17561
rect 11716 17524 11744 17555
rect 11164 17496 11744 17524
rect 12452 17524 12480 17555
rect 13078 17552 13084 17604
rect 13136 17552 13142 17604
rect 14182 17552 14188 17604
rect 14240 17552 14246 17604
rect 17586 17552 17592 17604
rect 17644 17552 17650 17604
rect 18046 17552 18052 17604
rect 18104 17552 18110 17604
rect 14642 17524 14648 17536
rect 12452 17496 14648 17524
rect 10928 17484 10934 17496
rect 14642 17484 14648 17496
rect 14700 17484 14706 17536
rect 16666 17484 16672 17536
rect 16724 17484 16730 17536
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 17862 17524 17868 17536
rect 17184 17496 17868 17524
rect 17184 17484 17190 17496
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 18892 17524 18920 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19518 17620 19524 17672
rect 19576 17620 19582 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19702 17660 19708 17672
rect 19659 17632 19708 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 19702 17620 19708 17632
rect 19760 17620 19766 17672
rect 19794 17620 19800 17672
rect 19852 17620 19858 17672
rect 22278 17620 22284 17672
rect 22336 17620 22342 17672
rect 22646 17620 22652 17672
rect 22704 17660 22710 17672
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 22704 17632 22753 17660
rect 22704 17620 22710 17632
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 23290 17620 23296 17672
rect 23348 17620 23354 17672
rect 23492 17669 23520 17700
rect 23750 17688 23756 17700
rect 23808 17688 23814 17740
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17629 23535 17663
rect 23860 17660 23888 17768
rect 25041 17765 25053 17799
rect 25087 17765 25099 17799
rect 25041 17759 25099 17765
rect 23937 17731 23995 17737
rect 23937 17697 23949 17731
rect 23983 17728 23995 17731
rect 24854 17728 24860 17740
rect 23983 17700 24860 17728
rect 23983 17697 23995 17700
rect 23937 17691 23995 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25792 17737 25820 17836
rect 25958 17824 25964 17876
rect 26016 17864 26022 17876
rect 27157 17867 27215 17873
rect 26016 17836 27016 17864
rect 26016 17824 26022 17836
rect 25869 17799 25927 17805
rect 25869 17765 25881 17799
rect 25915 17796 25927 17799
rect 26234 17796 26240 17808
rect 25915 17768 26240 17796
rect 25915 17765 25927 17768
rect 25869 17759 25927 17765
rect 26234 17756 26240 17768
rect 26292 17756 26298 17808
rect 26436 17768 26924 17796
rect 26436 17740 26464 17768
rect 25777 17731 25835 17737
rect 25240 17700 25682 17728
rect 24394 17660 24400 17672
rect 23860 17632 24400 17660
rect 23477 17623 23535 17629
rect 24394 17620 24400 17632
rect 24452 17620 24458 17672
rect 25240 17660 25268 17700
rect 25654 17669 25682 17700
rect 25777 17697 25789 17731
rect 25823 17697 25835 17731
rect 25777 17691 25835 17697
rect 26050 17688 26056 17740
rect 26108 17688 26114 17740
rect 26142 17688 26148 17740
rect 26200 17688 26206 17740
rect 26418 17688 26424 17740
rect 26476 17688 26482 17740
rect 26510 17688 26516 17740
rect 26568 17688 26574 17740
rect 24990 17632 25268 17660
rect 25501 17663 25559 17669
rect 18966 17552 18972 17604
rect 19024 17592 19030 17604
rect 19024 17564 20838 17592
rect 19024 17552 19030 17564
rect 23566 17552 23572 17604
rect 23624 17552 23630 17604
rect 23661 17595 23719 17601
rect 23661 17561 23673 17595
rect 23707 17561 23719 17595
rect 23661 17555 23719 17561
rect 23799 17595 23857 17601
rect 23799 17561 23811 17595
rect 23845 17592 23857 17595
rect 24026 17592 24032 17604
rect 23845 17564 24032 17592
rect 23845 17561 23857 17564
rect 23799 17555 23857 17561
rect 18472 17496 18920 17524
rect 18472 17484 18478 17496
rect 19058 17484 19064 17536
rect 19116 17484 19122 17536
rect 22557 17527 22615 17533
rect 22557 17493 22569 17527
rect 22603 17524 22615 17527
rect 23106 17524 23112 17536
rect 22603 17496 23112 17524
rect 22603 17493 22615 17496
rect 22557 17487 22615 17493
rect 23106 17484 23112 17496
rect 23164 17484 23170 17536
rect 23676 17524 23704 17555
rect 24026 17552 24032 17564
rect 24084 17592 24090 17604
rect 24990 17592 25018 17632
rect 25314 17598 25320 17650
rect 25372 17598 25378 17650
rect 25501 17629 25513 17663
rect 25547 17629 25559 17663
rect 25501 17623 25559 17629
rect 25639 17663 25697 17669
rect 25639 17629 25651 17663
rect 25685 17660 25697 17663
rect 25958 17660 25964 17672
rect 25685 17632 25964 17660
rect 25685 17629 25697 17632
rect 25639 17623 25697 17629
rect 24084 17564 25018 17592
rect 25056 17564 25268 17592
rect 24084 17552 24090 17564
rect 25056 17524 25084 17564
rect 25240 17536 25268 17564
rect 25406 17552 25412 17604
rect 25464 17552 25470 17604
rect 25516 17592 25544 17623
rect 25958 17620 25964 17632
rect 26016 17620 26022 17672
rect 26602 17620 26608 17672
rect 26660 17620 26666 17672
rect 26896 17669 26924 17768
rect 26988 17669 27016 17836
rect 27157 17833 27169 17867
rect 27203 17864 27215 17867
rect 27246 17864 27252 17876
rect 27203 17836 27252 17864
rect 27203 17833 27215 17836
rect 27157 17827 27215 17833
rect 27246 17824 27252 17836
rect 27304 17824 27310 17876
rect 27338 17756 27344 17808
rect 27396 17796 27402 17808
rect 27985 17799 28043 17805
rect 27985 17796 27997 17799
rect 27396 17768 27997 17796
rect 27396 17756 27402 17768
rect 27985 17765 27997 17768
rect 28031 17765 28043 17799
rect 27985 17759 28043 17765
rect 27632 17700 28304 17728
rect 26881 17663 26939 17669
rect 26881 17629 26893 17663
rect 26927 17629 26939 17663
rect 26881 17623 26939 17629
rect 26973 17663 27031 17669
rect 26973 17629 26985 17663
rect 27019 17629 27031 17663
rect 26973 17623 27031 17629
rect 27522 17620 27528 17672
rect 27580 17660 27586 17672
rect 27632 17669 27660 17700
rect 27617 17663 27675 17669
rect 27617 17660 27629 17663
rect 27580 17632 27629 17660
rect 27580 17620 27586 17632
rect 27617 17629 27629 17632
rect 27663 17660 27675 17663
rect 27663 17632 27717 17660
rect 27663 17629 27675 17632
rect 27617 17623 27675 17629
rect 27890 17620 27896 17672
rect 27948 17620 27954 17672
rect 28169 17663 28227 17669
rect 28169 17660 28181 17663
rect 28000 17632 28181 17660
rect 26789 17595 26847 17601
rect 26789 17592 26801 17595
rect 25516 17564 26801 17592
rect 23676 17496 25084 17524
rect 25130 17484 25136 17536
rect 25188 17484 25194 17536
rect 25222 17484 25228 17536
rect 25280 17524 25286 17536
rect 25516 17524 25544 17564
rect 26789 17561 26801 17564
rect 26835 17561 26847 17595
rect 26789 17555 26847 17561
rect 27154 17552 27160 17604
rect 27212 17592 27218 17604
rect 27433 17595 27491 17601
rect 27433 17592 27445 17595
rect 27212 17564 27445 17592
rect 27212 17552 27218 17564
rect 27433 17561 27445 17564
rect 27479 17561 27491 17595
rect 28000 17592 28028 17632
rect 28169 17629 28181 17632
rect 28215 17629 28227 17663
rect 28169 17623 28227 17629
rect 27433 17555 27491 17561
rect 27816 17564 28028 17592
rect 28276 17592 28304 17700
rect 28353 17663 28411 17669
rect 28353 17629 28365 17663
rect 28399 17660 28411 17663
rect 28399 17632 28488 17660
rect 28399 17629 28411 17632
rect 28353 17623 28411 17629
rect 28460 17604 28488 17632
rect 28276 17564 28396 17592
rect 25280 17496 25544 17524
rect 25280 17484 25286 17496
rect 25590 17484 25596 17536
rect 25648 17524 25654 17536
rect 26142 17524 26148 17536
rect 25648 17496 26148 17524
rect 25648 17484 25654 17496
rect 26142 17484 26148 17496
rect 26200 17524 26206 17536
rect 26237 17527 26295 17533
rect 26237 17524 26249 17527
rect 26200 17496 26249 17524
rect 26200 17484 26206 17496
rect 26237 17493 26249 17496
rect 26283 17493 26295 17527
rect 26237 17487 26295 17493
rect 26421 17527 26479 17533
rect 26421 17493 26433 17527
rect 26467 17524 26479 17527
rect 26510 17524 26516 17536
rect 26467 17496 26516 17524
rect 26467 17493 26479 17496
rect 26421 17487 26479 17493
rect 26510 17484 26516 17496
rect 26568 17484 26574 17536
rect 27614 17484 27620 17536
rect 27672 17524 27678 17536
rect 27816 17533 27844 17564
rect 28368 17536 28396 17564
rect 28442 17552 28448 17604
rect 28500 17552 28506 17604
rect 27801 17527 27859 17533
rect 27801 17524 27813 17527
rect 27672 17496 27813 17524
rect 27672 17484 27678 17496
rect 27801 17493 27813 17496
rect 27847 17493 27859 17527
rect 27801 17487 27859 17493
rect 28074 17484 28080 17536
rect 28132 17524 28138 17536
rect 28261 17527 28319 17533
rect 28261 17524 28273 17527
rect 28132 17496 28273 17524
rect 28132 17484 28138 17496
rect 28261 17493 28273 17496
rect 28307 17493 28319 17527
rect 28261 17487 28319 17493
rect 28350 17484 28356 17536
rect 28408 17484 28414 17536
rect 1104 17434 29440 17456
rect 1104 17382 5151 17434
rect 5203 17382 5215 17434
rect 5267 17382 5279 17434
rect 5331 17382 5343 17434
rect 5395 17382 5407 17434
rect 5459 17382 12234 17434
rect 12286 17382 12298 17434
rect 12350 17382 12362 17434
rect 12414 17382 12426 17434
rect 12478 17382 12490 17434
rect 12542 17382 19317 17434
rect 19369 17382 19381 17434
rect 19433 17382 19445 17434
rect 19497 17382 19509 17434
rect 19561 17382 19573 17434
rect 19625 17382 26400 17434
rect 26452 17382 26464 17434
rect 26516 17382 26528 17434
rect 26580 17382 26592 17434
rect 26644 17382 26656 17434
rect 26708 17382 29440 17434
rect 1104 17360 29440 17382
rect 4062 17320 4068 17332
rect 3712 17292 4068 17320
rect 3234 17212 3240 17264
rect 3292 17252 3298 17264
rect 3513 17255 3571 17261
rect 3513 17252 3525 17255
rect 3292 17224 3525 17252
rect 3292 17212 3298 17224
rect 3513 17221 3525 17224
rect 3559 17221 3571 17255
rect 3513 17215 3571 17221
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17184 3387 17187
rect 3375 17156 3464 17184
rect 3375 17153 3387 17156
rect 3329 17147 3387 17153
rect 3436 17128 3464 17156
rect 3418 17076 3424 17128
rect 3476 17076 3482 17128
rect 3528 17116 3556 17215
rect 3602 17144 3608 17196
rect 3660 17144 3666 17196
rect 3712 17193 3740 17292
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4522 17280 4528 17332
rect 4580 17280 4586 17332
rect 4982 17320 4988 17332
rect 4632 17292 4988 17320
rect 4249 17255 4307 17261
rect 4249 17221 4261 17255
rect 4295 17252 4307 17255
rect 4632 17252 4660 17292
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5169 17323 5227 17329
rect 5169 17320 5181 17323
rect 5132 17292 5181 17320
rect 5132 17280 5138 17292
rect 5169 17289 5181 17292
rect 5215 17289 5227 17323
rect 5169 17283 5227 17289
rect 5258 17280 5264 17332
rect 5316 17280 5322 17332
rect 5368 17292 7420 17320
rect 4801 17255 4859 17261
rect 4801 17252 4813 17255
rect 4295 17224 4660 17252
rect 4295 17221 4307 17224
rect 4249 17215 4307 17221
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 3970 17144 3976 17196
rect 4028 17144 4034 17196
rect 4632 17193 4660 17224
rect 4724 17224 4813 17252
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17153 4215 17187
rect 4157 17147 4215 17153
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17153 4399 17187
rect 4341 17147 4399 17153
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 4172 17116 4200 17147
rect 3528 17088 4200 17116
rect 3988 17060 4016 17088
rect 3970 17008 3976 17060
rect 4028 17008 4034 17060
rect 4356 17048 4384 17147
rect 4080 17020 4384 17048
rect 4724 17048 4752 17224
rect 4801 17221 4813 17224
rect 4847 17221 4859 17255
rect 5276 17252 5304 17280
rect 4801 17215 4859 17221
rect 5092 17224 5304 17252
rect 4893 17187 4951 17193
rect 4893 17184 4905 17187
rect 4816 17156 4905 17184
rect 4816 17128 4844 17156
rect 4893 17153 4905 17156
rect 4939 17153 4951 17187
rect 4893 17147 4951 17153
rect 4985 17187 5043 17193
rect 4985 17153 4997 17187
rect 5031 17184 5043 17187
rect 5092 17184 5120 17224
rect 5031 17156 5120 17184
rect 5031 17153 5043 17156
rect 4985 17147 5043 17153
rect 5166 17144 5172 17196
rect 5224 17184 5230 17196
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 5224 17156 5273 17184
rect 5224 17144 5230 17156
rect 5261 17153 5273 17156
rect 5307 17184 5319 17187
rect 5368 17184 5396 17292
rect 5445 17255 5503 17261
rect 5445 17221 5457 17255
rect 5491 17252 5503 17255
rect 5994 17252 6000 17264
rect 5491 17224 6000 17252
rect 5491 17221 5503 17224
rect 5445 17215 5503 17221
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 7392 17196 7420 17292
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 12802 17320 12808 17332
rect 10008 17292 12204 17320
rect 10008 17280 10014 17292
rect 9968 17252 9996 17280
rect 9600 17224 9996 17252
rect 5534 17193 5540 17196
rect 5307 17156 5396 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 5533 17147 5540 17193
rect 5534 17144 5540 17147
rect 5592 17144 5598 17196
rect 5626 17144 5632 17196
rect 5684 17184 5690 17196
rect 5684 17156 6224 17184
rect 5684 17144 5690 17156
rect 4798 17076 4804 17128
rect 4856 17076 4862 17128
rect 4724 17020 6040 17048
rect 4080 16992 4108 17020
rect 6012 16992 6040 17020
rect 6196 16992 6224 17156
rect 7374 17144 7380 17196
rect 7432 17144 7438 17196
rect 9600 17193 9628 17224
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 10870 17144 10876 17196
rect 10928 17184 10934 17196
rect 12176 17193 12204 17292
rect 12452 17292 12808 17320
rect 12452 17261 12480 17292
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 13909 17323 13967 17329
rect 13909 17320 13921 17323
rect 13872 17292 13921 17320
rect 13872 17280 13878 17292
rect 13909 17289 13921 17292
rect 13955 17289 13967 17323
rect 16666 17320 16672 17332
rect 13909 17283 13967 17289
rect 15028 17292 16672 17320
rect 12437 17255 12495 17261
rect 12437 17221 12449 17255
rect 12483 17221 12495 17255
rect 12437 17215 12495 17221
rect 12161 17187 12219 17193
rect 10928 17170 10994 17184
rect 10928 17156 11008 17170
rect 10928 17144 10934 17156
rect 9858 17076 9864 17128
rect 9916 17076 9922 17128
rect 10980 17116 11008 17156
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 13078 17116 13084 17128
rect 10980 17088 13084 17116
rect 13078 17076 13084 17088
rect 13136 17116 13142 17128
rect 13556 17116 13584 17170
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 15028 17193 15056 17292
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 16758 17280 16764 17332
rect 16816 17320 16822 17332
rect 16816 17292 17356 17320
rect 16816 17280 16822 17292
rect 15102 17212 15108 17264
rect 15160 17212 15166 17264
rect 15197 17255 15255 17261
rect 15197 17221 15209 17255
rect 15243 17252 15255 17255
rect 15746 17252 15752 17264
rect 15243 17224 15752 17252
rect 15243 17221 15255 17224
rect 15197 17215 15255 17221
rect 15746 17212 15752 17224
rect 15804 17212 15810 17264
rect 16114 17212 16120 17264
rect 16172 17252 16178 17264
rect 16172 17224 17080 17252
rect 16172 17212 16178 17224
rect 14001 17187 14059 17193
rect 14001 17184 14013 17187
rect 13964 17156 14013 17184
rect 13964 17144 13970 17156
rect 14001 17153 14013 17156
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 15120 17184 15148 17212
rect 15289 17187 15347 17193
rect 15289 17184 15301 17187
rect 15120 17156 15301 17184
rect 13136 17088 13584 17116
rect 13136 17076 13142 17088
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14366 17116 14372 17128
rect 14148 17088 14372 17116
rect 14148 17076 14154 17088
rect 14366 17076 14372 17088
rect 14424 17116 14430 17128
rect 15120 17116 15148 17156
rect 15289 17153 15301 17156
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 14424 17088 15148 17116
rect 14424 17076 14430 17088
rect 11238 17008 11244 17060
rect 11296 17048 11302 17060
rect 11333 17051 11391 17057
rect 11333 17048 11345 17051
rect 11296 17020 11345 17048
rect 11296 17008 11302 17020
rect 11333 17017 11345 17020
rect 11379 17017 11391 17051
rect 11333 17011 11391 17017
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 3881 16983 3939 16989
rect 3881 16980 3893 16983
rect 3384 16952 3893 16980
rect 3384 16940 3390 16952
rect 3881 16949 3893 16952
rect 3927 16949 3939 16983
rect 3881 16943 3939 16949
rect 4062 16940 4068 16992
rect 4120 16940 4126 16992
rect 5810 16940 5816 16992
rect 5868 16940 5874 16992
rect 5994 16940 6000 16992
rect 6052 16940 6058 16992
rect 6178 16940 6184 16992
rect 6236 16940 6242 16992
rect 14090 16940 14096 16992
rect 14148 16980 14154 16992
rect 14645 16983 14703 16989
rect 14645 16980 14657 16983
rect 14148 16952 14657 16980
rect 14148 16940 14154 16952
rect 14645 16949 14657 16952
rect 14691 16949 14703 16983
rect 15396 16980 15424 17147
rect 16942 17144 16948 17196
rect 17000 17144 17006 17196
rect 17052 17193 17080 17224
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17126 17144 17132 17196
rect 17184 17144 17190 17196
rect 17328 17193 17356 17292
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 18785 17323 18843 17329
rect 18785 17320 18797 17323
rect 17644 17292 18797 17320
rect 17644 17280 17650 17292
rect 18785 17289 18797 17292
rect 18831 17289 18843 17323
rect 19058 17320 19064 17332
rect 18785 17283 18843 17289
rect 18892 17292 19064 17320
rect 18892 17261 18920 17292
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19242 17280 19248 17332
rect 19300 17280 19306 17332
rect 20346 17280 20352 17332
rect 20404 17320 20410 17332
rect 20809 17323 20867 17329
rect 20809 17320 20821 17323
rect 20404 17292 20821 17320
rect 20404 17280 20410 17292
rect 20809 17289 20821 17292
rect 20855 17289 20867 17323
rect 20809 17283 20867 17289
rect 21821 17323 21879 17329
rect 21821 17289 21833 17323
rect 21867 17289 21879 17323
rect 21821 17283 21879 17289
rect 23385 17323 23443 17329
rect 23385 17289 23397 17323
rect 23431 17320 23443 17323
rect 23566 17320 23572 17332
rect 23431 17292 23572 17320
rect 23431 17289 23443 17292
rect 23385 17283 23443 17289
rect 18877 17255 18935 17261
rect 18877 17252 18889 17255
rect 17604 17224 18889 17252
rect 17604 17193 17632 17224
rect 18877 17221 18889 17224
rect 18923 17221 18935 17255
rect 18877 17215 18935 17221
rect 19150 17212 19156 17264
rect 19208 17212 19214 17264
rect 21836 17252 21864 17283
rect 23566 17280 23572 17292
rect 23624 17280 23630 17332
rect 25130 17320 25136 17332
rect 23768 17292 25136 17320
rect 21008 17224 21864 17252
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 18141 17187 18199 17193
rect 18141 17153 18153 17187
rect 18187 17184 18199 17187
rect 18233 17187 18291 17193
rect 18233 17184 18245 17187
rect 18187 17156 18245 17184
rect 18187 17153 18199 17156
rect 18141 17147 18199 17153
rect 18233 17153 18245 17156
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17153 18475 17187
rect 18417 17147 18475 17153
rect 15470 17076 15476 17128
rect 15528 17076 15534 17128
rect 16669 17119 16727 17125
rect 16669 17085 16681 17119
rect 16715 17116 16727 17119
rect 18340 17116 18368 17144
rect 16715 17088 18368 17116
rect 16715 17085 16727 17088
rect 16669 17079 16727 17085
rect 15488 17048 15516 17076
rect 15565 17051 15623 17057
rect 15565 17048 15577 17051
rect 15488 17020 15577 17048
rect 15565 17017 15577 17020
rect 15611 17017 15623 17051
rect 15565 17011 15623 17017
rect 17494 17008 17500 17060
rect 17552 17048 17558 17060
rect 18432 17048 18460 17147
rect 18506 17144 18512 17196
rect 18564 17144 18570 17196
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19168 17184 19196 17212
rect 21008 17193 21036 17224
rect 22002 17212 22008 17264
rect 22060 17252 22066 17264
rect 23768 17261 23796 17292
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 25406 17280 25412 17332
rect 25464 17320 25470 17332
rect 25869 17323 25927 17329
rect 25869 17320 25881 17323
rect 25464 17292 25881 17320
rect 25464 17280 25470 17292
rect 25869 17289 25881 17292
rect 25915 17289 25927 17323
rect 25869 17283 25927 17289
rect 26050 17280 26056 17332
rect 26108 17280 26114 17332
rect 26142 17280 26148 17332
rect 26200 17320 26206 17332
rect 26418 17320 26424 17332
rect 26200 17292 26424 17320
rect 26200 17280 26206 17292
rect 26418 17280 26424 17292
rect 26476 17280 26482 17332
rect 26789 17323 26847 17329
rect 26789 17320 26801 17323
rect 26528 17292 26801 17320
rect 22281 17255 22339 17261
rect 22281 17252 22293 17255
rect 22060 17224 22293 17252
rect 22060 17212 22066 17224
rect 22281 17221 22293 17224
rect 22327 17221 22339 17255
rect 22281 17215 22339 17221
rect 23753 17255 23811 17261
rect 23753 17221 23765 17255
rect 23799 17221 23811 17255
rect 23753 17215 23811 17221
rect 25038 17212 25044 17264
rect 25096 17252 25102 17264
rect 26068 17252 26096 17280
rect 26237 17255 26295 17261
rect 26237 17252 26249 17255
rect 25096 17224 25452 17252
rect 25096 17212 25102 17224
rect 19107 17156 19196 17184
rect 20993 17187 21051 17193
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 22020 17184 22048 17212
rect 25424 17196 25452 17224
rect 25700 17224 26249 17252
rect 21315 17156 22048 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 17552 17020 18460 17048
rect 17552 17008 17558 17020
rect 16114 16980 16120 16992
rect 15396 16952 16120 16980
rect 14645 16943 14703 16949
rect 16114 16940 16120 16952
rect 16172 16980 16178 16992
rect 18616 16980 18644 17147
rect 22186 17144 22192 17196
rect 22244 17144 22250 17196
rect 22830 17144 22836 17196
rect 22888 17144 22894 17196
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17116 21419 17119
rect 22370 17116 22376 17128
rect 21407 17088 22376 17116
rect 21407 17085 21419 17088
rect 21361 17079 21419 17085
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 22465 17119 22523 17125
rect 22465 17085 22477 17119
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17116 23167 17119
rect 23198 17116 23204 17128
rect 23155 17088 23204 17116
rect 23155 17085 23167 17088
rect 23109 17079 23167 17085
rect 21637 17051 21695 17057
rect 21637 17017 21649 17051
rect 21683 17048 21695 17051
rect 22278 17048 22284 17060
rect 21683 17020 22284 17048
rect 21683 17017 21695 17020
rect 21637 17011 21695 17017
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 22480 17048 22508 17079
rect 23198 17076 23204 17088
rect 23256 17076 23262 17128
rect 23474 17076 23480 17128
rect 23532 17076 23538 17128
rect 24872 17116 24900 17170
rect 25406 17144 25412 17196
rect 25464 17144 25470 17196
rect 25498 17144 25504 17196
rect 25556 17184 25562 17196
rect 25593 17187 25651 17193
rect 25593 17184 25605 17187
rect 25556 17156 25605 17184
rect 25556 17144 25562 17156
rect 25593 17153 25605 17156
rect 25639 17153 25651 17187
rect 25593 17147 25651 17153
rect 24946 17116 24952 17128
rect 24872 17088 24952 17116
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 25700 17116 25728 17224
rect 26237 17221 26249 17224
rect 26283 17221 26295 17255
rect 26528 17252 26556 17292
rect 26789 17289 26801 17292
rect 26835 17320 26847 17323
rect 27890 17320 27896 17332
rect 26835 17292 27896 17320
rect 26835 17289 26847 17292
rect 26789 17283 26847 17289
rect 27890 17280 27896 17292
rect 27948 17280 27954 17332
rect 27522 17252 27528 17264
rect 26237 17215 26295 17221
rect 26344 17224 26556 17252
rect 26712 17224 27528 17252
rect 26344 17193 26372 17224
rect 26712 17196 26740 17224
rect 27522 17212 27528 17224
rect 27580 17212 27586 17264
rect 27706 17212 27712 17264
rect 27764 17252 27770 17264
rect 28261 17255 28319 17261
rect 28261 17252 28273 17255
rect 27764 17224 28273 17252
rect 27764 17212 27770 17224
rect 28261 17221 28273 17224
rect 28307 17221 28319 17255
rect 28261 17215 28319 17221
rect 26053 17187 26111 17193
rect 26053 17153 26065 17187
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17153 26387 17187
rect 26329 17147 26387 17153
rect 26421 17187 26479 17193
rect 26421 17153 26433 17187
rect 26467 17184 26479 17187
rect 26510 17184 26516 17196
rect 26467 17156 26516 17184
rect 26467 17153 26479 17156
rect 26421 17147 26479 17153
rect 25240 17088 25728 17116
rect 26068 17116 26096 17147
rect 26510 17144 26516 17156
rect 26568 17144 26574 17196
rect 26605 17187 26663 17193
rect 26605 17153 26617 17187
rect 26651 17184 26663 17187
rect 26694 17184 26700 17196
rect 26651 17156 26700 17184
rect 26651 17153 26663 17156
rect 26605 17147 26663 17153
rect 26694 17144 26700 17156
rect 26752 17144 26758 17196
rect 26988 17184 27108 17188
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 26804 17160 27169 17184
rect 26804 17156 27016 17160
rect 27080 17156 27169 17160
rect 26804 17116 26832 17156
rect 27157 17153 27169 17156
rect 27203 17184 27215 17187
rect 27617 17187 27675 17193
rect 27203 17156 27568 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27540 17128 27568 17156
rect 27617 17153 27629 17187
rect 27663 17184 27675 17187
rect 27798 17184 27804 17196
rect 27663 17156 27804 17184
rect 27663 17153 27675 17156
rect 27617 17147 27675 17153
rect 27798 17144 27804 17156
rect 27856 17144 27862 17196
rect 27890 17144 27896 17196
rect 27948 17184 27954 17196
rect 28442 17184 28448 17196
rect 27948 17156 28448 17184
rect 27948 17144 27954 17156
rect 28442 17144 28448 17156
rect 28500 17144 28506 17196
rect 26068 17088 26832 17116
rect 22480 17020 23612 17048
rect 23584 16992 23612 17020
rect 16172 16952 18644 16980
rect 16172 16940 16178 16952
rect 23106 16940 23112 16992
rect 23164 16940 23170 16992
rect 23566 16940 23572 16992
rect 23624 16940 23630 16992
rect 24394 16940 24400 16992
rect 24452 16980 24458 16992
rect 25240 16989 25268 17088
rect 27246 17076 27252 17128
rect 27304 17076 27310 17128
rect 27341 17119 27399 17125
rect 27341 17085 27353 17119
rect 27387 17085 27399 17119
rect 27341 17079 27399 17085
rect 25777 17051 25835 17057
rect 25777 17017 25789 17051
rect 25823 17048 25835 17051
rect 26510 17048 26516 17060
rect 25823 17020 26516 17048
rect 25823 17017 25835 17020
rect 25777 17011 25835 17017
rect 26510 17008 26516 17020
rect 26568 17008 26574 17060
rect 26970 17008 26976 17060
rect 27028 17008 27034 17060
rect 27356 17048 27384 17079
rect 27430 17076 27436 17128
rect 27488 17076 27494 17128
rect 27522 17076 27528 17128
rect 27580 17076 27586 17128
rect 28169 17119 28227 17125
rect 28169 17085 28181 17119
rect 28215 17116 28227 17119
rect 28350 17116 28356 17128
rect 28215 17088 28356 17116
rect 28215 17085 28227 17088
rect 28169 17079 28227 17085
rect 28350 17076 28356 17088
rect 28408 17076 28414 17128
rect 27709 17051 27767 17057
rect 27709 17048 27721 17051
rect 27356 17020 27721 17048
rect 27709 17017 27721 17020
rect 27755 17017 27767 17051
rect 27709 17011 27767 17017
rect 25225 16983 25283 16989
rect 25225 16980 25237 16983
rect 24452 16952 25237 16980
rect 24452 16940 24458 16952
rect 25225 16949 25237 16952
rect 25271 16949 25283 16983
rect 25225 16943 25283 16949
rect 26326 16940 26332 16992
rect 26384 16980 26390 16992
rect 26421 16983 26479 16989
rect 26421 16980 26433 16983
rect 26384 16952 26433 16980
rect 26384 16940 26390 16952
rect 26421 16949 26433 16952
rect 26467 16949 26479 16983
rect 26421 16943 26479 16949
rect 26602 16940 26608 16992
rect 26660 16980 26666 16992
rect 27246 16980 27252 16992
rect 26660 16952 27252 16980
rect 26660 16940 26666 16952
rect 27246 16940 27252 16952
rect 27304 16980 27310 16992
rect 28077 16983 28135 16989
rect 28077 16980 28089 16983
rect 27304 16952 28089 16980
rect 27304 16940 27310 16952
rect 28077 16949 28089 16952
rect 28123 16949 28135 16983
rect 28077 16943 28135 16949
rect 28626 16940 28632 16992
rect 28684 16940 28690 16992
rect 1104 16890 29440 16912
rect 1104 16838 4491 16890
rect 4543 16838 4555 16890
rect 4607 16838 4619 16890
rect 4671 16838 4683 16890
rect 4735 16838 4747 16890
rect 4799 16838 11574 16890
rect 11626 16838 11638 16890
rect 11690 16838 11702 16890
rect 11754 16838 11766 16890
rect 11818 16838 11830 16890
rect 11882 16838 18657 16890
rect 18709 16838 18721 16890
rect 18773 16838 18785 16890
rect 18837 16838 18849 16890
rect 18901 16838 18913 16890
rect 18965 16838 25740 16890
rect 25792 16838 25804 16890
rect 25856 16838 25868 16890
rect 25920 16838 25932 16890
rect 25984 16838 25996 16890
rect 26048 16838 29440 16890
rect 1104 16816 29440 16838
rect 3602 16736 3608 16788
rect 3660 16776 3666 16788
rect 5166 16776 5172 16788
rect 3660 16748 5172 16776
rect 3660 16736 3666 16748
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 5592 16748 6285 16776
rect 5592 16736 5598 16748
rect 6273 16745 6285 16748
rect 6319 16745 6331 16779
rect 6273 16739 6331 16745
rect 14642 16736 14648 16788
rect 14700 16736 14706 16788
rect 16942 16736 16948 16788
rect 17000 16776 17006 16788
rect 19150 16776 19156 16788
rect 17000 16748 19156 16776
rect 17000 16736 17006 16748
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 22005 16779 22063 16785
rect 22005 16745 22017 16779
rect 22051 16776 22063 16779
rect 22186 16776 22192 16788
rect 22051 16748 22192 16776
rect 22051 16745 22063 16748
rect 22005 16739 22063 16745
rect 22186 16736 22192 16748
rect 22244 16736 22250 16788
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 22373 16779 22431 16785
rect 22373 16776 22385 16779
rect 22336 16748 22385 16776
rect 22336 16736 22342 16748
rect 22373 16745 22385 16748
rect 22419 16745 22431 16779
rect 22373 16739 22431 16745
rect 22646 16736 22652 16788
rect 22704 16776 22710 16788
rect 22741 16779 22799 16785
rect 22741 16776 22753 16779
rect 22704 16748 22753 16776
rect 22704 16736 22710 16748
rect 22741 16745 22753 16748
rect 22787 16745 22799 16779
rect 22741 16739 22799 16745
rect 3418 16668 3424 16720
rect 3476 16708 3482 16720
rect 4982 16708 4988 16720
rect 3476 16680 4988 16708
rect 3476 16668 3482 16680
rect 4982 16668 4988 16680
rect 5040 16668 5046 16720
rect 7190 16708 7196 16720
rect 5276 16680 7196 16708
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3191 16612 3801 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 5276 16640 5304 16680
rect 7190 16668 7196 16680
rect 7248 16668 7254 16720
rect 10502 16668 10508 16720
rect 10560 16708 10566 16720
rect 16850 16708 16856 16720
rect 10560 16680 16856 16708
rect 10560 16668 10566 16680
rect 16850 16668 16856 16680
rect 16908 16668 16914 16720
rect 3789 16603 3847 16609
rect 4908 16612 5304 16640
rect 4908 16584 4936 16612
rect 1394 16532 1400 16584
rect 1452 16532 1458 16584
rect 4890 16532 4896 16584
rect 4948 16532 4954 16584
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 1670 16464 1676 16516
rect 1728 16464 1734 16516
rect 3878 16504 3884 16516
rect 2898 16476 3884 16504
rect 3878 16464 3884 16476
rect 3936 16464 3942 16516
rect 4430 16396 4436 16448
rect 4488 16396 4494 16448
rect 5000 16436 5028 16535
rect 5074 16532 5080 16584
rect 5132 16532 5138 16584
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16572 5227 16575
rect 5276 16572 5304 16612
rect 5460 16612 7512 16640
rect 5215 16544 5304 16572
rect 5353 16575 5411 16581
rect 5215 16541 5227 16544
rect 5169 16535 5227 16541
rect 5353 16541 5365 16575
rect 5399 16572 5411 16575
rect 5460 16572 5488 16612
rect 7484 16584 7512 16612
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10134 16640 10140 16652
rect 9824 16612 10140 16640
rect 9824 16600 9830 16612
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 10962 16640 10968 16652
rect 10735 16612 10968 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 16960 16640 16988 16736
rect 22756 16708 22784 16739
rect 22830 16736 22836 16788
rect 22888 16776 22894 16788
rect 23109 16779 23167 16785
rect 23109 16776 23121 16779
rect 22888 16748 23121 16776
rect 22888 16736 22894 16748
rect 23109 16745 23121 16748
rect 23155 16745 23167 16779
rect 23382 16776 23388 16788
rect 23109 16739 23167 16745
rect 23216 16748 23388 16776
rect 23216 16708 23244 16748
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 23753 16779 23811 16785
rect 23753 16745 23765 16779
rect 23799 16776 23811 16779
rect 23842 16776 23848 16788
rect 23799 16748 23848 16776
rect 23799 16745 23811 16748
rect 23753 16739 23811 16745
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 24397 16779 24455 16785
rect 24397 16745 24409 16779
rect 24443 16776 24455 16779
rect 25314 16776 25320 16788
rect 24443 16748 25320 16776
rect 24443 16745 24455 16748
rect 24397 16739 24455 16745
rect 25314 16736 25320 16748
rect 25372 16736 25378 16788
rect 26234 16736 26240 16788
rect 26292 16736 26298 16788
rect 26510 16736 26516 16788
rect 26568 16776 26574 16788
rect 27154 16776 27160 16788
rect 26568 16748 27160 16776
rect 26568 16736 26574 16748
rect 27154 16736 27160 16748
rect 27212 16736 27218 16788
rect 27798 16736 27804 16788
rect 27856 16736 27862 16788
rect 22756 16680 23244 16708
rect 23290 16668 23296 16720
rect 23348 16708 23354 16720
rect 23661 16711 23719 16717
rect 23661 16708 23673 16711
rect 23348 16680 23673 16708
rect 23348 16668 23354 16680
rect 23661 16677 23673 16680
rect 23707 16677 23719 16711
rect 26252 16708 26280 16736
rect 23661 16671 23719 16677
rect 24964 16680 27016 16708
rect 14292 16612 14872 16640
rect 5399 16544 5488 16572
rect 5399 16541 5411 16544
rect 5353 16535 5411 16541
rect 5718 16532 5724 16584
rect 5776 16532 5782 16584
rect 7466 16532 7472 16584
rect 7524 16532 7530 16584
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16572 9919 16575
rect 9950 16572 9956 16584
rect 9907 16544 9956 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 10152 16572 10180 16600
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 10152 16544 10241 16572
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 14090 16532 14096 16584
rect 14148 16532 14154 16584
rect 14292 16581 14320 16612
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14461 16575 14519 16581
rect 14461 16541 14473 16575
rect 14507 16572 14519 16575
rect 14734 16572 14740 16584
rect 14507 16544 14740 16572
rect 14507 16541 14519 16544
rect 14461 16535 14519 16541
rect 5092 16504 5120 16532
rect 5253 16507 5311 16513
rect 5253 16504 5265 16507
rect 5092 16476 5265 16504
rect 5253 16473 5265 16476
rect 5299 16473 5311 16507
rect 5253 16467 5311 16473
rect 10045 16507 10103 16513
rect 10045 16473 10057 16507
rect 10091 16473 10103 16507
rect 10045 16467 10103 16473
rect 10137 16507 10195 16513
rect 10137 16473 10149 16507
rect 10183 16504 10195 16507
rect 11241 16507 11299 16513
rect 11241 16504 11253 16507
rect 10183 16476 11253 16504
rect 10183 16473 10195 16476
rect 10137 16467 10195 16473
rect 11241 16473 11253 16476
rect 11287 16473 11299 16507
rect 11241 16467 11299 16473
rect 5074 16436 5080 16448
rect 5000 16408 5080 16436
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5534 16396 5540 16448
rect 5592 16396 5598 16448
rect 10060 16436 10088 16467
rect 14366 16464 14372 16516
rect 14424 16464 14430 16516
rect 10318 16436 10324 16448
rect 10060 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 10410 16396 10416 16448
rect 10468 16396 10474 16448
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 14476 16436 14504 16535
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 14844 16504 14872 16612
rect 15120 16612 16988 16640
rect 14918 16532 14924 16584
rect 14976 16572 14982 16584
rect 15120 16581 15148 16612
rect 22002 16600 22008 16652
rect 22060 16640 22066 16652
rect 22833 16643 22891 16649
rect 22833 16640 22845 16643
rect 22060 16612 22845 16640
rect 22060 16600 22066 16612
rect 22833 16609 22845 16612
rect 22879 16640 22891 16643
rect 23845 16643 23903 16649
rect 22879 16612 23520 16640
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 15105 16575 15163 16581
rect 15105 16572 15117 16575
rect 14976 16544 15117 16572
rect 14976 16532 14982 16544
rect 15105 16541 15117 16544
rect 15151 16541 15163 16575
rect 15105 16535 15163 16541
rect 15197 16575 15255 16581
rect 15197 16541 15209 16575
rect 15243 16541 15255 16575
rect 15197 16535 15255 16541
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16572 15347 16575
rect 15335 16544 15424 16572
rect 15335 16541 15347 16544
rect 15289 16535 15347 16541
rect 15010 16504 15016 16516
rect 14844 16476 15016 16504
rect 15010 16464 15016 16476
rect 15068 16464 15074 16516
rect 15212 16504 15240 16535
rect 15396 16504 15424 16544
rect 15470 16532 15476 16584
rect 15528 16532 15534 16584
rect 22189 16575 22247 16581
rect 22189 16541 22201 16575
rect 22235 16572 22247 16575
rect 22278 16572 22284 16584
rect 22235 16544 22284 16572
rect 22235 16541 22247 16544
rect 22189 16535 22247 16541
rect 22278 16532 22284 16544
rect 22336 16532 22342 16584
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 15654 16504 15660 16516
rect 15212 16476 15332 16504
rect 15396 16476 15660 16504
rect 15304 16448 15332 16476
rect 15654 16464 15660 16476
rect 15712 16504 15718 16516
rect 17126 16504 17132 16516
rect 15712 16476 17132 16504
rect 15712 16464 15718 16476
rect 17126 16464 17132 16476
rect 17184 16464 17190 16516
rect 22480 16504 22508 16535
rect 22738 16532 22744 16584
rect 22796 16532 22802 16584
rect 23201 16575 23259 16581
rect 23201 16541 23213 16575
rect 23247 16572 23259 16575
rect 23247 16544 23336 16572
rect 23247 16541 23259 16544
rect 23201 16535 23259 16541
rect 22480 16476 23244 16504
rect 23216 16448 23244 16476
rect 12216 16408 14504 16436
rect 14829 16439 14887 16445
rect 12216 16396 12222 16408
rect 14829 16405 14841 16439
rect 14875 16436 14887 16439
rect 15102 16436 15108 16448
rect 14875 16408 15108 16436
rect 14875 16405 14887 16408
rect 14829 16399 14887 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 15286 16396 15292 16448
rect 15344 16396 15350 16448
rect 23198 16396 23204 16448
rect 23256 16396 23262 16448
rect 23308 16436 23336 16544
rect 23382 16532 23388 16584
rect 23440 16532 23446 16584
rect 23492 16581 23520 16612
rect 23845 16609 23857 16643
rect 23891 16609 23903 16643
rect 23845 16603 23903 16609
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16541 23627 16575
rect 23860 16572 23888 16603
rect 23934 16572 23940 16584
rect 23860 16544 23940 16572
rect 23569 16535 23627 16541
rect 23400 16504 23428 16532
rect 23584 16504 23612 16535
rect 23934 16532 23940 16544
rect 23992 16532 23998 16584
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16572 24639 16575
rect 24670 16572 24676 16584
rect 24627 16544 24676 16572
rect 24627 16541 24639 16544
rect 24581 16535 24639 16541
rect 24670 16532 24676 16544
rect 24728 16532 24734 16584
rect 24964 16581 24992 16680
rect 25406 16600 25412 16652
rect 25464 16640 25470 16652
rect 25464 16612 25544 16640
rect 25464 16600 25470 16612
rect 25516 16581 25544 16612
rect 25590 16600 25596 16652
rect 25648 16640 25654 16652
rect 26145 16643 26203 16649
rect 25648 16612 25728 16640
rect 25648 16600 25654 16612
rect 25700 16581 25728 16612
rect 26145 16609 26157 16643
rect 26191 16640 26203 16643
rect 26234 16640 26240 16652
rect 26191 16612 26240 16640
rect 26191 16609 26203 16612
rect 26145 16603 26203 16609
rect 26234 16600 26240 16612
rect 26292 16600 26298 16652
rect 26344 16581 26372 16680
rect 26786 16640 26792 16652
rect 26436 16612 26792 16640
rect 26436 16584 26464 16612
rect 26786 16600 26792 16612
rect 26844 16640 26850 16652
rect 26844 16612 26924 16640
rect 26844 16600 26850 16612
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16541 25007 16575
rect 24949 16535 25007 16541
rect 25501 16575 25559 16581
rect 25501 16541 25513 16575
rect 25547 16541 25559 16575
rect 25501 16535 25559 16541
rect 25685 16575 25743 16581
rect 25685 16541 25697 16575
rect 25731 16541 25743 16575
rect 25685 16535 25743 16541
rect 26329 16575 26387 16581
rect 26329 16541 26341 16575
rect 26375 16541 26387 16575
rect 26329 16535 26387 16541
rect 23400 16476 23612 16504
rect 23750 16464 23756 16516
rect 23808 16504 23814 16516
rect 24872 16504 24900 16535
rect 26418 16532 26424 16584
rect 26476 16532 26482 16584
rect 26510 16532 26516 16584
rect 26568 16532 26574 16584
rect 26896 16581 26924 16612
rect 26605 16575 26663 16581
rect 26605 16541 26617 16575
rect 26651 16541 26663 16575
rect 26605 16535 26663 16541
rect 26881 16575 26939 16581
rect 26881 16541 26893 16575
rect 26927 16541 26939 16575
rect 26988 16572 27016 16680
rect 27172 16640 27200 16736
rect 27172 16612 28212 16640
rect 27433 16575 27491 16581
rect 27433 16572 27445 16575
rect 26988 16544 27445 16572
rect 26881 16535 26939 16541
rect 27433 16541 27445 16544
rect 27479 16541 27491 16575
rect 27433 16535 27491 16541
rect 25041 16507 25099 16513
rect 25041 16504 25053 16507
rect 23808 16476 25053 16504
rect 23808 16464 23814 16476
rect 25041 16473 25053 16476
rect 25087 16473 25099 16507
rect 25041 16467 25099 16473
rect 25593 16507 25651 16513
rect 25593 16473 25605 16507
rect 25639 16504 25651 16507
rect 26620 16504 26648 16535
rect 25639 16476 26648 16504
rect 26697 16507 26755 16513
rect 25639 16473 25651 16476
rect 25593 16467 25651 16473
rect 26697 16473 26709 16507
rect 26743 16504 26755 16507
rect 26786 16504 26792 16516
rect 26743 16476 26792 16504
rect 26743 16473 26755 16476
rect 26697 16467 26755 16473
rect 26786 16464 26792 16476
rect 26844 16464 26850 16516
rect 27448 16504 27476 16535
rect 27614 16532 27620 16584
rect 27672 16532 27678 16584
rect 27709 16575 27767 16581
rect 27709 16541 27721 16575
rect 27755 16572 27767 16575
rect 27755 16544 28028 16572
rect 27755 16541 27767 16544
rect 27709 16535 27767 16541
rect 27801 16507 27859 16513
rect 27801 16504 27813 16507
rect 26988 16476 27384 16504
rect 27448 16476 27813 16504
rect 24765 16439 24823 16445
rect 24765 16436 24777 16439
rect 23308 16408 24777 16436
rect 24765 16405 24777 16408
rect 24811 16436 24823 16439
rect 26988 16436 27016 16476
rect 24811 16408 27016 16436
rect 27065 16439 27123 16445
rect 24811 16405 24823 16408
rect 24765 16399 24823 16405
rect 27065 16405 27077 16439
rect 27111 16436 27123 16439
rect 27154 16436 27160 16448
rect 27111 16408 27160 16436
rect 27111 16405 27123 16408
rect 27065 16399 27123 16405
rect 27154 16396 27160 16408
rect 27212 16396 27218 16448
rect 27246 16396 27252 16448
rect 27304 16396 27310 16448
rect 27356 16436 27384 16476
rect 27801 16473 27813 16476
rect 27847 16473 27859 16507
rect 28000 16504 28028 16544
rect 28074 16532 28080 16584
rect 28132 16532 28138 16584
rect 28184 16581 28212 16612
rect 28169 16575 28227 16581
rect 28169 16541 28181 16575
rect 28215 16541 28227 16575
rect 28169 16535 28227 16541
rect 28350 16532 28356 16584
rect 28408 16581 28414 16584
rect 28408 16572 28419 16581
rect 28408 16544 28453 16572
rect 28408 16535 28419 16544
rect 28408 16532 28414 16535
rect 28626 16532 28632 16584
rect 28684 16532 28690 16584
rect 28261 16507 28319 16513
rect 28261 16504 28273 16507
rect 28000 16476 28273 16504
rect 27801 16467 27859 16473
rect 28261 16473 28273 16476
rect 28307 16473 28319 16507
rect 28261 16467 28319 16473
rect 27985 16439 28043 16445
rect 27985 16436 27997 16439
rect 27356 16408 27997 16436
rect 27985 16405 27997 16408
rect 28031 16436 28043 16439
rect 28644 16436 28672 16532
rect 28031 16408 28672 16436
rect 28031 16405 28043 16408
rect 27985 16399 28043 16405
rect 1104 16346 29440 16368
rect 1104 16294 5151 16346
rect 5203 16294 5215 16346
rect 5267 16294 5279 16346
rect 5331 16294 5343 16346
rect 5395 16294 5407 16346
rect 5459 16294 12234 16346
rect 12286 16294 12298 16346
rect 12350 16294 12362 16346
rect 12414 16294 12426 16346
rect 12478 16294 12490 16346
rect 12542 16294 19317 16346
rect 19369 16294 19381 16346
rect 19433 16294 19445 16346
rect 19497 16294 19509 16346
rect 19561 16294 19573 16346
rect 19625 16294 26400 16346
rect 26452 16294 26464 16346
rect 26516 16294 26528 16346
rect 26580 16294 26592 16346
rect 26644 16294 26656 16346
rect 26708 16294 29440 16346
rect 1104 16272 29440 16294
rect 1397 16235 1455 16241
rect 1397 16201 1409 16235
rect 1443 16232 1455 16235
rect 1670 16232 1676 16244
rect 1443 16204 1676 16232
rect 1443 16201 1455 16204
rect 1397 16195 1455 16201
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 4430 16232 4436 16244
rect 2792 16204 4436 16232
rect 2792 16173 2820 16204
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 4982 16192 4988 16244
rect 5040 16192 5046 16244
rect 5074 16192 5080 16244
rect 5132 16232 5138 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5132 16204 6193 16232
rect 5132 16192 5138 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6181 16195 6239 16201
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 7432 16204 9536 16232
rect 7432 16192 7438 16204
rect 2777 16167 2835 16173
rect 2777 16133 2789 16167
rect 2823 16133 2835 16167
rect 2777 16127 2835 16133
rect 5736 16136 6500 16164
rect 5736 16108 5764 16136
rect 934 16056 940 16108
rect 992 16096 998 16108
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 992 16068 1593 16096
rect 992 16056 998 16068
rect 1581 16065 1593 16068
rect 1627 16065 1639 16099
rect 1581 16059 1639 16065
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 5166 16096 5172 16108
rect 3936 16068 5172 16096
rect 3936 16056 3942 16068
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 5718 16056 5724 16108
rect 5776 16056 5782 16108
rect 5902 16056 5908 16108
rect 5960 16096 5966 16108
rect 6472 16105 6500 16136
rect 6546 16124 6552 16176
rect 6604 16164 6610 16176
rect 9309 16167 9367 16173
rect 9309 16164 9321 16167
rect 6604 16136 6914 16164
rect 6604 16124 6610 16136
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 5960 16068 6377 16096
rect 5960 16056 5966 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 6458 16099 6516 16105
rect 6458 16065 6470 16099
rect 6504 16065 6516 16099
rect 6458 16059 6516 16065
rect 6638 16056 6644 16108
rect 6696 16056 6702 16108
rect 6886 16105 6914 16136
rect 7116 16136 9321 16164
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 6871 16099 6929 16105
rect 6871 16065 6883 16099
rect 6917 16096 6929 16099
rect 7006 16096 7012 16108
rect 6917 16068 7012 16096
rect 6917 16065 6929 16068
rect 6871 16059 6929 16065
rect 1394 15988 1400 16040
rect 1452 16028 1458 16040
rect 2501 16031 2559 16037
rect 2501 16028 2513 16031
rect 1452 16000 2513 16028
rect 1452 15988 1458 16000
rect 2501 15997 2513 16000
rect 2547 15997 2559 16031
rect 2501 15991 2559 15997
rect 4433 16031 4491 16037
rect 4433 15997 4445 16031
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 4338 15920 4344 15972
rect 4396 15960 4402 15972
rect 4448 15960 4476 15991
rect 5626 15988 5632 16040
rect 5684 15988 5690 16040
rect 6748 15960 6776 16059
rect 7006 16056 7012 16068
rect 7064 16056 7070 16108
rect 7116 16105 7144 16136
rect 9309 16133 9321 16136
rect 9355 16133 9367 16167
rect 9309 16127 9367 16133
rect 9508 16108 9536 16204
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 11330 16232 11336 16244
rect 10008 16204 11336 16232
rect 10008 16192 10014 16204
rect 10042 16124 10048 16176
rect 10100 16124 10106 16176
rect 10152 16173 10180 16204
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 17954 16232 17960 16244
rect 12360 16204 17960 16232
rect 10137 16167 10195 16173
rect 10137 16133 10149 16167
rect 10183 16133 10195 16167
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 10137 16127 10195 16133
rect 10428 16136 12173 16164
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 7248 16068 7297 16096
rect 7248 16056 7254 16068
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7374 16056 7380 16108
rect 7432 16056 7438 16108
rect 7466 16056 7472 16108
rect 7524 16056 7530 16108
rect 7926 16056 7932 16108
rect 7984 16056 7990 16108
rect 8110 16056 8116 16108
rect 8168 16096 8174 16108
rect 8297 16099 8355 16105
rect 8297 16096 8309 16099
rect 8168 16068 8309 16096
rect 8168 16056 8174 16068
rect 8297 16065 8309 16068
rect 8343 16065 8355 16099
rect 8297 16059 8355 16065
rect 9490 16056 9496 16108
rect 9548 16056 9554 16108
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 4396 15932 6776 15960
rect 6932 16000 8616 16028
rect 4396 15920 4402 15932
rect 4249 15895 4307 15901
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 6932 15892 6960 16000
rect 7009 15963 7067 15969
rect 7009 15929 7021 15963
rect 7055 15960 7067 15963
rect 8294 15960 8300 15972
rect 7055 15932 8300 15960
rect 7055 15929 7067 15932
rect 7009 15923 7067 15929
rect 8294 15920 8300 15932
rect 8352 15920 8358 15972
rect 8588 15960 8616 16000
rect 8662 15988 8668 16040
rect 8720 15988 8726 16040
rect 9876 16028 9904 16059
rect 10226 16056 10232 16108
rect 10284 16056 10290 16108
rect 10428 16028 10456 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 12161 16127 12219 16133
rect 12360 16096 12388 16204
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 22830 16192 22836 16244
rect 22888 16232 22894 16244
rect 26786 16232 26792 16244
rect 22888 16204 26792 16232
rect 22888 16192 22894 16204
rect 12894 16124 12900 16176
rect 12952 16164 12958 16176
rect 13265 16167 13323 16173
rect 12952 16136 13216 16164
rect 12952 16124 12958 16136
rect 13188 16108 13216 16136
rect 13265 16133 13277 16167
rect 13311 16164 13323 16167
rect 13311 16136 13952 16164
rect 13311 16133 13323 16136
rect 13265 16127 13323 16133
rect 13924 16108 13952 16136
rect 14090 16124 14096 16176
rect 14148 16164 14154 16176
rect 14918 16164 14924 16176
rect 14148 16136 14924 16164
rect 14148 16124 14154 16136
rect 14918 16124 14924 16136
rect 14976 16164 14982 16176
rect 16025 16167 16083 16173
rect 16025 16164 16037 16167
rect 14976 16136 16037 16164
rect 14976 16124 14982 16136
rect 16025 16133 16037 16136
rect 16071 16133 16083 16167
rect 16025 16127 16083 16133
rect 23198 16124 23204 16176
rect 23256 16164 23262 16176
rect 23293 16167 23351 16173
rect 23293 16164 23305 16167
rect 23256 16136 23305 16164
rect 23256 16124 23262 16136
rect 23293 16133 23305 16136
rect 23339 16133 23351 16167
rect 23293 16127 23351 16133
rect 25406 16124 25412 16176
rect 25464 16124 25470 16176
rect 10520 16068 12388 16096
rect 10520 16037 10548 16068
rect 12986 16056 12992 16108
rect 13044 16056 13050 16108
rect 13170 16056 13176 16108
rect 13228 16056 13234 16108
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16096 13415 16099
rect 13446 16096 13452 16108
rect 13403 16068 13452 16096
rect 13403 16065 13415 16068
rect 13357 16059 13415 16065
rect 13446 16056 13452 16068
rect 13504 16056 13510 16108
rect 13906 16056 13912 16108
rect 13964 16056 13970 16108
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15703 16068 15761 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15838 16056 15844 16108
rect 15896 16096 15902 16108
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 15896 16068 15945 16096
rect 15896 16056 15902 16068
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 16114 16056 16120 16108
rect 16172 16096 16178 16108
rect 17034 16096 17040 16108
rect 16172 16068 17040 16096
rect 16172 16056 16178 16068
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23934 16096 23940 16108
rect 23523 16068 23940 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 23934 16056 23940 16068
rect 23992 16056 23998 16108
rect 9876 16000 10456 16028
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 10520 15960 10548 15991
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 10928 16000 11529 16028
rect 10928 15988 10934 16000
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 16028 15163 16031
rect 15286 16028 15292 16040
rect 15151 16000 15292 16028
rect 15151 15997 15163 16000
rect 15105 15991 15163 15997
rect 15286 15988 15292 16000
rect 15344 16028 15350 16040
rect 25424 16028 25452 16124
rect 25700 16105 25728 16204
rect 26786 16192 26792 16204
rect 26844 16192 26850 16244
rect 25685 16099 25743 16105
rect 25685 16065 25697 16099
rect 25731 16065 25743 16099
rect 25685 16059 25743 16065
rect 25869 16099 25927 16105
rect 25869 16065 25881 16099
rect 25915 16096 25927 16099
rect 26326 16096 26332 16108
rect 25915 16068 26332 16096
rect 25915 16065 25927 16068
rect 25869 16059 25927 16065
rect 25884 16028 25912 16059
rect 26326 16056 26332 16068
rect 26384 16056 26390 16108
rect 27522 16028 27528 16040
rect 15344 16000 16160 16028
rect 25424 16000 25912 16028
rect 25976 16000 27528 16028
rect 15344 15988 15350 16000
rect 8588 15932 10548 15960
rect 13464 15932 16068 15960
rect 4295 15864 6960 15892
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 7650 15852 7656 15904
rect 7708 15852 7714 15904
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 10008 15864 10425 15892
rect 10008 15852 10014 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 13464 15892 13492 15932
rect 16040 15904 16068 15932
rect 16132 15904 16160 16000
rect 23290 15920 23296 15972
rect 23348 15960 23354 15972
rect 23658 15960 23664 15972
rect 23348 15932 23664 15960
rect 23348 15920 23354 15932
rect 23658 15920 23664 15932
rect 23716 15960 23722 15972
rect 25976 15960 26004 16000
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 23716 15932 26004 15960
rect 23716 15920 23722 15932
rect 26234 15920 26240 15972
rect 26292 15960 26298 15972
rect 26786 15960 26792 15972
rect 26292 15932 26792 15960
rect 26292 15920 26298 15932
rect 26786 15920 26792 15932
rect 26844 15920 26850 15972
rect 11195 15864 13492 15892
rect 13541 15895 13599 15901
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 13541 15861 13553 15895
rect 13587 15892 13599 15895
rect 13814 15892 13820 15904
rect 13587 15864 13820 15892
rect 13587 15861 13599 15864
rect 13541 15855 13599 15861
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 15654 15892 15660 15904
rect 15344 15864 15660 15892
rect 15344 15852 15350 15864
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 16022 15852 16028 15904
rect 16080 15852 16086 15904
rect 16114 15852 16120 15904
rect 16172 15852 16178 15904
rect 16298 15852 16304 15904
rect 16356 15852 16362 15904
rect 25777 15895 25835 15901
rect 25777 15861 25789 15895
rect 25823 15892 25835 15895
rect 26142 15892 26148 15904
rect 25823 15864 26148 15892
rect 25823 15861 25835 15864
rect 25777 15855 25835 15861
rect 26142 15852 26148 15864
rect 26200 15852 26206 15904
rect 1104 15802 29440 15824
rect 1104 15750 4491 15802
rect 4543 15750 4555 15802
rect 4607 15750 4619 15802
rect 4671 15750 4683 15802
rect 4735 15750 4747 15802
rect 4799 15750 11574 15802
rect 11626 15750 11638 15802
rect 11690 15750 11702 15802
rect 11754 15750 11766 15802
rect 11818 15750 11830 15802
rect 11882 15750 18657 15802
rect 18709 15750 18721 15802
rect 18773 15750 18785 15802
rect 18837 15750 18849 15802
rect 18901 15750 18913 15802
rect 18965 15750 25740 15802
rect 25792 15750 25804 15802
rect 25856 15750 25868 15802
rect 25920 15750 25932 15802
rect 25984 15750 25996 15802
rect 26048 15750 29440 15802
rect 1104 15728 29440 15750
rect 3605 15691 3663 15697
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 4338 15688 4344 15700
rect 3651 15660 4344 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 5997 15691 6055 15697
rect 5997 15688 6009 15691
rect 5776 15660 6009 15688
rect 5776 15648 5782 15660
rect 5997 15657 6009 15660
rect 6043 15657 6055 15691
rect 7926 15688 7932 15700
rect 5997 15651 6055 15657
rect 6380 15660 7932 15688
rect 5810 15580 5816 15632
rect 5868 15580 5874 15632
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 1857 15555 1915 15561
rect 1857 15552 1869 15555
rect 1452 15524 1869 15552
rect 1452 15512 1458 15524
rect 1857 15521 1869 15524
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 3326 15552 3332 15564
rect 2179 15524 3332 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 5828 15552 5856 15580
rect 4571 15524 5856 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 3234 15444 3240 15496
rect 3292 15484 3298 15496
rect 3878 15484 3884 15496
rect 3292 15456 3884 15484
rect 3292 15444 3298 15456
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4172 15456 4261 15484
rect 4172 15360 4200 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 6086 15484 6092 15496
rect 5658 15456 6092 15484
rect 4249 15447 4307 15453
rect 6086 15444 6092 15456
rect 6144 15484 6150 15496
rect 6380 15484 6408 15660
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 8389 15691 8447 15697
rect 8389 15657 8401 15691
rect 8435 15688 8447 15691
rect 8662 15688 8668 15700
rect 8435 15660 8668 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 9480 15691 9538 15697
rect 9480 15657 9492 15691
rect 9526 15688 9538 15691
rect 9950 15688 9956 15700
rect 9526 15660 9956 15688
rect 9526 15657 9538 15660
rect 9480 15651 9538 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10870 15648 10876 15700
rect 10928 15688 10934 15700
rect 10965 15691 11023 15697
rect 10965 15688 10977 15691
rect 10928 15660 10977 15688
rect 10928 15648 10934 15660
rect 10965 15657 10977 15660
rect 11011 15657 11023 15691
rect 15010 15688 15016 15700
rect 10965 15651 11023 15657
rect 12176 15660 15016 15688
rect 12176 15620 12204 15660
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 16114 15648 16120 15700
rect 16172 15648 16178 15700
rect 16298 15648 16304 15700
rect 16356 15648 16362 15700
rect 23566 15648 23572 15700
rect 23624 15648 23630 15700
rect 24026 15648 24032 15700
rect 24084 15688 24090 15700
rect 24946 15688 24952 15700
rect 24084 15660 24952 15688
rect 24084 15648 24090 15660
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 26142 15648 26148 15700
rect 26200 15688 26206 15700
rect 26237 15691 26295 15697
rect 26237 15688 26249 15691
rect 26200 15660 26249 15688
rect 26200 15648 26206 15660
rect 26237 15657 26249 15660
rect 26283 15657 26295 15691
rect 26237 15651 26295 15657
rect 26694 15648 26700 15700
rect 26752 15688 26758 15700
rect 26973 15691 27031 15697
rect 26973 15688 26985 15691
rect 26752 15660 26985 15688
rect 26752 15648 26758 15660
rect 26973 15657 26985 15660
rect 27019 15688 27031 15691
rect 27154 15688 27160 15700
rect 27019 15660 27160 15688
rect 27019 15657 27031 15660
rect 26973 15651 27031 15657
rect 27154 15648 27160 15660
rect 27212 15688 27218 15700
rect 27614 15688 27620 15700
rect 27212 15660 27620 15688
rect 27212 15648 27218 15660
rect 27614 15648 27620 15660
rect 27672 15648 27678 15700
rect 11164 15592 12204 15620
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15552 6975 15555
rect 7650 15552 7656 15564
rect 6963 15524 7656 15552
rect 6963 15521 6975 15524
rect 6917 15515 6975 15521
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 8110 15552 8116 15564
rect 8036 15524 8116 15552
rect 6144 15456 6408 15484
rect 6144 15444 6150 15456
rect 6546 15444 6552 15496
rect 6604 15484 6610 15496
rect 6641 15487 6699 15493
rect 6641 15484 6653 15487
rect 6604 15456 6653 15484
rect 6604 15444 6610 15456
rect 6641 15453 6653 15456
rect 6687 15453 6699 15487
rect 8036 15470 8064 15524
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 9490 15512 9496 15564
rect 9548 15552 9554 15564
rect 10502 15552 10508 15564
rect 9548 15524 10508 15552
rect 9548 15512 9554 15524
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 6641 15447 6699 15453
rect 9214 15444 9220 15496
rect 9272 15444 9278 15496
rect 10042 15376 10048 15428
rect 10100 15376 10106 15428
rect 4154 15308 4160 15360
rect 4212 15308 4218 15360
rect 5166 15308 5172 15360
rect 5224 15348 5230 15360
rect 5810 15348 5816 15360
rect 5224 15320 5816 15348
rect 5224 15308 5230 15320
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 11164 15348 11192 15592
rect 11882 15444 11888 15496
rect 11940 15444 11946 15496
rect 12176 15494 12204 15592
rect 12342 15512 12348 15564
rect 12400 15552 12406 15564
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 12400 15524 13185 15552
rect 12400 15512 12406 15524
rect 13173 15521 13185 15524
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 14366 15512 14372 15564
rect 14424 15512 14430 15564
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15552 14703 15555
rect 16316 15552 16344 15648
rect 18785 15623 18843 15629
rect 18785 15589 18797 15623
rect 18831 15620 18843 15623
rect 19058 15620 19064 15632
rect 18831 15592 19064 15620
rect 18831 15589 18843 15592
rect 18785 15583 18843 15589
rect 19058 15580 19064 15592
rect 19116 15620 19122 15632
rect 23201 15623 23259 15629
rect 19116 15592 20208 15620
rect 19116 15580 19122 15592
rect 14691 15524 16344 15552
rect 16485 15555 16543 15561
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 16485 15521 16497 15555
rect 16531 15552 16543 15555
rect 17402 15552 17408 15564
rect 16531 15524 17408 15552
rect 16531 15521 16543 15524
rect 16485 15515 16543 15521
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18693 15555 18751 15561
rect 18693 15552 18705 15555
rect 18012 15524 18705 15552
rect 18012 15512 18018 15524
rect 18693 15521 18705 15524
rect 18739 15521 18751 15555
rect 18693 15515 18751 15521
rect 19720 15524 20024 15552
rect 12084 15493 12204 15494
rect 12069 15487 12204 15493
rect 12069 15453 12081 15487
rect 12115 15466 12204 15487
rect 12115 15453 12127 15466
rect 12069 15447 12127 15453
rect 12250 15444 12256 15496
rect 12308 15444 12314 15496
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13906 15484 13912 15496
rect 13403 15456 13912 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 11330 15376 11336 15428
rect 11388 15416 11394 15428
rect 11790 15416 11796 15428
rect 11388 15388 11796 15416
rect 11388 15376 11394 15388
rect 11790 15376 11796 15388
rect 11848 15416 11854 15428
rect 12161 15419 12219 15425
rect 12161 15416 12173 15419
rect 11848 15388 12173 15416
rect 11848 15376 11854 15388
rect 12161 15385 12173 15388
rect 12207 15385 12219 15419
rect 12161 15379 12219 15385
rect 7248 15320 11192 15348
rect 7248 15308 7254 15320
rect 11238 15308 11244 15360
rect 11296 15348 11302 15360
rect 12268 15348 12296 15444
rect 12636 15416 12664 15447
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 19720 15493 19748 15524
rect 18417 15487 18475 15493
rect 18417 15484 18429 15487
rect 18196 15456 18429 15484
rect 18196 15444 18202 15456
rect 18417 15453 18429 15456
rect 18463 15453 18475 15487
rect 18417 15447 18475 15453
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19659 15456 19717 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19794 15444 19800 15496
rect 19852 15444 19858 15496
rect 19996 15493 20024 15524
rect 20180 15493 20208 15592
rect 23201 15589 23213 15623
rect 23247 15620 23259 15623
rect 23290 15620 23296 15632
rect 23247 15592 23296 15620
rect 23247 15589 23259 15592
rect 23201 15583 23259 15589
rect 23290 15580 23296 15592
rect 23348 15580 23354 15632
rect 23676 15592 24716 15620
rect 22278 15512 22284 15564
rect 22336 15552 22342 15564
rect 22336 15524 23428 15552
rect 22336 15512 22342 15524
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15453 19947 15487
rect 19889 15447 19947 15453
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 12986 15416 12992 15428
rect 12636 15388 12992 15416
rect 12986 15376 12992 15388
rect 13044 15416 13050 15428
rect 13044 15388 13400 15416
rect 13044 15376 13050 15388
rect 13372 15360 13400 15388
rect 15654 15376 15660 15428
rect 15712 15376 15718 15428
rect 16022 15376 16028 15428
rect 16080 15416 16086 15428
rect 16761 15419 16819 15425
rect 16761 15416 16773 15419
rect 16080 15388 16773 15416
rect 16080 15376 16086 15388
rect 16761 15385 16773 15388
rect 16807 15385 16819 15419
rect 16761 15379 16819 15385
rect 16850 15376 16856 15428
rect 16908 15376 16914 15428
rect 17218 15376 17224 15428
rect 17276 15376 17282 15428
rect 18506 15416 18512 15428
rect 18064 15388 18512 15416
rect 11296 15320 12296 15348
rect 12437 15351 12495 15357
rect 11296 15308 11302 15320
rect 12437 15317 12449 15351
rect 12483 15348 12495 15351
rect 12618 15348 12624 15360
rect 12483 15320 12624 15348
rect 12483 15317 12495 15320
rect 12437 15311 12495 15317
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 13354 15308 13360 15360
rect 13412 15308 13418 15360
rect 13538 15308 13544 15360
rect 13596 15348 13602 15360
rect 13909 15351 13967 15357
rect 13909 15348 13921 15351
rect 13596 15320 13921 15348
rect 13596 15308 13602 15320
rect 13909 15317 13921 15320
rect 13955 15317 13967 15351
rect 16868 15348 16896 15376
rect 18064 15348 18092 15388
rect 18506 15376 18512 15388
rect 18564 15416 18570 15428
rect 19245 15419 19303 15425
rect 19245 15416 19257 15419
rect 18564 15388 19257 15416
rect 18564 15376 18570 15388
rect 19245 15385 19257 15388
rect 19291 15385 19303 15419
rect 19245 15379 19303 15385
rect 19429 15419 19487 15425
rect 19429 15385 19441 15419
rect 19475 15416 19487 15419
rect 19904 15416 19932 15447
rect 23198 15444 23204 15496
rect 23256 15444 23262 15496
rect 23400 15493 23428 15524
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15484 23443 15487
rect 23676 15484 23704 15592
rect 24688 15564 24716 15592
rect 24762 15580 24768 15632
rect 24820 15620 24826 15632
rect 26513 15623 26571 15629
rect 26513 15620 26525 15623
rect 24820 15592 26525 15620
rect 24820 15580 24826 15592
rect 26513 15589 26525 15592
rect 26559 15589 26571 15623
rect 27430 15620 27436 15632
rect 26513 15583 26571 15589
rect 26620 15592 27436 15620
rect 23750 15512 23756 15564
rect 23808 15512 23814 15564
rect 24026 15512 24032 15564
rect 24084 15512 24090 15564
rect 24670 15512 24676 15564
rect 24728 15552 24734 15564
rect 26620 15552 26648 15592
rect 27430 15580 27436 15592
rect 27488 15580 27494 15632
rect 24728 15524 26648 15552
rect 27160 15560 27218 15561
rect 27160 15555 27384 15560
rect 24728 15512 24734 15524
rect 23431 15456 23704 15484
rect 23845 15487 23903 15493
rect 23431 15453 23443 15456
rect 23385 15447 23443 15453
rect 23845 15453 23857 15487
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 23860 15416 23888 15447
rect 23934 15444 23940 15496
rect 23992 15484 23998 15496
rect 23992 15456 24716 15484
rect 23992 15444 23998 15456
rect 24210 15416 24216 15428
rect 19475 15388 19840 15416
rect 19904 15388 24216 15416
rect 19475 15385 19487 15388
rect 19429 15379 19487 15385
rect 16868 15320 18092 15348
rect 13909 15311 13967 15317
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 18196 15320 18245 15348
rect 18196 15308 18202 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 19812 15348 19840 15388
rect 24210 15376 24216 15388
rect 24268 15376 24274 15428
rect 19978 15348 19984 15360
rect 19812 15320 19984 15348
rect 18233 15311 18291 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20070 15308 20076 15360
rect 20128 15308 20134 15360
rect 24688 15348 24716 15456
rect 24854 15376 24860 15428
rect 24912 15416 24918 15428
rect 25222 15416 25228 15428
rect 24912 15388 25228 15416
rect 24912 15376 24918 15388
rect 25222 15376 25228 15388
rect 25280 15376 25286 15428
rect 26068 15425 26096 15524
rect 27160 15521 27172 15555
rect 27206 15552 27384 15555
rect 27706 15552 27712 15564
rect 27206 15532 27712 15552
rect 27206 15521 27218 15532
rect 27356 15524 27712 15532
rect 27160 15515 27218 15521
rect 27706 15512 27712 15524
rect 27764 15512 27770 15564
rect 26694 15484 26700 15496
rect 26284 15459 26700 15484
rect 26283 15456 26700 15459
rect 26283 15453 26341 15456
rect 26053 15419 26111 15425
rect 26053 15385 26065 15419
rect 26099 15385 26111 15419
rect 26283 15419 26295 15453
rect 26329 15419 26341 15453
rect 26694 15444 26700 15456
rect 26752 15444 26758 15496
rect 26786 15444 26792 15496
rect 26844 15444 26850 15496
rect 26881 15487 26939 15493
rect 26881 15453 26893 15487
rect 26927 15453 26939 15487
rect 26881 15447 26939 15453
rect 26283 15413 26341 15419
rect 26513 15419 26571 15425
rect 26053 15379 26111 15385
rect 26513 15385 26525 15419
rect 26559 15385 26571 15419
rect 26896 15416 26924 15447
rect 27246 15444 27252 15496
rect 27304 15444 27310 15496
rect 27338 15444 27344 15496
rect 27396 15444 27402 15496
rect 27433 15487 27491 15493
rect 27433 15453 27445 15487
rect 27479 15453 27491 15487
rect 27433 15447 27491 15453
rect 27356 15416 27384 15444
rect 26896 15388 27384 15416
rect 27448 15416 27476 15447
rect 27890 15416 27896 15428
rect 27448 15388 27896 15416
rect 26513 15379 26571 15385
rect 26326 15348 26332 15360
rect 24688 15320 26332 15348
rect 26326 15308 26332 15320
rect 26384 15308 26390 15360
rect 26421 15351 26479 15357
rect 26421 15317 26433 15351
rect 26467 15348 26479 15351
rect 26528 15348 26556 15379
rect 27890 15376 27896 15388
rect 27948 15376 27954 15428
rect 26467 15320 26556 15348
rect 26467 15317 26479 15320
rect 26421 15311 26479 15317
rect 26602 15308 26608 15360
rect 26660 15348 26666 15360
rect 26697 15351 26755 15357
rect 26697 15348 26709 15351
rect 26660 15320 26709 15348
rect 26660 15308 26666 15320
rect 26697 15317 26709 15320
rect 26743 15317 26755 15351
rect 26697 15311 26755 15317
rect 26970 15308 26976 15360
rect 27028 15348 27034 15360
rect 27157 15351 27215 15357
rect 27157 15348 27169 15351
rect 27028 15320 27169 15348
rect 27028 15308 27034 15320
rect 27157 15317 27169 15320
rect 27203 15317 27215 15351
rect 27157 15311 27215 15317
rect 27246 15308 27252 15360
rect 27304 15348 27310 15360
rect 27341 15351 27399 15357
rect 27341 15348 27353 15351
rect 27304 15320 27353 15348
rect 27304 15308 27310 15320
rect 27341 15317 27353 15320
rect 27387 15317 27399 15351
rect 27341 15311 27399 15317
rect 1104 15258 29440 15280
rect 1104 15206 5151 15258
rect 5203 15206 5215 15258
rect 5267 15206 5279 15258
rect 5331 15206 5343 15258
rect 5395 15206 5407 15258
rect 5459 15206 12234 15258
rect 12286 15206 12298 15258
rect 12350 15206 12362 15258
rect 12414 15206 12426 15258
rect 12478 15206 12490 15258
rect 12542 15206 19317 15258
rect 19369 15206 19381 15258
rect 19433 15206 19445 15258
rect 19497 15206 19509 15258
rect 19561 15206 19573 15258
rect 19625 15206 26400 15258
rect 26452 15206 26464 15258
rect 26516 15206 26528 15258
rect 26580 15206 26592 15258
rect 26644 15206 26656 15258
rect 26708 15206 29440 15258
rect 1104 15184 29440 15206
rect 4154 15144 4160 15156
rect 4080 15116 4160 15144
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 4080 14949 4108 15116
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 5350 15144 5356 15156
rect 4356 15116 5356 15144
rect 4356 15085 4384 15116
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5684 15116 5825 15144
rect 5684 15104 5690 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 5813 15107 5871 15113
rect 5920 15116 8156 15144
rect 4341 15079 4399 15085
rect 4341 15045 4353 15079
rect 4387 15045 4399 15079
rect 5920 15076 5948 15116
rect 8128 15088 8156 15116
rect 8662 15104 8668 15156
rect 8720 15104 8726 15156
rect 9398 15104 9404 15156
rect 9456 15104 9462 15156
rect 10410 15144 10416 15156
rect 9508 15116 10416 15144
rect 8110 15076 8116 15088
rect 5566 15048 5948 15076
rect 8050 15048 8116 15076
rect 4341 15039 4399 15045
rect 5828 15020 5856 15048
rect 8110 15036 8116 15048
rect 8168 15036 8174 15088
rect 8202 15036 8208 15088
rect 8260 15076 8266 15088
rect 8680 15076 8708 15104
rect 8757 15079 8815 15085
rect 8757 15076 8769 15079
rect 8260 15048 8616 15076
rect 8680 15048 8769 15076
rect 8260 15036 8266 15048
rect 5810 14968 5816 15020
rect 5868 14968 5874 15020
rect 8294 14968 8300 15020
rect 8352 15008 8358 15020
rect 8389 15011 8447 15017
rect 8389 15008 8401 15011
rect 8352 14980 8401 15008
rect 8352 14968 8358 14980
rect 8389 14977 8401 14980
rect 8435 14977 8447 15011
rect 8389 14971 8447 14977
rect 8482 15011 8540 15017
rect 8482 14977 8494 15011
rect 8528 14977 8540 15011
rect 8588 15008 8616 15048
rect 8757 15045 8769 15048
rect 8803 15045 8815 15079
rect 9416 15076 9444 15104
rect 9508 15085 9536 15116
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 11514 15104 11520 15156
rect 11572 15144 11578 15156
rect 12158 15144 12164 15156
rect 11572 15116 12164 15144
rect 11572 15104 11578 15116
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 12618 15144 12624 15156
rect 12452 15116 12624 15144
rect 8757 15039 8815 15045
rect 9232 15048 9444 15076
rect 9493 15079 9551 15085
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 8588 14980 8677 15008
rect 8482 14971 8540 14977
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 8895 15011 8953 15017
rect 8895 14977 8907 15011
rect 8941 15008 8953 15011
rect 9232 15008 9260 15048
rect 9493 15045 9505 15079
rect 9539 15045 9551 15079
rect 9493 15039 9551 15045
rect 10042 15036 10048 15088
rect 10100 15036 10106 15088
rect 12342 15076 12348 15088
rect 11440 15048 12348 15076
rect 8941 14980 9260 15008
rect 8941 14977 8953 14980
rect 8895 14971 8953 14977
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 1452 14912 4077 14940
rect 1452 14900 1458 14912
rect 4065 14909 4077 14912
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 6546 14940 6552 14952
rect 5592 14912 6552 14940
rect 5592 14900 5598 14912
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 8497 14940 8525 14971
rect 8312 14912 8525 14940
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 8312 14813 8340 14912
rect 9214 14900 9220 14952
rect 9272 14900 9278 14952
rect 11440 14940 11468 15048
rect 12342 15036 12348 15048
rect 12400 15036 12406 15088
rect 12452 15085 12480 15116
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 12728 15116 13768 15144
rect 12437 15079 12495 15085
rect 12437 15045 12449 15079
rect 12483 15045 12495 15079
rect 12437 15039 12495 15045
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 12728 15076 12756 15116
rect 12584 15048 12756 15076
rect 13740 15076 13768 15116
rect 13906 15104 13912 15156
rect 13964 15104 13970 15156
rect 15470 15144 15476 15156
rect 14016 15116 15476 15144
rect 14016 15076 14044 15116
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 15654 15104 15660 15156
rect 15712 15144 15718 15156
rect 15712 15116 15884 15144
rect 15712 15104 15718 15116
rect 13740 15048 14044 15076
rect 12584 15036 12590 15048
rect 11514 14968 11520 15020
rect 11572 14968 11578 15020
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 9324 14912 11468 14940
rect 11716 14940 11744 14971
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 12066 15008 12072 15020
rect 11931 14980 12072 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 12066 14968 12072 14980
rect 12124 14968 12130 15020
rect 13538 14968 13544 15020
rect 13596 14968 13602 15020
rect 15856 15008 15884 15116
rect 16022 15104 16028 15156
rect 16080 15104 16086 15156
rect 16114 15104 16120 15156
rect 16172 15144 16178 15156
rect 19613 15147 19671 15153
rect 19613 15144 19625 15147
rect 16172 15116 19625 15144
rect 16172 15104 16178 15116
rect 19613 15113 19625 15116
rect 19659 15144 19671 15147
rect 19978 15144 19984 15156
rect 19659 15116 19984 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 19978 15104 19984 15116
rect 20036 15144 20042 15156
rect 20036 15116 21588 15144
rect 20036 15104 20042 15116
rect 16040 15076 16068 15104
rect 16390 15076 16396 15088
rect 16040 15048 16396 15076
rect 16390 15036 16396 15048
rect 16448 15076 16454 15088
rect 16669 15079 16727 15085
rect 16669 15076 16681 15079
rect 16448 15048 16681 15076
rect 16448 15036 16454 15048
rect 16669 15045 16681 15048
rect 16715 15045 16727 15079
rect 16669 15039 16727 15045
rect 16022 15008 16028 15020
rect 15856 14994 16028 15008
rect 15870 14980 16028 14994
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16206 14968 16212 15020
rect 16264 15008 16270 15020
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 16264 14980 16313 15008
rect 16264 14968 16270 14980
rect 16301 14977 16313 14980
rect 16347 14977 16359 15011
rect 16684 15008 16712 15039
rect 17402 15036 17408 15088
rect 17460 15036 17466 15088
rect 17681 15079 17739 15085
rect 17681 15045 17693 15079
rect 17727 15076 17739 15079
rect 18138 15076 18144 15088
rect 17727 15048 18144 15076
rect 17727 15045 17739 15048
rect 17681 15039 17739 15045
rect 18138 15036 18144 15048
rect 18196 15036 18202 15088
rect 19061 15079 19119 15085
rect 19061 15045 19073 15079
rect 19107 15076 19119 15079
rect 20162 15076 20168 15088
rect 19107 15048 20168 15076
rect 19107 15045 19119 15048
rect 19061 15039 19119 15045
rect 18233 15011 18291 15017
rect 18233 15008 18245 15011
rect 16684 14980 18245 15008
rect 16301 14971 16359 14977
rect 18233 14977 18245 14980
rect 18279 14977 18291 15011
rect 18233 14971 18291 14977
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 12161 14943 12219 14949
rect 11716 14912 12112 14940
rect 9033 14875 9091 14881
rect 9033 14841 9045 14875
rect 9079 14872 9091 14875
rect 9324 14872 9352 14912
rect 9079 14844 9352 14872
rect 9079 14841 9091 14844
rect 9033 14835 9091 14841
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 8168 14776 8309 14804
rect 8168 14764 8174 14776
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 8297 14767 8355 14773
rect 8570 14764 8576 14816
rect 8628 14804 8634 14816
rect 11716 14804 11744 14912
rect 12084 14872 12112 14912
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12434 14940 12440 14952
rect 12207 14912 12440 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14424 14912 14473 14940
rect 14424 14900 14430 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14940 14795 14943
rect 15470 14940 15476 14952
rect 14783 14912 15476 14940
rect 14783 14909 14795 14912
rect 14737 14903 14795 14909
rect 12084 14844 12193 14872
rect 8628 14776 11744 14804
rect 8628 14764 8634 14776
rect 12066 14764 12072 14816
rect 12124 14764 12130 14816
rect 12165 14804 12193 14844
rect 12618 14804 12624 14816
rect 12165 14776 12624 14804
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 14476 14804 14504 14903
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 16040 14940 16068 14968
rect 17218 14940 17224 14952
rect 16040 14912 17224 14940
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 17126 14872 17132 14884
rect 16132 14844 17132 14872
rect 14734 14804 14740 14816
rect 14476 14776 14740 14804
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 14826 14764 14832 14816
rect 14884 14804 14890 14816
rect 16132 14804 16160 14844
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 17954 14832 17960 14884
rect 18012 14832 18018 14884
rect 18248 14872 18276 14971
rect 19444 14940 19472 14971
rect 19610 14968 19616 15020
rect 19668 15008 19674 15020
rect 19705 15011 19763 15017
rect 19705 15008 19717 15011
rect 19668 14980 19717 15008
rect 19668 14968 19674 14980
rect 19705 14977 19717 14980
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 19794 14968 19800 15020
rect 19852 14968 19858 15020
rect 19904 15017 19932 15048
rect 20162 15036 20168 15048
rect 20220 15036 20226 15088
rect 19889 15011 19947 15017
rect 19889 14977 19901 15011
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 21232 14980 21298 15008
rect 21232 14968 21238 14980
rect 19812 14940 19840 14968
rect 21560 14952 21588 15116
rect 25222 15104 25228 15156
rect 25280 15144 25286 15156
rect 26234 15144 26240 15156
rect 25280 15116 26240 15144
rect 25280 15104 25286 15116
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 26344 15116 27502 15144
rect 24026 15036 24032 15088
rect 24084 15036 24090 15088
rect 24670 15036 24676 15088
rect 24728 15036 24734 15088
rect 24762 15036 24768 15088
rect 24820 15036 24826 15088
rect 24854 15036 24860 15088
rect 24912 15036 24918 15088
rect 24946 15036 24952 15088
rect 25004 15085 25010 15088
rect 25004 15079 25033 15085
rect 25021 15076 25033 15079
rect 26344 15076 26372 15116
rect 25021 15048 26372 15076
rect 25021 15045 25033 15048
rect 25004 15039 25033 15045
rect 25004 15036 25010 15039
rect 24674 15033 24732 15036
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 19444 14912 19840 14940
rect 20162 14900 20168 14952
rect 20220 14900 20226 14952
rect 21542 14900 21548 14952
rect 21600 14900 21606 14952
rect 21637 14943 21695 14949
rect 21637 14909 21649 14943
rect 21683 14940 21695 14943
rect 22112 14940 22140 14971
rect 22370 14968 22376 15020
rect 22428 15008 22434 15020
rect 22925 15011 22983 15017
rect 22925 15008 22937 15011
rect 22428 14980 22937 15008
rect 22428 14968 22434 14980
rect 22925 14977 22937 14980
rect 22971 14977 22983 15011
rect 22925 14971 22983 14977
rect 23198 14968 23204 15020
rect 23256 15008 23262 15020
rect 23293 15011 23351 15017
rect 23293 15008 23305 15011
rect 23256 14980 23305 15008
rect 23256 14968 23262 14980
rect 23293 14977 23305 14980
rect 23339 14977 23351 15011
rect 23293 14971 23351 14977
rect 21683 14912 22140 14940
rect 22281 14943 22339 14949
rect 21683 14909 21695 14912
rect 21637 14903 21695 14909
rect 22281 14909 22293 14943
rect 22327 14909 22339 14943
rect 23308 14940 23336 14971
rect 23382 14968 23388 15020
rect 23440 15008 23446 15020
rect 23753 15011 23811 15017
rect 23753 15008 23765 15011
rect 23440 14980 23765 15008
rect 23440 14968 23446 14980
rect 23753 14977 23765 14980
rect 23799 14977 23811 15011
rect 24674 14999 24686 15033
rect 24720 14999 24732 15033
rect 24674 14993 24732 14999
rect 25133 15011 25191 15017
rect 23753 14971 23811 14977
rect 25133 14977 25145 15011
rect 25179 15008 25191 15011
rect 26053 15011 26111 15017
rect 26053 15008 26065 15011
rect 25179 14980 26065 15008
rect 25179 14977 25191 14980
rect 25133 14971 25191 14977
rect 26053 14977 26065 14980
rect 26099 14977 26111 15011
rect 26053 14971 26111 14977
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 24854 14940 24860 14952
rect 23308 14912 24860 14940
rect 22281 14903 22339 14909
rect 21560 14872 21588 14900
rect 22296 14872 22324 14903
rect 24854 14900 24860 14912
rect 24912 14900 24918 14952
rect 25406 14900 25412 14952
rect 25464 14900 25470 14952
rect 18248 14844 20024 14872
rect 21560 14844 22324 14872
rect 14884 14776 16160 14804
rect 14884 14764 14890 14776
rect 16206 14764 16212 14816
rect 16264 14764 16270 14816
rect 16393 14807 16451 14813
rect 16393 14773 16405 14807
rect 16439 14804 16451 14807
rect 16574 14804 16580 14816
rect 16439 14776 16580 14804
rect 16439 14773 16451 14776
rect 16393 14767 16451 14773
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 18138 14764 18144 14816
rect 18196 14764 18202 14816
rect 19242 14764 19248 14816
rect 19300 14764 19306 14816
rect 19996 14804 20024 14844
rect 23842 14832 23848 14884
rect 23900 14872 23906 14884
rect 26160 14872 26188 14971
rect 26234 14968 26240 15020
rect 26292 14968 26298 15020
rect 26344 15017 26372 15048
rect 26970 15036 26976 15088
rect 27028 15076 27034 15088
rect 27474 15085 27502 15116
rect 27614 15104 27620 15156
rect 27672 15104 27678 15156
rect 27893 15147 27951 15153
rect 27893 15113 27905 15147
rect 27939 15144 27951 15147
rect 28350 15144 28356 15156
rect 27939 15116 28356 15144
rect 27939 15113 27951 15116
rect 27893 15107 27951 15113
rect 27249 15079 27307 15085
rect 27249 15076 27261 15079
rect 27028 15048 27261 15076
rect 27028 15036 27034 15048
rect 27249 15045 27261 15048
rect 27295 15045 27307 15079
rect 27249 15039 27307 15045
rect 27459 15079 27517 15085
rect 27459 15045 27471 15079
rect 27505 15045 27517 15079
rect 27632 15076 27660 15104
rect 27632 15048 28028 15076
rect 27459 15039 27517 15045
rect 28000 15017 28028 15048
rect 26329 15011 26387 15017
rect 26329 14977 26341 15011
rect 26375 14977 26387 15011
rect 26329 14971 26387 14977
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 14977 27399 15011
rect 27709 15011 27767 15017
rect 27709 15008 27721 15011
rect 27341 14971 27399 14977
rect 27540 14980 27721 15008
rect 23900 14844 26188 14872
rect 26252 14872 26280 14968
rect 27172 14940 27200 14971
rect 27246 14940 27252 14952
rect 27172 14912 27252 14940
rect 27246 14900 27252 14912
rect 27304 14900 27310 14952
rect 27356 14872 27384 14971
rect 27540 14952 27568 14980
rect 27709 14977 27721 14980
rect 27755 14977 27767 15011
rect 27709 14971 27767 14977
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 27522 14900 27528 14952
rect 27580 14900 27586 14952
rect 27617 14943 27675 14949
rect 27617 14909 27629 14943
rect 27663 14940 27675 14943
rect 28092 14940 28120 15116
rect 28350 15104 28356 15116
rect 28408 15144 28414 15156
rect 28408 15116 28856 15144
rect 28408 15104 28414 15116
rect 28828 15020 28856 15116
rect 28810 14968 28816 15020
rect 28868 14968 28874 15020
rect 27663 14912 28120 14940
rect 27663 14909 27675 14912
rect 27617 14903 27675 14909
rect 27632 14872 27660 14903
rect 26252 14844 27384 14872
rect 27448 14844 27660 14872
rect 23900 14832 23906 14844
rect 20714 14804 20720 14816
rect 19996 14776 20720 14804
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 24486 14764 24492 14816
rect 24544 14764 24550 14816
rect 26973 14807 27031 14813
rect 26973 14773 26985 14807
rect 27019 14804 27031 14807
rect 27062 14804 27068 14816
rect 27019 14776 27068 14804
rect 27019 14773 27031 14776
rect 26973 14767 27031 14773
rect 27062 14764 27068 14776
rect 27120 14764 27126 14816
rect 27338 14764 27344 14816
rect 27396 14804 27402 14816
rect 27448 14804 27476 14844
rect 27706 14832 27712 14884
rect 27764 14832 27770 14884
rect 27396 14776 27476 14804
rect 27396 14764 27402 14776
rect 1104 14714 29440 14736
rect 1104 14662 4491 14714
rect 4543 14662 4555 14714
rect 4607 14662 4619 14714
rect 4671 14662 4683 14714
rect 4735 14662 4747 14714
rect 4799 14662 11574 14714
rect 11626 14662 11638 14714
rect 11690 14662 11702 14714
rect 11754 14662 11766 14714
rect 11818 14662 11830 14714
rect 11882 14662 18657 14714
rect 18709 14662 18721 14714
rect 18773 14662 18785 14714
rect 18837 14662 18849 14714
rect 18901 14662 18913 14714
rect 18965 14662 25740 14714
rect 25792 14662 25804 14714
rect 25856 14662 25868 14714
rect 25920 14662 25932 14714
rect 25984 14662 25996 14714
rect 26048 14662 29440 14714
rect 1104 14640 29440 14662
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 6880 14572 7665 14600
rect 6880 14560 6886 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 10410 14560 10416 14612
rect 10468 14600 10474 14612
rect 11330 14600 11336 14612
rect 10468 14572 11336 14600
rect 10468 14560 10474 14572
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 11872 14603 11930 14609
rect 11872 14569 11884 14603
rect 11918 14600 11930 14603
rect 12066 14600 12072 14612
rect 11918 14572 12072 14600
rect 11918 14569 11930 14572
rect 11872 14563 11930 14569
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 13354 14560 13360 14612
rect 13412 14560 13418 14612
rect 16025 14603 16083 14609
rect 16025 14569 16037 14603
rect 16071 14600 16083 14603
rect 16114 14600 16120 14612
rect 16071 14572 16120 14600
rect 16071 14569 16083 14572
rect 16025 14563 16083 14569
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 16206 14560 16212 14612
rect 16264 14560 16270 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18785 14603 18843 14609
rect 18785 14600 18797 14603
rect 18196 14572 18797 14600
rect 18196 14560 18202 14572
rect 18785 14569 18797 14572
rect 18831 14569 18843 14603
rect 18785 14563 18843 14569
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 19300 14572 20085 14600
rect 19300 14560 19306 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 20073 14563 20131 14569
rect 20162 14560 20168 14612
rect 20220 14600 20226 14612
rect 20717 14603 20775 14609
rect 20717 14600 20729 14603
rect 20220 14572 20729 14600
rect 20220 14560 20226 14572
rect 20717 14569 20729 14572
rect 20763 14569 20775 14603
rect 20717 14563 20775 14569
rect 20898 14560 20904 14612
rect 20956 14600 20962 14612
rect 23109 14603 23167 14609
rect 20956 14572 23060 14600
rect 20956 14560 20962 14572
rect 10502 14532 10508 14544
rect 7852 14504 10508 14532
rect 7852 14408 7880 14504
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 10594 14492 10600 14544
rect 10652 14532 10658 14544
rect 10870 14532 10876 14544
rect 10652 14504 10876 14532
rect 10652 14492 10658 14504
rect 10870 14492 10876 14504
rect 10928 14492 10934 14544
rect 8110 14424 8116 14476
rect 8168 14424 8174 14476
rect 11609 14467 11667 14473
rect 11609 14464 11621 14467
rect 9232 14436 11621 14464
rect 9232 14408 9260 14436
rect 11609 14433 11621 14436
rect 11655 14464 11667 14467
rect 12434 14464 12440 14476
rect 11655 14436 12440 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 15105 14467 15163 14473
rect 15105 14464 15117 14467
rect 14424 14436 15117 14464
rect 14424 14424 14430 14436
rect 15105 14433 15117 14436
rect 15151 14464 15163 14467
rect 16224 14464 16252 14560
rect 18506 14492 18512 14544
rect 18564 14492 18570 14544
rect 18690 14492 18696 14544
rect 18748 14532 18754 14544
rect 22281 14535 22339 14541
rect 22281 14532 22293 14535
rect 18748 14504 20208 14532
rect 18748 14492 18754 14504
rect 15151 14436 16252 14464
rect 18524 14464 18552 14492
rect 19076 14476 19104 14504
rect 18524 14436 18920 14464
rect 15151 14433 15163 14436
rect 15105 14427 15163 14433
rect 18892 14408 18920 14436
rect 19058 14424 19064 14476
rect 19116 14424 19122 14476
rect 20070 14464 20076 14476
rect 19444 14436 20076 14464
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14365 7159 14399
rect 7101 14359 7159 14365
rect 7116 14260 7144 14359
rect 7374 14356 7380 14408
rect 7432 14356 7438 14408
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14396 7527 14399
rect 7834 14396 7840 14408
rect 7515 14368 7840 14396
rect 7515 14365 7527 14368
rect 7469 14359 7527 14365
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 9214 14356 9220 14408
rect 9272 14356 9278 14408
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 10561 14399 10619 14405
rect 10561 14365 10573 14399
rect 10607 14396 10619 14399
rect 10607 14365 10640 14396
rect 10561 14359 10640 14365
rect 7285 14331 7343 14337
rect 7285 14297 7297 14331
rect 7331 14328 7343 14331
rect 7558 14328 7564 14340
rect 7331 14300 7564 14328
rect 7331 14297 7343 14300
rect 7285 14291 7343 14297
rect 7558 14288 7564 14300
rect 7616 14328 7622 14340
rect 8570 14328 8576 14340
rect 7616 14300 8576 14328
rect 7616 14288 7622 14300
rect 8570 14288 8576 14300
rect 8628 14288 8634 14340
rect 8665 14263 8723 14269
rect 8665 14260 8677 14263
rect 7116 14232 8677 14260
rect 8665 14229 8677 14232
rect 8711 14229 8723 14263
rect 10612 14260 10640 14359
rect 10778 14356 10784 14408
rect 10836 14356 10842 14408
rect 10870 14356 10876 14408
rect 10928 14405 10934 14408
rect 10928 14396 10936 14405
rect 14185 14399 14243 14405
rect 10928 14368 10973 14396
rect 10928 14359 10936 14368
rect 14185 14365 14197 14399
rect 14231 14396 14243 14399
rect 14274 14396 14280 14408
rect 14231 14368 14280 14396
rect 14231 14365 14243 14368
rect 14185 14359 14243 14365
rect 10928 14356 10934 14359
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 16022 14396 16028 14408
rect 15795 14368 16028 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16298 14356 16304 14408
rect 16356 14356 16362 14408
rect 16482 14356 16488 14408
rect 16540 14356 16546 14408
rect 16574 14356 16580 14408
rect 16632 14396 16638 14408
rect 18509 14399 18567 14405
rect 18509 14396 18521 14399
rect 16632 14368 18521 14396
rect 16632 14356 16638 14368
rect 18509 14365 18521 14368
rect 18555 14365 18567 14399
rect 18509 14359 18567 14365
rect 18598 14356 18604 14408
rect 18656 14356 18662 14408
rect 18874 14356 18880 14408
rect 18932 14356 18938 14408
rect 19444 14405 19472 14436
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 20180 14408 20208 14504
rect 20272 14504 22293 14532
rect 20272 14473 20300 14504
rect 22281 14501 22293 14504
rect 22327 14501 22339 14535
rect 22281 14495 22339 14501
rect 20257 14467 20315 14473
rect 20257 14433 20269 14467
rect 20303 14433 20315 14467
rect 20257 14427 20315 14433
rect 20364 14436 21036 14464
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19610 14356 19616 14408
rect 19668 14356 19674 14408
rect 19794 14405 19800 14408
rect 19751 14399 19800 14405
rect 19751 14365 19763 14399
rect 19797 14365 19800 14399
rect 19751 14359 19800 14365
rect 19794 14356 19800 14359
rect 19852 14356 19858 14408
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20162 14396 20168 14408
rect 19935 14368 20168 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 20162 14356 20168 14368
rect 20220 14396 20226 14408
rect 20364 14396 20392 14436
rect 20220 14368 20392 14396
rect 20441 14399 20499 14405
rect 20220 14356 20226 14368
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 20530 14396 20536 14408
rect 20487 14368 20536 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 20901 14399 20959 14405
rect 20640 14394 20760 14396
rect 20901 14394 20913 14399
rect 20640 14368 20913 14394
rect 10686 14288 10692 14340
rect 10744 14288 10750 14340
rect 13538 14328 13544 14340
rect 13110 14300 13544 14328
rect 13538 14288 13544 14300
rect 13596 14328 13602 14340
rect 14553 14331 14611 14337
rect 14553 14328 14565 14331
rect 13596 14300 14565 14328
rect 13596 14288 13602 14300
rect 14553 14297 14565 14300
rect 14599 14297 14611 14331
rect 14553 14291 14611 14297
rect 10962 14260 10968 14272
rect 10612 14232 10968 14260
rect 8665 14223 8723 14229
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 11054 14220 11060 14272
rect 11112 14220 11118 14272
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 15562 14260 15568 14272
rect 12032 14232 15568 14260
rect 12032 14220 12038 14232
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 15654 14220 15660 14272
rect 15712 14220 15718 14272
rect 16209 14263 16267 14269
rect 16209 14229 16221 14263
rect 16255 14260 16267 14263
rect 16316 14260 16344 14356
rect 19521 14331 19579 14337
rect 19521 14297 19533 14331
rect 19567 14297 19579 14331
rect 19628 14328 19656 14356
rect 19628 14300 19932 14328
rect 19521 14291 19579 14297
rect 16255 14232 16344 14260
rect 16255 14229 16267 14232
rect 16209 14223 16267 14229
rect 16758 14220 16764 14272
rect 16816 14220 16822 14272
rect 18322 14220 18328 14272
rect 18380 14220 18386 14272
rect 19242 14220 19248 14272
rect 19300 14220 19306 14272
rect 19536 14260 19564 14291
rect 19904 14272 19932 14300
rect 19978 14288 19984 14340
rect 20036 14288 20042 14340
rect 19610 14260 19616 14272
rect 19536 14232 19616 14260
rect 19610 14220 19616 14232
rect 19668 14220 19674 14272
rect 19886 14220 19892 14272
rect 19944 14220 19950 14272
rect 20640 14269 20668 14368
rect 20732 14366 20913 14368
rect 20901 14365 20913 14366
rect 20947 14365 20959 14399
rect 21008 14396 21036 14436
rect 21082 14424 21088 14476
rect 21140 14464 21146 14476
rect 22741 14467 22799 14473
rect 21140 14436 22600 14464
rect 21140 14424 21146 14436
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 21008 14368 21373 14396
rect 20901 14359 20959 14365
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21542 14356 21548 14408
rect 21600 14356 21606 14408
rect 21634 14356 21640 14408
rect 21692 14356 21698 14408
rect 21730 14399 21788 14405
rect 21730 14365 21742 14399
rect 21776 14365 21788 14399
rect 21730 14359 21788 14365
rect 22143 14399 22201 14405
rect 22143 14365 22155 14399
rect 22189 14396 22201 14399
rect 22278 14396 22284 14408
rect 22189 14368 22284 14396
rect 22189 14365 22201 14368
rect 22143 14359 22201 14365
rect 21453 14331 21511 14337
rect 21453 14297 21465 14331
rect 21499 14328 21511 14331
rect 21744 14328 21772 14359
rect 22278 14356 22284 14368
rect 22336 14356 22342 14408
rect 22370 14356 22376 14408
rect 22428 14356 22434 14408
rect 22572 14405 22600 14436
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 23032 14464 23060 14572
rect 23109 14569 23121 14603
rect 23155 14600 23167 14603
rect 23382 14600 23388 14612
rect 23155 14572 23388 14600
rect 23155 14569 23167 14572
rect 23109 14563 23167 14569
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 23566 14560 23572 14612
rect 23624 14560 23630 14612
rect 24486 14560 24492 14612
rect 24544 14600 24550 14612
rect 24746 14603 24804 14609
rect 24746 14600 24758 14603
rect 24544 14572 24758 14600
rect 24544 14560 24550 14572
rect 24746 14569 24758 14572
rect 24792 14569 24804 14603
rect 24746 14563 24804 14569
rect 26878 14560 26884 14612
rect 26936 14560 26942 14612
rect 23842 14464 23848 14476
rect 22787 14436 23848 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 23842 14424 23848 14436
rect 23900 14424 23906 14476
rect 24486 14424 24492 14476
rect 24544 14464 24550 14476
rect 26789 14467 26847 14473
rect 26789 14464 26801 14467
rect 24544 14436 26801 14464
rect 24544 14424 24550 14436
rect 26789 14433 26801 14436
rect 26835 14464 26847 14467
rect 26896 14464 26924 14560
rect 26835 14436 26924 14464
rect 26835 14433 26847 14436
rect 26789 14427 26847 14433
rect 27062 14424 27068 14476
rect 27120 14424 27126 14476
rect 28810 14424 28816 14476
rect 28868 14424 28874 14476
rect 22557 14399 22615 14405
rect 22557 14365 22569 14399
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 22646 14356 22652 14408
rect 22704 14356 22710 14408
rect 22830 14356 22836 14408
rect 22888 14396 22894 14408
rect 22925 14399 22983 14405
rect 22925 14396 22937 14399
rect 22888 14368 22937 14396
rect 22888 14356 22894 14368
rect 22925 14365 22937 14368
rect 22971 14365 22983 14399
rect 22925 14359 22983 14365
rect 23477 14399 23535 14405
rect 23477 14365 23489 14399
rect 23523 14396 23535 14399
rect 23658 14396 23664 14408
rect 23523 14368 23664 14396
rect 23523 14365 23535 14368
rect 23477 14359 23535 14365
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 21499 14300 21772 14328
rect 21913 14331 21971 14337
rect 21499 14297 21511 14300
rect 21453 14291 21511 14297
rect 21913 14297 21925 14331
rect 21959 14297 21971 14331
rect 21913 14291 21971 14297
rect 22005 14331 22063 14337
rect 22005 14297 22017 14331
rect 22051 14328 22063 14331
rect 25038 14328 25044 14340
rect 22051 14300 25044 14328
rect 22051 14297 22063 14300
rect 22005 14291 22063 14297
rect 20625 14263 20683 14269
rect 20625 14229 20637 14263
rect 20671 14229 20683 14263
rect 21928 14260 21956 14291
rect 25038 14288 25044 14300
rect 25096 14288 25102 14340
rect 25314 14288 25320 14340
rect 25372 14288 25378 14340
rect 26513 14331 26571 14337
rect 26513 14297 26525 14331
rect 26559 14297 26571 14331
rect 26513 14291 26571 14297
rect 22094 14260 22100 14272
rect 21928 14232 22100 14260
rect 20625 14223 20683 14229
rect 22094 14220 22100 14232
rect 22152 14220 22158 14272
rect 23934 14220 23940 14272
rect 23992 14220 23998 14272
rect 25406 14220 25412 14272
rect 25464 14260 25470 14272
rect 26528 14260 26556 14291
rect 27522 14288 27528 14340
rect 27580 14288 27586 14340
rect 25464 14232 26556 14260
rect 25464 14220 25470 14232
rect 1104 14170 29440 14192
rect 1104 14118 5151 14170
rect 5203 14118 5215 14170
rect 5267 14118 5279 14170
rect 5331 14118 5343 14170
rect 5395 14118 5407 14170
rect 5459 14118 12234 14170
rect 12286 14118 12298 14170
rect 12350 14118 12362 14170
rect 12414 14118 12426 14170
rect 12478 14118 12490 14170
rect 12542 14118 19317 14170
rect 19369 14118 19381 14170
rect 19433 14118 19445 14170
rect 19497 14118 19509 14170
rect 19561 14118 19573 14170
rect 19625 14118 26400 14170
rect 26452 14118 26464 14170
rect 26516 14118 26528 14170
rect 26580 14118 26592 14170
rect 26644 14118 26656 14170
rect 26708 14118 29440 14170
rect 1104 14096 29440 14118
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10962 14056 10968 14068
rect 10376 14028 10968 14056
rect 10376 14016 10382 14028
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11054 14016 11060 14068
rect 11112 14016 11118 14068
rect 13814 14016 13820 14068
rect 13872 14016 13878 14068
rect 14366 14016 14372 14068
rect 14424 14016 14430 14068
rect 15654 14056 15660 14068
rect 14936 14028 15660 14056
rect 3234 13988 3240 14000
rect 3082 13960 3240 13988
rect 3234 13948 3240 13960
rect 3292 13948 3298 14000
rect 3602 13948 3608 14000
rect 3660 13948 3666 14000
rect 9876 13960 10916 13988
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1452 13892 1593 13920
rect 1452 13880 1458 13892
rect 1581 13889 1593 13892
rect 1627 13889 1639 13923
rect 1581 13883 1639 13889
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 9876 13929 9904 13960
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 5684 13892 6561 13920
rect 5684 13880 5690 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 9861 13923 9919 13929
rect 6779 13892 7328 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7300 13864 7328 13892
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 10045 13923 10103 13929
rect 10045 13920 10057 13923
rect 10008 13892 10057 13920
rect 10008 13880 10014 13892
rect 10045 13889 10057 13892
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 1854 13812 1860 13864
rect 1912 13812 1918 13864
rect 5902 13812 5908 13864
rect 5960 13812 5966 13864
rect 6638 13812 6644 13864
rect 6696 13812 6702 13864
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 5920 13784 5948 13812
rect 6546 13784 6552 13796
rect 5920 13756 6552 13784
rect 6546 13744 6552 13756
rect 6604 13784 6610 13796
rect 6840 13784 6868 13815
rect 7282 13812 7288 13864
rect 7340 13812 7346 13864
rect 10152 13852 10180 13883
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 10502 13920 10508 13932
rect 10284 13892 10508 13920
rect 10284 13880 10290 13892
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 10152 13824 10732 13852
rect 7098 13784 7104 13796
rect 6604 13756 7104 13784
rect 6604 13744 6610 13756
rect 7098 13744 7104 13756
rect 7156 13744 7162 13796
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 10704 13784 10732 13824
rect 10778 13812 10784 13864
rect 10836 13812 10842 13864
rect 10888 13852 10916 13960
rect 11072 13920 11100 14016
rect 13832 13988 13860 14016
rect 13832 13960 14228 13988
rect 14200 13929 14228 13960
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 11072 13892 14105 13920
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14384 13861 14412 14016
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13920 14519 13923
rect 14826 13920 14832 13932
rect 14507 13892 14832 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 14936 13929 14964 14028
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 18414 14016 18420 14068
rect 18472 14056 18478 14068
rect 19058 14056 19064 14068
rect 18472 14028 19064 14056
rect 18472 14016 18478 14028
rect 19058 14016 19064 14028
rect 19116 14056 19122 14068
rect 19116 14028 19288 14056
rect 19116 14016 19122 14028
rect 15197 13991 15255 13997
rect 15197 13957 15209 13991
rect 15243 13988 15255 13991
rect 15562 13988 15568 14000
rect 15243 13960 15568 13988
rect 15243 13957 15255 13960
rect 15197 13951 15255 13957
rect 15562 13948 15568 13960
rect 15620 13948 15626 14000
rect 18340 13988 18368 14016
rect 18340 13960 18920 13988
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13920 15163 13923
rect 15289 13923 15347 13929
rect 15151 13892 15240 13920
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 10888 13824 11345 13852
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 11422 13784 11428 13796
rect 7248 13756 10548 13784
rect 10704 13756 11428 13784
rect 7248 13744 7254 13756
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 6362 13716 6368 13728
rect 6236 13688 6368 13716
rect 6236 13676 6242 13688
rect 6362 13676 6368 13688
rect 6420 13716 6426 13728
rect 10134 13716 10140 13728
rect 6420 13688 10140 13716
rect 6420 13676 6426 13688
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10410 13676 10416 13728
rect 10468 13676 10474 13728
rect 10520 13716 10548 13756
rect 11422 13744 11428 13756
rect 11480 13744 11486 13796
rect 13909 13787 13967 13793
rect 13909 13753 13921 13787
rect 13955 13784 13967 13787
rect 15102 13784 15108 13796
rect 13955 13756 15108 13784
rect 13955 13753 13967 13756
rect 13909 13747 13967 13753
rect 15102 13744 15108 13756
rect 15160 13744 15166 13796
rect 11146 13716 11152 13728
rect 10520 13688 11152 13716
rect 11146 13676 11152 13688
rect 11204 13716 11210 13728
rect 14090 13716 14096 13728
rect 11204 13688 14096 13716
rect 11204 13676 11210 13688
rect 14090 13676 14096 13688
rect 14148 13676 14154 13728
rect 15212 13716 15240 13892
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 17034 13920 17040 13932
rect 15335 13892 17040 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 18616 13852 18644 13883
rect 18690 13880 18696 13932
rect 18748 13880 18754 13932
rect 18892 13929 18920 13960
rect 19150 13948 19156 14000
rect 19208 13948 19214 14000
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 18969 13923 19027 13929
rect 18969 13889 18981 13923
rect 19015 13920 19027 13923
rect 19061 13923 19119 13929
rect 19061 13920 19073 13923
rect 19015 13892 19073 13920
rect 19015 13889 19027 13892
rect 18969 13883 19027 13889
rect 19061 13889 19073 13892
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 19168 13852 19196 13948
rect 19260 13929 19288 14028
rect 19352 14028 19932 14056
rect 19352 13929 19380 14028
rect 19702 13948 19708 14000
rect 19760 13948 19766 14000
rect 19904 13997 19932 14028
rect 19978 14016 19984 14068
rect 20036 14056 20042 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 20036 14028 20545 14056
rect 20036 14016 20042 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 20533 14019 20591 14025
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 20680 14028 21557 14056
rect 20680 14016 20686 14028
rect 21545 14025 21557 14028
rect 21591 14025 21603 14059
rect 21545 14019 21603 14025
rect 22370 14016 22376 14068
rect 22428 14056 22434 14068
rect 23382 14056 23388 14068
rect 22428 14028 23388 14056
rect 22428 14016 22434 14028
rect 23382 14016 23388 14028
rect 23440 14056 23446 14068
rect 23661 14059 23719 14065
rect 23661 14056 23673 14059
rect 23440 14028 23673 14056
rect 23440 14016 23446 14028
rect 23661 14025 23673 14028
rect 23707 14025 23719 14059
rect 26237 14059 26295 14065
rect 26237 14056 26249 14059
rect 23661 14019 23719 14025
rect 25056 14028 26249 14056
rect 25056 14000 25084 14028
rect 26237 14025 26249 14028
rect 26283 14056 26295 14059
rect 27614 14056 27620 14068
rect 26283 14028 27620 14056
rect 26283 14025 26295 14028
rect 26237 14019 26295 14025
rect 27614 14016 27620 14028
rect 27672 14016 27678 14068
rect 19889 13991 19947 13997
rect 19889 13957 19901 13991
rect 19935 13988 19947 13991
rect 21450 13988 21456 14000
rect 19935 13960 21456 13988
rect 19935 13957 19947 13960
rect 19889 13951 19947 13957
rect 21450 13948 21456 13960
rect 21508 13988 21514 14000
rect 21726 13988 21732 14000
rect 21508 13960 21732 13988
rect 21508 13948 21514 13960
rect 21726 13948 21732 13960
rect 21784 13948 21790 14000
rect 23566 13948 23572 14000
rect 23624 13988 23630 14000
rect 24210 13988 24216 14000
rect 23624 13960 24216 13988
rect 23624 13948 23630 13960
rect 24210 13948 24216 13960
rect 24268 13948 24274 14000
rect 25038 13948 25044 14000
rect 25096 13948 25102 14000
rect 25314 13948 25320 14000
rect 25372 13948 25378 14000
rect 19245 13923 19303 13929
rect 19245 13889 19257 13923
rect 19291 13889 19303 13923
rect 19245 13883 19303 13889
rect 19337 13923 19395 13929
rect 19337 13889 19349 13923
rect 19383 13889 19395 13923
rect 19337 13883 19395 13889
rect 19518 13880 19524 13932
rect 19576 13880 19582 13932
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13920 19671 13923
rect 20070 13920 20076 13932
rect 19659 13892 20076 13920
rect 19659 13889 19671 13892
rect 19613 13883 19671 13889
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20165 13923 20223 13929
rect 20165 13889 20177 13923
rect 20211 13920 20223 13923
rect 20211 13892 20668 13920
rect 20211 13889 20223 13892
rect 20165 13883 20223 13889
rect 20180 13852 20208 13883
rect 18616 13824 19196 13852
rect 19260 13824 20208 13852
rect 15470 13744 15476 13796
rect 15528 13744 15534 13796
rect 16850 13744 16856 13796
rect 16908 13744 16914 13796
rect 18138 13744 18144 13796
rect 18196 13784 18202 13796
rect 19260 13784 19288 13824
rect 20254 13812 20260 13864
rect 20312 13812 20318 13864
rect 20640 13852 20668 13892
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 20772 13892 22661 13920
rect 20772 13880 20778 13892
rect 22649 13889 22661 13892
rect 22695 13889 22707 13923
rect 22649 13883 22707 13889
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 24486 13920 24492 13932
rect 23532 13892 24492 13920
rect 23532 13880 23538 13892
rect 24486 13880 24492 13892
rect 24544 13880 24550 13932
rect 27982 13880 27988 13932
rect 28040 13880 28046 13932
rect 20990 13852 20996 13864
rect 20640 13824 20996 13852
rect 20990 13812 20996 13824
rect 21048 13812 21054 13864
rect 21085 13855 21143 13861
rect 21085 13821 21097 13855
rect 21131 13852 21143 13855
rect 22186 13852 22192 13864
rect 21131 13824 22192 13852
rect 21131 13821 21143 13824
rect 21085 13815 21143 13821
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 24029 13855 24087 13861
rect 24029 13821 24041 13855
rect 24075 13821 24087 13855
rect 24029 13815 24087 13821
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24210 13852 24216 13864
rect 24167 13824 24216 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 18196 13756 19288 13784
rect 18196 13744 18202 13756
rect 19794 13744 19800 13796
rect 19852 13784 19858 13796
rect 20073 13787 20131 13793
rect 20073 13784 20085 13787
rect 19852 13756 20085 13784
rect 19852 13744 19858 13756
rect 20073 13753 20085 13756
rect 20119 13753 20131 13787
rect 21358 13784 21364 13796
rect 20073 13747 20131 13753
rect 20180 13756 21364 13784
rect 15746 13716 15752 13728
rect 15212 13688 15752 13716
rect 15746 13676 15752 13688
rect 15804 13716 15810 13728
rect 16868 13716 16896 13744
rect 15804 13688 16896 13716
rect 15804 13676 15810 13688
rect 18414 13676 18420 13728
rect 18472 13676 18478 13728
rect 18874 13676 18880 13728
rect 18932 13716 18938 13728
rect 20180 13725 20208 13756
rect 21358 13744 21364 13756
rect 21416 13744 21422 13796
rect 20165 13719 20223 13725
rect 20165 13716 20177 13719
rect 18932 13688 20177 13716
rect 18932 13676 18938 13688
rect 20165 13685 20177 13688
rect 20211 13685 20223 13719
rect 24044 13716 24072 13815
rect 24210 13812 24216 13824
rect 24268 13812 24274 13864
rect 24305 13855 24363 13861
rect 24305 13821 24317 13855
rect 24351 13852 24363 13855
rect 24765 13855 24823 13861
rect 24765 13852 24777 13855
rect 24351 13824 24777 13852
rect 24351 13821 24363 13824
rect 24305 13815 24363 13821
rect 24765 13821 24777 13824
rect 24811 13821 24823 13855
rect 24765 13815 24823 13821
rect 25314 13812 25320 13864
rect 25372 13852 25378 13864
rect 27522 13852 27528 13864
rect 25372 13824 27528 13852
rect 25372 13812 25378 13824
rect 27522 13812 27528 13824
rect 27580 13852 27586 13864
rect 28353 13855 28411 13861
rect 28353 13852 28365 13855
rect 27580 13824 28365 13852
rect 27580 13812 27586 13824
rect 28353 13821 28365 13824
rect 28399 13821 28411 13855
rect 28353 13815 28411 13821
rect 24946 13716 24952 13728
rect 24044 13688 24952 13716
rect 20165 13679 20223 13685
rect 24946 13676 24952 13688
rect 25004 13676 25010 13728
rect 1104 13626 29440 13648
rect 1104 13574 4491 13626
rect 4543 13574 4555 13626
rect 4607 13574 4619 13626
rect 4671 13574 4683 13626
rect 4735 13574 4747 13626
rect 4799 13574 11574 13626
rect 11626 13574 11638 13626
rect 11690 13574 11702 13626
rect 11754 13574 11766 13626
rect 11818 13574 11830 13626
rect 11882 13574 18657 13626
rect 18709 13574 18721 13626
rect 18773 13574 18785 13626
rect 18837 13574 18849 13626
rect 18901 13574 18913 13626
rect 18965 13574 25740 13626
rect 25792 13574 25804 13626
rect 25856 13574 25868 13626
rect 25920 13574 25932 13626
rect 25984 13574 25996 13626
rect 26048 13574 29440 13626
rect 1104 13552 29440 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 2225 13515 2283 13521
rect 2225 13512 2237 13515
rect 1912 13484 2237 13512
rect 1912 13472 1918 13484
rect 2225 13481 2237 13484
rect 2271 13481 2283 13515
rect 2225 13475 2283 13481
rect 3602 13472 3608 13524
rect 3660 13472 3666 13524
rect 6273 13515 6331 13521
rect 6273 13481 6285 13515
rect 6319 13512 6331 13515
rect 6638 13512 6644 13524
rect 6319 13484 6644 13512
rect 6319 13481 6331 13484
rect 6273 13475 6331 13481
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 7190 13472 7196 13524
rect 7248 13472 7254 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 13262 13512 13268 13524
rect 8527 13484 13268 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 16942 13512 16948 13524
rect 15304 13484 16948 13512
rect 2593 13447 2651 13453
rect 2593 13413 2605 13447
rect 2639 13413 2651 13447
rect 2593 13407 2651 13413
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2608 13308 2636 13407
rect 3237 13379 3295 13385
rect 3237 13345 3249 13379
rect 3283 13376 3295 13379
rect 3620 13376 3648 13472
rect 7208 13444 7236 13472
rect 15304 13456 15332 13484
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18785 13515 18843 13521
rect 18785 13512 18797 13515
rect 18564 13484 18797 13512
rect 18564 13472 18570 13484
rect 18785 13481 18797 13484
rect 18831 13481 18843 13515
rect 18785 13475 18843 13481
rect 3283 13348 3648 13376
rect 6104 13416 7236 13444
rect 3283 13345 3295 13348
rect 3237 13339 3295 13345
rect 2455 13280 2636 13308
rect 2961 13311 3019 13317
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 3050 13308 3056 13320
rect 3007 13280 3056 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 3050 13268 3056 13280
rect 3108 13308 3114 13320
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 3108 13280 3433 13308
rect 3108 13268 3114 13280
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13308 3663 13311
rect 6104 13308 6132 13416
rect 9766 13404 9772 13456
rect 9824 13444 9830 13456
rect 12069 13447 12127 13453
rect 12069 13444 12081 13447
rect 9824 13416 12081 13444
rect 9824 13404 9830 13416
rect 12069 13413 12081 13416
rect 12115 13413 12127 13447
rect 12069 13407 12127 13413
rect 15286 13404 15292 13456
rect 15344 13404 15350 13456
rect 15841 13447 15899 13453
rect 15841 13413 15853 13447
rect 15887 13444 15899 13447
rect 17586 13444 17592 13456
rect 15887 13416 17592 13444
rect 15887 13413 15899 13416
rect 15841 13407 15899 13413
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 6196 13348 9168 13376
rect 6196 13317 6224 13348
rect 7208 13320 7236 13348
rect 3651 13280 6132 13308
rect 6181 13311 6239 13317
rect 3651 13277 3663 13280
rect 3605 13271 3663 13277
rect 6181 13277 6193 13311
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13308 6607 13311
rect 6914 13308 6920 13320
rect 6595 13280 6920 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 6914 13268 6920 13280
rect 6972 13268 6978 13320
rect 7098 13268 7104 13320
rect 7156 13268 7162 13320
rect 7190 13268 7196 13320
rect 7248 13268 7254 13320
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 8128 13317 8156 13348
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 7116 13240 7144 13268
rect 7576 13240 7604 13271
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 9140 13317 9168 13348
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 13446 13376 13452 13388
rect 9456 13348 13452 13376
rect 9456 13336 9462 13348
rect 13446 13336 13452 13348
rect 13504 13376 13510 13388
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 13504 13348 14504 13376
rect 13504 13336 13510 13348
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 8260 13280 8401 13308
rect 8260 13268 8266 13280
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 10318 13308 10324 13320
rect 9723 13280 10324 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 7116 13212 7604 13240
rect 7837 13243 7895 13249
rect 7837 13209 7849 13243
rect 7883 13240 7895 13243
rect 8220 13240 8248 13268
rect 7883 13212 8248 13240
rect 8956 13240 8984 13271
rect 10318 13268 10324 13280
rect 10376 13308 10382 13320
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 10376 13280 10425 13308
rect 10376 13268 10382 13280
rect 10413 13277 10425 13280
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 10560 13280 10605 13308
rect 10560 13268 10566 13280
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 10870 13268 10876 13320
rect 10928 13317 10934 13320
rect 10928 13271 10936 13317
rect 10928 13268 10934 13271
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11480 13280 11529 13308
rect 11480 13268 11486 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11664 13280 11897 13308
rect 11664 13268 11670 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12710 13308 12716 13320
rect 12216 13280 12716 13308
rect 12216 13268 12222 13280
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 9858 13240 9864 13252
rect 8956 13212 9864 13240
rect 7883 13209 7895 13212
rect 7837 13203 7895 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 10686 13200 10692 13252
rect 10744 13200 10750 13252
rect 3053 13175 3111 13181
rect 3053 13141 3065 13175
rect 3099 13172 3111 13175
rect 3234 13172 3240 13184
rect 3099 13144 3240 13172
rect 3099 13141 3111 13144
rect 3053 13135 3111 13141
rect 3234 13132 3240 13144
rect 3292 13172 3298 13184
rect 3513 13175 3571 13181
rect 3513 13172 3525 13175
rect 3292 13144 3525 13172
rect 3292 13132 3298 13144
rect 3513 13141 3525 13144
rect 3559 13141 3571 13175
rect 3513 13135 3571 13141
rect 7098 13132 7104 13184
rect 7156 13132 7162 13184
rect 9125 13175 9183 13181
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 9398 13172 9404 13184
rect 9171 13144 9404 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 10888 13172 10916 13268
rect 14476 13252 14504 13348
rect 15580 13348 17325 13376
rect 15580 13317 15608 13348
rect 17313 13345 17325 13348
rect 17359 13345 17371 13379
rect 18800 13376 18828 13475
rect 19518 13472 19524 13524
rect 19576 13512 19582 13524
rect 20622 13512 20628 13524
rect 19576 13484 20628 13512
rect 19576 13472 19582 13484
rect 20622 13472 20628 13484
rect 20680 13472 20686 13524
rect 21358 13472 21364 13524
rect 21416 13472 21422 13524
rect 24946 13472 24952 13524
rect 25004 13512 25010 13524
rect 25777 13515 25835 13521
rect 25777 13512 25789 13515
rect 25004 13484 25789 13512
rect 25004 13472 25010 13484
rect 25777 13481 25789 13484
rect 25823 13481 25835 13515
rect 25777 13475 25835 13481
rect 28902 13472 28908 13524
rect 28960 13512 28966 13524
rect 28997 13515 29055 13521
rect 28997 13512 29009 13515
rect 28960 13484 29009 13512
rect 28960 13472 28966 13484
rect 28997 13481 29009 13484
rect 29043 13481 29055 13515
rect 28997 13475 29055 13481
rect 19337 13379 19395 13385
rect 19337 13376 19349 13379
rect 18800 13348 19349 13376
rect 17313 13339 17371 13345
rect 19337 13345 19349 13348
rect 19383 13345 19395 13379
rect 19337 13339 19395 13345
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15746 13268 15752 13320
rect 15804 13268 15810 13320
rect 16301 13311 16359 13317
rect 16040 13280 16252 13308
rect 10962 13200 10968 13252
rect 11020 13240 11026 13252
rect 11701 13243 11759 13249
rect 11701 13240 11713 13243
rect 11020 13212 11713 13240
rect 11020 13200 11026 13212
rect 11701 13209 11713 13212
rect 11747 13209 11759 13243
rect 11701 13203 11759 13209
rect 11790 13200 11796 13252
rect 11848 13200 11854 13252
rect 11992 13212 12434 13240
rect 10284 13144 10916 13172
rect 11057 13175 11115 13181
rect 10284 13132 10290 13144
rect 11057 13141 11069 13175
rect 11103 13172 11115 13175
rect 11992 13172 12020 13212
rect 11103 13144 12020 13172
rect 12406 13172 12434 13212
rect 14458 13200 14464 13252
rect 14516 13200 14522 13252
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 16040 13240 16068 13280
rect 15160 13212 16068 13240
rect 16117 13243 16175 13249
rect 15160 13200 15166 13212
rect 16117 13209 16129 13243
rect 16163 13209 16175 13243
rect 16224 13240 16252 13280
rect 16301 13277 16313 13311
rect 16347 13308 16359 13311
rect 16482 13308 16488 13320
rect 16347 13280 16488 13308
rect 16347 13277 16359 13280
rect 16301 13271 16359 13277
rect 16482 13268 16488 13280
rect 16540 13308 16546 13320
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16540 13280 16957 13308
rect 16540 13268 16546 13280
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 17126 13268 17132 13320
rect 17184 13308 17190 13320
rect 17954 13308 17960 13320
rect 17184 13280 17960 13308
rect 17184 13268 17190 13280
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 18138 13268 18144 13320
rect 18196 13308 18202 13320
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 18196 13280 18797 13308
rect 18196 13268 18202 13280
rect 18785 13277 18797 13280
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 18969 13311 19027 13317
rect 18969 13277 18981 13311
rect 19015 13277 19027 13311
rect 18969 13271 19027 13277
rect 16758 13240 16764 13252
rect 16224 13212 16764 13240
rect 16117 13203 16175 13209
rect 16132 13172 16160 13203
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 18984 13240 19012 13271
rect 19242 13268 19248 13320
rect 19300 13268 19306 13320
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13308 19579 13311
rect 19978 13308 19984 13320
rect 19567 13280 19984 13308
rect 19567 13277 19579 13280
rect 19521 13271 19579 13277
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20254 13268 20260 13320
rect 20312 13268 20318 13320
rect 21376 13308 21404 13472
rect 22465 13447 22523 13453
rect 22465 13444 22477 13447
rect 21468 13416 22477 13444
rect 21468 13388 21496 13416
rect 22465 13413 22477 13416
rect 22511 13444 22523 13447
rect 22830 13444 22836 13456
rect 22511 13416 22836 13444
rect 22511 13413 22523 13416
rect 22465 13407 22523 13413
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 21450 13336 21456 13388
rect 21508 13336 21514 13388
rect 22186 13376 22192 13388
rect 22066 13348 22192 13376
rect 21729 13311 21787 13317
rect 21729 13308 21741 13311
rect 21376 13280 21741 13308
rect 21729 13277 21741 13280
rect 21775 13277 21787 13311
rect 21729 13271 21787 13277
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13308 21971 13311
rect 22066 13308 22094 13348
rect 22186 13336 22192 13348
rect 22244 13376 22250 13388
rect 22646 13376 22652 13388
rect 22244 13348 22652 13376
rect 22244 13336 22250 13348
rect 22646 13336 22652 13348
rect 22704 13376 22710 13388
rect 22704 13348 23336 13376
rect 22704 13336 22710 13348
rect 23308 13320 23336 13348
rect 25038 13336 25044 13388
rect 25096 13376 25102 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 25096 13348 25145 13376
rect 25096 13336 25102 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 21959 13280 22094 13308
rect 22833 13311 22891 13317
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 22833 13277 22845 13311
rect 22879 13277 22891 13311
rect 22833 13271 22891 13277
rect 20272 13240 20300 13268
rect 18984 13212 20300 13240
rect 12406 13144 16160 13172
rect 11103 13141 11115 13144
rect 11057 13135 11115 13141
rect 16574 13132 16580 13184
rect 16632 13172 16638 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 16632 13144 16865 13172
rect 16632 13132 16638 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 16853 13135 16911 13141
rect 19705 13175 19763 13181
rect 19705 13141 19717 13175
rect 19751 13172 19763 13175
rect 19794 13172 19800 13184
rect 19751 13144 19800 13172
rect 19751 13141 19763 13144
rect 19705 13135 19763 13141
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 21818 13132 21824 13184
rect 21876 13132 21882 13184
rect 22848 13172 22876 13271
rect 23290 13268 23296 13320
rect 23348 13268 23354 13320
rect 27614 13268 27620 13320
rect 27672 13308 27678 13320
rect 28813 13311 28871 13317
rect 28813 13308 28825 13311
rect 27672 13280 28825 13308
rect 27672 13268 27678 13280
rect 28813 13277 28825 13280
rect 28859 13277 28871 13311
rect 28813 13271 28871 13277
rect 23750 13172 23756 13184
rect 22848 13144 23756 13172
rect 23750 13132 23756 13144
rect 23808 13172 23814 13184
rect 24026 13172 24032 13184
rect 23808 13144 24032 13172
rect 23808 13132 23814 13144
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 1104 13082 29440 13104
rect 1104 13030 5151 13082
rect 5203 13030 5215 13082
rect 5267 13030 5279 13082
rect 5331 13030 5343 13082
rect 5395 13030 5407 13082
rect 5459 13030 12234 13082
rect 12286 13030 12298 13082
rect 12350 13030 12362 13082
rect 12414 13030 12426 13082
rect 12478 13030 12490 13082
rect 12542 13030 19317 13082
rect 19369 13030 19381 13082
rect 19433 13030 19445 13082
rect 19497 13030 19509 13082
rect 19561 13030 19573 13082
rect 19625 13030 26400 13082
rect 26452 13030 26464 13082
rect 26516 13030 26528 13082
rect 26580 13030 26592 13082
rect 26644 13030 26656 13082
rect 26708 13030 29440 13082
rect 1104 13008 29440 13030
rect 5166 12968 5172 12980
rect 1780 12940 5172 12968
rect 1394 12792 1400 12844
rect 1452 12832 1458 12844
rect 1780 12841 1808 12940
rect 5166 12928 5172 12940
rect 5224 12968 5230 12980
rect 5534 12968 5540 12980
rect 5224 12940 5540 12968
rect 5224 12928 5230 12940
rect 3602 12860 3608 12912
rect 3660 12860 3666 12912
rect 5368 12909 5396 12940
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 7098 12968 7104 12980
rect 5920 12940 7104 12968
rect 5920 12909 5948 12940
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 10410 12968 10416 12980
rect 9508 12940 10416 12968
rect 5353 12903 5411 12909
rect 5353 12869 5365 12903
rect 5399 12869 5411 12903
rect 5353 12863 5411 12869
rect 5905 12903 5963 12909
rect 5905 12869 5917 12903
rect 5951 12869 5963 12903
rect 5905 12863 5963 12869
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 9508 12909 9536 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 10778 12928 10784 12980
rect 10836 12968 10842 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10836 12940 10977 12968
rect 10836 12928 10842 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11848 12940 12173 12968
rect 11848 12928 11854 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 14645 12971 14703 12977
rect 13320 12940 14320 12968
rect 13320 12928 13326 12940
rect 7469 12903 7527 12909
rect 7469 12900 7481 12903
rect 6788 12872 7481 12900
rect 6788 12860 6794 12872
rect 7469 12869 7481 12872
rect 7515 12900 7527 12903
rect 9493 12903 9551 12909
rect 7515 12872 7972 12900
rect 7515 12869 7527 12872
rect 7469 12863 7527 12869
rect 1765 12835 1823 12841
rect 1765 12832 1777 12835
rect 1452 12804 1777 12832
rect 1452 12792 1458 12804
rect 1765 12801 1777 12804
rect 1811 12801 1823 12835
rect 1765 12795 1823 12801
rect 3142 12792 3148 12844
rect 3200 12792 3206 12844
rect 3620 12832 3648 12860
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 3620 12804 3893 12832
rect 3881 12801 3893 12804
rect 3927 12801 3939 12835
rect 3881 12795 3939 12801
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4890 12832 4896 12844
rect 4663 12804 4896 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 2038 12724 2044 12776
rect 2096 12724 2102 12776
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12764 3847 12767
rect 4080 12764 4108 12795
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 6362 12832 6368 12844
rect 6043 12804 6368 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 5644 12764 5672 12795
rect 3835 12736 5672 12764
rect 5828 12764 5856 12795
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 5828 12736 6040 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 3804 12628 3832 12727
rect 6012 12708 6040 12736
rect 5994 12656 6000 12708
rect 6052 12656 6058 12708
rect 6932 12696 6960 12795
rect 7190 12792 7196 12844
rect 7248 12792 7254 12844
rect 7558 12792 7564 12844
rect 7616 12792 7622 12844
rect 7944 12776 7972 12872
rect 9493 12869 9505 12903
rect 9539 12869 9551 12903
rect 9493 12863 9551 12869
rect 10042 12860 10048 12912
rect 10100 12860 10106 12912
rect 11422 12860 11428 12912
rect 11480 12860 11486 12912
rect 14292 12909 14320 12940
rect 14645 12937 14657 12971
rect 14691 12968 14703 12971
rect 15746 12968 15752 12980
rect 14691 12940 15752 12968
rect 14691 12937 14703 12940
rect 14645 12931 14703 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16482 12928 16488 12980
rect 16540 12928 16546 12980
rect 17126 12968 17132 12980
rect 16960 12940 17132 12968
rect 16960 12909 16988 12940
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 18414 12968 18420 12980
rect 18340 12940 18420 12968
rect 18340 12909 18368 12940
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 21177 12971 21235 12977
rect 21177 12937 21189 12971
rect 21223 12968 21235 12971
rect 21634 12968 21640 12980
rect 21223 12940 21640 12968
rect 21223 12937 21235 12940
rect 21177 12931 21235 12937
rect 21634 12928 21640 12940
rect 21692 12928 21698 12980
rect 22278 12928 22284 12980
rect 22336 12928 22342 12980
rect 14001 12903 14059 12909
rect 14001 12900 14013 12903
rect 12268 12872 14013 12900
rect 10502 12792 10508 12844
rect 10560 12792 10566 12844
rect 11440 12832 11468 12860
rect 12268 12841 12296 12872
rect 14001 12869 14013 12872
rect 14047 12869 14059 12903
rect 14001 12863 14059 12869
rect 14277 12903 14335 12909
rect 14277 12869 14289 12903
rect 14323 12869 14335 12903
rect 14277 12863 14335 12869
rect 16945 12903 17003 12909
rect 16945 12869 16957 12903
rect 16991 12869 17003 12903
rect 16945 12863 17003 12869
rect 18325 12903 18383 12909
rect 18325 12869 18337 12903
rect 18371 12869 18383 12903
rect 18325 12863 18383 12869
rect 20714 12860 20720 12912
rect 20772 12900 20778 12912
rect 22005 12903 22063 12909
rect 22005 12900 22017 12903
rect 20772 12872 22017 12900
rect 20772 12860 20778 12872
rect 22005 12869 22017 12872
rect 22051 12869 22063 12903
rect 22296 12900 22324 12928
rect 22922 12900 22928 12912
rect 22296 12872 22928 12900
rect 22005 12863 22063 12869
rect 22922 12860 22928 12872
rect 22980 12900 22986 12912
rect 22980 12872 23152 12900
rect 22980 12860 22986 12872
rect 12253 12835 12311 12841
rect 11440 12804 12204 12832
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 7282 12696 7288 12708
rect 6932 12668 7288 12696
rect 7282 12656 7288 12668
rect 7340 12656 7346 12708
rect 7852 12696 7880 12727
rect 7926 12724 7932 12776
rect 7984 12724 7990 12776
rect 9214 12724 9220 12776
rect 9272 12724 9278 12776
rect 10226 12764 10232 12776
rect 9324 12736 10232 12764
rect 9324 12696 9352 12736
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10520 12764 10548 12792
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 10520 12736 11529 12764
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 12176 12764 12204 12804
rect 12253 12801 12265 12835
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 12434 12792 12440 12844
rect 12492 12792 12498 12844
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 12621 12835 12679 12841
rect 12621 12801 12633 12835
rect 12667 12832 12679 12835
rect 12710 12832 12716 12844
rect 12667 12804 12716 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 12544 12764 12572 12795
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12832 13507 12835
rect 13814 12832 13820 12844
rect 13495 12804 13820 12832
rect 13495 12801 13507 12804
rect 13449 12795 13507 12801
rect 13814 12792 13820 12804
rect 13872 12832 13878 12844
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13872 12804 14105 12832
rect 13872 12792 13878 12804
rect 14093 12801 14105 12804
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14366 12792 14372 12844
rect 14424 12792 14430 12844
rect 14458 12792 14464 12844
rect 14516 12792 14522 12844
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16632 12804 16681 12832
rect 16632 12792 16638 12804
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 17034 12792 17040 12844
rect 17092 12792 17098 12844
rect 17402 12792 17408 12844
rect 17460 12832 17466 12844
rect 18049 12835 18107 12841
rect 18049 12832 18061 12835
rect 17460 12804 18061 12832
rect 17460 12792 17466 12804
rect 18049 12801 18061 12804
rect 18095 12801 18107 12835
rect 19458 12818 21036 12832
rect 18049 12795 18107 12801
rect 19444 12804 21036 12818
rect 14550 12764 14556 12776
rect 12176 12736 14556 12764
rect 11517 12727 11575 12733
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 14734 12724 14740 12776
rect 14792 12724 14798 12776
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 15059 12736 17264 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 7852 12668 9352 12696
rect 3878 12628 3884 12640
rect 3804 12600 3884 12628
rect 3878 12588 3884 12600
rect 3936 12588 3942 12640
rect 4246 12588 4252 12640
rect 4304 12588 4310 12640
rect 6178 12588 6184 12640
rect 6236 12588 6242 12640
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7852 12628 7880 12668
rect 10686 12656 10692 12708
rect 10744 12656 10750 12708
rect 7064 12600 7880 12628
rect 7064 12588 7070 12600
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 10704 12628 10732 12656
rect 7984 12600 10732 12628
rect 7984 12588 7990 12600
rect 12802 12588 12808 12640
rect 12860 12588 12866 12640
rect 14568 12628 14596 12724
rect 17236 12705 17264 12736
rect 17221 12699 17279 12705
rect 17221 12665 17233 12699
rect 17267 12665 17279 12699
rect 17221 12659 17279 12665
rect 17126 12628 17132 12640
rect 14568 12600 17132 12628
rect 17126 12588 17132 12600
rect 17184 12588 17190 12640
rect 19058 12588 19064 12640
rect 19116 12628 19122 12640
rect 19444 12628 19472 12804
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12764 20131 12767
rect 20530 12764 20536 12776
rect 20119 12736 20536 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 21008 12764 21036 12804
rect 21082 12792 21088 12844
rect 21140 12832 21146 12844
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 21140 12804 21465 12832
rect 21140 12792 21146 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 21453 12795 21511 12801
rect 21818 12792 21824 12844
rect 21876 12832 21882 12844
rect 23124 12841 23152 12872
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 21876 12804 23029 12832
rect 21876 12792 21882 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 23109 12835 23167 12841
rect 23109 12801 23121 12835
rect 23155 12801 23167 12835
rect 23109 12795 23167 12801
rect 21174 12764 21180 12776
rect 21008 12736 21180 12764
rect 21174 12724 21180 12736
rect 21232 12724 21238 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12733 21419 12767
rect 21361 12727 21419 12733
rect 21545 12767 21603 12773
rect 21545 12733 21557 12767
rect 21591 12764 21603 12767
rect 21726 12764 21732 12776
rect 21591 12736 21732 12764
rect 21591 12733 21603 12736
rect 21545 12727 21603 12733
rect 21376 12696 21404 12727
rect 21726 12724 21732 12736
rect 21784 12764 21790 12776
rect 22186 12764 22192 12776
rect 21784 12736 22192 12764
rect 21784 12724 21790 12736
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 22738 12724 22744 12776
rect 22796 12724 22802 12776
rect 22646 12696 22652 12708
rect 21376 12668 22652 12696
rect 22646 12656 22652 12668
rect 22704 12656 22710 12708
rect 19116 12600 19472 12628
rect 19116 12588 19122 12600
rect 21634 12588 21640 12640
rect 21692 12628 21698 12640
rect 23017 12631 23075 12637
rect 23017 12628 23029 12631
rect 21692 12600 23029 12628
rect 21692 12588 21698 12600
rect 23017 12597 23029 12600
rect 23063 12597 23075 12631
rect 23017 12591 23075 12597
rect 23385 12631 23443 12637
rect 23385 12597 23397 12631
rect 23431 12628 23443 12631
rect 23474 12628 23480 12640
rect 23431 12600 23480 12628
rect 23431 12597 23443 12600
rect 23385 12591 23443 12597
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 1104 12538 29440 12560
rect 1104 12486 4491 12538
rect 4543 12486 4555 12538
rect 4607 12486 4619 12538
rect 4671 12486 4683 12538
rect 4735 12486 4747 12538
rect 4799 12486 11574 12538
rect 11626 12486 11638 12538
rect 11690 12486 11702 12538
rect 11754 12486 11766 12538
rect 11818 12486 11830 12538
rect 11882 12486 18657 12538
rect 18709 12486 18721 12538
rect 18773 12486 18785 12538
rect 18837 12486 18849 12538
rect 18901 12486 18913 12538
rect 18965 12486 25740 12538
rect 25792 12486 25804 12538
rect 25856 12486 25868 12538
rect 25920 12486 25932 12538
rect 25984 12486 25996 12538
rect 26048 12486 29440 12538
rect 1104 12464 29440 12486
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 2685 12427 2743 12433
rect 2685 12424 2697 12427
rect 2096 12396 2697 12424
rect 2096 12384 2102 12396
rect 2685 12393 2697 12396
rect 2731 12393 2743 12427
rect 3513 12427 3571 12433
rect 3513 12424 3525 12427
rect 2685 12387 2743 12393
rect 2884 12396 3525 12424
rect 2884 12229 2912 12396
rect 3513 12393 3525 12396
rect 3559 12393 3571 12427
rect 5902 12424 5908 12436
rect 3513 12387 3571 12393
rect 4632 12396 5908 12424
rect 4246 12356 4252 12368
rect 2976 12328 4252 12356
rect 2976 12229 3004 12328
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 4632 12297 4660 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6144 12396 6684 12424
rect 6144 12384 6150 12396
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 4617 12291 4675 12297
rect 3375 12260 3648 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 2961 12183 3019 12189
rect 3050 12180 3056 12232
rect 3108 12180 3114 12232
rect 3234 12229 3240 12232
rect 3191 12223 3240 12229
rect 3191 12189 3203 12223
rect 3237 12189 3240 12223
rect 3191 12183 3240 12189
rect 3234 12180 3240 12183
rect 3292 12180 3298 12232
rect 3620 12229 3648 12260
rect 4617 12257 4629 12291
rect 4663 12257 4675 12291
rect 4617 12251 4675 12257
rect 5166 12248 5172 12300
rect 5224 12248 5230 12300
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 6178 12288 6184 12300
rect 5491 12260 6184 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 3651 12192 3924 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 3436 12152 3464 12183
rect 3436 12124 3648 12152
rect 3620 12096 3648 12124
rect 3896 12096 3924 12192
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 5074 12220 5080 12232
rect 4755 12192 5080 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4540 12152 4568 12183
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 6656 12152 6684 12396
rect 6914 12384 6920 12436
rect 6972 12384 6978 12436
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7248 12396 7512 12424
rect 7248 12384 7254 12396
rect 6932 12356 6960 12384
rect 6932 12328 7328 12356
rect 7300 12288 7328 12328
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 7300 12260 7389 12288
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 7484 12288 7512 12396
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 7616 12396 7941 12424
rect 7616 12384 7622 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 10560 12396 10977 12424
rect 10560 12384 10566 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 10965 12387 11023 12393
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 16574 12424 16580 12436
rect 14792 12396 16580 12424
rect 14792 12384 14798 12396
rect 16574 12384 16580 12396
rect 16632 12424 16638 12436
rect 17402 12424 17408 12436
rect 16632 12396 17408 12424
rect 16632 12384 16638 12396
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 15381 12359 15439 12365
rect 15381 12356 15393 12359
rect 13740 12328 15393 12356
rect 7484 12260 7788 12288
rect 7377 12251 7435 12257
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7650 12220 7656 12232
rect 7340 12192 7656 12220
rect 7340 12180 7346 12192
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 7760 12229 7788 12260
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 9272 12260 11805 12288
rect 9272 12248 9278 12260
rect 11793 12257 11805 12260
rect 11839 12288 11851 12291
rect 12066 12288 12072 12300
rect 11839 12260 12072 12288
rect 11839 12257 11851 12260
rect 11793 12251 11851 12257
rect 12066 12248 12072 12260
rect 12124 12288 12130 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 12124 12260 12173 12288
rect 12124 12248 12130 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12288 12495 12291
rect 13740 12288 13768 12328
rect 15381 12325 15393 12328
rect 15427 12325 15439 12359
rect 15381 12319 15439 12325
rect 16209 12359 16267 12365
rect 16209 12325 16221 12359
rect 16255 12356 16267 12359
rect 17218 12356 17224 12368
rect 16255 12328 17224 12356
rect 16255 12325 16267 12328
rect 16209 12319 16267 12325
rect 17218 12316 17224 12328
rect 17276 12316 17282 12368
rect 22922 12316 22928 12368
rect 22980 12356 22986 12368
rect 22980 12328 23060 12356
rect 22980 12316 22986 12328
rect 16390 12288 16396 12300
rect 12483 12260 13768 12288
rect 13832 12260 16396 12288
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 9493 12155 9551 12161
rect 4540 12124 5672 12152
rect 6656 12138 9076 12152
rect 6670 12124 9076 12138
rect 5644 12096 5672 12124
rect 3602 12044 3608 12096
rect 3660 12044 3666 12096
rect 3878 12044 3884 12096
rect 3936 12044 3942 12096
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 5534 12084 5540 12096
rect 4295 12056 5540 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 5626 12044 5632 12096
rect 5684 12044 5690 12096
rect 7006 12044 7012 12096
rect 7064 12044 7070 12096
rect 9048 12084 9076 12124
rect 9493 12121 9505 12155
rect 9539 12152 9551 12155
rect 9766 12152 9772 12164
rect 9539 12124 9772 12152
rect 9539 12121 9551 12124
rect 9493 12115 9551 12121
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 9950 12152 9956 12164
rect 9876 12124 9956 12152
rect 9674 12084 9680 12096
rect 9048 12056 9680 12084
rect 9674 12044 9680 12056
rect 9732 12084 9738 12096
rect 9876 12084 9904 12124
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 11057 12155 11115 12161
rect 11057 12121 11069 12155
rect 11103 12121 11115 12155
rect 11057 12115 11115 12121
rect 9732 12056 9904 12084
rect 9732 12044 9738 12056
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 11072 12084 11100 12115
rect 13446 12112 13452 12164
rect 13504 12112 13510 12164
rect 13832 12084 13860 12260
rect 16390 12248 16396 12260
rect 16448 12248 16454 12300
rect 16758 12248 16764 12300
rect 16816 12248 16822 12300
rect 23032 12297 23060 12328
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12257 23075 12291
rect 23017 12251 23075 12257
rect 14185 12223 14243 12229
rect 14185 12189 14197 12223
rect 14231 12220 14243 12223
rect 14366 12220 14372 12232
rect 14231 12192 14372 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 10192 12056 13860 12084
rect 13909 12087 13967 12093
rect 10192 12044 10198 12056
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14200 12084 14228 12183
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14783 12192 14841 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 15010 12180 15016 12232
rect 15068 12180 15074 12232
rect 15194 12180 15200 12232
rect 15252 12180 15258 12232
rect 16114 12180 16120 12232
rect 16172 12180 16178 12232
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 16942 12220 16948 12232
rect 16724 12192 16948 12220
rect 16724 12180 16730 12192
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 19978 12180 19984 12232
rect 20036 12180 20042 12232
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22465 12223 22523 12229
rect 22465 12220 22477 12223
rect 22244 12192 22477 12220
rect 22244 12180 22250 12192
rect 22465 12189 22477 12192
rect 22511 12189 22523 12223
rect 22465 12183 22523 12189
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 22925 12223 22983 12229
rect 22925 12220 22937 12223
rect 22704 12192 22937 12220
rect 22704 12180 22710 12192
rect 22925 12189 22937 12192
rect 22971 12220 22983 12223
rect 23106 12220 23112 12232
rect 22971 12192 23112 12220
rect 22971 12189 22983 12192
rect 22925 12183 22983 12189
rect 23106 12180 23112 12192
rect 23164 12180 23170 12232
rect 23474 12180 23480 12232
rect 23532 12220 23538 12232
rect 24029 12223 24087 12229
rect 24029 12220 24041 12223
rect 23532 12192 24041 12220
rect 23532 12180 23538 12192
rect 24029 12189 24041 12192
rect 24075 12189 24087 12223
rect 24029 12183 24087 12189
rect 14568 12152 14596 12180
rect 15105 12155 15163 12161
rect 15105 12152 15117 12155
rect 14568 12124 15117 12152
rect 15105 12121 15117 12124
rect 15151 12121 15163 12155
rect 22278 12152 22284 12164
rect 15105 12115 15163 12121
rect 16224 12124 22284 12152
rect 16224 12096 16252 12124
rect 22278 12112 22284 12124
rect 22336 12112 22342 12164
rect 23014 12112 23020 12164
rect 23072 12152 23078 12164
rect 23385 12155 23443 12161
rect 23385 12152 23397 12155
rect 23072 12124 23397 12152
rect 23072 12112 23078 12124
rect 23385 12121 23397 12124
rect 23431 12121 23443 12155
rect 23385 12115 23443 12121
rect 13955 12056 14228 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 16206 12044 16212 12096
rect 16264 12044 16270 12096
rect 19794 12044 19800 12096
rect 19852 12044 19858 12096
rect 23661 12087 23719 12093
rect 23661 12053 23673 12087
rect 23707 12084 23719 12087
rect 23750 12084 23756 12096
rect 23707 12056 23756 12084
rect 23707 12053 23719 12056
rect 23661 12047 23719 12053
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 23842 12044 23848 12096
rect 23900 12044 23906 12096
rect 1104 11994 29440 12016
rect 1104 11942 5151 11994
rect 5203 11942 5215 11994
rect 5267 11942 5279 11994
rect 5331 11942 5343 11994
rect 5395 11942 5407 11994
rect 5459 11942 12234 11994
rect 12286 11942 12298 11994
rect 12350 11942 12362 11994
rect 12414 11942 12426 11994
rect 12478 11942 12490 11994
rect 12542 11942 19317 11994
rect 19369 11942 19381 11994
rect 19433 11942 19445 11994
rect 19497 11942 19509 11994
rect 19561 11942 19573 11994
rect 19625 11942 26400 11994
rect 26452 11942 26464 11994
rect 26516 11942 26528 11994
rect 26580 11942 26592 11994
rect 26644 11942 26656 11994
rect 26708 11942 29440 11994
rect 1104 11920 29440 11942
rect 4065 11883 4123 11889
rect 4065 11849 4077 11883
rect 4111 11880 4123 11883
rect 4430 11880 4436 11892
rect 4111 11852 4436 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4430 11840 4436 11852
rect 4488 11840 4494 11892
rect 5626 11840 5632 11892
rect 5684 11880 5690 11892
rect 7009 11883 7067 11889
rect 7009 11880 7021 11883
rect 5684 11852 7021 11880
rect 5684 11840 5690 11852
rect 7009 11849 7021 11852
rect 7055 11880 7067 11883
rect 7190 11880 7196 11892
rect 7055 11852 7196 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 9858 11880 9864 11892
rect 7708 11852 9864 11880
rect 7708 11840 7714 11852
rect 9858 11840 9864 11852
rect 9916 11880 9922 11892
rect 12710 11880 12716 11892
rect 9916 11852 10916 11880
rect 9916 11840 9922 11852
rect 3142 11772 3148 11824
rect 3200 11772 3206 11824
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11744 1823 11747
rect 2222 11744 2228 11756
rect 1811 11716 2228 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4448 11744 4476 11840
rect 5074 11772 5080 11824
rect 5132 11812 5138 11824
rect 5718 11812 5724 11824
rect 5132 11784 5724 11812
rect 5132 11772 5138 11784
rect 5718 11772 5724 11784
rect 5776 11812 5782 11824
rect 6457 11815 6515 11821
rect 6457 11812 6469 11815
rect 5776 11784 6469 11812
rect 5776 11772 5782 11784
rect 6457 11781 6469 11784
rect 6503 11812 6515 11815
rect 6546 11812 6552 11824
rect 6503 11784 6552 11812
rect 6503 11781 6515 11784
rect 6457 11775 6515 11781
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 4295 11716 4476 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 6362 11744 6368 11756
rect 4948 11716 6368 11744
rect 4948 11704 4954 11716
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7282 11744 7288 11756
rect 6963 11716 7288 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7282 11704 7288 11716
rect 7340 11744 7346 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7340 11716 7573 11744
rect 7340 11704 7346 11716
rect 7561 11713 7573 11716
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 4338 11676 4344 11688
rect 2639 11648 4344 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 2222 11500 2228 11552
rect 2280 11540 2286 11552
rect 2332 11540 2360 11639
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 5442 11676 5448 11688
rect 4632 11648 5448 11676
rect 4632 11608 4660 11648
rect 5442 11636 5448 11648
rect 5500 11676 5506 11688
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 5500 11648 5641 11676
rect 5500 11636 5506 11648
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 5629 11639 5687 11645
rect 4172 11580 4660 11608
rect 4172 11540 4200 11580
rect 5994 11568 6000 11620
rect 6052 11608 6058 11620
rect 6457 11611 6515 11617
rect 6457 11608 6469 11611
rect 6052 11580 6469 11608
rect 6052 11568 6058 11580
rect 6457 11577 6469 11580
rect 6503 11608 6515 11611
rect 7668 11608 7696 11840
rect 9766 11772 9772 11824
rect 9824 11772 9830 11824
rect 10888 11821 10916 11852
rect 12360 11852 12716 11880
rect 12360 11821 12388 11852
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 13814 11840 13820 11892
rect 13872 11840 13878 11892
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 16485 11883 16543 11889
rect 16485 11880 16497 11883
rect 16172 11852 16497 11880
rect 16172 11840 16178 11852
rect 16485 11849 16497 11852
rect 16531 11849 16543 11883
rect 16485 11843 16543 11849
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 19981 11883 20039 11889
rect 19981 11880 19993 11883
rect 19116 11852 19993 11880
rect 19116 11840 19122 11852
rect 19981 11849 19993 11852
rect 20027 11880 20039 11883
rect 20162 11880 20168 11892
rect 20027 11852 20168 11880
rect 20027 11849 20039 11852
rect 19981 11843 20039 11849
rect 20162 11840 20168 11852
rect 20220 11840 20226 11892
rect 20254 11840 20260 11892
rect 20312 11840 20318 11892
rect 22278 11840 22284 11892
rect 22336 11880 22342 11892
rect 22336 11852 23060 11880
rect 22336 11840 22342 11852
rect 10873 11815 10931 11821
rect 10873 11781 10885 11815
rect 10919 11781 10931 11815
rect 10873 11775 10931 11781
rect 12345 11815 12403 11821
rect 12345 11781 12357 11815
rect 12391 11781 12403 11815
rect 12345 11775 12403 11781
rect 13909 11815 13967 11821
rect 13909 11781 13921 11815
rect 13955 11812 13967 11815
rect 14274 11812 14280 11824
rect 13955 11784 14280 11812
rect 13955 11781 13967 11784
rect 13909 11775 13967 11781
rect 14274 11772 14280 11784
rect 14332 11772 14338 11824
rect 16206 11772 16212 11824
rect 16264 11772 16270 11824
rect 20272 11812 20300 11840
rect 23032 11812 23060 11852
rect 23106 11840 23112 11892
rect 23164 11880 23170 11892
rect 23753 11883 23811 11889
rect 23753 11880 23765 11883
rect 23164 11852 23765 11880
rect 23164 11840 23170 11852
rect 23753 11849 23765 11852
rect 23799 11849 23811 11883
rect 23753 11843 23811 11849
rect 24397 11883 24455 11889
rect 24397 11849 24409 11883
rect 24443 11880 24455 11883
rect 25498 11880 25504 11892
rect 24443 11852 25504 11880
rect 24443 11849 24455 11852
rect 24397 11843 24455 11849
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 19536 11784 20300 11812
rect 20456 11784 21864 11812
rect 9784 11744 9812 11772
rect 10459 11747 10517 11753
rect 9784 11716 9904 11744
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11676 8723 11679
rect 8938 11676 8944 11688
rect 8711 11648 8944 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9033 11679 9091 11685
rect 9033 11645 9045 11679
rect 9079 11676 9091 11679
rect 9766 11676 9772 11688
rect 9079 11648 9772 11676
rect 9079 11645 9091 11648
rect 9033 11639 9091 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 9876 11676 9904 11716
rect 10459 11713 10471 11747
rect 10505 11744 10517 11747
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10505 11716 10609 11744
rect 10505 11713 10517 11716
rect 10459 11707 10517 11713
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 12066 11704 12072 11756
rect 12124 11704 12130 11756
rect 13446 11704 13452 11756
rect 13504 11704 13510 11756
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 14642 11744 14648 11756
rect 14148 11716 14648 11744
rect 14148 11704 14154 11716
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15712 11716 15945 11744
rect 15712 11704 15718 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16482 11744 16488 11756
rect 16347 11716 16488 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 13464 11676 13492 11704
rect 13630 11676 13636 11688
rect 9876 11648 13636 11676
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 16132 11676 16160 11707
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 18506 11704 18512 11756
rect 18564 11704 18570 11756
rect 19536 11753 19564 11784
rect 20456 11756 20484 11784
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11713 19579 11747
rect 19521 11707 19579 11713
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11744 19855 11747
rect 20070 11744 20076 11756
rect 19843 11716 20076 11744
rect 19843 11713 19855 11716
rect 19797 11707 19855 11713
rect 20070 11704 20076 11716
rect 20128 11704 20134 11756
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20438 11744 20444 11756
rect 20303 11716 20444 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 20530 11704 20536 11756
rect 20588 11744 20594 11756
rect 21836 11753 21864 11784
rect 22204 11784 22876 11812
rect 23032 11784 25728 11812
rect 22204 11756 22232 11784
rect 21821 11747 21879 11753
rect 20588 11716 21404 11744
rect 20588 11704 20594 11716
rect 16206 11676 16212 11688
rect 16132 11648 16212 11676
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 17037 11679 17095 11685
rect 17037 11645 17049 11679
rect 17083 11676 17095 11679
rect 18046 11676 18052 11688
rect 17083 11648 18052 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 19978 11676 19984 11688
rect 19392 11648 19984 11676
rect 19392 11636 19398 11648
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 6503 11580 7696 11608
rect 6503 11577 6515 11580
rect 6457 11571 6515 11577
rect 16666 11568 16672 11620
rect 16724 11608 16730 11620
rect 18417 11611 18475 11617
rect 18417 11608 18429 11611
rect 16724 11580 18429 11608
rect 16724 11568 16730 11580
rect 18417 11577 18429 11580
rect 18463 11577 18475 11611
rect 18417 11571 18475 11577
rect 2280 11512 4200 11540
rect 2280 11500 2286 11512
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4304 11512 4813 11540
rect 4304 11500 4310 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 4801 11503 4859 11509
rect 7190 11500 7196 11552
rect 7248 11500 7254 11552
rect 7374 11500 7380 11552
rect 7432 11540 7438 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7432 11512 8217 11540
rect 7432 11500 7438 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 14277 11543 14335 11549
rect 14277 11509 14289 11543
rect 14323 11540 14335 11543
rect 14550 11540 14556 11552
rect 14323 11512 14556 11540
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 17586 11500 17592 11552
rect 17644 11500 17650 11552
rect 21376 11540 21404 11716
rect 21821 11713 21833 11747
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 21836 11676 21864 11707
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 22646 11704 22652 11756
rect 22704 11704 22710 11756
rect 22848 11753 22876 11784
rect 22833 11747 22891 11753
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 22922 11704 22928 11756
rect 22980 11744 22986 11756
rect 23477 11747 23535 11753
rect 23477 11744 23489 11747
rect 22980 11716 23489 11744
rect 22980 11704 22986 11716
rect 23477 11713 23489 11716
rect 23523 11744 23535 11747
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23523 11716 23949 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 24026 11704 24032 11756
rect 24084 11744 24090 11756
rect 25700 11753 25728 11784
rect 24213 11747 24271 11753
rect 24213 11744 24225 11747
rect 24084 11716 24225 11744
rect 24084 11704 24090 11716
rect 24213 11713 24225 11716
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11744 25743 11747
rect 26694 11744 26700 11756
rect 25731 11716 26700 11744
rect 25731 11713 25743 11716
rect 25685 11707 25743 11713
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 21836 11648 22232 11676
rect 22204 11608 22232 11648
rect 23290 11636 23296 11688
rect 23348 11636 23354 11688
rect 23569 11679 23627 11685
rect 23569 11645 23581 11679
rect 23615 11645 23627 11679
rect 23569 11639 23627 11645
rect 22462 11608 22468 11620
rect 22204 11580 22468 11608
rect 22462 11568 22468 11580
rect 22520 11608 22526 11620
rect 23584 11608 23612 11639
rect 23750 11636 23756 11688
rect 23808 11676 23814 11688
rect 25593 11679 25651 11685
rect 25593 11676 25605 11679
rect 23808 11648 25605 11676
rect 23808 11636 23814 11648
rect 25593 11645 25605 11648
rect 25639 11645 25651 11679
rect 25593 11639 25651 11645
rect 22520 11580 24624 11608
rect 22520 11568 22526 11580
rect 24596 11552 24624 11580
rect 22370 11540 22376 11552
rect 21376 11512 22376 11540
rect 22370 11500 22376 11512
rect 22428 11540 22434 11552
rect 22646 11540 22652 11552
rect 22428 11512 22652 11540
rect 22428 11500 22434 11512
rect 22646 11500 22652 11512
rect 22704 11540 22710 11552
rect 24118 11540 24124 11552
rect 22704 11512 24124 11540
rect 22704 11500 22710 11512
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 24578 11500 24584 11552
rect 24636 11500 24642 11552
rect 26053 11543 26111 11549
rect 26053 11509 26065 11543
rect 26099 11540 26111 11543
rect 26142 11540 26148 11552
rect 26099 11512 26148 11540
rect 26099 11509 26111 11512
rect 26053 11503 26111 11509
rect 26142 11500 26148 11512
rect 26200 11500 26206 11552
rect 1104 11450 29440 11472
rect 1104 11398 4491 11450
rect 4543 11398 4555 11450
rect 4607 11398 4619 11450
rect 4671 11398 4683 11450
rect 4735 11398 4747 11450
rect 4799 11398 11574 11450
rect 11626 11398 11638 11450
rect 11690 11398 11702 11450
rect 11754 11398 11766 11450
rect 11818 11398 11830 11450
rect 11882 11398 18657 11450
rect 18709 11398 18721 11450
rect 18773 11398 18785 11450
rect 18837 11398 18849 11450
rect 18901 11398 18913 11450
rect 18965 11398 25740 11450
rect 25792 11398 25804 11450
rect 25856 11398 25868 11450
rect 25920 11398 25932 11450
rect 25984 11398 25996 11450
rect 26048 11398 29440 11450
rect 1104 11376 29440 11398
rect 4338 11296 4344 11348
rect 4396 11296 4402 11348
rect 5708 11339 5766 11345
rect 5708 11305 5720 11339
rect 5754 11336 5766 11339
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 5754 11308 7849 11336
rect 5754 11305 5766 11308
rect 5708 11299 5766 11305
rect 7837 11305 7849 11308
rect 7883 11305 7895 11339
rect 7837 11299 7895 11305
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 12158 11336 12164 11348
rect 11296 11308 12164 11336
rect 11296 11296 11302 11308
rect 12158 11296 12164 11308
rect 12216 11336 12222 11348
rect 15194 11336 15200 11348
rect 12216 11308 15200 11336
rect 12216 11296 12222 11308
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 17586 11336 17592 11348
rect 15948 11308 17592 11336
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 7193 11271 7251 11277
rect 4120 11240 4200 11268
rect 4120 11228 4126 11240
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11200 1915 11203
rect 2222 11200 2228 11212
rect 1903 11172 2228 11200
rect 1903 11169 1915 11172
rect 1857 11163 1915 11169
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 3878 11160 3884 11212
rect 3936 11160 3942 11212
rect 3142 11092 3148 11144
rect 3200 11132 3206 11144
rect 3200 11104 3266 11132
rect 3200 11092 3206 11104
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3752 11104 3801 11132
rect 3752 11092 3758 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 2130 11024 2136 11076
rect 2188 11024 2194 11076
rect 3896 11064 3924 11160
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 4172 11141 4200 11240
rect 7193 11237 7205 11271
rect 7239 11268 7251 11271
rect 7282 11268 7288 11280
rect 7239 11240 7288 11268
rect 7239 11237 7251 11240
rect 7193 11231 7251 11237
rect 7282 11228 7288 11240
rect 7340 11228 7346 11280
rect 4356 11172 4660 11200
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4356 11132 4384 11172
rect 4632 11144 4660 11172
rect 5442 11160 5448 11212
rect 5500 11160 5506 11212
rect 6362 11160 6368 11212
rect 6420 11200 6426 11212
rect 10134 11200 10140 11212
rect 6420 11172 10140 11200
rect 6420 11160 6426 11172
rect 4203 11104 4384 11132
rect 4525 11135 4583 11141
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 3896 11036 4077 11064
rect 4065 11033 4077 11036
rect 4111 11033 4123 11067
rect 4540 11064 4568 11095
rect 4614 11092 4620 11144
rect 4672 11092 4678 11144
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7374 11132 7380 11144
rect 7331 11104 7380 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7653 11135 7711 11141
rect 7653 11101 7665 11135
rect 7699 11132 7711 11135
rect 7834 11132 7840 11144
rect 7699 11104 7840 11132
rect 7699 11101 7711 11104
rect 7653 11095 7711 11101
rect 7834 11092 7840 11104
rect 7892 11132 7898 11144
rect 8110 11132 8116 11144
rect 7892 11104 8116 11132
rect 7892 11092 7898 11104
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 9968 11141 9996 11172
rect 10134 11160 10140 11172
rect 10192 11160 10198 11212
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 15948 11132 15976 11308
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 18046 11296 18052 11348
rect 18104 11296 18110 11348
rect 19794 11296 19800 11348
rect 19852 11336 19858 11348
rect 20238 11339 20296 11345
rect 20238 11336 20250 11339
rect 19852 11308 20250 11336
rect 19852 11296 19858 11308
rect 20238 11305 20250 11308
rect 20284 11305 20296 11339
rect 20238 11299 20296 11305
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22646 11336 22652 11348
rect 22152 11308 22652 11336
rect 22152 11296 22158 11308
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 26694 11296 26700 11348
rect 26752 11296 26758 11348
rect 16209 11271 16267 11277
rect 16209 11237 16221 11271
rect 16255 11237 16267 11271
rect 16209 11231 16267 11237
rect 15703 11104 15976 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 6178 11064 6184 11076
rect 4065 11027 4123 11033
rect 4172 11036 5948 11064
rect 3605 10999 3663 11005
rect 3605 10965 3617 10999
rect 3651 10996 3663 10999
rect 4172 10996 4200 11036
rect 5920 11008 5948 11036
rect 6104 11036 6184 11064
rect 3651 10968 4200 10996
rect 3651 10965 3663 10968
rect 3605 10959 3663 10965
rect 4706 10956 4712 11008
rect 4764 10996 4770 11008
rect 5077 10999 5135 11005
rect 5077 10996 5089 10999
rect 4764 10968 5089 10996
rect 4764 10956 4770 10968
rect 5077 10965 5089 10968
rect 5123 10965 5135 10999
rect 5077 10959 5135 10965
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 6104 10996 6132 11036
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 7466 11024 7472 11076
rect 7524 11024 7530 11076
rect 7558 11024 7564 11076
rect 7616 11024 7622 11076
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 10689 11067 10747 11073
rect 10689 11064 10701 11067
rect 8996 11036 10701 11064
rect 8996 11024 9002 11036
rect 10689 11033 10701 11036
rect 10735 11033 10747 11067
rect 10689 11027 10747 11033
rect 15841 11067 15899 11073
rect 15841 11033 15853 11067
rect 15887 11033 15899 11067
rect 15841 11027 15899 11033
rect 7098 10996 7104 11008
rect 6104 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7576 10996 7604 11024
rect 13538 10996 13544 11008
rect 7576 10968 13544 10996
rect 13538 10956 13544 10968
rect 13596 10956 13602 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14550 10996 14556 11008
rect 13872 10968 14556 10996
rect 13872 10956 13878 10968
rect 14550 10956 14556 10968
rect 14608 10956 14614 11008
rect 15856 10996 15884 11027
rect 15930 11024 15936 11076
rect 15988 11024 15994 11076
rect 16224 11064 16252 11231
rect 18874 11228 18880 11280
rect 18932 11268 18938 11280
rect 19334 11268 19340 11280
rect 18932 11240 19340 11268
rect 18932 11228 18938 11240
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 22462 11228 22468 11280
rect 22520 11228 22526 11280
rect 22664 11268 22692 11296
rect 24673 11271 24731 11277
rect 24673 11268 24685 11271
rect 22664 11240 24685 11268
rect 24673 11237 24685 11240
rect 24719 11237 24731 11271
rect 24673 11231 24731 11237
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11200 16359 11203
rect 16574 11200 16580 11212
rect 16347 11172 16580 11200
rect 16347 11169 16359 11172
rect 16301 11163 16359 11169
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 19058 11160 19064 11212
rect 19116 11160 19122 11212
rect 19981 11203 20039 11209
rect 19981 11200 19993 11203
rect 19260 11172 19993 11200
rect 18138 11132 18144 11144
rect 17710 11104 18144 11132
rect 18138 11092 18144 11104
rect 18196 11092 18202 11144
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 18509 11135 18567 11141
rect 18509 11132 18521 11135
rect 18288 11104 18521 11132
rect 18288 11092 18294 11104
rect 18509 11101 18521 11104
rect 18555 11101 18567 11135
rect 18509 11095 18567 11101
rect 18690 11092 18696 11144
rect 18748 11132 18754 11144
rect 19076 11132 19104 11160
rect 19260 11144 19288 11172
rect 19981 11169 19993 11172
rect 20027 11200 20039 11203
rect 22738 11200 22744 11212
rect 20027 11172 22744 11200
rect 20027 11169 20039 11172
rect 19981 11163 20039 11169
rect 22738 11160 22744 11172
rect 22796 11200 22802 11212
rect 24946 11200 24952 11212
rect 22796 11172 24952 11200
rect 22796 11160 22802 11172
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 26712 11200 26740 11296
rect 26881 11203 26939 11209
rect 26881 11200 26893 11203
rect 26712 11172 26893 11200
rect 26881 11169 26893 11172
rect 26927 11169 26939 11203
rect 26881 11163 26939 11169
rect 28902 11160 28908 11212
rect 28960 11200 28966 11212
rect 28997 11203 29055 11209
rect 28997 11200 29009 11203
rect 28960 11172 29009 11200
rect 28960 11160 28966 11172
rect 28997 11169 29009 11172
rect 29043 11169 29055 11203
rect 28997 11163 29055 11169
rect 18748 11104 19104 11132
rect 18748 11092 18754 11104
rect 19242 11092 19248 11144
rect 19300 11092 19306 11144
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 19475 11104 19840 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 16577 11067 16635 11073
rect 16577 11064 16589 11067
rect 16224 11036 16589 11064
rect 16577 11033 16589 11036
rect 16623 11033 16635 11067
rect 16850 11064 16856 11076
rect 16577 11027 16635 11033
rect 16684 11036 16856 11064
rect 16684 10996 16712 11036
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 19444 11064 19472 11095
rect 17880 11036 18460 11064
rect 15856 10968 16712 10996
rect 16758 10956 16764 11008
rect 16816 10996 16822 11008
rect 17880 10996 17908 11036
rect 16816 10968 17908 10996
rect 18432 10996 18460 11036
rect 19076 11036 19472 11064
rect 19076 10996 19104 11036
rect 19702 11024 19708 11076
rect 19760 11024 19766 11076
rect 19812 11064 19840 11104
rect 22094 11092 22100 11144
rect 22152 11092 22158 11144
rect 22281 11135 22339 11141
rect 22281 11101 22293 11135
rect 22327 11101 22339 11135
rect 22281 11095 22339 11101
rect 20346 11064 20352 11076
rect 19812 11036 20352 11064
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 22005 11067 22063 11073
rect 21482 11036 21956 11064
rect 18432 10968 19104 10996
rect 16816 10956 16822 10968
rect 21174 10956 21180 11008
rect 21232 10996 21238 11008
rect 21560 10996 21588 11036
rect 21232 10968 21588 10996
rect 21928 10996 21956 11036
rect 22005 11033 22017 11067
rect 22051 11064 22063 11067
rect 22296 11064 22324 11095
rect 22370 11092 22376 11144
rect 22428 11092 22434 11144
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11132 22707 11135
rect 22922 11132 22928 11144
rect 22695 11104 22928 11132
rect 22695 11101 22707 11104
rect 22649 11095 22707 11101
rect 22462 11064 22468 11076
rect 22051 11036 22468 11064
rect 22051 11033 22063 11036
rect 22005 11027 22063 11033
rect 22462 11024 22468 11036
rect 22520 11064 22526 11076
rect 22664 11064 22692 11095
rect 22922 11092 22928 11104
rect 22980 11092 22986 11144
rect 23385 11135 23443 11141
rect 23385 11101 23397 11135
rect 23431 11132 23443 11135
rect 23431 11104 24900 11132
rect 23431 11101 23443 11104
rect 23385 11095 23443 11101
rect 22520 11036 22692 11064
rect 22520 11024 22526 11036
rect 23106 11024 23112 11076
rect 23164 11064 23170 11076
rect 23566 11064 23572 11076
rect 23164 11036 23572 11064
rect 23164 11024 23170 11036
rect 23566 11024 23572 11036
rect 23624 11024 23630 11076
rect 23658 11024 23664 11076
rect 23716 11064 23722 11076
rect 24029 11067 24087 11073
rect 24029 11064 24041 11067
rect 23716 11036 24041 11064
rect 23716 11024 23722 11036
rect 24029 11033 24041 11036
rect 24075 11033 24087 11067
rect 24029 11027 24087 11033
rect 23934 10996 23940 11008
rect 21928 10968 23940 10996
rect 21232 10956 21238 10968
rect 23934 10956 23940 10968
rect 23992 10956 23998 11008
rect 24044 10996 24072 11027
rect 24118 11024 24124 11076
rect 24176 11064 24182 11076
rect 24397 11067 24455 11073
rect 24397 11064 24409 11067
rect 24176 11036 24409 11064
rect 24176 11024 24182 11036
rect 24397 11033 24409 11036
rect 24443 11033 24455 11067
rect 24397 11027 24455 11033
rect 24302 10996 24308 11008
rect 24044 10968 24308 10996
rect 24302 10956 24308 10968
rect 24360 10956 24366 11008
rect 24872 11005 24900 11104
rect 28718 11092 28724 11144
rect 28776 11092 28782 11144
rect 25222 11024 25228 11076
rect 25280 11024 25286 11076
rect 27062 11064 27068 11076
rect 26450 11036 27068 11064
rect 24857 10999 24915 11005
rect 24857 10965 24869 10999
rect 24903 10965 24915 10999
rect 24857 10959 24915 10965
rect 25038 10956 25044 11008
rect 25096 10996 25102 11008
rect 25314 10996 25320 11008
rect 25096 10968 25320 10996
rect 25096 10956 25102 10968
rect 25314 10956 25320 10968
rect 25372 10996 25378 11008
rect 26528 10996 26556 11036
rect 27062 11024 27068 11036
rect 27120 11024 27126 11076
rect 25372 10968 26556 10996
rect 25372 10956 25378 10968
rect 26786 10956 26792 11008
rect 26844 10996 26850 11008
rect 27525 10999 27583 11005
rect 27525 10996 27537 10999
rect 26844 10968 27537 10996
rect 26844 10956 26850 10968
rect 27525 10965 27537 10968
rect 27571 10965 27583 10999
rect 27525 10959 27583 10965
rect 1104 10906 29440 10928
rect 1104 10854 5151 10906
rect 5203 10854 5215 10906
rect 5267 10854 5279 10906
rect 5331 10854 5343 10906
rect 5395 10854 5407 10906
rect 5459 10854 12234 10906
rect 12286 10854 12298 10906
rect 12350 10854 12362 10906
rect 12414 10854 12426 10906
rect 12478 10854 12490 10906
rect 12542 10854 19317 10906
rect 19369 10854 19381 10906
rect 19433 10854 19445 10906
rect 19497 10854 19509 10906
rect 19561 10854 19573 10906
rect 19625 10854 26400 10906
rect 26452 10854 26464 10906
rect 26516 10854 26528 10906
rect 26580 10854 26592 10906
rect 26644 10854 26656 10906
rect 26708 10854 29440 10906
rect 1104 10832 29440 10854
rect 4062 10752 4068 10804
rect 4120 10752 4126 10804
rect 4154 10752 4160 10804
rect 4212 10752 4218 10804
rect 4706 10792 4712 10804
rect 4632 10764 4712 10792
rect 3973 10727 4031 10733
rect 3973 10693 3985 10727
rect 4019 10724 4031 10727
rect 4080 10724 4108 10752
rect 4019 10696 4108 10724
rect 4019 10693 4031 10696
rect 3973 10687 4031 10693
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3804 10452 3832 10619
rect 4062 10616 4068 10668
rect 4120 10616 4126 10668
rect 4172 10665 4200 10752
rect 4632 10665 4660 10764
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5718 10792 5724 10804
rect 5215 10764 5304 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5276 10736 5304 10764
rect 5460 10764 5724 10792
rect 4801 10727 4859 10733
rect 4801 10724 4813 10727
rect 4724 10696 4813 10724
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 4172 10520 4200 10619
rect 4724 10588 4752 10696
rect 4801 10693 4813 10696
rect 4847 10693 4859 10727
rect 4801 10687 4859 10693
rect 4890 10684 4896 10736
rect 4948 10684 4954 10736
rect 5258 10684 5264 10736
rect 5316 10684 5322 10736
rect 5460 10733 5488 10764
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 5902 10752 5908 10804
rect 5960 10752 5966 10804
rect 5994 10752 6000 10804
rect 6052 10752 6058 10804
rect 9677 10795 9735 10801
rect 9677 10761 9689 10795
rect 9723 10792 9735 10795
rect 9766 10792 9772 10804
rect 9723 10764 9772 10792
rect 9723 10761 9735 10764
rect 9677 10755 9735 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 13998 10752 14004 10804
rect 14056 10792 14062 10804
rect 14461 10795 14519 10801
rect 14461 10792 14473 10795
rect 14056 10764 14473 10792
rect 14056 10752 14062 10764
rect 14461 10761 14473 10764
rect 14507 10761 14519 10795
rect 14461 10755 14519 10761
rect 14550 10752 14556 10804
rect 14608 10752 14614 10804
rect 17865 10795 17923 10801
rect 17865 10761 17877 10795
rect 17911 10792 17923 10795
rect 18506 10792 18512 10804
rect 17911 10764 18512 10792
rect 17911 10761 17923 10764
rect 17865 10755 17923 10761
rect 18506 10752 18512 10764
rect 18564 10792 18570 10804
rect 19981 10795 20039 10801
rect 19981 10792 19993 10795
rect 18564 10764 19993 10792
rect 18564 10752 18570 10764
rect 19981 10761 19993 10764
rect 20027 10761 20039 10795
rect 19981 10755 20039 10761
rect 20346 10752 20352 10804
rect 20404 10752 20410 10804
rect 22741 10795 22799 10801
rect 22741 10761 22753 10795
rect 22787 10792 22799 10795
rect 23014 10792 23020 10804
rect 22787 10764 23020 10792
rect 22787 10761 22799 10764
rect 22741 10755 22799 10761
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 23842 10792 23848 10804
rect 23124 10764 23848 10792
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10693 5503 10727
rect 5445 10687 5503 10693
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 5592 10696 6377 10724
rect 5592 10684 5598 10696
rect 6365 10693 6377 10696
rect 6411 10693 6423 10727
rect 17129 10727 17187 10733
rect 17129 10724 17141 10727
rect 6365 10687 6423 10693
rect 9600 10696 17141 10724
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7190 10656 7196 10668
rect 6687 10628 7196 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 4798 10588 4804 10600
rect 4724 10560 4804 10588
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5000 10588 5028 10619
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 4908 10560 5028 10588
rect 6181 10591 6239 10597
rect 4172 10492 4660 10520
rect 4062 10452 4068 10464
rect 3804 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4341 10455 4399 10461
rect 4341 10452 4353 10455
rect 4212 10424 4353 10452
rect 4212 10412 4218 10424
rect 4341 10421 4353 10424
rect 4387 10421 4399 10455
rect 4632 10452 4660 10492
rect 4908 10452 4936 10560
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 6227 10560 6469 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 6457 10557 6469 10560
rect 6503 10557 6515 10591
rect 7006 10588 7012 10600
rect 6457 10551 6515 10557
rect 6564 10560 7012 10588
rect 5258 10480 5264 10532
rect 5316 10520 5322 10532
rect 5445 10523 5503 10529
rect 5445 10520 5457 10523
rect 5316 10492 5457 10520
rect 5316 10480 5322 10492
rect 5445 10489 5457 10492
rect 5491 10520 5503 10523
rect 5626 10520 5632 10532
rect 5491 10492 5632 10520
rect 5491 10489 5503 10492
rect 5445 10483 5503 10489
rect 5626 10480 5632 10492
rect 5684 10480 5690 10532
rect 5534 10452 5540 10464
rect 4632 10424 5540 10452
rect 4341 10415 4399 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6564 10461 6592 10560
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 6825 10523 6883 10529
rect 6825 10489 6837 10523
rect 6871 10520 6883 10523
rect 9600 10520 9628 10696
rect 17129 10693 17141 10696
rect 17175 10693 17187 10727
rect 17129 10687 17187 10693
rect 17221 10727 17279 10733
rect 17221 10693 17233 10727
rect 17267 10724 17279 10727
rect 19794 10724 19800 10736
rect 17267 10696 19800 10724
rect 17267 10693 17279 10696
rect 17221 10687 17279 10693
rect 19794 10684 19800 10696
rect 19852 10684 19858 10736
rect 20070 10684 20076 10736
rect 20128 10724 20134 10736
rect 23124 10733 23152 10764
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 23934 10752 23940 10804
rect 23992 10792 23998 10804
rect 23992 10764 24256 10792
rect 23992 10752 23998 10764
rect 23109 10727 23167 10733
rect 20128 10696 22508 10724
rect 20128 10684 20134 10696
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 9876 10588 9904 10619
rect 9950 10616 9956 10668
rect 10008 10616 10014 10668
rect 10134 10616 10140 10668
rect 10192 10616 10198 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 9876 10560 9996 10588
rect 6871 10492 9628 10520
rect 6871 10489 6883 10492
rect 6825 10483 6883 10489
rect 9968 10464 9996 10560
rect 10244 10520 10272 10619
rect 10318 10616 10324 10668
rect 10376 10616 10382 10668
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 10428 10628 10517 10656
rect 10428 10600 10456 10628
rect 10505 10625 10517 10628
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 13538 10616 13544 10668
rect 13596 10616 13602 10668
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 13863 10628 14381 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 14369 10625 14381 10628
rect 14415 10656 14427 10659
rect 14918 10656 14924 10668
rect 14415 10628 14924 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 14918 10616 14924 10628
rect 14976 10656 14982 10668
rect 15470 10656 15476 10668
rect 14976 10628 15476 10656
rect 14976 10616 14982 10628
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 16206 10656 16212 10668
rect 15764 10628 16212 10656
rect 10410 10548 10416 10600
rect 10468 10588 10474 10600
rect 11422 10588 11428 10600
rect 10468 10560 11428 10588
rect 10468 10548 10474 10560
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 10594 10520 10600 10532
rect 10244 10492 10600 10520
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 13556 10520 13584 10616
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 13925 10520 13953 10551
rect 13998 10548 14004 10600
rect 14056 10548 14062 10600
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 15764 10588 15792 10628
rect 16206 10616 16212 10628
rect 16264 10656 16270 10668
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 16264 10628 16313 10656
rect 16264 10616 16270 10628
rect 16301 10625 16313 10628
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10656 16543 10659
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16531 10628 16865 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17001 10659 17059 10665
rect 17001 10625 17013 10659
rect 17047 10656 17059 10659
rect 17047 10625 17080 10656
rect 17001 10619 17080 10625
rect 15344 10560 15792 10588
rect 16117 10591 16175 10597
rect 15344 10548 15350 10560
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16316 10588 16344 10619
rect 16758 10588 16764 10600
rect 16316 10560 16764 10588
rect 16117 10551 16175 10557
rect 14185 10523 14243 10529
rect 14185 10520 14197 10523
rect 13556 10492 14197 10520
rect 14185 10489 14197 10492
rect 14231 10520 14243 10523
rect 15930 10520 15936 10532
rect 14231 10492 15936 10520
rect 14231 10489 14243 10492
rect 14185 10483 14243 10489
rect 15930 10480 15936 10492
rect 15988 10520 15994 10532
rect 16132 10520 16160 10551
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 17052 10588 17080 10619
rect 17310 10616 17316 10668
rect 17368 10665 17374 10668
rect 17368 10656 17376 10665
rect 17770 10656 17776 10668
rect 17368 10628 17776 10656
rect 17368 10619 17376 10628
rect 17368 10616 17374 10619
rect 17770 10616 17776 10628
rect 17828 10616 17834 10668
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 17920 10628 17962 10656
rect 17920 10616 17926 10628
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 18104 10628 18245 10656
rect 18104 10616 18110 10628
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10625 18843 10659
rect 18785 10619 18843 10625
rect 18325 10591 18383 10597
rect 17052 10560 17724 10588
rect 17696 10529 17724 10560
rect 18325 10557 18337 10591
rect 18371 10588 18383 10591
rect 18414 10588 18420 10600
rect 18371 10560 18420 10588
rect 18371 10557 18383 10560
rect 18325 10551 18383 10557
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 15988 10492 16160 10520
rect 17681 10523 17739 10529
rect 15988 10480 15994 10492
rect 17681 10489 17693 10523
rect 17727 10489 17739 10523
rect 17681 10483 17739 10489
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10421 6607 10455
rect 6549 10415 6607 10421
rect 9950 10412 9956 10464
rect 10008 10412 10014 10464
rect 10042 10412 10048 10464
rect 10100 10452 10106 10464
rect 10410 10452 10416 10464
rect 10100 10424 10416 10452
rect 10100 10412 10106 10424
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10689 10455 10747 10461
rect 10689 10452 10701 10455
rect 10560 10424 10701 10452
rect 10560 10412 10566 10424
rect 10689 10421 10701 10424
rect 10735 10421 10747 10455
rect 10689 10415 10747 10421
rect 13538 10412 13544 10464
rect 13596 10412 13602 10464
rect 14734 10412 14740 10464
rect 14792 10412 14798 10464
rect 17402 10412 17408 10464
rect 17460 10452 17466 10464
rect 17497 10455 17555 10461
rect 17497 10452 17509 10455
rect 17460 10424 17509 10452
rect 17460 10412 17466 10424
rect 17497 10421 17509 10424
rect 17543 10421 17555 10455
rect 18616 10452 18644 10619
rect 18800 10588 18828 10619
rect 18966 10616 18972 10668
rect 19024 10616 19030 10668
rect 19058 10616 19064 10668
rect 19116 10656 19122 10668
rect 19153 10659 19211 10665
rect 19153 10656 19165 10659
rect 19116 10628 19165 10656
rect 19116 10616 19122 10628
rect 19153 10625 19165 10628
rect 19199 10625 19211 10659
rect 19153 10619 19211 10625
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 20088 10656 20116 10684
rect 19291 10628 20116 10656
rect 20165 10659 20223 10665
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 20165 10625 20177 10659
rect 20211 10656 20223 10659
rect 20530 10656 20536 10668
rect 20211 10628 20536 10656
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 20640 10665 20668 10696
rect 22480 10668 22508 10696
rect 23109 10693 23121 10727
rect 23155 10693 23167 10727
rect 23109 10687 23167 10693
rect 20625 10659 20683 10665
rect 20625 10625 20637 10659
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10656 20867 10659
rect 22002 10656 22008 10668
rect 20855 10628 22008 10656
rect 20855 10625 20867 10628
rect 20809 10619 20867 10625
rect 19705 10591 19763 10597
rect 18800 10560 19104 10588
rect 19076 10520 19104 10560
rect 19705 10557 19717 10591
rect 19751 10588 19763 10591
rect 20438 10588 20444 10600
rect 19751 10560 20444 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 19720 10520 19748 10551
rect 20438 10548 20444 10560
rect 20496 10588 20502 10600
rect 20824 10588 20852 10619
rect 22002 10616 22008 10628
rect 22060 10656 22066 10668
rect 22097 10659 22155 10665
rect 22097 10656 22109 10659
rect 22060 10628 22109 10656
rect 22060 10616 22066 10628
rect 22097 10625 22109 10628
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 22462 10616 22468 10668
rect 22520 10656 22526 10668
rect 22557 10659 22615 10665
rect 22557 10656 22569 10659
rect 22520 10628 22569 10656
rect 22520 10616 22526 10628
rect 22557 10625 22569 10628
rect 22603 10625 22615 10659
rect 22557 10619 22615 10625
rect 22738 10616 22744 10668
rect 22796 10656 22802 10668
rect 22833 10659 22891 10665
rect 22833 10656 22845 10659
rect 22796 10628 22845 10656
rect 22796 10616 22802 10628
rect 22833 10625 22845 10628
rect 22879 10625 22891 10659
rect 24228 10656 24256 10764
rect 25222 10752 25228 10804
rect 25280 10792 25286 10804
rect 25409 10795 25467 10801
rect 25409 10792 25421 10795
rect 25280 10764 25421 10792
rect 25280 10752 25286 10764
rect 25409 10761 25421 10764
rect 25455 10761 25467 10795
rect 26145 10795 26203 10801
rect 26145 10792 26157 10795
rect 25409 10755 25467 10761
rect 25608 10764 26157 10792
rect 24578 10684 24584 10736
rect 24636 10724 24642 10736
rect 24857 10727 24915 10733
rect 24857 10724 24869 10727
rect 24636 10696 24869 10724
rect 24636 10684 24642 10696
rect 24857 10693 24869 10696
rect 24903 10693 24915 10727
rect 24857 10687 24915 10693
rect 25038 10684 25044 10736
rect 25096 10684 25102 10736
rect 25056 10656 25084 10684
rect 24228 10642 25084 10656
rect 24242 10628 25084 10642
rect 25608 10656 25636 10764
rect 26145 10761 26157 10764
rect 26191 10761 26203 10795
rect 26145 10755 26203 10761
rect 25774 10684 25780 10736
rect 25832 10724 25838 10736
rect 25961 10727 26019 10733
rect 25961 10724 25973 10727
rect 25832 10696 25973 10724
rect 25832 10684 25838 10696
rect 25961 10693 25973 10696
rect 26007 10724 26019 10727
rect 26007 10696 26740 10724
rect 26007 10693 26019 10696
rect 25961 10687 26019 10693
rect 25685 10659 25743 10665
rect 25685 10656 25697 10659
rect 25608 10628 25697 10656
rect 22833 10619 22891 10625
rect 25685 10625 25697 10628
rect 25731 10625 25743 10659
rect 25685 10619 25743 10625
rect 26142 10616 26148 10668
rect 26200 10656 26206 10668
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 26200 10628 26341 10656
rect 26200 10616 26206 10628
rect 26329 10625 26341 10628
rect 26375 10625 26387 10659
rect 26329 10619 26387 10625
rect 26418 10616 26424 10668
rect 26476 10616 26482 10668
rect 26510 10616 26516 10668
rect 26568 10616 26574 10668
rect 26602 10616 26608 10668
rect 26660 10616 26666 10668
rect 26712 10665 26740 10696
rect 26697 10659 26755 10665
rect 26697 10625 26709 10659
rect 26743 10625 26755 10659
rect 26697 10619 26755 10625
rect 26789 10659 26847 10665
rect 26789 10625 26801 10659
rect 26835 10625 26847 10659
rect 26789 10619 26847 10625
rect 20496 10560 20852 10588
rect 20496 10548 20502 10560
rect 20898 10548 20904 10600
rect 20956 10588 20962 10600
rect 22186 10588 22192 10600
rect 20956 10560 22192 10588
rect 20956 10548 20962 10560
rect 22186 10548 22192 10560
rect 22244 10588 22250 10600
rect 22373 10591 22431 10597
rect 22373 10588 22385 10591
rect 22244 10560 22385 10588
rect 22244 10548 22250 10560
rect 22373 10557 22385 10560
rect 22419 10557 22431 10591
rect 22373 10551 22431 10557
rect 25590 10548 25596 10600
rect 25648 10548 25654 10600
rect 26053 10591 26111 10597
rect 26053 10557 26065 10591
rect 26099 10588 26111 10591
rect 26620 10588 26648 10616
rect 26099 10560 26648 10588
rect 26099 10557 26111 10560
rect 26053 10551 26111 10557
rect 19076 10492 19748 10520
rect 20530 10480 20536 10532
rect 20588 10480 20594 10532
rect 24302 10480 24308 10532
rect 24360 10520 24366 10532
rect 26804 10520 26832 10619
rect 24360 10492 26832 10520
rect 24360 10480 24366 10492
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 18616 10424 19625 10452
rect 17497 10415 17555 10421
rect 19613 10421 19625 10424
rect 19659 10452 19671 10455
rect 19886 10452 19892 10464
rect 19659 10424 19892 10452
rect 19659 10421 19671 10424
rect 19613 10415 19671 10421
rect 19886 10412 19892 10424
rect 19944 10452 19950 10464
rect 20548 10452 20576 10480
rect 19944 10424 20576 10452
rect 19944 10412 19950 10424
rect 22370 10412 22376 10464
rect 22428 10412 22434 10464
rect 1104 10362 29440 10384
rect 1104 10310 4491 10362
rect 4543 10310 4555 10362
rect 4607 10310 4619 10362
rect 4671 10310 4683 10362
rect 4735 10310 4747 10362
rect 4799 10310 11574 10362
rect 11626 10310 11638 10362
rect 11690 10310 11702 10362
rect 11754 10310 11766 10362
rect 11818 10310 11830 10362
rect 11882 10310 18657 10362
rect 18709 10310 18721 10362
rect 18773 10310 18785 10362
rect 18837 10310 18849 10362
rect 18901 10310 18913 10362
rect 18965 10310 25740 10362
rect 25792 10310 25804 10362
rect 25856 10310 25868 10362
rect 25920 10310 25932 10362
rect 25984 10310 25996 10362
rect 26048 10310 29440 10362
rect 1104 10288 29440 10310
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 4120 10220 4721 10248
rect 4120 10208 4126 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 10042 10248 10048 10260
rect 9824 10220 10048 10248
rect 9824 10208 9830 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10192 10220 10609 10248
rect 10192 10208 10198 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 12618 10248 12624 10260
rect 11020 10220 12624 10248
rect 11020 10208 11026 10220
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13538 10208 13544 10260
rect 13596 10257 13602 10260
rect 13596 10251 13621 10257
rect 13609 10217 13621 10251
rect 13596 10211 13621 10217
rect 13596 10208 13602 10211
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 17310 10248 17316 10260
rect 16540 10220 17316 10248
rect 16540 10208 16546 10220
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 19150 10248 19156 10260
rect 18196 10220 19156 10248
rect 18196 10208 18202 10220
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 20254 10208 20260 10260
rect 20312 10248 20318 10260
rect 20717 10251 20775 10257
rect 20717 10248 20729 10251
rect 20312 10220 20729 10248
rect 20312 10208 20318 10220
rect 20717 10217 20729 10220
rect 20763 10217 20775 10251
rect 20717 10211 20775 10217
rect 22646 10208 22652 10260
rect 22704 10208 22710 10260
rect 22833 10251 22891 10257
rect 22833 10217 22845 10251
rect 22879 10217 22891 10251
rect 22833 10211 22891 10217
rect 9416 10152 12664 10180
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 9416 10053 9444 10152
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10284 10084 10640 10112
rect 10284 10072 10290 10084
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9858 10004 9864 10056
rect 9916 10004 9922 10056
rect 10042 10004 10048 10056
rect 10100 10004 10106 10056
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10044 10195 10047
rect 10318 10044 10324 10056
rect 10183 10016 10324 10044
rect 10183 10013 10195 10016
rect 10137 10007 10195 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10612 10044 10640 10084
rect 10686 10072 10692 10124
rect 10744 10072 10750 10124
rect 11333 10115 11391 10121
rect 11333 10112 11345 10115
rect 10796 10084 11345 10112
rect 10796 10044 10824 10084
rect 11333 10081 11345 10084
rect 11379 10081 11391 10115
rect 11333 10075 11391 10081
rect 11974 10072 11980 10124
rect 12032 10072 12038 10124
rect 12636 10112 12664 10152
rect 13262 10140 13268 10192
rect 13320 10140 13326 10192
rect 13648 10152 16712 10180
rect 13280 10112 13308 10140
rect 12636 10084 13308 10112
rect 10612 10016 10824 10044
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10044 10931 10047
rect 10962 10044 10968 10056
rect 10919 10016 10968 10044
rect 10919 10013 10931 10016
rect 10873 10007 10931 10013
rect 9493 9979 9551 9985
rect 9493 9945 9505 9979
rect 9539 9976 9551 9979
rect 9950 9976 9956 9988
rect 9539 9948 9956 9976
rect 9539 9945 9551 9948
rect 9493 9939 9551 9945
rect 9950 9936 9956 9948
rect 10008 9976 10014 9988
rect 10888 9976 10916 10007
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11149 10047 11207 10053
rect 11149 10044 11161 10047
rect 11112 10016 11161 10044
rect 11112 10004 11118 10016
rect 11149 10013 11161 10016
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11247 10047 11305 10053
rect 11247 10013 11259 10047
rect 11293 10013 11305 10047
rect 11247 10007 11305 10013
rect 11256 9976 11284 10007
rect 11422 10004 11428 10056
rect 11480 10046 11486 10056
rect 12636 10053 12664 10084
rect 11701 10047 11759 10053
rect 11480 10018 11523 10046
rect 11480 10004 11486 10018
rect 11701 10013 11713 10047
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10013 12679 10047
rect 12621 10007 12679 10013
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 13648 10044 13676 10152
rect 16574 10072 16580 10124
rect 16632 10072 16638 10124
rect 16684 10112 16712 10152
rect 17862 10140 17868 10192
rect 17920 10180 17926 10192
rect 20272 10180 20300 10208
rect 17920 10152 20300 10180
rect 20349 10183 20407 10189
rect 17920 10140 17926 10152
rect 20349 10149 20361 10183
rect 20395 10180 20407 10183
rect 20898 10180 20904 10192
rect 20395 10152 20904 10180
rect 20395 10149 20407 10152
rect 20349 10143 20407 10149
rect 18230 10112 18236 10124
rect 16684 10084 18236 10112
rect 18230 10072 18236 10084
rect 18288 10112 18294 10124
rect 19058 10112 19064 10124
rect 18288 10084 19064 10112
rect 18288 10072 18294 10084
rect 19058 10072 19064 10084
rect 19116 10112 19122 10124
rect 20364 10112 20392 10143
rect 20898 10140 20904 10152
rect 20956 10140 20962 10192
rect 19116 10084 20392 10112
rect 19116 10072 19122 10084
rect 20438 10072 20444 10124
rect 20496 10072 20502 10124
rect 22664 10112 22692 10208
rect 22296 10084 22692 10112
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 12851 10016 13676 10044
rect 13740 10016 14289 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 10008 9948 10916 9976
rect 10980 9948 11284 9976
rect 10008 9936 10014 9948
rect 9030 9868 9036 9920
rect 9088 9868 9094 9920
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 10870 9908 10876 9920
rect 10376 9880 10876 9908
rect 10376 9868 10382 9880
rect 10870 9868 10876 9880
rect 10928 9908 10934 9920
rect 10980 9908 11008 9948
rect 11330 9936 11336 9988
rect 11388 9936 11394 9988
rect 11716 9976 11744 10007
rect 12820 9976 12848 10007
rect 11716 9948 12848 9976
rect 13354 9936 13360 9988
rect 13412 9936 13418 9988
rect 10928 9880 11008 9908
rect 11057 9911 11115 9917
rect 10928 9868 10934 9880
rect 11057 9877 11069 9911
rect 11103 9908 11115 9911
rect 11348 9908 11376 9936
rect 11103 9880 11376 9908
rect 11103 9877 11115 9880
rect 11057 9871 11115 9877
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 12124 9880 12817 9908
rect 12124 9868 12130 9880
rect 12805 9877 12817 9880
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13740 9917 13768 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 15286 10004 15292 10056
rect 15344 10004 15350 10056
rect 15378 10004 15384 10056
rect 15436 10004 15442 10056
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 15657 10047 15715 10053
rect 15528 10016 15573 10044
rect 15528 10004 15534 10016
rect 15657 10013 15669 10047
rect 15703 10013 15715 10047
rect 15657 10007 15715 10013
rect 15887 10047 15945 10053
rect 15887 10013 15899 10047
rect 15933 10044 15945 10047
rect 16482 10044 16488 10056
rect 15933 10016 16488 10044
rect 15933 10013 15945 10016
rect 15887 10007 15945 10013
rect 15304 9976 15332 10004
rect 15672 9976 15700 10007
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 18138 10044 18144 10056
rect 17986 10016 18144 10044
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18417 10047 18475 10053
rect 18417 10044 18429 10047
rect 18380 10016 18429 10044
rect 18380 10004 18386 10016
rect 18417 10013 18429 10016
rect 18463 10013 18475 10047
rect 18417 10007 18475 10013
rect 19886 10004 19892 10056
rect 19944 10004 19950 10056
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20070 10044 20076 10056
rect 20027 10016 20076 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 22296 10053 22324 10084
rect 22281 10047 22339 10053
rect 22281 10013 22293 10047
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10044 22523 10047
rect 22848 10044 22876 10211
rect 22922 10208 22928 10260
rect 22980 10208 22986 10260
rect 23293 10251 23351 10257
rect 23293 10217 23305 10251
rect 23339 10248 23351 10251
rect 23382 10248 23388 10260
rect 23339 10220 23388 10248
rect 23339 10217 23351 10220
rect 23293 10211 23351 10217
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 25590 10208 25596 10260
rect 25648 10248 25654 10260
rect 25869 10251 25927 10257
rect 25869 10248 25881 10251
rect 25648 10220 25881 10248
rect 25648 10208 25654 10220
rect 25869 10217 25881 10220
rect 25915 10217 25927 10251
rect 25869 10211 25927 10217
rect 22940 10056 22968 10208
rect 23017 10115 23075 10121
rect 23017 10081 23029 10115
rect 23063 10112 23075 10115
rect 23198 10112 23204 10124
rect 23063 10084 23204 10112
rect 23063 10081 23075 10084
rect 23017 10075 23075 10081
rect 23198 10072 23204 10084
rect 23256 10072 23262 10124
rect 26510 10112 26516 10124
rect 26068 10084 26516 10112
rect 22511 10016 22876 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 15304 9948 15700 9976
rect 15749 9979 15807 9985
rect 15749 9945 15761 9979
rect 15795 9976 15807 9979
rect 15795 9948 16804 9976
rect 15795 9945 15807 9948
rect 15749 9939 15807 9945
rect 13557 9911 13615 9917
rect 13557 9908 13569 9911
rect 13136 9880 13569 9908
rect 13136 9868 13142 9880
rect 13557 9877 13569 9880
rect 13603 9877 13615 9911
rect 13557 9871 13615 9877
rect 13725 9911 13783 9917
rect 13725 9877 13737 9911
rect 13771 9877 13783 9911
rect 13725 9871 13783 9877
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13872 9880 14105 9908
rect 13872 9868 13878 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 15252 9880 16037 9908
rect 15252 9868 15258 9880
rect 16025 9877 16037 9880
rect 16071 9877 16083 9911
rect 16776 9908 16804 9948
rect 16850 9936 16856 9988
rect 16908 9936 16914 9988
rect 22186 9976 22192 9988
rect 18248 9948 22192 9976
rect 18248 9908 18276 9948
rect 22186 9936 22192 9948
rect 22244 9976 22250 9988
rect 22480 9976 22508 10007
rect 22922 10004 22928 10056
rect 22980 10044 22986 10056
rect 26068 10053 26096 10084
rect 26510 10072 26516 10084
rect 26568 10112 26574 10124
rect 26878 10112 26884 10124
rect 26568 10084 26884 10112
rect 26568 10072 26574 10084
rect 26878 10072 26884 10084
rect 26936 10072 26942 10124
rect 23109 10047 23167 10053
rect 23109 10044 23121 10047
rect 22980 10016 23121 10044
rect 22980 10004 22986 10016
rect 23109 10013 23121 10016
rect 23155 10013 23167 10047
rect 23109 10007 23167 10013
rect 26053 10047 26111 10053
rect 26053 10013 26065 10047
rect 26099 10013 26111 10047
rect 26053 10007 26111 10013
rect 26145 10047 26203 10053
rect 26145 10013 26157 10047
rect 26191 10044 26203 10047
rect 26418 10044 26424 10056
rect 26191 10016 26424 10044
rect 26191 10013 26203 10016
rect 26145 10007 26203 10013
rect 22244 9948 22508 9976
rect 22244 9936 22250 9948
rect 22830 9936 22836 9988
rect 22888 9936 22894 9988
rect 25869 9979 25927 9985
rect 25869 9945 25881 9979
rect 25915 9945 25927 9979
rect 25869 9939 25927 9945
rect 16776 9880 18276 9908
rect 16025 9871 16083 9877
rect 18322 9868 18328 9920
rect 18380 9868 18386 9920
rect 19058 9868 19064 9920
rect 19116 9868 19122 9920
rect 22370 9868 22376 9920
rect 22428 9868 22434 9920
rect 25884 9908 25912 9939
rect 26252 9920 26280 10016
rect 26418 10004 26424 10016
rect 26476 10004 26482 10056
rect 26142 9908 26148 9920
rect 25884 9880 26148 9908
rect 26142 9868 26148 9880
rect 26200 9868 26206 9920
rect 26234 9868 26240 9920
rect 26292 9868 26298 9920
rect 1104 9818 29440 9840
rect 1104 9766 5151 9818
rect 5203 9766 5215 9818
rect 5267 9766 5279 9818
rect 5331 9766 5343 9818
rect 5395 9766 5407 9818
rect 5459 9766 12234 9818
rect 12286 9766 12298 9818
rect 12350 9766 12362 9818
rect 12414 9766 12426 9818
rect 12478 9766 12490 9818
rect 12542 9766 19317 9818
rect 19369 9766 19381 9818
rect 19433 9766 19445 9818
rect 19497 9766 19509 9818
rect 19561 9766 19573 9818
rect 19625 9766 26400 9818
rect 26452 9766 26464 9818
rect 26516 9766 26528 9818
rect 26580 9766 26592 9818
rect 26644 9766 26656 9818
rect 26708 9766 29440 9818
rect 1104 9744 29440 9766
rect 3697 9707 3755 9713
rect 3697 9673 3709 9707
rect 3743 9704 3755 9707
rect 3743 9676 4108 9704
rect 3743 9673 3755 9676
rect 3697 9667 3755 9673
rect 4080 9648 4108 9676
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 9677 9707 9735 9713
rect 6052 9676 6914 9704
rect 6052 9664 6058 9676
rect 2222 9636 2228 9648
rect 1964 9608 2228 9636
rect 1964 9577 1992 9608
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 4120 9608 5580 9636
rect 4120 9596 4126 9608
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 4890 9528 4896 9580
rect 4948 9528 4954 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 5031 9540 5089 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 4154 9500 4160 9512
rect 2271 9472 4160 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 4908 9500 4936 9528
rect 5276 9500 5304 9531
rect 4908 9472 5304 9500
rect 5368 9500 5396 9531
rect 5442 9528 5448 9580
rect 5500 9528 5506 9580
rect 5552 9568 5580 9608
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 6457 9639 6515 9645
rect 6457 9636 6469 9639
rect 6328 9608 6469 9636
rect 6328 9596 6334 9608
rect 6457 9605 6469 9608
rect 6503 9605 6515 9639
rect 6886 9636 6914 9676
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 9950 9704 9956 9716
rect 9723 9676 9956 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 7009 9639 7067 9645
rect 7009 9636 7021 9639
rect 6886 9608 7021 9636
rect 6457 9599 6515 9605
rect 7009 9605 7021 9608
rect 7055 9605 7067 9639
rect 9692 9636 9720 9667
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10502 9704 10508 9716
rect 10152 9676 10508 9704
rect 10152 9645 10180 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 10594 9664 10600 9716
rect 10652 9664 10658 9716
rect 10686 9664 10692 9716
rect 10744 9664 10750 9716
rect 10870 9664 10876 9716
rect 10928 9664 10934 9716
rect 16850 9664 16856 9716
rect 16908 9704 16914 9716
rect 17221 9707 17279 9713
rect 17221 9704 17233 9707
rect 16908 9676 17233 9704
rect 16908 9664 16914 9676
rect 17221 9673 17233 9676
rect 17267 9673 17279 9707
rect 17221 9667 17279 9673
rect 17773 9707 17831 9713
rect 17773 9673 17785 9707
rect 17819 9704 17831 9707
rect 18506 9704 18512 9716
rect 17819 9676 18512 9704
rect 17819 9673 17831 9676
rect 17773 9667 17831 9673
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 18966 9664 18972 9716
rect 19024 9704 19030 9716
rect 21450 9704 21456 9716
rect 19024 9676 21456 9704
rect 19024 9664 19030 9676
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 7009 9599 7067 9605
rect 8772 9608 9720 9636
rect 10137 9639 10195 9645
rect 8772 9577 8800 9608
rect 10137 9605 10149 9639
rect 10183 9605 10195 9639
rect 10137 9599 10195 9605
rect 10226 9596 10232 9648
rect 10284 9596 10290 9648
rect 10367 9639 10425 9645
rect 10367 9605 10379 9639
rect 10413 9636 10425 9639
rect 10704 9636 10732 9664
rect 10413 9608 10732 9636
rect 10888 9636 10916 9664
rect 11149 9639 11207 9645
rect 10888 9608 11100 9636
rect 10413 9605 10425 9608
rect 10367 9599 10425 9605
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 5552 9540 6929 9568
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9030 9528 9036 9580
rect 9088 9568 9094 9580
rect 9309 9571 9367 9577
rect 9309 9568 9321 9571
rect 9088 9540 9321 9568
rect 9088 9528 9094 9540
rect 9309 9537 9321 9540
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9539 9571 9597 9577
rect 9539 9537 9551 9571
rect 9585 9568 9597 9571
rect 9858 9568 9864 9580
rect 9585 9540 9864 9568
rect 9585 9537 9597 9540
rect 9539 9531 9597 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10045 9571 10103 9577
rect 10045 9568 10057 9571
rect 10008 9540 10057 9568
rect 10008 9528 10014 9540
rect 10045 9537 10057 9540
rect 10091 9537 10103 9571
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 10045 9531 10103 9537
rect 10428 9540 10517 9568
rect 6178 9500 6184 9512
rect 5368 9472 6184 9500
rect 4341 9463 4399 9469
rect 4356 9376 4384 9463
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 8711 9472 8800 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 6457 9435 6515 9441
rect 6457 9432 6469 9435
rect 5552 9404 6469 9432
rect 4338 9324 4344 9376
rect 4396 9324 4402 9376
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5552 9364 5580 9404
rect 6457 9401 6469 9404
rect 6503 9401 6515 9435
rect 6457 9395 6515 9401
rect 5132 9336 5580 9364
rect 5132 9324 5138 9336
rect 5626 9324 5632 9376
rect 5684 9324 5690 9376
rect 6472 9364 6500 9395
rect 6546 9392 6552 9444
rect 6604 9432 6610 9444
rect 8481 9435 8539 9441
rect 8481 9432 8493 9435
rect 6604 9404 8493 9432
rect 6604 9392 6610 9404
rect 8481 9401 8493 9404
rect 8527 9401 8539 9435
rect 8481 9395 8539 9401
rect 6638 9364 6644 9376
rect 6472 9336 6644 9364
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7190 9324 7196 9376
rect 7248 9324 7254 9376
rect 8772 9364 8800 9472
rect 8846 9460 8852 9512
rect 8904 9460 8910 9512
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 8956 9432 8984 9463
rect 9122 9460 9128 9512
rect 9180 9460 9186 9512
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9674 9500 9680 9512
rect 9447 9472 9680 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9500 9827 9503
rect 10318 9500 10324 9512
rect 9815 9472 10324 9500
rect 9815 9469 9827 9472
rect 9769 9463 9827 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 9861 9435 9919 9441
rect 9861 9432 9873 9435
rect 8956 9404 9873 9432
rect 9861 9401 9873 9404
rect 9907 9401 9919 9435
rect 9861 9395 9919 9401
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10428 9432 10456 9540
rect 10505 9537 10517 9540
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10643 9540 10824 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 10192 9404 10456 9432
rect 10192 9392 10198 9404
rect 10686 9392 10692 9444
rect 10744 9392 10750 9444
rect 10042 9364 10048 9376
rect 8772 9336 10048 9364
rect 10042 9324 10048 9336
rect 10100 9364 10106 9376
rect 10704 9364 10732 9392
rect 10100 9336 10732 9364
rect 10796 9364 10824 9540
rect 10888 9509 10916 9608
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 11072 9568 11100 9608
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 11330 9636 11336 9648
rect 11195 9608 11336 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 11330 9596 11336 9608
rect 11388 9636 11394 9648
rect 11388 9608 11928 9636
rect 11388 9596 11394 9608
rect 11900 9577 11928 9608
rect 13170 9596 13176 9648
rect 13228 9596 13234 9648
rect 13446 9636 13452 9648
rect 13280 9608 13452 9636
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 11072 9540 11253 9568
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 11974 9528 11980 9580
rect 12032 9568 12038 9580
rect 13280 9577 13308 9608
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 13541 9639 13599 9645
rect 13541 9605 13553 9639
rect 13587 9636 13599 9639
rect 13814 9636 13820 9648
rect 13587 9608 13820 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14274 9596 14280 9648
rect 14332 9596 14338 9648
rect 16684 9608 19104 9636
rect 16684 9577 16712 9608
rect 19076 9580 19104 9608
rect 26878 9596 26884 9648
rect 26936 9636 26942 9648
rect 26936 9608 28028 9636
rect 26936 9596 26942 9608
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12032 9540 12541 9568
rect 12032 9528 12038 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 16669 9571 16727 9577
rect 16669 9537 16681 9571
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16850 9528 16856 9580
rect 16908 9528 16914 9580
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 11054 9460 11060 9512
rect 11112 9460 11118 9512
rect 10965 9435 11023 9441
rect 10965 9401 10977 9435
rect 11011 9432 11023 9435
rect 11072 9432 11100 9460
rect 11011 9404 11100 9432
rect 11011 9401 11023 9404
rect 10965 9395 11023 9401
rect 11992 9364 12020 9528
rect 13998 9460 14004 9512
rect 14056 9500 14062 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 14056 9472 15301 9500
rect 14056 9460 14062 9472
rect 15289 9469 15301 9472
rect 15335 9500 15347 9503
rect 16574 9500 16580 9512
rect 15335 9472 16580 9500
rect 15335 9469 15347 9472
rect 15289 9463 15347 9469
rect 16574 9460 16580 9472
rect 16632 9500 16638 9512
rect 16960 9500 16988 9531
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 17770 9571 17828 9577
rect 17770 9537 17782 9571
rect 17816 9568 17828 9571
rect 18141 9571 18199 9577
rect 17816 9540 17908 9568
rect 17816 9537 17828 9540
rect 17770 9531 17828 9537
rect 16632 9472 16988 9500
rect 16632 9460 16638 9472
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 17052 9432 17080 9528
rect 17880 9444 17908 9540
rect 18141 9537 18153 9571
rect 18187 9568 18199 9571
rect 18322 9568 18328 9580
rect 18187 9540 18328 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 18506 9571 18564 9577
rect 18506 9568 18518 9571
rect 18432 9540 18518 9568
rect 18230 9460 18236 9512
rect 18288 9460 18294 9512
rect 16080 9404 17080 9432
rect 16080 9392 16086 9404
rect 17862 9392 17868 9444
rect 17920 9432 17926 9444
rect 18432 9432 18460 9540
rect 18506 9537 18518 9540
rect 18552 9537 18564 9571
rect 18506 9531 18564 9537
rect 19058 9528 19064 9580
rect 19116 9528 19122 9580
rect 22554 9528 22560 9580
rect 22612 9528 22618 9580
rect 26326 9528 26332 9580
rect 26384 9528 26390 9580
rect 26421 9571 26479 9577
rect 26421 9537 26433 9571
rect 26467 9568 26479 9571
rect 26973 9571 27031 9577
rect 26973 9568 26985 9571
rect 26467 9540 26985 9568
rect 26467 9537 26479 9540
rect 26421 9531 26479 9537
rect 26973 9537 26985 9540
rect 27019 9568 27031 9571
rect 27798 9568 27804 9580
rect 27019 9540 27804 9568
rect 27019 9537 27031 9540
rect 26973 9531 27031 9537
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 17920 9404 18460 9432
rect 18616 9472 18981 9500
rect 17920 9392 17926 9404
rect 10796 9336 12020 9364
rect 10100 9324 10106 9336
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 14274 9364 14280 9376
rect 13688 9336 14280 9364
rect 13688 9324 13694 9336
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 17586 9324 17592 9376
rect 17644 9324 17650 9376
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 18012 9336 18337 9364
rect 18012 9324 18018 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 18414 9324 18420 9376
rect 18472 9364 18478 9376
rect 18616 9364 18644 9472
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 22572 9500 22600 9528
rect 26436 9500 26464 9531
rect 27798 9528 27804 9540
rect 27856 9528 27862 9580
rect 28000 9577 28028 9608
rect 28074 9596 28080 9648
rect 28132 9636 28138 9648
rect 28132 9608 28304 9636
rect 28132 9596 28138 9608
rect 27893 9571 27951 9577
rect 27893 9537 27905 9571
rect 27939 9537 27951 9571
rect 27893 9531 27951 9537
rect 27985 9571 28043 9577
rect 27985 9537 27997 9571
rect 28031 9537 28043 9571
rect 27985 9531 28043 9537
rect 22572 9472 26464 9500
rect 26605 9503 26663 9509
rect 18969 9463 19027 9469
rect 26605 9469 26617 9503
rect 26651 9500 26663 9503
rect 26878 9500 26884 9512
rect 26651 9472 26884 9500
rect 26651 9469 26663 9472
rect 26605 9463 26663 9469
rect 26878 9460 26884 9472
rect 26936 9460 26942 9512
rect 27908 9500 27936 9531
rect 28166 9528 28172 9580
rect 28224 9528 28230 9580
rect 28276 9577 28304 9608
rect 28261 9571 28319 9577
rect 28261 9537 28273 9571
rect 28307 9537 28319 9571
rect 28261 9531 28319 9537
rect 27908 9472 28488 9500
rect 26142 9392 26148 9444
rect 26200 9432 26206 9444
rect 27617 9435 27675 9441
rect 27617 9432 27629 9435
rect 26200 9404 27629 9432
rect 26200 9392 26206 9404
rect 27617 9401 27629 9404
rect 27663 9401 27675 9435
rect 27617 9395 27675 9401
rect 28460 9376 28488 9472
rect 18472 9336 18644 9364
rect 18877 9367 18935 9373
rect 18472 9324 18478 9336
rect 18877 9333 18889 9367
rect 18923 9364 18935 9367
rect 19334 9364 19340 9376
rect 18923 9336 19340 9364
rect 18923 9333 18935 9336
rect 18877 9327 18935 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 25590 9324 25596 9376
rect 25648 9364 25654 9376
rect 27709 9367 27767 9373
rect 27709 9364 27721 9367
rect 25648 9336 27721 9364
rect 25648 9324 25654 9336
rect 27709 9333 27721 9336
rect 27755 9333 27767 9367
rect 27709 9327 27767 9333
rect 28442 9324 28448 9376
rect 28500 9324 28506 9376
rect 1104 9274 29440 9296
rect 1104 9222 4491 9274
rect 4543 9222 4555 9274
rect 4607 9222 4619 9274
rect 4671 9222 4683 9274
rect 4735 9222 4747 9274
rect 4799 9222 11574 9274
rect 11626 9222 11638 9274
rect 11690 9222 11702 9274
rect 11754 9222 11766 9274
rect 11818 9222 11830 9274
rect 11882 9222 18657 9274
rect 18709 9222 18721 9274
rect 18773 9222 18785 9274
rect 18837 9222 18849 9274
rect 18901 9222 18913 9274
rect 18965 9222 25740 9274
rect 25792 9222 25804 9274
rect 25856 9222 25868 9274
rect 25920 9222 25932 9274
rect 25984 9222 25996 9274
rect 26048 9222 29440 9274
rect 1104 9200 29440 9222
rect 2120 9163 2178 9169
rect 2120 9129 2132 9163
rect 2166 9160 2178 9163
rect 5626 9160 5632 9172
rect 2166 9132 5632 9160
rect 2166 9129 2178 9132
rect 2120 9123 2178 9129
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 5736 9132 13032 9160
rect 3326 9052 3332 9104
rect 3384 9052 3390 9104
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 5353 9095 5411 9101
rect 5353 9092 5365 9095
rect 5132 9064 5365 9092
rect 5132 9052 5138 9064
rect 5353 9061 5365 9064
rect 5399 9061 5411 9095
rect 5353 9055 5411 9061
rect 5534 9052 5540 9104
rect 5592 9092 5598 9104
rect 5736 9092 5764 9132
rect 5592 9064 5764 9092
rect 5592 9052 5598 9064
rect 10410 9052 10416 9104
rect 10468 9092 10474 9104
rect 13004 9092 13032 9132
rect 13078 9120 13084 9172
rect 13136 9120 13142 9172
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 22557 9163 22615 9169
rect 22557 9160 22569 9163
rect 17552 9132 22569 9160
rect 17552 9120 17558 9132
rect 22557 9129 22569 9132
rect 22603 9129 22615 9163
rect 22557 9123 22615 9129
rect 17310 9092 17316 9104
rect 10468 9064 10548 9092
rect 13004 9064 17316 9092
rect 10468 9052 10474 9064
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 2222 9024 2228 9036
rect 1903 8996 2228 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 3344 8956 3372 9052
rect 3605 9027 3663 9033
rect 3605 8993 3617 9027
rect 3651 9024 3663 9027
rect 4338 9024 4344 9036
rect 3651 8996 4344 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 4396 8996 5825 9024
rect 4396 8984 4402 8996
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 5994 9024 6000 9036
rect 5951 8996 6000 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6227 8996 8984 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 8956 8968 8984 8996
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 9309 9027 9367 9033
rect 9309 9024 9321 9027
rect 9180 8996 9321 9024
rect 9180 8984 9186 8996
rect 9309 8993 9321 8996
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 9858 8984 9864 9036
rect 9916 9024 9922 9036
rect 10134 9024 10140 9036
rect 9916 8996 10140 9024
rect 9916 8984 9922 8996
rect 10134 8984 10140 8996
rect 10192 9024 10198 9036
rect 10520 9024 10548 9064
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 18322 9052 18328 9104
rect 18380 9052 18386 9104
rect 22572 9092 22600 9123
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 23017 9163 23075 9169
rect 23017 9160 23029 9163
rect 22888 9132 23029 9160
rect 22888 9120 22894 9132
rect 23017 9129 23029 9132
rect 23063 9129 23075 9163
rect 23017 9123 23075 9129
rect 24946 9120 24952 9172
rect 25004 9160 25010 9172
rect 25004 9132 26280 9160
rect 25004 9120 25010 9132
rect 24026 9092 24032 9104
rect 22572 9064 24032 9092
rect 24026 9052 24032 9064
rect 24084 9052 24090 9104
rect 25590 9052 25596 9104
rect 25648 9052 25654 9104
rect 25682 9052 25688 9104
rect 25740 9092 25746 9104
rect 25740 9064 26030 9092
rect 25740 9052 25746 9064
rect 11054 9024 11060 9036
rect 10192 8996 10456 9024
rect 10520 8996 11060 9024
rect 10192 8984 10198 8996
rect 3266 8928 3372 8956
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4295 8928 4384 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4356 8832 4384 8928
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 10428 8956 10456 8996
rect 11054 8984 11060 8996
rect 11112 9024 11118 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 11112 8996 11161 9024
rect 11112 8984 11118 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 11358 9027 11416 9033
rect 11358 9024 11370 9027
rect 11296 8996 11370 9024
rect 11296 8984 11302 8996
rect 11358 8993 11370 8996
rect 11404 9024 11416 9027
rect 12066 9024 12072 9036
rect 11404 8996 12072 9024
rect 11404 8993 11416 8996
rect 11358 8987 11416 8993
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 9024 14703 9027
rect 15654 9024 15660 9036
rect 14691 8996 15660 9024
rect 14691 8993 14703 8996
rect 14645 8987 14703 8993
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 18138 9024 18144 9036
rect 16408 8996 18144 9024
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10428 8928 10885 8956
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 10873 8919 10931 8925
rect 11532 8928 11621 8956
rect 5353 8891 5411 8897
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 6270 8888 6276 8900
rect 5399 8860 6276 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 7098 8848 7104 8900
rect 7156 8848 7162 8900
rect 9674 8848 9680 8900
rect 9732 8848 9738 8900
rect 11241 8891 11299 8897
rect 11241 8857 11253 8891
rect 11287 8888 11299 8891
rect 11330 8888 11336 8900
rect 11287 8860 11336 8888
rect 11287 8857 11299 8860
rect 11241 8851 11299 8857
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 4338 8780 4344 8832
rect 4396 8780 4402 8832
rect 4890 8780 4896 8832
rect 4948 8780 4954 8832
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 5132 8792 6101 8820
rect 5132 8780 5138 8792
rect 6089 8789 6101 8792
rect 6135 8789 6147 8823
rect 6288 8820 6316 8848
rect 7975 8823 8033 8829
rect 7975 8820 7987 8823
rect 6288 8792 7987 8820
rect 6089 8783 6147 8789
rect 7975 8789 7987 8792
rect 8021 8789 8033 8823
rect 7975 8783 8033 8789
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 11532 8829 11560 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 12158 8956 12164 8968
rect 11931 8928 12164 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13722 8956 13728 8968
rect 13035 8928 13728 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 13817 8959 13875 8965
rect 13817 8925 13829 8959
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 13541 8891 13599 8897
rect 13541 8888 13553 8891
rect 13320 8860 13553 8888
rect 13320 8848 13326 8860
rect 13541 8857 13553 8860
rect 13587 8857 13599 8891
rect 13832 8888 13860 8919
rect 16408 8900 16436 8996
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18046 8956 18052 8968
rect 18003 8928 18052 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18340 8965 18368 9052
rect 22186 8984 22192 9036
rect 22244 8984 22250 9036
rect 22278 8984 22284 9036
rect 22336 8984 22342 9036
rect 22462 8984 22468 9036
rect 22520 9024 22526 9036
rect 22649 9027 22707 9033
rect 22649 9024 22661 9027
rect 22520 8996 22661 9024
rect 22520 8984 22526 8996
rect 22649 8993 22661 8996
rect 22695 8993 22707 9027
rect 22649 8987 22707 8993
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 22097 8959 22155 8965
rect 19392 8928 20668 8956
rect 19392 8916 19398 8928
rect 13906 8888 13912 8900
rect 13832 8860 13912 8888
rect 13541 8851 13599 8857
rect 13906 8848 13912 8860
rect 13964 8848 13970 8900
rect 16390 8848 16396 8900
rect 16448 8848 16454 8900
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 18141 8891 18199 8897
rect 18141 8888 18153 8891
rect 16908 8860 18153 8888
rect 16908 8848 16914 8860
rect 18141 8857 18153 8860
rect 18187 8857 18199 8891
rect 18141 8851 18199 8857
rect 18230 8848 18236 8900
rect 18288 8848 18294 8900
rect 19889 8891 19947 8897
rect 19889 8888 19901 8891
rect 18432 8860 19901 8888
rect 10735 8823 10793 8829
rect 10735 8820 10747 8823
rect 10008 8792 10747 8820
rect 10008 8780 10014 8792
rect 10735 8789 10747 8792
rect 10781 8789 10793 8823
rect 10735 8783 10793 8789
rect 11517 8823 11575 8829
rect 11517 8789 11529 8823
rect 11563 8789 11575 8823
rect 13630 8820 13636 8832
rect 13688 8829 13694 8832
rect 13597 8792 13636 8820
rect 11517 8783 11575 8789
rect 13630 8780 13636 8792
rect 13688 8783 13697 8829
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 15197 8823 15255 8829
rect 15197 8820 15209 8823
rect 13771 8792 15209 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 15197 8789 15209 8792
rect 15243 8789 15255 8823
rect 15197 8783 15255 8789
rect 13688 8780 13694 8783
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 18432 8820 18460 8860
rect 19889 8857 19901 8860
rect 19935 8857 19947 8891
rect 19889 8851 19947 8857
rect 20640 8832 20668 8928
rect 22097 8925 22109 8959
rect 22143 8956 22155 8959
rect 22370 8956 22376 8968
rect 22143 8928 22376 8956
rect 22143 8925 22155 8928
rect 22097 8919 22155 8925
rect 22370 8916 22376 8928
rect 22428 8916 22434 8968
rect 22833 8959 22891 8965
rect 22833 8956 22845 8959
rect 22664 8928 22845 8956
rect 22554 8848 22560 8900
rect 22612 8848 22618 8900
rect 18104 8792 18460 8820
rect 18104 8780 18110 8792
rect 18506 8780 18512 8832
rect 18564 8780 18570 8832
rect 20622 8780 20628 8832
rect 20680 8780 20686 8832
rect 21726 8780 21732 8832
rect 21784 8780 21790 8832
rect 22094 8780 22100 8832
rect 22152 8820 22158 8832
rect 22572 8820 22600 8848
rect 22664 8832 22692 8928
rect 22833 8925 22845 8928
rect 22879 8956 22891 8959
rect 23382 8956 23388 8968
rect 22879 8928 23388 8956
rect 22879 8925 22891 8928
rect 22833 8919 22891 8925
rect 23382 8916 23388 8928
rect 23440 8916 23446 8968
rect 25608 8956 25636 9052
rect 26002 8965 26030 9064
rect 26252 9033 26280 9132
rect 27798 9120 27804 9172
rect 27856 9160 27862 9172
rect 27985 9163 28043 9169
rect 27985 9160 27997 9163
rect 27856 9132 27997 9160
rect 27856 9120 27862 9132
rect 27985 9129 27997 9132
rect 28031 9129 28043 9163
rect 27985 9123 28043 9129
rect 26237 9027 26295 9033
rect 26237 8993 26249 9027
rect 26283 8993 26295 9027
rect 26237 8987 26295 8993
rect 25686 8959 25744 8965
rect 25686 8956 25698 8959
rect 25608 8928 25698 8956
rect 25686 8925 25698 8928
rect 25732 8925 25744 8959
rect 25686 8919 25744 8925
rect 25987 8959 26045 8965
rect 25987 8925 25999 8959
rect 26033 8925 26045 8959
rect 25987 8919 26045 8925
rect 26142 8916 26148 8968
rect 26200 8916 26206 8968
rect 28000 8956 28028 9123
rect 28353 8959 28411 8965
rect 28353 8956 28365 8959
rect 28000 8928 28365 8956
rect 28353 8925 28365 8928
rect 28399 8925 28411 8959
rect 28353 8919 28411 8925
rect 25774 8848 25780 8900
rect 25832 8848 25838 8900
rect 25866 8848 25872 8900
rect 25924 8848 25930 8900
rect 26513 8891 26571 8897
rect 26513 8857 26525 8891
rect 26559 8857 26571 8891
rect 26513 8851 26571 8857
rect 22152 8792 22600 8820
rect 22152 8780 22158 8792
rect 22646 8780 22652 8832
rect 22704 8780 22710 8832
rect 25501 8823 25559 8829
rect 25501 8789 25513 8823
rect 25547 8820 25559 8823
rect 26528 8820 26556 8851
rect 26786 8848 26792 8900
rect 26844 8848 26850 8900
rect 27062 8848 27068 8900
rect 27120 8848 27126 8900
rect 28169 8891 28227 8897
rect 28169 8857 28181 8891
rect 28215 8857 28227 8891
rect 28169 8851 28227 8857
rect 25547 8792 26556 8820
rect 26804 8820 26832 8848
rect 28184 8820 28212 8851
rect 28442 8848 28448 8900
rect 28500 8888 28506 8900
rect 28537 8891 28595 8897
rect 28537 8888 28549 8891
rect 28500 8860 28549 8888
rect 28500 8848 28506 8860
rect 28537 8857 28549 8860
rect 28583 8857 28595 8891
rect 28537 8851 28595 8857
rect 26804 8792 28212 8820
rect 25547 8789 25559 8792
rect 25501 8783 25559 8789
rect 1104 8730 29440 8752
rect 1104 8678 5151 8730
rect 5203 8678 5215 8730
rect 5267 8678 5279 8730
rect 5331 8678 5343 8730
rect 5395 8678 5407 8730
rect 5459 8678 12234 8730
rect 12286 8678 12298 8730
rect 12350 8678 12362 8730
rect 12414 8678 12426 8730
rect 12478 8678 12490 8730
rect 12542 8678 19317 8730
rect 19369 8678 19381 8730
rect 19433 8678 19445 8730
rect 19497 8678 19509 8730
rect 19561 8678 19573 8730
rect 19625 8678 26400 8730
rect 26452 8678 26464 8730
rect 26516 8678 26528 8730
rect 26580 8678 26592 8730
rect 26644 8678 26656 8730
rect 26708 8678 29440 8730
rect 1104 8656 29440 8678
rect 2222 8576 2228 8628
rect 2280 8576 2286 8628
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 3384 8588 3556 8616
rect 3384 8576 3390 8588
rect 2240 8548 2268 8576
rect 2682 8548 2688 8560
rect 2148 8520 2688 8548
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 2148 8489 2176 8520
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 2133 8483 2191 8489
rect 2133 8480 2145 8483
rect 1728 8452 2145 8480
rect 1728 8440 1734 8452
rect 2133 8449 2145 8452
rect 2179 8449 2191 8483
rect 3528 8466 3556 8588
rect 4890 8576 4896 8628
rect 4948 8576 4954 8628
rect 5445 8619 5503 8625
rect 5445 8585 5457 8619
rect 5491 8616 5503 8619
rect 5534 8616 5540 8628
rect 5491 8588 5540 8616
rect 5491 8585 5503 8588
rect 5445 8579 5503 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8585 5687 8619
rect 5629 8579 5687 8585
rect 4908 8548 4936 8576
rect 3988 8520 4936 8548
rect 4985 8551 5043 8557
rect 3988 8489 4016 8520
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 5644 8548 5672 8579
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6730 8616 6736 8628
rect 6052 8588 6736 8616
rect 6052 8576 6058 8588
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 9950 8616 9956 8628
rect 7668 8588 9168 8616
rect 5031 8520 5672 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 5810 8508 5816 8560
rect 5868 8548 5874 8560
rect 6012 8548 6040 8576
rect 7668 8557 7696 8588
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 5868 8520 6040 8548
rect 5868 8508 5874 8520
rect 3973 8483 4031 8489
rect 2133 8443 2191 8449
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4246 8440 4252 8492
rect 4304 8440 4310 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4430 8480 4436 8492
rect 4387 8452 4436 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4430 8440 4436 8452
rect 4488 8480 4494 8492
rect 5261 8483 5319 8489
rect 4488 8452 5028 8480
rect 4488 8440 4494 8452
rect 5000 8424 5028 8452
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5442 8480 5448 8492
rect 5307 8452 5448 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5736 8452 5948 8480
rect 5736 8424 5764 8452
rect 2409 8415 2467 8421
rect 2409 8381 2421 8415
rect 2455 8412 2467 8415
rect 2455 8384 4568 8412
rect 2455 8381 2467 8384
rect 2409 8375 2467 8381
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4338 8344 4344 8356
rect 3927 8316 4344 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4338 8304 4344 8316
rect 4396 8344 4402 8356
rect 4540 8353 4568 8384
rect 4982 8372 4988 8424
rect 5040 8372 5046 8424
rect 5074 8372 5080 8424
rect 5132 8372 5138 8424
rect 5718 8372 5724 8424
rect 5776 8372 5782 8424
rect 5920 8421 5948 8452
rect 6012 8421 6040 8520
rect 6104 8520 7665 8548
rect 6104 8421 6132 8520
rect 7653 8517 7665 8520
rect 7699 8517 7711 8551
rect 7653 8511 7711 8517
rect 8297 8551 8355 8557
rect 8297 8517 8309 8551
rect 8343 8517 8355 8551
rect 8297 8511 8355 8517
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6822 8480 6828 8492
rect 6328 8452 6828 8480
rect 6328 8440 6334 8452
rect 6822 8440 6828 8452
rect 6880 8480 6886 8492
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 6880 8452 7297 8480
rect 6880 8440 6886 8452
rect 7285 8449 7297 8452
rect 7331 8480 7343 8483
rect 8312 8480 8340 8511
rect 9030 8508 9036 8560
rect 9088 8508 9094 8560
rect 7331 8452 8340 8480
rect 9140 8480 9168 8588
rect 9232 8588 9956 8616
rect 9232 8557 9260 8588
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 13320 8588 13369 8616
rect 13320 8576 13326 8588
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 13556 8588 15516 8616
rect 9217 8551 9275 8557
rect 9217 8517 9229 8551
rect 9263 8517 9275 8551
rect 13556 8548 13584 8588
rect 9217 8511 9275 8517
rect 13096 8520 13584 8548
rect 9766 8480 9772 8492
rect 9140 8452 9772 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 13096 8489 13124 8520
rect 13630 8508 13636 8560
rect 13688 8548 13694 8560
rect 13725 8551 13783 8557
rect 13725 8548 13737 8551
rect 13688 8520 13737 8548
rect 13688 8508 13694 8520
rect 13725 8517 13737 8520
rect 13771 8517 13783 8551
rect 13725 8511 13783 8517
rect 14274 8508 14280 8560
rect 14332 8508 14338 8560
rect 15488 8557 15516 8588
rect 16758 8576 16764 8628
rect 16816 8576 16822 8628
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 18506 8576 18512 8628
rect 18564 8576 18570 8628
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 19208 8588 19564 8616
rect 19208 8576 19214 8588
rect 15473 8551 15531 8557
rect 15473 8517 15485 8551
rect 15519 8548 15531 8551
rect 15654 8548 15660 8560
rect 15519 8520 15660 8548
rect 15519 8517 15531 8520
rect 15473 8511 15531 8517
rect 15654 8508 15660 8520
rect 15712 8508 15718 8560
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 16574 8440 16580 8492
rect 16632 8480 16638 8492
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 16632 8452 16681 8480
rect 16632 8440 16638 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16776 8480 16804 8576
rect 17604 8548 17632 8576
rect 17328 8520 17632 8548
rect 17328 8489 17356 8520
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16776 8452 16865 8480
rect 16669 8443 16727 8449
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17129 8483 17187 8489
rect 17129 8480 17141 8483
rect 17083 8452 17141 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 17129 8449 17141 8452
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 17277 8483 17356 8489
rect 17277 8449 17289 8483
rect 17323 8452 17356 8483
rect 17405 8483 17463 8489
rect 17323 8449 17335 8452
rect 17277 8443 17335 8449
rect 17405 8449 17417 8483
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8381 5871 8415
rect 5813 8375 5871 8381
rect 5905 8415 5963 8421
rect 5905 8381 5917 8415
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 5997 8415 6055 8421
rect 5997 8381 6009 8415
rect 6043 8381 6055 8415
rect 5997 8375 6055 8381
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 4525 8347 4583 8353
rect 4396 8316 4476 8344
rect 4396 8304 4402 8316
rect 4448 8276 4476 8316
rect 4525 8313 4537 8347
rect 4571 8313 4583 8347
rect 5828 8344 5856 8375
rect 6564 8344 6592 8375
rect 6638 8372 6644 8424
rect 6696 8372 6702 8424
rect 6730 8372 6736 8424
rect 6788 8372 6794 8424
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8260 8384 8769 8412
rect 8260 8372 8266 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 9490 8412 9496 8424
rect 8895 8384 9496 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 4525 8307 4583 8313
rect 4632 8316 5856 8344
rect 5920 8316 6592 8344
rect 4632 8276 4660 8316
rect 4448 8248 4660 8276
rect 5074 8236 5080 8288
rect 5132 8236 5138 8288
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 5920 8276 5948 8316
rect 5592 8248 5948 8276
rect 5592 8236 5598 8248
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 6236 8248 6377 8276
rect 6236 8236 6242 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 6656 8276 6684 8372
rect 6748 8344 6776 8372
rect 8297 8347 8355 8353
rect 8297 8344 8309 8347
rect 6748 8316 8309 8344
rect 8297 8313 8309 8316
rect 8343 8313 8355 8347
rect 8864 8344 8892 8375
rect 9490 8372 9496 8384
rect 9548 8412 9554 8424
rect 9953 8415 10011 8421
rect 9953 8412 9965 8415
rect 9548 8384 9965 8412
rect 9548 8372 9554 8384
rect 9953 8381 9965 8384
rect 9999 8381 10011 8415
rect 13354 8412 13360 8424
rect 9953 8375 10011 8381
rect 12176 8384 13360 8412
rect 12176 8356 12204 8384
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 13446 8372 13452 8424
rect 13504 8372 13510 8424
rect 8297 8307 8355 8313
rect 8404 8316 8892 8344
rect 8404 8276 8432 8316
rect 12158 8304 12164 8356
rect 12216 8304 12222 8356
rect 13173 8347 13231 8353
rect 13173 8313 13185 8347
rect 13219 8344 13231 8347
rect 13219 8316 13584 8344
rect 13219 8313 13231 8316
rect 13173 8307 13231 8313
rect 6656 8248 8432 8276
rect 13556 8276 13584 8316
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 17420 8344 17448 8443
rect 17494 8440 17500 8492
rect 17552 8440 17558 8492
rect 17635 8483 17693 8489
rect 17635 8449 17647 8483
rect 17681 8480 17693 8483
rect 17770 8480 17776 8492
rect 17681 8452 17776 8480
rect 17681 8449 17693 8452
rect 17635 8443 17693 8449
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 18524 8412 18552 8576
rect 19242 8548 19248 8560
rect 18892 8520 19248 8548
rect 18892 8489 18920 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 19536 8548 19564 8588
rect 20622 8576 20628 8628
rect 20680 8576 20686 8628
rect 21726 8576 21732 8628
rect 21784 8576 21790 8628
rect 23014 8576 23020 8628
rect 23072 8616 23078 8628
rect 23072 8588 23796 8616
rect 23072 8576 23078 8588
rect 19536 8520 19642 8548
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8449 18935 8483
rect 18877 8443 18935 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8480 21143 8483
rect 21744 8480 21772 8576
rect 23385 8551 23443 8557
rect 23385 8548 23397 8551
rect 22572 8520 23397 8548
rect 22572 8492 22600 8520
rect 23385 8517 23397 8520
rect 23431 8548 23443 8551
rect 23658 8548 23664 8560
rect 23431 8520 23664 8548
rect 23431 8517 23443 8520
rect 23385 8511 23443 8517
rect 23658 8508 23664 8520
rect 23716 8508 23722 8560
rect 23768 8548 23796 8588
rect 24210 8548 24216 8560
rect 23768 8520 24216 8548
rect 21131 8452 21772 8480
rect 21131 8449 21143 8452
rect 21085 8443 21143 8449
rect 22554 8440 22560 8492
rect 22612 8440 22618 8492
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 18524 8384 19165 8412
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 22848 8412 22876 8443
rect 22922 8440 22928 8492
rect 22980 8480 22986 8492
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 22980 8452 23029 8480
rect 22980 8440 22986 8452
rect 23017 8449 23029 8452
rect 23063 8480 23075 8483
rect 23198 8480 23204 8492
rect 23063 8452 23204 8480
rect 23063 8449 23075 8452
rect 23017 8443 23075 8449
rect 23198 8440 23204 8452
rect 23256 8440 23262 8492
rect 23474 8440 23480 8492
rect 23532 8480 23538 8492
rect 23952 8489 23980 8520
rect 24210 8508 24216 8520
rect 24268 8508 24274 8560
rect 25774 8508 25780 8560
rect 25832 8548 25838 8560
rect 26234 8548 26240 8560
rect 25832 8520 26240 8548
rect 25832 8508 25838 8520
rect 26234 8508 26240 8520
rect 26292 8548 26298 8560
rect 27065 8551 27123 8557
rect 27065 8548 27077 8551
rect 26292 8520 27077 8548
rect 26292 8508 26298 8520
rect 27065 8517 27077 8520
rect 27111 8517 27123 8551
rect 28442 8548 28448 8560
rect 27065 8511 27123 8517
rect 27264 8520 28448 8548
rect 23569 8483 23627 8489
rect 23569 8480 23581 8483
rect 23532 8452 23581 8480
rect 23532 8440 23538 8452
rect 23569 8449 23581 8452
rect 23615 8449 23627 8483
rect 23937 8483 23995 8489
rect 23569 8443 23627 8449
rect 23676 8452 23888 8480
rect 22848 8384 23060 8412
rect 19153 8375 19211 8381
rect 23032 8356 23060 8384
rect 23382 8372 23388 8424
rect 23440 8412 23446 8424
rect 23676 8412 23704 8452
rect 23440 8384 23704 8412
rect 23440 8372 23446 8384
rect 23750 8372 23756 8424
rect 23808 8372 23814 8424
rect 23860 8412 23888 8452
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 24026 8440 24032 8492
rect 24084 8480 24090 8492
rect 24121 8483 24179 8489
rect 24121 8480 24133 8483
rect 24084 8452 24133 8480
rect 24084 8440 24090 8452
rect 24121 8449 24133 8452
rect 24167 8449 24179 8483
rect 24228 8480 24256 8508
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 24228 8452 26065 8480
rect 24121 8443 24179 8449
rect 26053 8449 26065 8452
rect 26099 8480 26111 8483
rect 26418 8480 26424 8492
rect 26099 8452 26424 8480
rect 26099 8449 26111 8452
rect 26053 8443 26111 8449
rect 26418 8440 26424 8452
rect 26476 8480 26482 8492
rect 26476 8452 26740 8480
rect 26476 8440 26482 8452
rect 25869 8415 25927 8421
rect 25869 8412 25881 8415
rect 23860 8384 25881 8412
rect 25869 8381 25881 8384
rect 25915 8381 25927 8415
rect 25869 8375 25927 8381
rect 16632 8316 17448 8344
rect 16632 8304 16638 8316
rect 23014 8304 23020 8356
rect 23072 8304 23078 8356
rect 23658 8304 23664 8356
rect 23716 8344 23722 8356
rect 23937 8347 23995 8353
rect 23937 8344 23949 8347
rect 23716 8316 23949 8344
rect 23716 8304 23722 8316
rect 23937 8313 23949 8316
rect 23983 8313 23995 8347
rect 25884 8344 25912 8375
rect 26326 8372 26332 8424
rect 26384 8372 26390 8424
rect 26510 8344 26516 8356
rect 25884 8316 26516 8344
rect 23937 8307 23995 8313
rect 26510 8304 26516 8316
rect 26568 8304 26574 8356
rect 26602 8304 26608 8356
rect 26660 8304 26666 8356
rect 26712 8344 26740 8452
rect 26878 8440 26884 8492
rect 26936 8480 26942 8492
rect 27264 8489 27292 8520
rect 28442 8508 28448 8520
rect 28500 8508 28506 8560
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26936 8452 26985 8480
rect 26936 8440 26942 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 27525 8483 27583 8489
rect 27525 8449 27537 8483
rect 27571 8449 27583 8483
rect 27525 8443 27583 8449
rect 26789 8415 26847 8421
rect 26789 8381 26801 8415
rect 26835 8412 26847 8415
rect 27540 8412 27568 8443
rect 27614 8440 27620 8492
rect 27672 8480 27678 8492
rect 27801 8483 27859 8489
rect 27801 8480 27813 8483
rect 27672 8452 27813 8480
rect 27672 8440 27678 8452
rect 27801 8449 27813 8452
rect 27847 8480 27859 8483
rect 28074 8480 28080 8492
rect 27847 8452 28080 8480
rect 27847 8449 27859 8452
rect 27801 8443 27859 8449
rect 28074 8440 28080 8452
rect 28132 8440 28138 8492
rect 28166 8440 28172 8492
rect 28224 8440 28230 8492
rect 28184 8412 28212 8440
rect 26835 8384 28212 8412
rect 26835 8381 26847 8384
rect 26789 8375 26847 8381
rect 26878 8344 26884 8356
rect 26712 8316 26884 8344
rect 26878 8304 26884 8316
rect 26936 8304 26942 8356
rect 27522 8304 27528 8356
rect 27580 8304 27586 8356
rect 13906 8276 13912 8288
rect 13556 8248 13912 8276
rect 6365 8239 6423 8245
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 17034 8236 17040 8288
rect 17092 8276 17098 8288
rect 17773 8279 17831 8285
rect 17773 8276 17785 8279
rect 17092 8248 17785 8276
rect 17092 8236 17098 8248
rect 17773 8245 17785 8248
rect 17819 8245 17831 8279
rect 17773 8239 17831 8245
rect 20898 8236 20904 8288
rect 20956 8236 20962 8288
rect 22462 8236 22468 8288
rect 22520 8276 22526 8288
rect 22922 8276 22928 8288
rect 22520 8248 22928 8276
rect 22520 8236 22526 8248
rect 22922 8236 22928 8248
rect 22980 8276 22986 8288
rect 23201 8279 23259 8285
rect 23201 8276 23213 8279
rect 22980 8248 23213 8276
rect 22980 8236 22986 8248
rect 23201 8245 23213 8248
rect 23247 8245 23259 8279
rect 23201 8239 23259 8245
rect 23845 8279 23903 8285
rect 23845 8245 23857 8279
rect 23891 8276 23903 8279
rect 24670 8276 24676 8288
rect 23891 8248 24676 8276
rect 23891 8245 23903 8248
rect 23845 8239 23903 8245
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 26237 8279 26295 8285
rect 26237 8245 26249 8279
rect 26283 8276 26295 8279
rect 27540 8276 27568 8304
rect 26283 8248 27568 8276
rect 26283 8245 26295 8248
rect 26237 8239 26295 8245
rect 1104 8186 29440 8208
rect 1104 8134 4491 8186
rect 4543 8134 4555 8186
rect 4607 8134 4619 8186
rect 4671 8134 4683 8186
rect 4735 8134 4747 8186
rect 4799 8134 11574 8186
rect 11626 8134 11638 8186
rect 11690 8134 11702 8186
rect 11754 8134 11766 8186
rect 11818 8134 11830 8186
rect 11882 8134 18657 8186
rect 18709 8134 18721 8186
rect 18773 8134 18785 8186
rect 18837 8134 18849 8186
rect 18901 8134 18913 8186
rect 18965 8134 25740 8186
rect 25792 8134 25804 8186
rect 25856 8134 25868 8186
rect 25920 8134 25932 8186
rect 25984 8134 25996 8186
rect 26048 8134 29440 8186
rect 1104 8112 29440 8134
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 3988 8044 5181 8072
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 3988 7936 4016 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 6089 8075 6147 8081
rect 6089 8072 6101 8075
rect 5583 8044 6101 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 6089 8041 6101 8044
rect 6135 8041 6147 8075
rect 13725 8075 13783 8081
rect 6089 8035 6147 8041
rect 6196 8044 12434 8072
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 6196 8004 6224 8044
rect 4120 7976 6224 8004
rect 4120 7964 4126 7976
rect 6730 7964 6736 8016
rect 6788 7964 6794 8016
rect 12406 8004 12434 8044
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 14090 8072 14096 8084
rect 13771 8044 14096 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 14090 8032 14096 8044
rect 14148 8072 14154 8084
rect 14458 8072 14464 8084
rect 14148 8044 14464 8072
rect 14148 8032 14154 8044
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 14734 8032 14740 8084
rect 14792 8032 14798 8084
rect 18046 8072 18052 8084
rect 17328 8044 18052 8072
rect 14182 8004 14188 8016
rect 12406 7976 14188 8004
rect 14182 7964 14188 7976
rect 14240 7964 14246 8016
rect 5442 7936 5448 7948
rect 1995 7908 4016 7936
rect 4448 7908 5448 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 1670 7828 1676 7880
rect 1728 7828 1734 7880
rect 3326 7868 3332 7880
rect 3082 7840 3332 7868
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4448 7868 4476 7908
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 6273 7939 6331 7945
rect 5776 7908 6040 7936
rect 5776 7896 5782 7908
rect 4019 7840 4476 7868
rect 4525 7871 4583 7877
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4571 7840 4629 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 3988 7732 4016 7831
rect 4982 7828 4988 7880
rect 5040 7828 5046 7880
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5902 7828 5908 7880
rect 5960 7828 5966 7880
rect 6012 7868 6040 7908
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 7190 7936 7196 7948
rect 6319 7908 7196 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 13998 7936 14004 7948
rect 10008 7908 14004 7936
rect 10008 7896 10014 7908
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 14752 7936 14780 8032
rect 17328 8016 17356 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 21821 8075 21879 8081
rect 21821 8041 21833 8075
rect 21867 8072 21879 8075
rect 22186 8072 22192 8084
rect 21867 8044 22192 8072
rect 21867 8041 21879 8044
rect 21821 8035 21879 8041
rect 22186 8032 22192 8044
rect 22244 8032 22250 8084
rect 22278 8032 22284 8084
rect 22336 8032 22342 8084
rect 23842 8072 23848 8084
rect 22664 8044 23848 8072
rect 17310 7964 17316 8016
rect 17368 7964 17374 8016
rect 17770 7964 17776 8016
rect 17828 7964 17834 8016
rect 22296 8004 22324 8032
rect 22664 8004 22692 8044
rect 23842 8032 23848 8044
rect 23900 8032 23906 8084
rect 25225 8075 25283 8081
rect 25225 8041 25237 8075
rect 25271 8072 25283 8075
rect 26602 8072 26608 8084
rect 25271 8044 26608 8072
rect 25271 8041 25283 8044
rect 25225 8035 25283 8041
rect 26602 8032 26608 8044
rect 26660 8032 26666 8084
rect 27338 8032 27344 8084
rect 27396 8072 27402 8084
rect 27522 8072 27528 8084
rect 27396 8044 27528 8072
rect 27396 8032 27402 8044
rect 27522 8032 27528 8044
rect 27580 8032 27586 8084
rect 22296 7976 22692 8004
rect 17788 7936 17816 7964
rect 20349 7939 20407 7945
rect 14292 7908 14780 7936
rect 16776 7908 17080 7936
rect 6365 7871 6423 7877
rect 6012 7840 6316 7868
rect 4154 7760 4160 7812
rect 4212 7800 4218 7812
rect 4801 7803 4859 7809
rect 4801 7800 4813 7803
rect 4212 7772 4813 7800
rect 4212 7760 4218 7772
rect 4801 7769 4813 7772
rect 4847 7769 4859 7803
rect 4801 7763 4859 7769
rect 4890 7760 4896 7812
rect 4948 7760 4954 7812
rect 6089 7803 6147 7809
rect 6089 7769 6101 7803
rect 6135 7800 6147 7803
rect 6178 7800 6184 7812
rect 6135 7772 6184 7800
rect 6135 7769 6147 7772
rect 6089 7763 6147 7769
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6288 7800 6316 7840
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 6411 7840 7481 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 7469 7837 7481 7840
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 14090 7828 14096 7880
rect 14148 7828 14154 7880
rect 14292 7877 14320 7908
rect 16776 7880 16804 7908
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 6638 7800 6644 7812
rect 6288 7772 6644 7800
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 6733 7803 6791 7809
rect 6733 7769 6745 7803
rect 6779 7800 6791 7803
rect 6822 7800 6828 7812
rect 6779 7772 6828 7800
rect 6779 7769 6791 7772
rect 6733 7763 6791 7769
rect 6822 7760 6828 7772
rect 6880 7760 6886 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 6932 7772 7297 7800
rect 3467 7704 4016 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 6270 7732 6276 7744
rect 4304 7704 6276 7732
rect 4304 7692 4310 7704
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 6656 7732 6684 7760
rect 6932 7732 6960 7772
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7285 7763 7343 7769
rect 9858 7760 9864 7812
rect 9916 7800 9922 7812
rect 13541 7803 13599 7809
rect 13541 7800 13553 7803
rect 9916 7772 13553 7800
rect 9916 7760 9922 7772
rect 13541 7769 13553 7772
rect 13587 7800 13599 7803
rect 13630 7800 13636 7812
rect 13587 7772 13636 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 13722 7760 13728 7812
rect 13780 7809 13786 7812
rect 13780 7803 13815 7809
rect 13803 7800 13815 7803
rect 14292 7800 14320 7831
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 14516 7840 14565 7868
rect 14516 7828 14522 7840
rect 14553 7837 14565 7840
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 14642 7828 14648 7880
rect 14700 7868 14706 7880
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 14700 7840 14749 7868
rect 14700 7828 14706 7840
rect 14737 7837 14749 7840
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 14752 7800 14780 7831
rect 15102 7828 15108 7880
rect 15160 7828 15166 7880
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 16390 7868 16396 7880
rect 15528 7840 16396 7868
rect 15528 7828 15534 7840
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 16758 7868 16764 7880
rect 16623 7840 16764 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 17052 7877 17080 7908
rect 17696 7908 18184 7936
rect 16853 7871 16911 7877
rect 16853 7837 16865 7871
rect 16899 7837 16911 7871
rect 16853 7831 16911 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 13803 7772 14320 7800
rect 14384 7772 14780 7800
rect 15120 7800 15148 7828
rect 16868 7800 16896 7831
rect 17402 7828 17408 7880
rect 17460 7828 17466 7880
rect 17696 7877 17724 7908
rect 17954 7877 17960 7880
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 17921 7871 17960 7877
rect 17921 7837 17933 7871
rect 17921 7831 17960 7837
rect 15120 7772 16896 7800
rect 13803 7769 13815 7772
rect 13780 7763 13815 7769
rect 13780 7760 13786 7763
rect 6656 7704 6960 7732
rect 7190 7692 7196 7744
rect 7248 7692 7254 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 13740 7732 13768 7760
rect 13412 7704 13768 7732
rect 13412 7692 13418 7704
rect 13906 7692 13912 7744
rect 13964 7692 13970 7744
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 14384 7732 14412 7772
rect 17218 7760 17224 7812
rect 17276 7760 17282 7812
rect 17788 7800 17816 7831
rect 17954 7828 17960 7831
rect 18012 7828 18018 7880
rect 18046 7828 18052 7880
rect 18104 7828 18110 7880
rect 18156 7868 18184 7908
rect 20349 7905 20361 7939
rect 20395 7936 20407 7939
rect 20898 7936 20904 7948
rect 20395 7908 20904 7936
rect 20395 7905 20407 7908
rect 20349 7899 20407 7905
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 22462 7936 22468 7948
rect 22204 7908 22468 7936
rect 18238 7871 18296 7877
rect 18238 7868 18250 7871
rect 18156 7840 18250 7868
rect 18238 7837 18250 7840
rect 18284 7837 18296 7871
rect 18238 7831 18296 7837
rect 20070 7828 20076 7880
rect 20128 7828 20134 7880
rect 22002 7828 22008 7880
rect 22060 7828 22066 7880
rect 22204 7877 22232 7908
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 22278 7828 22284 7880
rect 22336 7828 22342 7880
rect 22554 7865 22560 7880
rect 22388 7837 22560 7865
rect 17420 7772 17816 7800
rect 18141 7803 18199 7809
rect 14056 7704 14412 7732
rect 14056 7692 14062 7704
rect 14458 7692 14464 7744
rect 14516 7692 14522 7744
rect 14642 7692 14648 7744
rect 14700 7692 14706 7744
rect 16758 7692 16764 7744
rect 16816 7732 16822 7744
rect 17420 7732 17448 7772
rect 18141 7769 18153 7803
rect 18187 7800 18199 7803
rect 21910 7800 21916 7812
rect 18187 7772 19288 7800
rect 21574 7772 21916 7800
rect 18187 7769 18199 7772
rect 18141 7763 18199 7769
rect 16816 7704 17448 7732
rect 16816 7692 16822 7704
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 18156 7732 18184 7763
rect 17552 7704 18184 7732
rect 17552 7692 17558 7704
rect 18414 7692 18420 7744
rect 18472 7692 18478 7744
rect 19260 7732 19288 7772
rect 21910 7760 21916 7772
rect 21968 7760 21974 7812
rect 22388 7800 22416 7837
rect 22554 7828 22560 7837
rect 22612 7828 22618 7880
rect 22664 7865 22692 7976
rect 23014 7964 23020 8016
rect 23072 8004 23078 8016
rect 24026 8004 24032 8016
rect 23072 7976 23158 8004
rect 23072 7964 23078 7976
rect 22859 7871 22917 7877
rect 22859 7868 22871 7871
rect 22848 7865 22871 7868
rect 22664 7837 22871 7865
rect 22905 7837 22917 7871
rect 22859 7831 22917 7837
rect 23014 7828 23020 7880
rect 23072 7828 23078 7880
rect 23130 7877 23158 7976
rect 23216 7976 24032 8004
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7837 23167 7871
rect 23109 7831 23167 7837
rect 22296 7772 22416 7800
rect 22649 7803 22707 7809
rect 22094 7732 22100 7744
rect 19260 7704 22100 7732
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22296 7741 22324 7772
rect 22649 7769 22661 7803
rect 22695 7769 22707 7803
rect 22649 7763 22707 7769
rect 22741 7803 22799 7809
rect 22741 7769 22753 7803
rect 22787 7800 22799 7803
rect 23216 7800 23244 7976
rect 24026 7964 24032 7976
rect 24084 8004 24090 8016
rect 26142 8004 26148 8016
rect 24084 7976 26148 8004
rect 24084 7964 24090 7976
rect 26142 7964 26148 7976
rect 26200 7964 26206 8016
rect 26326 7964 26332 8016
rect 26384 8004 26390 8016
rect 26384 7976 27568 8004
rect 26384 7964 26390 7976
rect 27540 7948 27568 7976
rect 23492 7908 23888 7936
rect 23492 7880 23520 7908
rect 23293 7871 23351 7877
rect 23293 7837 23305 7871
rect 23339 7868 23351 7871
rect 23382 7868 23388 7880
rect 23339 7840 23388 7868
rect 23339 7837 23351 7840
rect 23293 7831 23351 7837
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 23566 7828 23572 7880
rect 23624 7828 23630 7880
rect 23658 7828 23664 7880
rect 23716 7828 23722 7880
rect 23750 7828 23756 7880
rect 23808 7828 23814 7880
rect 23860 7877 23888 7908
rect 24210 7896 24216 7948
rect 24268 7936 24274 7948
rect 25498 7936 25504 7948
rect 24268 7908 24624 7936
rect 24268 7896 24274 7908
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7837 23903 7871
rect 23845 7831 23903 7837
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 22787 7772 23244 7800
rect 23584 7800 23612 7828
rect 24044 7800 24072 7831
rect 24118 7828 24124 7880
rect 24176 7868 24182 7880
rect 24596 7877 24624 7908
rect 24964 7908 25504 7936
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 24176 7840 24409 7868
rect 24176 7828 24182 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24728 7840 24869 7868
rect 24728 7828 24734 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 23584 7772 24072 7800
rect 22787 7769 22799 7772
rect 22741 7763 22799 7769
rect 22281 7735 22339 7741
rect 22281 7701 22293 7735
rect 22327 7701 22339 7735
rect 22281 7695 22339 7701
rect 22370 7692 22376 7744
rect 22428 7692 22434 7744
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 22664 7732 22692 7763
rect 24210 7760 24216 7812
rect 24268 7800 24274 7812
rect 24964 7800 24992 7908
rect 25498 7896 25504 7908
rect 25556 7936 25562 7948
rect 26237 7939 26295 7945
rect 25556 7908 26122 7936
rect 25556 7896 25562 7908
rect 26094 7877 26122 7908
rect 26237 7905 26249 7939
rect 26283 7936 26295 7939
rect 27157 7939 27215 7945
rect 27157 7936 27169 7939
rect 26283 7908 27169 7936
rect 26283 7905 26295 7908
rect 26237 7899 26295 7905
rect 27157 7905 27169 7908
rect 27203 7905 27215 7939
rect 27157 7899 27215 7905
rect 27522 7896 27528 7948
rect 27580 7896 27586 7948
rect 25041 7871 25099 7877
rect 25041 7837 25053 7871
rect 25087 7868 25099 7871
rect 25777 7871 25835 7877
rect 25087 7840 25176 7868
rect 25087 7837 25099 7840
rect 25041 7831 25099 7837
rect 24268 7772 24992 7800
rect 24268 7760 24274 7772
rect 22520 7704 22692 7732
rect 22520 7692 22526 7704
rect 23290 7692 23296 7744
rect 23348 7692 23354 7744
rect 23385 7735 23443 7741
rect 23385 7701 23397 7735
rect 23431 7732 23443 7735
rect 23658 7732 23664 7744
rect 23431 7704 23664 7732
rect 23431 7701 23443 7704
rect 23385 7695 23443 7701
rect 23658 7692 23664 7704
rect 23716 7692 23722 7744
rect 23750 7692 23756 7744
rect 23808 7732 23814 7744
rect 24765 7735 24823 7741
rect 24765 7732 24777 7735
rect 23808 7704 24777 7732
rect 23808 7692 23814 7704
rect 24765 7701 24777 7704
rect 24811 7732 24823 7735
rect 25148 7732 25176 7840
rect 25777 7837 25789 7871
rect 25823 7837 25835 7871
rect 25777 7831 25835 7837
rect 26079 7871 26137 7877
rect 26079 7837 26091 7871
rect 26125 7837 26137 7871
rect 26079 7831 26137 7837
rect 24811 7704 25176 7732
rect 24811 7701 24823 7704
rect 24765 7695 24823 7701
rect 25590 7692 25596 7744
rect 25648 7692 25654 7744
rect 25792 7732 25820 7831
rect 26510 7828 26516 7880
rect 26568 7828 26574 7880
rect 26602 7828 26608 7880
rect 26660 7868 26666 7880
rect 26970 7868 26976 7880
rect 26660 7840 26976 7868
rect 26660 7828 26666 7840
rect 26970 7828 26976 7840
rect 27028 7868 27034 7880
rect 27249 7871 27307 7877
rect 27249 7868 27261 7871
rect 27028 7840 27261 7868
rect 27028 7828 27034 7840
rect 27249 7837 27261 7840
rect 27295 7837 27307 7871
rect 27249 7831 27307 7837
rect 25866 7760 25872 7812
rect 25924 7760 25930 7812
rect 25961 7803 26019 7809
rect 25961 7769 25973 7803
rect 26007 7800 26019 7803
rect 26234 7800 26240 7812
rect 26007 7772 26240 7800
rect 26007 7769 26019 7772
rect 25961 7763 26019 7769
rect 26234 7760 26240 7772
rect 26292 7760 26298 7812
rect 26528 7800 26556 7828
rect 26786 7800 26792 7812
rect 26528 7772 26792 7800
rect 26786 7760 26792 7772
rect 26844 7760 26850 7812
rect 27801 7735 27859 7741
rect 27801 7732 27813 7735
rect 25792 7704 27813 7732
rect 27801 7701 27813 7704
rect 27847 7701 27859 7735
rect 27801 7695 27859 7701
rect 1104 7642 29440 7664
rect 1104 7590 5151 7642
rect 5203 7590 5215 7642
rect 5267 7590 5279 7642
rect 5331 7590 5343 7642
rect 5395 7590 5407 7642
rect 5459 7590 12234 7642
rect 12286 7590 12298 7642
rect 12350 7590 12362 7642
rect 12414 7590 12426 7642
rect 12478 7590 12490 7642
rect 12542 7590 19317 7642
rect 19369 7590 19381 7642
rect 19433 7590 19445 7642
rect 19497 7590 19509 7642
rect 19561 7590 19573 7642
rect 19625 7590 26400 7642
rect 26452 7590 26464 7642
rect 26516 7590 26528 7642
rect 26580 7590 26592 7642
rect 26644 7590 26656 7642
rect 26708 7590 29440 7642
rect 1104 7568 29440 7590
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 5132 7500 5641 7528
rect 5132 7488 5138 7500
rect 5629 7497 5641 7500
rect 5675 7497 5687 7531
rect 5629 7491 5687 7497
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 12342 7528 12348 7540
rect 6604 7500 12348 7528
rect 6604 7488 6610 7500
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 14642 7528 14648 7540
rect 12912 7500 14648 7528
rect 5828 7460 5856 7488
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 5828 7432 6132 7460
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5736 7364 6009 7392
rect 5736 7336 5764 7364
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 5810 7284 5816 7336
rect 5868 7284 5874 7336
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6104 7324 6132 7432
rect 10336 7432 11529 7460
rect 10336 7401 10364 7432
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 11517 7423 11575 7429
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10594 7352 10600 7404
rect 10652 7352 10658 7404
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7392 10931 7395
rect 11330 7392 11336 7404
rect 10919 7364 11336 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11422 7352 11428 7404
rect 11480 7352 11486 7404
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 12158 7392 12164 7404
rect 11839 7364 12164 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 12158 7352 12164 7364
rect 12216 7352 12222 7404
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7361 12311 7395
rect 12912 7392 12940 7500
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 16758 7488 16764 7540
rect 16816 7488 16822 7540
rect 16945 7531 17003 7537
rect 16945 7497 16957 7531
rect 16991 7528 17003 7531
rect 17126 7528 17132 7540
rect 16991 7500 17132 7528
rect 16991 7497 17003 7500
rect 16945 7491 17003 7497
rect 17126 7488 17132 7500
rect 17184 7488 17190 7540
rect 17402 7528 17408 7540
rect 17292 7500 17408 7528
rect 12989 7463 13047 7469
rect 12989 7429 13001 7463
rect 13035 7460 13047 7463
rect 13817 7463 13875 7469
rect 13817 7460 13829 7463
rect 13035 7432 13829 7460
rect 13035 7429 13047 7432
rect 12989 7423 13047 7429
rect 13817 7429 13829 7432
rect 13863 7429 13875 7463
rect 13817 7423 13875 7429
rect 14274 7420 14280 7472
rect 14332 7420 14338 7472
rect 16776 7460 16804 7488
rect 16776 7432 17172 7460
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 12912 7364 13185 7392
rect 12253 7355 12311 7361
rect 13173 7361 13185 7364
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 5951 7296 6132 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10612 7324 10640 7352
rect 9732 7296 10640 7324
rect 9732 7284 9738 7296
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10836 7296 11069 7324
rect 10836 7284 10842 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 11440 7324 11468 7352
rect 12268 7324 12296 7355
rect 13354 7352 13360 7404
rect 13412 7352 13418 7404
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 16761 7395 16819 7401
rect 16761 7361 16773 7395
rect 16807 7361 16819 7395
rect 16761 7355 16819 7361
rect 11440 7296 12296 7324
rect 13449 7327 13507 7333
rect 11057 7287 11115 7293
rect 13449 7293 13461 7327
rect 13495 7324 13507 7327
rect 14182 7324 14188 7336
rect 13495 7296 14188 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 14182 7284 14188 7296
rect 14240 7324 14246 7336
rect 15102 7324 15108 7336
rect 14240 7296 15108 7324
rect 14240 7284 14246 7296
rect 15102 7284 15108 7296
rect 15160 7324 15166 7336
rect 15565 7327 15623 7333
rect 15565 7324 15577 7327
rect 15160 7296 15577 7324
rect 15160 7284 15166 7296
rect 15565 7293 15577 7296
rect 15611 7293 15623 7327
rect 16776 7324 16804 7355
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 17144 7401 17172 7432
rect 17292 7401 17320 7500
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 17678 7488 17684 7540
rect 17736 7528 17742 7540
rect 18046 7528 18052 7540
rect 17736 7500 18052 7528
rect 17736 7488 17742 7500
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 22554 7488 22560 7540
rect 22612 7488 22618 7540
rect 22922 7488 22928 7540
rect 22980 7488 22986 7540
rect 23014 7488 23020 7540
rect 23072 7488 23078 7540
rect 23658 7488 23664 7540
rect 23716 7528 23722 7540
rect 23716 7500 24716 7528
rect 23716 7488 23722 7500
rect 17770 7420 17776 7472
rect 17828 7420 17834 7472
rect 22465 7463 22523 7469
rect 18248 7432 18552 7460
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 17277 7395 17335 7401
rect 17277 7361 17289 7395
rect 17323 7361 17335 7395
rect 17277 7355 17335 7361
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 17494 7352 17500 7404
rect 17552 7352 17558 7404
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17788 7392 17816 7420
rect 17635 7364 17816 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 17862 7352 17868 7404
rect 17920 7352 17926 7404
rect 18046 7352 18052 7404
rect 18104 7352 18110 7404
rect 18248 7401 18276 7432
rect 18524 7404 18552 7432
rect 22465 7429 22477 7463
rect 22511 7460 22523 7463
rect 23032 7460 23060 7488
rect 22511 7432 23060 7460
rect 23753 7463 23811 7469
rect 22511 7429 22523 7432
rect 22465 7423 22523 7429
rect 23753 7429 23765 7463
rect 23799 7460 23811 7463
rect 24121 7463 24179 7469
rect 24121 7460 24133 7463
rect 23799 7432 24133 7460
rect 23799 7429 23811 7432
rect 23753 7423 23811 7429
rect 24121 7429 24133 7432
rect 24167 7429 24179 7463
rect 24121 7423 24179 7429
rect 24578 7420 24584 7472
rect 24636 7420 24642 7472
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 18414 7352 18420 7404
rect 18472 7352 18478 7404
rect 18506 7352 18512 7404
rect 18564 7352 18570 7404
rect 22278 7352 22284 7404
rect 22336 7392 22342 7404
rect 22741 7395 22799 7401
rect 22741 7392 22753 7395
rect 22336 7364 22753 7392
rect 22336 7352 22342 7364
rect 22741 7361 22753 7364
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 22830 7352 22836 7404
rect 22888 7352 22894 7404
rect 23017 7395 23075 7401
rect 23017 7361 23029 7395
rect 23063 7392 23075 7395
rect 23290 7392 23296 7404
rect 23063 7364 23296 7392
rect 23063 7361 23075 7364
rect 23017 7355 23075 7361
rect 18325 7327 18383 7333
rect 18325 7324 18337 7327
rect 16776 7296 18337 7324
rect 15565 7287 15623 7293
rect 18325 7293 18337 7296
rect 18371 7293 18383 7327
rect 18325 7287 18383 7293
rect 21913 7327 21971 7333
rect 21913 7293 21925 7327
rect 21959 7324 21971 7327
rect 22186 7324 22192 7336
rect 21959 7296 22192 7324
rect 21959 7293 21971 7296
rect 21913 7287 21971 7293
rect 22186 7284 22192 7296
rect 22244 7324 22250 7336
rect 22848 7324 22876 7352
rect 22244 7296 22876 7324
rect 22244 7284 22250 7296
rect 12069 7259 12127 7265
rect 12069 7256 12081 7259
rect 11072 7228 12081 7256
rect 11072 7200 11100 7228
rect 12069 7225 12081 7228
rect 12115 7225 12127 7259
rect 12069 7219 12127 7225
rect 22002 7216 22008 7268
rect 22060 7256 22066 7268
rect 23032 7256 23060 7355
rect 23290 7352 23296 7364
rect 23348 7352 23354 7404
rect 23845 7395 23903 7401
rect 23845 7361 23857 7395
rect 23891 7361 23903 7395
rect 23845 7355 23903 7361
rect 23201 7327 23259 7333
rect 23201 7293 23213 7327
rect 23247 7293 23259 7327
rect 23860 7324 23888 7355
rect 24026 7352 24032 7404
rect 24084 7352 24090 7404
rect 24210 7352 24216 7404
rect 24268 7352 24274 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 24596 7392 24624 7420
rect 24688 7401 24716 7500
rect 25590 7488 25596 7540
rect 25648 7488 25654 7540
rect 25866 7488 25872 7540
rect 25924 7528 25930 7540
rect 27157 7531 27215 7537
rect 27157 7528 27169 7531
rect 25924 7500 27169 7528
rect 25924 7488 25930 7500
rect 27157 7497 27169 7500
rect 27203 7497 27215 7531
rect 27157 7491 27215 7497
rect 25225 7463 25283 7469
rect 25225 7429 25237 7463
rect 25271 7460 25283 7463
rect 25608 7460 25636 7488
rect 25271 7432 25636 7460
rect 26896 7432 27568 7460
rect 25271 7429 25283 7432
rect 25225 7423 25283 7429
rect 26896 7404 26924 7432
rect 24535 7364 24624 7392
rect 24673 7395 24731 7401
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 24673 7361 24685 7395
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 24946 7352 24952 7404
rect 25004 7352 25010 7404
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 23860 7296 24593 7324
rect 23201 7287 23259 7293
rect 24581 7293 24593 7296
rect 24627 7293 24639 7327
rect 24581 7287 24639 7293
rect 22060 7228 23060 7256
rect 23216 7256 23244 7287
rect 25314 7284 25320 7336
rect 25372 7324 25378 7336
rect 26344 7324 26372 7378
rect 26878 7352 26884 7404
rect 26936 7352 26942 7404
rect 26970 7352 26976 7404
rect 27028 7352 27034 7404
rect 27062 7352 27068 7404
rect 27120 7352 27126 7404
rect 27249 7395 27307 7401
rect 27249 7361 27261 7395
rect 27295 7392 27307 7395
rect 27338 7392 27344 7404
rect 27295 7364 27344 7392
rect 27295 7361 27307 7364
rect 27249 7355 27307 7361
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 27540 7401 27568 7432
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 27525 7395 27583 7401
rect 27525 7361 27537 7395
rect 27571 7361 27583 7395
rect 27709 7395 27767 7401
rect 27709 7392 27721 7395
rect 27525 7355 27583 7361
rect 27632 7364 27721 7392
rect 27080 7324 27108 7352
rect 25372 7296 27108 7324
rect 27448 7324 27476 7355
rect 27448 7296 27568 7324
rect 25372 7284 25378 7296
rect 27540 7268 27568 7296
rect 24118 7256 24124 7268
rect 23216 7228 24124 7256
rect 22060 7216 22066 7228
rect 24118 7216 24124 7228
rect 24176 7216 24182 7268
rect 26697 7259 26755 7265
rect 26697 7225 26709 7259
rect 26743 7256 26755 7259
rect 26786 7256 26792 7268
rect 26743 7228 26792 7256
rect 26743 7225 26755 7228
rect 26697 7219 26755 7225
rect 26786 7216 26792 7228
rect 26844 7216 26850 7268
rect 27522 7216 27528 7268
rect 27580 7216 27586 7268
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 7742 7188 7748 7200
rect 6328 7160 7748 7188
rect 6328 7148 6334 7160
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 11054 7148 11060 7200
rect 11112 7148 11118 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11882 7188 11888 7200
rect 11204 7160 11888 7188
rect 11204 7148 11210 7160
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 11974 7148 11980 7200
rect 12032 7148 12038 7200
rect 16758 7148 16764 7200
rect 16816 7148 16822 7200
rect 17129 7191 17187 7197
rect 17129 7157 17141 7191
rect 17175 7188 17187 7191
rect 17402 7188 17408 7200
rect 17175 7160 17408 7188
rect 17175 7157 17187 7160
rect 17129 7151 17187 7157
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 17862 7148 17868 7200
rect 17920 7148 17926 7200
rect 24394 7148 24400 7200
rect 24452 7148 24458 7200
rect 26804 7188 26832 7216
rect 27632 7188 27660 7364
rect 27709 7361 27721 7364
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 28718 7352 28724 7404
rect 28776 7352 28782 7404
rect 26804 7160 27660 7188
rect 28902 7148 28908 7200
rect 28960 7188 28966 7200
rect 28997 7191 29055 7197
rect 28997 7188 29009 7191
rect 28960 7160 29009 7188
rect 28960 7148 28966 7160
rect 28997 7157 29009 7160
rect 29043 7157 29055 7191
rect 28997 7151 29055 7157
rect 1104 7098 29440 7120
rect 1104 7046 4491 7098
rect 4543 7046 4555 7098
rect 4607 7046 4619 7098
rect 4671 7046 4683 7098
rect 4735 7046 4747 7098
rect 4799 7046 11574 7098
rect 11626 7046 11638 7098
rect 11690 7046 11702 7098
rect 11754 7046 11766 7098
rect 11818 7046 11830 7098
rect 11882 7046 18657 7098
rect 18709 7046 18721 7098
rect 18773 7046 18785 7098
rect 18837 7046 18849 7098
rect 18901 7046 18913 7098
rect 18965 7046 25740 7098
rect 25792 7046 25804 7098
rect 25856 7046 25868 7098
rect 25920 7046 25932 7098
rect 25984 7046 25996 7098
rect 26048 7046 29440 7098
rect 1104 7024 29440 7046
rect 4890 6984 4896 6996
rect 4816 6956 4896 6984
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4816 6780 4844 6956
rect 4890 6944 4896 6956
rect 4948 6984 4954 6996
rect 8110 6984 8116 6996
rect 4948 6956 7052 6984
rect 4948 6944 4954 6956
rect 5074 6876 5080 6928
rect 5132 6876 5138 6928
rect 5276 6888 6408 6916
rect 4571 6752 4844 6780
rect 4893 6783 4951 6789
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 4893 6749 4905 6783
rect 4939 6780 4951 6783
rect 5276 6780 5304 6888
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5902 6848 5908 6860
rect 5399 6820 5908 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 6270 6848 6276 6860
rect 6012 6820 6276 6848
rect 6012 6789 6040 6820
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 4939 6752 5304 6780
rect 5997 6783 6055 6789
rect 4939 6749 4951 6752
rect 4893 6743 4951 6749
rect 5997 6749 6009 6783
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6086 6740 6092 6792
rect 6144 6740 6150 6792
rect 6380 6789 6408 6888
rect 7024 6860 7052 6956
rect 7576 6956 8116 6984
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 7377 6919 7435 6925
rect 7377 6916 7389 6919
rect 7340 6888 7389 6916
rect 7340 6876 7346 6888
rect 7377 6885 7389 6888
rect 7423 6885 7435 6919
rect 7377 6879 7435 6885
rect 7006 6808 7012 6860
rect 7064 6848 7070 6860
rect 7576 6848 7604 6956
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 11149 6987 11207 6993
rect 11149 6984 11161 6987
rect 10468 6956 11161 6984
rect 10468 6944 10474 6956
rect 11149 6953 11161 6956
rect 11195 6984 11207 6987
rect 11238 6984 11244 6996
rect 11195 6956 11244 6984
rect 11195 6953 11207 6956
rect 11149 6947 11207 6953
rect 11238 6944 11244 6956
rect 11296 6984 11302 6996
rect 11698 6984 11704 6996
rect 11296 6956 11704 6984
rect 11296 6944 11302 6956
rect 11698 6944 11704 6956
rect 11756 6984 11762 6996
rect 12161 6987 12219 6993
rect 12161 6984 12173 6987
rect 11756 6956 12173 6984
rect 11756 6944 11762 6956
rect 12161 6953 12173 6956
rect 12207 6953 12219 6987
rect 12161 6947 12219 6953
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12400 6956 14412 6984
rect 12400 6944 12406 6956
rect 10134 6876 10140 6928
rect 10192 6916 10198 6928
rect 10192 6888 11284 6916
rect 10192 6876 10198 6888
rect 9858 6848 9864 6860
rect 7064 6820 7144 6848
rect 7064 6808 7070 6820
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6730 6780 6736 6792
rect 6411 6752 6736 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7116 6789 7144 6820
rect 7392 6820 7604 6848
rect 8220 6820 9864 6848
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7239 6783 7297 6789
rect 7239 6749 7251 6783
rect 7285 6780 7297 6783
rect 7392 6780 7420 6820
rect 7285 6752 7420 6780
rect 7285 6749 7297 6752
rect 7239 6743 7297 6749
rect 4709 6715 4767 6721
rect 4709 6681 4721 6715
rect 4755 6681 4767 6715
rect 4709 6675 4767 6681
rect 4801 6715 4859 6721
rect 4801 6681 4813 6715
rect 4847 6712 4859 6715
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 4847 6684 5917 6712
rect 4847 6681 4859 6684
rect 4801 6675 4859 6681
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 5905 6675 5963 6681
rect 6104 6712 6132 6740
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 6104 6684 6193 6712
rect 4724 6644 4752 6675
rect 6104 6644 6132 6684
rect 6181 6681 6193 6684
rect 6227 6681 6239 6715
rect 6181 6675 6239 6681
rect 6270 6672 6276 6724
rect 6328 6672 6334 6724
rect 6840 6656 6868 6743
rect 7466 6740 7472 6792
rect 7524 6740 7530 6792
rect 7650 6740 7656 6792
rect 7708 6740 7714 6792
rect 7883 6783 7941 6789
rect 7883 6749 7895 6783
rect 7929 6780 7941 6783
rect 8110 6780 8116 6792
rect 7929 6752 8116 6780
rect 7929 6749 7941 6752
rect 7883 6743 7941 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 7009 6715 7067 6721
rect 7009 6681 7021 6715
rect 7055 6712 7067 6715
rect 7055 6684 7420 6712
rect 7055 6681 7067 6684
rect 7009 6675 7067 6681
rect 4724 6616 6132 6644
rect 6546 6604 6552 6656
rect 6604 6604 6610 6656
rect 6822 6604 6828 6656
rect 6880 6604 6886 6656
rect 7392 6644 7420 6684
rect 7742 6672 7748 6724
rect 7800 6712 7806 6724
rect 8220 6712 8248 6820
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 11146 6848 11152 6860
rect 9968 6820 11152 6848
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 9968 6789 9996 6820
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11256 6848 11284 6888
rect 11330 6876 11336 6928
rect 11388 6876 11394 6928
rect 12066 6876 12072 6928
rect 12124 6876 12130 6928
rect 13906 6916 13912 6928
rect 13740 6888 13912 6916
rect 11422 6848 11428 6860
rect 11256 6820 11428 6848
rect 11422 6808 11428 6820
rect 11480 6808 11486 6860
rect 12084 6848 12112 6876
rect 12084 6820 12204 6848
rect 9953 6783 10011 6789
rect 8352 6752 9904 6780
rect 8352 6740 8358 6752
rect 9876 6724 9904 6752
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 11054 6780 11060 6792
rect 10827 6752 11060 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11974 6780 11980 6792
rect 11388 6752 11980 6780
rect 11388 6740 11394 6752
rect 11974 6740 11980 6752
rect 12032 6780 12038 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 12032 6752 12081 6780
rect 12032 6740 12038 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 7800 6684 8248 6712
rect 7800 6672 7806 6684
rect 9766 6672 9772 6724
rect 9824 6672 9830 6724
rect 9858 6672 9864 6724
rect 9916 6672 9922 6724
rect 10042 6672 10048 6724
rect 10100 6672 10106 6724
rect 10505 6715 10563 6721
rect 10505 6681 10517 6715
rect 10551 6681 10563 6715
rect 10505 6675 10563 6681
rect 7650 6644 7656 6656
rect 7392 6616 7656 6644
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 8018 6604 8024 6656
rect 8076 6604 8082 6656
rect 9784 6644 9812 6672
rect 10520 6644 10548 6675
rect 10594 6672 10600 6724
rect 10652 6712 10658 6724
rect 11609 6715 11667 6721
rect 11609 6712 11621 6715
rect 10652 6684 11621 6712
rect 10652 6672 10658 6684
rect 11609 6681 11621 6684
rect 11655 6681 11667 6715
rect 11609 6675 11667 6681
rect 11698 6672 11704 6724
rect 11756 6672 11762 6724
rect 11793 6715 11851 6721
rect 11793 6681 11805 6715
rect 11839 6712 11851 6715
rect 12176 6712 12204 6820
rect 13630 6808 13636 6860
rect 13688 6808 13694 6860
rect 11839 6684 12204 6712
rect 13648 6712 13676 6808
rect 13740 6789 13768 6888
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 14384 6916 14412 6956
rect 14458 6944 14464 6996
rect 14516 6944 14522 6996
rect 16574 6944 16580 6996
rect 16632 6944 16638 6996
rect 16758 6944 16764 6996
rect 16816 6984 16822 6996
rect 17770 6984 17776 6996
rect 16816 6956 17776 6984
rect 16816 6944 16822 6956
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 20796 6987 20854 6993
rect 20796 6953 20808 6987
rect 20842 6984 20854 6987
rect 22370 6984 22376 6996
rect 20842 6956 22376 6984
rect 20842 6953 20854 6956
rect 20796 6947 20854 6953
rect 22370 6944 22376 6956
rect 22428 6944 22434 6996
rect 22728 6987 22786 6993
rect 22728 6953 22740 6987
rect 22774 6984 22786 6987
rect 24394 6984 24400 6996
rect 22774 6956 24400 6984
rect 22774 6953 22786 6956
rect 22728 6947 22786 6953
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 16592 6916 16620 6944
rect 14384 6888 16620 6916
rect 17586 6876 17592 6928
rect 17644 6916 17650 6928
rect 17644 6888 18092 6916
rect 17644 6876 17650 6888
rect 13817 6851 13875 6857
rect 13817 6817 13829 6851
rect 13863 6848 13875 6851
rect 13863 6820 14320 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13906 6740 13912 6792
rect 13964 6740 13970 6792
rect 14292 6789 14320 6820
rect 17144 6820 17632 6848
rect 17144 6792 17172 6820
rect 17604 6792 17632 6820
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 14568 6712 14596 6743
rect 15470 6712 15476 6724
rect 13648 6684 15476 6712
rect 11839 6681 11851 6684
rect 11793 6675 11851 6681
rect 9784 6616 10548 6644
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11808 6644 11836 6675
rect 15470 6672 15476 6684
rect 15528 6672 15534 6724
rect 17052 6712 17080 6743
rect 17126 6740 17132 6792
rect 17184 6740 17190 6792
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 17276 6752 17325 6780
rect 17276 6740 17282 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17402 6740 17408 6792
rect 17460 6740 17466 6792
rect 17586 6740 17592 6792
rect 17644 6740 17650 6792
rect 17678 6740 17684 6792
rect 17736 6740 17742 6792
rect 17770 6740 17776 6792
rect 17828 6780 17834 6792
rect 18064 6789 18092 6888
rect 22186 6876 22192 6928
rect 22244 6916 22250 6928
rect 22281 6919 22339 6925
rect 22281 6916 22293 6919
rect 22244 6888 22293 6916
rect 22244 6876 22250 6888
rect 22281 6885 22293 6888
rect 22327 6885 22339 6919
rect 22281 6879 22339 6885
rect 23842 6876 23848 6928
rect 23900 6876 23906 6928
rect 24026 6876 24032 6928
rect 24084 6876 24090 6928
rect 24118 6876 24124 6928
rect 24176 6916 24182 6928
rect 24213 6919 24271 6925
rect 24213 6916 24225 6919
rect 24176 6888 24225 6916
rect 24176 6876 24182 6888
rect 24213 6885 24225 6888
rect 24259 6885 24271 6919
rect 24213 6879 24271 6885
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20533 6851 20591 6857
rect 20533 6848 20545 6851
rect 20128 6820 20545 6848
rect 20128 6808 20134 6820
rect 20533 6817 20545 6820
rect 20579 6848 20591 6851
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 20579 6820 22477 6848
rect 20579 6817 20591 6820
rect 20533 6811 20591 6817
rect 22465 6817 22477 6820
rect 22511 6848 22523 6851
rect 22738 6848 22744 6860
rect 22511 6820 22744 6848
rect 22511 6817 22523 6820
rect 22465 6811 22523 6817
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 23860 6848 23888 6876
rect 24044 6848 24072 6876
rect 24489 6851 24547 6857
rect 24489 6848 24501 6851
rect 23860 6820 23980 6848
rect 24044 6820 24501 6848
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17828 6752 17877 6780
rect 17828 6740 17834 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 23952 6780 23980 6820
rect 24489 6817 24501 6820
rect 24535 6817 24547 6851
rect 24489 6811 24547 6817
rect 24210 6780 24216 6792
rect 21968 6752 22140 6780
rect 23952 6752 24216 6780
rect 21968 6740 21974 6752
rect 17420 6712 17448 6740
rect 17052 6684 17448 6712
rect 11204 6616 11836 6644
rect 11977 6647 12035 6653
rect 11204 6604 11210 6616
rect 11977 6613 11989 6647
rect 12023 6644 12035 6647
rect 12158 6644 12164 6656
rect 12023 6616 12164 6644
rect 12023 6613 12035 6616
rect 11977 6607 12035 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 17126 6644 17132 6656
rect 16899 6616 17132 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 17221 6647 17279 6653
rect 17221 6613 17233 6647
rect 17267 6644 17279 6647
rect 17696 6644 17724 6740
rect 17267 6616 17724 6644
rect 17267 6613 17279 6616
rect 17221 6607 17279 6613
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 17954 6604 17960 6656
rect 18012 6604 18018 6656
rect 22112 6644 22140 6752
rect 24210 6740 24216 6752
rect 24268 6780 24274 6792
rect 24397 6783 24455 6789
rect 24397 6780 24409 6783
rect 24268 6752 24409 6780
rect 24268 6740 24274 6752
rect 24397 6749 24409 6752
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 23966 6684 24256 6712
rect 24228 6644 24256 6684
rect 24302 6672 24308 6724
rect 24360 6712 24366 6724
rect 24596 6712 24624 6743
rect 24360 6684 24624 6712
rect 24360 6672 24366 6684
rect 25314 6672 25320 6724
rect 25372 6672 25378 6724
rect 25332 6644 25360 6672
rect 22112 6616 25360 6644
rect 1104 6554 29440 6576
rect 1104 6502 5151 6554
rect 5203 6502 5215 6554
rect 5267 6502 5279 6554
rect 5331 6502 5343 6554
rect 5395 6502 5407 6554
rect 5459 6502 12234 6554
rect 12286 6502 12298 6554
rect 12350 6502 12362 6554
rect 12414 6502 12426 6554
rect 12478 6502 12490 6554
rect 12542 6502 19317 6554
rect 19369 6502 19381 6554
rect 19433 6502 19445 6554
rect 19497 6502 19509 6554
rect 19561 6502 19573 6554
rect 19625 6502 26400 6554
rect 26452 6502 26464 6554
rect 26516 6502 26528 6554
rect 26580 6502 26592 6554
rect 26644 6502 26656 6554
rect 26708 6502 29440 6554
rect 1104 6480 29440 6502
rect 5074 6440 5080 6452
rect 4172 6412 5080 6440
rect 4172 6381 4200 6412
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 5902 6440 5908 6452
rect 5675 6412 5908 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6328 6412 7021 6440
rect 6328 6400 6334 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 7009 6403 7067 6409
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 7524 6412 8769 6440
rect 7524 6400 7530 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 8757 6403 8815 6409
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10284 6412 10885 6440
rect 10284 6400 10290 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 11057 6443 11115 6449
rect 11057 6409 11069 6443
rect 11103 6440 11115 6443
rect 11422 6440 11428 6452
rect 11103 6412 11428 6440
rect 11103 6409 11115 6412
rect 11057 6403 11115 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 12158 6400 12164 6452
rect 12216 6400 12222 6452
rect 14090 6440 14096 6452
rect 13740 6412 14096 6440
rect 4157 6375 4215 6381
rect 4157 6341 4169 6375
rect 4203 6341 4215 6375
rect 4157 6335 4215 6341
rect 6822 6332 6828 6384
rect 6880 6372 6886 6384
rect 8021 6375 8079 6381
rect 8021 6372 8033 6375
rect 6880 6344 8033 6372
rect 6880 6332 6886 6344
rect 8021 6341 8033 6344
rect 8067 6341 8079 6375
rect 8021 6335 8079 6341
rect 9858 6332 9864 6384
rect 9916 6372 9922 6384
rect 10045 6375 10103 6381
rect 10045 6372 10057 6375
rect 9916 6344 10057 6372
rect 9916 6332 9922 6344
rect 10045 6341 10057 6344
rect 10091 6372 10103 6375
rect 10505 6375 10563 6381
rect 10505 6372 10517 6375
rect 10091 6344 10517 6372
rect 10091 6341 10103 6344
rect 10045 6335 10103 6341
rect 10505 6341 10517 6344
rect 10551 6372 10563 6375
rect 10594 6372 10600 6384
rect 10551 6344 10600 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 3881 6307 3939 6313
rect 3881 6304 3893 6307
rect 2740 6276 3893 6304
rect 2740 6264 2746 6276
rect 3881 6273 3893 6276
rect 3927 6273 3939 6307
rect 7098 6304 7104 6316
rect 5290 6276 7104 6304
rect 3881 6267 3939 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7248 6276 7389 6304
rect 7248 6264 7254 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 8202 6264 8208 6316
rect 8260 6264 8266 6316
rect 9953 6307 10011 6313
rect 9953 6273 9965 6307
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5776 6208 6377 6236
rect 5776 6196 5782 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 9674 6236 9680 6248
rect 6788 6208 9680 6236
rect 6788 6196 6794 6208
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 9968 6236 9996 6267
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 10192 6276 10241 6304
rect 10192 6264 10198 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 10714 6307 10772 6313
rect 10468 6276 10640 6304
rect 10468 6264 10474 6276
rect 10502 6236 10508 6248
rect 9968 6208 10508 6236
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10612 6245 10640 6276
rect 10714 6273 10726 6307
rect 10760 6273 10772 6307
rect 10714 6267 10772 6273
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 6086 6128 6092 6180
rect 6144 6128 6150 6180
rect 8110 6128 8116 6180
rect 8168 6168 8174 6180
rect 10729 6168 10757 6267
rect 10962 6264 10968 6316
rect 11020 6313 11026 6316
rect 11020 6267 11029 6313
rect 11020 6264 11026 6267
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 12176 6304 12204 6400
rect 13740 6381 13768 6412
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16632 6412 17141 6440
rect 16632 6400 16638 6412
rect 17129 6409 17141 6412
rect 17175 6440 17187 6443
rect 17770 6440 17776 6452
rect 17175 6412 17776 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 17954 6400 17960 6452
rect 18012 6400 18018 6452
rect 20070 6400 20076 6452
rect 20128 6400 20134 6452
rect 20625 6443 20683 6449
rect 20625 6409 20637 6443
rect 20671 6440 20683 6443
rect 28718 6440 28724 6452
rect 20671 6412 28724 6440
rect 20671 6409 20683 6412
rect 20625 6403 20683 6409
rect 28718 6400 28724 6412
rect 28776 6400 28782 6452
rect 13725 6375 13783 6381
rect 13725 6341 13737 6375
rect 13771 6341 13783 6375
rect 13725 6335 13783 6341
rect 14182 6332 14188 6384
rect 14240 6332 14246 6384
rect 15470 6332 15476 6384
rect 15528 6332 15534 6384
rect 16850 6332 16856 6384
rect 16908 6372 16914 6384
rect 16945 6375 17003 6381
rect 16945 6372 16957 6375
rect 16908 6344 16957 6372
rect 16908 6332 16914 6344
rect 16945 6341 16957 6344
rect 16991 6372 17003 6375
rect 17862 6372 17868 6384
rect 16991 6344 17868 6372
rect 16991 6341 17003 6344
rect 16945 6335 17003 6341
rect 17862 6332 17868 6344
rect 17920 6332 17926 6384
rect 11563 6276 12204 6304
rect 17221 6307 17279 6313
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 17221 6273 17233 6307
rect 17267 6304 17279 6307
rect 17972 6304 18000 6400
rect 20272 6344 20852 6372
rect 20272 6316 20300 6344
rect 17267 6276 18000 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 20070 6264 20076 6316
rect 20128 6264 20134 6316
rect 20254 6264 20260 6316
rect 20312 6264 20318 6316
rect 20441 6307 20499 6313
rect 20441 6273 20453 6307
rect 20487 6273 20499 6307
rect 20441 6267 20499 6273
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11146 6168 11152 6180
rect 8168 6140 9904 6168
rect 10729 6140 11152 6168
rect 8168 6128 8174 6140
rect 6104 6100 6132 6128
rect 9766 6100 9772 6112
rect 6104 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 9876 6100 9904 6140
rect 11146 6128 11152 6140
rect 11204 6128 11210 6180
rect 11716 6100 11744 6199
rect 12618 6196 12624 6248
rect 12676 6236 12682 6248
rect 13446 6236 13452 6248
rect 12676 6208 13452 6236
rect 12676 6196 12682 6208
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 20088 6236 20116 6264
rect 20456 6236 20484 6267
rect 20530 6264 20536 6316
rect 20588 6264 20594 6316
rect 20824 6313 20852 6344
rect 20809 6307 20867 6313
rect 20809 6273 20821 6307
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 20993 6307 21051 6313
rect 20993 6273 21005 6307
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6273 21143 6307
rect 21085 6267 21143 6273
rect 21008 6236 21036 6267
rect 20088 6208 21036 6236
rect 9876 6072 11744 6100
rect 16945 6103 17003 6109
rect 16945 6069 16957 6103
rect 16991 6100 17003 6103
rect 17586 6100 17592 6112
rect 16991 6072 17592 6100
rect 16991 6069 17003 6072
rect 16945 6063 17003 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 21100 6100 21128 6267
rect 20496 6072 21128 6100
rect 20496 6060 20502 6072
rect 1104 6010 29440 6032
rect 1104 5958 4491 6010
rect 4543 5958 4555 6010
rect 4607 5958 4619 6010
rect 4671 5958 4683 6010
rect 4735 5958 4747 6010
rect 4799 5958 11574 6010
rect 11626 5958 11638 6010
rect 11690 5958 11702 6010
rect 11754 5958 11766 6010
rect 11818 5958 11830 6010
rect 11882 5958 18657 6010
rect 18709 5958 18721 6010
rect 18773 5958 18785 6010
rect 18837 5958 18849 6010
rect 18901 5958 18913 6010
rect 18965 5958 25740 6010
rect 25792 5958 25804 6010
rect 25856 5958 25868 6010
rect 25920 5958 25932 6010
rect 25984 5958 25996 6010
rect 26048 5958 29440 6010
rect 1104 5936 29440 5958
rect 4236 5899 4294 5905
rect 4236 5865 4248 5899
rect 4282 5896 4294 5899
rect 6546 5896 6552 5908
rect 4282 5868 6552 5896
rect 4282 5865 4294 5868
rect 4236 5859 4294 5865
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7248 5868 8033 5896
rect 7248 5856 7254 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 10042 5896 10048 5908
rect 8021 5859 8079 5865
rect 9416 5868 10048 5896
rect 5718 5788 5724 5840
rect 5776 5788 5782 5840
rect 2682 5720 2688 5772
rect 2740 5720 2746 5772
rect 6270 5760 6276 5772
rect 3988 5732 6276 5760
rect 2700 5692 2728 5720
rect 3988 5701 4016 5732
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 7282 5760 7288 5772
rect 6595 5732 7288 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 9416 5701 9444 5868
rect 10042 5856 10048 5868
rect 10100 5896 10106 5908
rect 10781 5899 10839 5905
rect 10781 5896 10793 5899
rect 10100 5868 10793 5896
rect 10100 5856 10106 5868
rect 10781 5865 10793 5868
rect 10827 5865 10839 5899
rect 10781 5859 10839 5865
rect 11054 5856 11060 5908
rect 11112 5856 11118 5908
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17000 5868 17693 5896
rect 17000 5856 17006 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 9692 5800 10364 5828
rect 9692 5701 9720 5800
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9916 5732 10057 5760
rect 9916 5720 9922 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 10134 5720 10140 5772
rect 10192 5720 10198 5772
rect 10336 5760 10364 5800
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 17865 5831 17923 5837
rect 17865 5828 17877 5831
rect 17276 5800 17877 5828
rect 17276 5788 17282 5800
rect 17865 5797 17877 5800
rect 17911 5797 17923 5831
rect 17865 5791 17923 5797
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 10336 5732 10885 5760
rect 10873 5729 10885 5732
rect 10919 5760 10931 5763
rect 11422 5760 11428 5772
rect 10919 5732 11428 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 11422 5720 11428 5732
rect 11480 5760 11486 5772
rect 11480 5732 11652 5760
rect 11480 5720 11486 5732
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 2700 5664 3985 5692
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5692 10287 5695
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10275 5664 10425 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 7006 5624 7012 5636
rect 5474 5596 7012 5624
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 7098 5584 7104 5636
rect 7156 5584 7162 5636
rect 9585 5627 9643 5633
rect 9585 5593 9597 5627
rect 9631 5593 9643 5627
rect 9968 5624 9996 5655
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 10560 5664 10609 5692
rect 10560 5652 10566 5664
rect 10597 5661 10609 5664
rect 10643 5692 10655 5695
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10643 5664 10977 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 11146 5652 11152 5704
rect 11204 5652 11210 5704
rect 11238 5652 11244 5704
rect 11296 5652 11302 5704
rect 11624 5701 11652 5732
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 18506 5760 18512 5772
rect 17460 5732 18512 5760
rect 17460 5720 17466 5732
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11348 5664 11529 5692
rect 11256 5624 11284 5652
rect 11348 5636 11376 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 17494 5652 17500 5704
rect 17552 5652 17558 5704
rect 17604 5701 17632 5732
rect 18248 5701 18276 5732
rect 18506 5720 18512 5732
rect 18564 5720 18570 5772
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5661 17647 5695
rect 18141 5695 18199 5701
rect 18141 5692 18153 5695
rect 17589 5655 17647 5661
rect 17972 5664 18153 5692
rect 9968 5596 11284 5624
rect 9585 5587 9643 5593
rect 9217 5559 9275 5565
rect 9217 5525 9229 5559
rect 9263 5556 9275 5559
rect 9306 5556 9312 5568
rect 9263 5528 9312 5556
rect 9263 5525 9275 5528
rect 9217 5519 9275 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 9600 5556 9628 5587
rect 11330 5584 11336 5636
rect 11388 5584 11394 5636
rect 11422 5584 11428 5636
rect 11480 5584 11486 5636
rect 16022 5584 16028 5636
rect 16080 5624 16086 5636
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 16080 5596 17417 5624
rect 16080 5584 16086 5596
rect 17405 5593 17417 5596
rect 17451 5624 17463 5627
rect 17512 5624 17540 5652
rect 17770 5624 17776 5636
rect 17451 5596 17776 5624
rect 17451 5593 17463 5596
rect 17405 5587 17463 5593
rect 17770 5584 17776 5596
rect 17828 5624 17834 5636
rect 17865 5627 17923 5633
rect 17865 5624 17877 5627
rect 17828 5596 17877 5624
rect 17828 5584 17834 5596
rect 17865 5593 17877 5596
rect 17911 5593 17923 5627
rect 17865 5587 17923 5593
rect 17972 5568 18000 5664
rect 18141 5661 18153 5664
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 18414 5652 18420 5704
rect 18472 5692 18478 5704
rect 18472 5664 18515 5692
rect 18472 5652 18478 5664
rect 9674 5556 9680 5568
rect 9600 5528 9680 5556
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 9766 5516 9772 5568
rect 9824 5516 9830 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 11146 5556 11152 5568
rect 10192 5528 11152 5556
rect 10192 5516 10198 5528
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 11790 5516 11796 5568
rect 11848 5516 11854 5568
rect 17954 5516 17960 5568
rect 18012 5516 18018 5568
rect 18049 5559 18107 5565
rect 18049 5525 18061 5559
rect 18095 5556 18107 5559
rect 18230 5556 18236 5568
rect 18095 5528 18236 5556
rect 18095 5525 18107 5528
rect 18049 5519 18107 5525
rect 18230 5516 18236 5528
rect 18288 5556 18294 5568
rect 18325 5559 18383 5565
rect 18325 5556 18337 5559
rect 18288 5528 18337 5556
rect 18288 5516 18294 5528
rect 18325 5525 18337 5528
rect 18371 5525 18383 5559
rect 18325 5519 18383 5525
rect 1104 5466 29440 5488
rect 1104 5414 5151 5466
rect 5203 5414 5215 5466
rect 5267 5414 5279 5466
rect 5331 5414 5343 5466
rect 5395 5414 5407 5466
rect 5459 5414 12234 5466
rect 12286 5414 12298 5466
rect 12350 5414 12362 5466
rect 12414 5414 12426 5466
rect 12478 5414 12490 5466
rect 12542 5414 19317 5466
rect 19369 5414 19381 5466
rect 19433 5414 19445 5466
rect 19497 5414 19509 5466
rect 19561 5414 19573 5466
rect 19625 5414 26400 5466
rect 26452 5414 26464 5466
rect 26516 5414 26528 5466
rect 26580 5414 26592 5466
rect 26644 5414 26656 5466
rect 26708 5414 29440 5466
rect 1104 5392 29440 5414
rect 8113 5355 8171 5361
rect 8113 5321 8125 5355
rect 8159 5352 8171 5355
rect 8202 5352 8208 5364
rect 8159 5324 8208 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 8938 5352 8944 5364
rect 8496 5324 8944 5352
rect 7098 5244 7104 5296
rect 7156 5244 7162 5296
rect 8018 5244 8024 5296
rect 8076 5244 8082 5296
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6328 5188 6377 5216
rect 6328 5176 6334 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5148 6699 5151
rect 8036 5148 8064 5244
rect 8496 5225 8524 5324
rect 8938 5312 8944 5324
rect 8996 5352 9002 5364
rect 12618 5352 12624 5364
rect 8996 5324 12624 5352
rect 8996 5312 9002 5324
rect 10321 5287 10379 5293
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 9766 5176 9772 5228
rect 9824 5176 9830 5228
rect 9876 5216 9904 5270
rect 10321 5253 10333 5287
rect 10367 5284 10379 5287
rect 10502 5284 10508 5296
rect 10367 5256 10508 5284
rect 10367 5253 10379 5256
rect 10321 5247 10379 5253
rect 10502 5244 10508 5256
rect 10560 5244 10566 5296
rect 10226 5216 10232 5228
rect 9876 5188 10232 5216
rect 10226 5176 10232 5188
rect 10284 5216 10290 5228
rect 11532 5225 11560 5324
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 16482 5352 16488 5364
rect 13872 5324 16488 5352
rect 13872 5312 13878 5324
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16879 5355 16937 5361
rect 16879 5321 16891 5355
rect 16925 5352 16937 5355
rect 17218 5352 17224 5364
rect 16925 5324 17224 5352
rect 16925 5321 16937 5324
rect 16879 5315 16937 5321
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 17368 5324 19656 5352
rect 17368 5312 17374 5324
rect 16669 5287 16727 5293
rect 11517 5219 11575 5225
rect 10284 5188 11192 5216
rect 10284 5176 10290 5188
rect 6687 5120 8064 5148
rect 8849 5151 8907 5157
rect 6687 5117 6699 5120
rect 6641 5111 6699 5117
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9784 5148 9812 5176
rect 8895 5120 9812 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10413 5151 10471 5157
rect 10413 5148 10425 5151
rect 10192 5120 10425 5148
rect 10192 5108 10198 5120
rect 10413 5117 10425 5120
rect 10459 5148 10471 5151
rect 10686 5148 10692 5160
rect 10459 5120 10692 5148
rect 10459 5117 10471 5120
rect 10413 5111 10471 5117
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 9674 5040 9680 5092
rect 9732 5080 9738 5092
rect 11057 5083 11115 5089
rect 11057 5080 11069 5083
rect 9732 5052 11069 5080
rect 9732 5040 9738 5052
rect 11057 5049 11069 5052
rect 11103 5049 11115 5083
rect 11057 5043 11115 5049
rect 11164 5012 11192 5188
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11848 5188 11897 5216
rect 11848 5176 11854 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12636 5216 12664 5270
rect 16669 5253 16681 5287
rect 16715 5284 16727 5287
rect 16715 5256 17724 5284
rect 16715 5253 16727 5256
rect 16669 5247 16727 5253
rect 17696 5228 17724 5256
rect 17880 5256 19012 5284
rect 17880 5228 17908 5256
rect 14182 5216 14188 5228
rect 12636 5188 14188 5216
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12434 5148 12440 5160
rect 11388 5120 12440 5148
rect 11388 5108 11394 5120
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12636 5012 12664 5188
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 16114 5176 16120 5228
rect 16172 5216 16178 5228
rect 17034 5216 17040 5228
rect 16172 5188 17040 5216
rect 16172 5176 16178 5188
rect 17034 5176 17040 5188
rect 17092 5216 17098 5228
rect 17129 5219 17187 5225
rect 17129 5216 17141 5219
rect 17092 5188 17141 5216
rect 17092 5176 17098 5188
rect 17129 5185 17141 5188
rect 17175 5216 17187 5219
rect 17402 5216 17408 5228
rect 17175 5188 17408 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17736 5188 17785 5216
rect 17736 5176 17742 5188
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 17862 5176 17868 5228
rect 17920 5176 17926 5228
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 13311 5151 13369 5157
rect 13311 5148 13323 5151
rect 12768 5120 13323 5148
rect 12768 5108 12774 5120
rect 13311 5117 13323 5120
rect 13357 5117 13369 5151
rect 13311 5111 13369 5117
rect 17497 5151 17555 5157
rect 17497 5117 17509 5151
rect 17543 5148 17555 5151
rect 17696 5148 17724 5176
rect 17543 5120 17724 5148
rect 17543 5117 17555 5120
rect 17497 5111 17555 5117
rect 18064 5092 18092 5179
rect 18230 5176 18236 5228
rect 18288 5176 18294 5228
rect 18506 5176 18512 5228
rect 18564 5176 18570 5228
rect 18984 5225 19012 5256
rect 19628 5225 19656 5324
rect 20254 5312 20260 5364
rect 20312 5352 20318 5364
rect 20349 5355 20407 5361
rect 20349 5352 20361 5355
rect 20312 5324 20361 5352
rect 20312 5312 20318 5324
rect 20349 5321 20361 5324
rect 20395 5321 20407 5355
rect 20349 5315 20407 5321
rect 28258 5312 28264 5364
rect 28316 5312 28322 5364
rect 18693 5219 18751 5225
rect 18693 5185 18705 5219
rect 18739 5185 18751 5219
rect 18693 5179 18751 5185
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 19153 5219 19211 5225
rect 19153 5185 19165 5219
rect 19199 5185 19211 5219
rect 19153 5179 19211 5185
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5185 19671 5219
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 19613 5179 19671 5185
rect 20088 5188 20269 5216
rect 18414 5148 18420 5160
rect 18248 5120 18420 5148
rect 18248 5092 18276 5120
rect 18414 5108 18420 5120
rect 18472 5148 18478 5160
rect 18708 5148 18736 5179
rect 19168 5148 19196 5179
rect 18472 5120 19196 5148
rect 18472 5108 18478 5120
rect 17037 5083 17095 5089
rect 17037 5049 17049 5083
rect 17083 5080 17095 5083
rect 17402 5080 17408 5092
rect 17083 5052 17408 5080
rect 17083 5049 17095 5052
rect 17037 5043 17095 5049
rect 17402 5040 17408 5052
rect 17460 5040 17466 5092
rect 18046 5080 18052 5092
rect 17512 5052 18052 5080
rect 11164 4984 12664 5012
rect 16850 4972 16856 5024
rect 16908 4972 16914 5024
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 17512 5021 17540 5052
rect 18046 5040 18052 5052
rect 18104 5040 18110 5092
rect 18230 5040 18236 5092
rect 18288 5040 18294 5092
rect 19628 5080 19656 5179
rect 20088 5157 20116 5188
rect 20257 5185 20269 5188
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 28074 5176 28080 5228
rect 28132 5176 28138 5228
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5117 20131 5151
rect 20073 5111 20131 5117
rect 19628 5052 20760 5080
rect 20732 5024 20760 5052
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17184 4984 17509 5012
rect 17184 4972 17190 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 17862 4972 17868 5024
rect 17920 4972 17926 5024
rect 17954 4972 17960 5024
rect 18012 5012 18018 5024
rect 18877 5015 18935 5021
rect 18877 5012 18889 5015
rect 18012 4984 18889 5012
rect 18012 4972 18018 4984
rect 18877 4981 18889 4984
rect 18923 4981 18935 5015
rect 18877 4975 18935 4981
rect 18969 5015 19027 5021
rect 18969 4981 18981 5015
rect 19015 5012 19027 5015
rect 19058 5012 19064 5024
rect 19015 4984 19064 5012
rect 19015 4981 19027 4984
rect 18969 4975 19027 4981
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19705 5015 19763 5021
rect 19705 5012 19717 5015
rect 19576 4984 19717 5012
rect 19576 4972 19582 4984
rect 19705 4981 19717 4984
rect 19751 4981 19763 5015
rect 19705 4975 19763 4981
rect 20714 4972 20720 5024
rect 20772 4972 20778 5024
rect 1104 4922 29440 4944
rect 1104 4870 4491 4922
rect 4543 4870 4555 4922
rect 4607 4870 4619 4922
rect 4671 4870 4683 4922
rect 4735 4870 4747 4922
rect 4799 4870 11574 4922
rect 11626 4870 11638 4922
rect 11690 4870 11702 4922
rect 11754 4870 11766 4922
rect 11818 4870 11830 4922
rect 11882 4870 18657 4922
rect 18709 4870 18721 4922
rect 18773 4870 18785 4922
rect 18837 4870 18849 4922
rect 18901 4870 18913 4922
rect 18965 4870 25740 4922
rect 25792 4870 25804 4922
rect 25856 4870 25868 4922
rect 25920 4870 25932 4922
rect 25984 4870 25996 4922
rect 26048 4870 29440 4922
rect 1104 4848 29440 4870
rect 10226 4768 10232 4820
rect 10284 4768 10290 4820
rect 10686 4768 10692 4820
rect 10744 4768 10750 4820
rect 11054 4768 11060 4820
rect 11112 4768 11118 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11422 4808 11428 4820
rect 11379 4780 11428 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 16025 4811 16083 4817
rect 16025 4777 16037 4811
rect 16071 4808 16083 4811
rect 16390 4808 16396 4820
rect 16071 4780 16396 4808
rect 16071 4777 16083 4780
rect 16025 4771 16083 4777
rect 16390 4768 16396 4780
rect 16448 4768 16454 4820
rect 16482 4768 16488 4820
rect 16540 4808 16546 4820
rect 16942 4808 16948 4820
rect 16540 4780 16948 4808
rect 16540 4768 16546 4780
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17586 4768 17592 4820
rect 17644 4768 17650 4820
rect 17770 4768 17776 4820
rect 17828 4768 17834 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 17920 4780 18920 4808
rect 17920 4768 17926 4780
rect 8938 4632 8944 4684
rect 8996 4632 9002 4684
rect 9306 4632 9312 4684
rect 9364 4632 9370 4684
rect 10244 4522 10272 4768
rect 11072 4672 11100 4768
rect 16114 4700 16120 4752
rect 16172 4700 16178 4752
rect 16209 4743 16267 4749
rect 16209 4709 16221 4743
rect 16255 4740 16267 4743
rect 18785 4743 18843 4749
rect 18785 4740 18797 4743
rect 16255 4712 18797 4740
rect 16255 4709 16267 4712
rect 16209 4703 16267 4709
rect 18785 4709 18797 4712
rect 18831 4709 18843 4743
rect 18785 4703 18843 4709
rect 18892 4740 18920 4780
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 19981 4811 20039 4817
rect 19981 4808 19993 4811
rect 19852 4780 19993 4808
rect 19852 4768 19858 4780
rect 19981 4777 19993 4780
rect 20027 4777 20039 4811
rect 19981 4771 20039 4777
rect 20441 4811 20499 4817
rect 20441 4777 20453 4811
rect 20487 4808 20499 4811
rect 28074 4808 28080 4820
rect 20487 4780 28080 4808
rect 20487 4777 20499 4780
rect 20441 4771 20499 4777
rect 28074 4768 28080 4780
rect 28132 4768 28138 4820
rect 20070 4740 20076 4752
rect 18892 4712 20076 4740
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 11072 4644 11161 4672
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 11149 4635 11207 4641
rect 13004 4644 13369 4672
rect 13004 4616 13032 4644
rect 13357 4641 13369 4644
rect 13403 4641 13415 4675
rect 13357 4635 13415 4641
rect 16022 4632 16028 4684
rect 16080 4632 16086 4684
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11330 4604 11336 4616
rect 11103 4576 11336 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 12986 4564 12992 4616
rect 13044 4564 13050 4616
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 13096 4536 13124 4567
rect 13262 4564 13268 4616
rect 13320 4564 13326 4616
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16040 4604 16068 4632
rect 16132 4613 16160 4700
rect 17494 4632 17500 4684
rect 17552 4672 17558 4684
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 17552 4644 17693 4672
rect 17552 4632 17558 4644
rect 17681 4641 17693 4644
rect 17727 4641 17739 4675
rect 17681 4635 17739 4641
rect 17770 4632 17776 4684
rect 17828 4632 17834 4684
rect 17862 4632 17868 4684
rect 17920 4672 17926 4684
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 17920 4644 18153 4672
rect 17920 4632 17926 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 18230 4632 18236 4684
rect 18288 4632 18294 4684
rect 18892 4681 18920 4712
rect 20070 4700 20076 4712
rect 20128 4700 20134 4752
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4672 18475 4675
rect 18877 4675 18935 4681
rect 18463 4644 18828 4672
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 15979 4576 16068 4604
rect 16117 4607 16175 4613
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16117 4573 16129 4607
rect 16163 4573 16175 4607
rect 16117 4567 16175 4573
rect 16482 4564 16488 4616
rect 16540 4564 16546 4616
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4573 16635 4607
rect 16577 4567 16635 4573
rect 13998 4536 14004 4548
rect 13096 4508 14004 4536
rect 13998 4496 14004 4508
rect 14056 4496 14062 4548
rect 16206 4496 16212 4548
rect 16264 4496 16270 4548
rect 16592 4536 16620 4567
rect 17402 4564 17408 4616
rect 17460 4564 17466 4616
rect 17785 4604 17813 4632
rect 17957 4607 18015 4613
rect 17785 4594 17816 4604
rect 17957 4594 17969 4607
rect 17785 4576 17969 4594
rect 17788 4573 17969 4576
rect 18003 4573 18015 4607
rect 17788 4567 18015 4573
rect 17788 4566 18000 4567
rect 18598 4564 18604 4616
rect 18656 4564 18662 4616
rect 16666 4536 16672 4548
rect 16592 4508 16672 4536
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 18616 4536 18644 4564
rect 18248 4508 18644 4536
rect 18800 4536 18828 4644
rect 18877 4641 18889 4675
rect 18923 4641 18935 4675
rect 19334 4672 19340 4684
rect 18877 4635 18935 4641
rect 19168 4644 19340 4672
rect 19168 4536 19196 4644
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 19426 4632 19432 4684
rect 19484 4632 19490 4684
rect 19518 4632 19524 4684
rect 19576 4632 19582 4684
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4672 19671 4675
rect 19659 4644 20208 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 20180 4616 20208 4644
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 19705 4607 19763 4613
rect 19352 4566 19564 4594
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 19794 4604 19800 4616
rect 19751 4576 19800 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 18800 4508 19196 4536
rect 19260 4536 19288 4564
rect 19352 4536 19380 4566
rect 19260 4508 19380 4536
rect 19536 4536 19564 4566
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4573 19947 4607
rect 19889 4567 19947 4573
rect 19904 4536 19932 4567
rect 20162 4564 20168 4616
rect 20220 4564 20226 4616
rect 20438 4564 20444 4616
rect 20496 4604 20502 4616
rect 20533 4607 20591 4613
rect 20533 4604 20545 4607
rect 20496 4576 20545 4604
rect 20496 4564 20502 4576
rect 20533 4573 20545 4576
rect 20579 4573 20591 4607
rect 20533 4567 20591 4573
rect 20714 4564 20720 4616
rect 20772 4564 20778 4616
rect 20625 4539 20683 4545
rect 20625 4536 20637 4539
rect 19536 4508 20637 4536
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 12897 4471 12955 4477
rect 12897 4468 12909 4471
rect 6512 4440 12909 4468
rect 6512 4428 6518 4440
rect 12897 4437 12909 4440
rect 12943 4437 12955 4471
rect 12897 4431 12955 4437
rect 16393 4471 16451 4477
rect 16393 4437 16405 4471
rect 16439 4468 16451 4471
rect 16850 4468 16856 4480
rect 16439 4440 16856 4468
rect 16439 4437 16451 4440
rect 16393 4431 16451 4437
rect 16850 4428 16856 4440
rect 16908 4468 16914 4480
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16908 4440 16957 4468
rect 16908 4428 16914 4440
rect 16945 4437 16957 4440
rect 16991 4437 17003 4471
rect 16945 4431 17003 4437
rect 17126 4428 17132 4480
rect 17184 4428 17190 4480
rect 17218 4428 17224 4480
rect 17276 4428 17282 4480
rect 18046 4428 18052 4480
rect 18104 4468 18110 4480
rect 18248 4468 18276 4508
rect 20625 4505 20637 4508
rect 20671 4505 20683 4539
rect 20625 4499 20683 4505
rect 18104 4440 18276 4468
rect 18104 4428 18110 4440
rect 18322 4428 18328 4480
rect 18380 4468 18386 4480
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 18380 4440 19257 4468
rect 18380 4428 18386 4440
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19794 4468 19800 4480
rect 19484 4440 19800 4468
rect 19484 4428 19490 4440
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 1104 4378 29440 4400
rect 1104 4326 5151 4378
rect 5203 4326 5215 4378
rect 5267 4326 5279 4378
rect 5331 4326 5343 4378
rect 5395 4326 5407 4378
rect 5459 4326 12234 4378
rect 12286 4326 12298 4378
rect 12350 4326 12362 4378
rect 12414 4326 12426 4378
rect 12478 4326 12490 4378
rect 12542 4326 19317 4378
rect 19369 4326 19381 4378
rect 19433 4326 19445 4378
rect 19497 4326 19509 4378
rect 19561 4326 19573 4378
rect 19625 4326 26400 4378
rect 26452 4326 26464 4378
rect 26516 4326 26528 4378
rect 26580 4326 26592 4378
rect 26644 4326 26656 4378
rect 26708 4326 29440 4378
rect 1104 4304 29440 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2464 4236 2774 4264
rect 2464 4224 2470 4236
rect 2746 4196 2774 4236
rect 12618 4224 12624 4276
rect 12676 4264 12682 4276
rect 13173 4267 13231 4273
rect 13173 4264 13185 4267
rect 12676 4236 13185 4264
rect 12676 4224 12682 4236
rect 13173 4233 13185 4236
rect 13219 4233 13231 4267
rect 13173 4227 13231 4233
rect 13909 4267 13967 4273
rect 13909 4233 13921 4267
rect 13955 4233 13967 4267
rect 13909 4227 13967 4233
rect 14461 4267 14519 4273
rect 14461 4233 14473 4267
rect 14507 4264 14519 4267
rect 14826 4264 14832 4276
rect 14507 4236 14832 4264
rect 14507 4233 14519 4236
rect 14461 4227 14519 4233
rect 13924 4196 13952 4227
rect 14826 4224 14832 4236
rect 14884 4224 14890 4276
rect 16390 4264 16396 4276
rect 15764 4236 16396 4264
rect 2746 4168 13952 4196
rect 14292 4168 14596 4196
rect 2406 4088 2412 4140
rect 2464 4088 2470 4140
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13111 4131 13169 4137
rect 13111 4128 13123 4131
rect 13044 4100 13123 4128
rect 13044 4088 13050 4100
rect 13111 4097 13123 4100
rect 13157 4097 13169 4131
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 13111 4091 13169 4097
rect 13280 4100 13645 4128
rect 13280 4060 13308 4100
rect 13633 4097 13645 4100
rect 13679 4097 13691 4131
rect 13633 4091 13691 4097
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 14292 4128 14320 4168
rect 14568 4137 14596 4168
rect 13771 4100 14320 4128
rect 14369 4131 14427 4137
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 14369 4097 14381 4131
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 14642 4128 14648 4140
rect 14599 4100 14648 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 13096 4032 13308 4060
rect 3510 3952 3516 4004
rect 3568 3992 3574 4004
rect 12989 3995 13047 4001
rect 12989 3992 13001 3995
rect 3568 3964 13001 3992
rect 3568 3952 3574 3964
rect 12989 3961 13001 3964
rect 13035 3961 13047 3995
rect 12989 3955 13047 3961
rect 13096 3936 13124 4032
rect 13354 4020 13360 4072
rect 13412 4060 13418 4072
rect 13740 4060 13768 4091
rect 13412 4032 13768 4060
rect 13412 4020 13418 4032
rect 14090 4020 14096 4072
rect 14148 4020 14154 4072
rect 14384 4060 14412 4091
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 15764 4137 15792 4236
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 16908 4236 17632 4264
rect 16908 4224 16914 4236
rect 16316 4168 16804 4196
rect 16316 4137 16344 4168
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 15212 4060 15240 4088
rect 14384 4032 15240 4060
rect 15580 4060 15608 4091
rect 15580 4032 15976 4060
rect 2222 3884 2228 3936
rect 2280 3884 2286 3936
rect 13078 3884 13084 3936
rect 13136 3884 13142 3936
rect 13538 3884 13544 3936
rect 13596 3884 13602 3936
rect 13906 3884 13912 3936
rect 13964 3924 13970 3936
rect 14277 3927 14335 3933
rect 14277 3924 14289 3927
rect 13964 3896 14289 3924
rect 13964 3884 13970 3896
rect 14277 3893 14289 3896
rect 14323 3924 14335 3927
rect 14384 3924 14412 4032
rect 14458 3952 14464 4004
rect 14516 3992 14522 4004
rect 15841 3995 15899 4001
rect 15841 3992 15853 3995
rect 14516 3964 15853 3992
rect 14516 3952 14522 3964
rect 15841 3961 15853 3964
rect 15887 3961 15899 3995
rect 15841 3955 15899 3961
rect 14323 3896 14412 3924
rect 14323 3893 14335 3896
rect 14277 3887 14335 3893
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 15948 3924 15976 4032
rect 16040 3992 16068 4091
rect 16574 4088 16580 4140
rect 16632 4128 16638 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16632 4100 16681 4128
rect 16632 4088 16638 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16776 4128 16804 4168
rect 16942 4156 16948 4208
rect 17000 4196 17006 4208
rect 17000 4168 17356 4196
rect 17000 4156 17006 4168
rect 17126 4128 17132 4140
rect 16776 4100 17132 4128
rect 16669 4091 16727 4097
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17218 4088 17224 4140
rect 17276 4088 17282 4140
rect 17328 4137 17356 4168
rect 17604 4137 17632 4236
rect 19702 4224 19708 4276
rect 19760 4224 19766 4276
rect 19981 4267 20039 4273
rect 19981 4233 19993 4267
rect 20027 4264 20039 4267
rect 20438 4264 20444 4276
rect 20027 4236 20444 4264
rect 20027 4233 20039 4236
rect 19981 4227 20039 4233
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 17589 4131 17647 4137
rect 17589 4097 17601 4131
rect 17635 4097 17647 4131
rect 17589 4091 17647 4097
rect 18414 4088 18420 4140
rect 18472 4128 18478 4140
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 18472 4100 18797 4128
rect 18472 4088 18478 4100
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 19242 4088 19248 4140
rect 19300 4088 19306 4140
rect 19720 4137 19748 4224
rect 19794 4156 19800 4208
rect 19852 4156 19858 4208
rect 24029 4199 24087 4205
rect 24029 4165 24041 4199
rect 24075 4196 24087 4199
rect 24213 4199 24271 4205
rect 24075 4168 24164 4196
rect 24075 4165 24087 4168
rect 24029 4159 24087 4165
rect 19705 4131 19763 4137
rect 19705 4097 19717 4131
rect 19751 4097 19763 4131
rect 19705 4091 19763 4097
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4060 16267 4063
rect 17236 4060 17264 4088
rect 16255 4032 17264 4060
rect 17405 4063 17463 4069
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 17405 4029 17417 4063
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 17310 3992 17316 4004
rect 16040 3964 17316 3992
rect 17310 3952 17316 3964
rect 17368 3952 17374 4004
rect 17420 3992 17448 4023
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 17552 4032 19533 4060
rect 17552 4020 17558 4032
rect 19521 4029 19533 4032
rect 19567 4029 19579 4063
rect 19521 4023 19579 4029
rect 19812 4060 19840 4156
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 24136 4128 24164 4168
rect 24213 4165 24225 4199
rect 24259 4196 24271 4199
rect 24302 4196 24308 4208
rect 24259 4168 24308 4196
rect 24259 4165 24271 4168
rect 24213 4159 24271 4165
rect 24302 4156 24308 4168
rect 24360 4196 24366 4208
rect 24765 4199 24823 4205
rect 24765 4196 24777 4199
rect 24360 4168 24777 4196
rect 24360 4156 24366 4168
rect 24765 4165 24777 4168
rect 24811 4165 24823 4199
rect 24765 4159 24823 4165
rect 24486 4128 24492 4140
rect 24136 4100 24492 4128
rect 24486 4088 24492 4100
rect 24544 4128 24550 4140
rect 24581 4131 24639 4137
rect 24581 4128 24593 4131
rect 24544 4100 24593 4128
rect 24544 4088 24550 4100
rect 24581 4097 24593 4100
rect 24627 4097 24639 4131
rect 24581 4091 24639 4097
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19812 4032 19993 4060
rect 19812 3992 19840 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 17420 3964 19840 3992
rect 17420 3936 17448 3964
rect 19886 3952 19892 4004
rect 19944 3952 19950 4004
rect 16482 3924 16488 3936
rect 15948 3896 16488 3924
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 17402 3884 17408 3936
rect 17460 3884 17466 3936
rect 19797 3927 19855 3933
rect 19797 3893 19809 3927
rect 19843 3924 19855 3927
rect 19904 3924 19932 3952
rect 19843 3896 19932 3924
rect 19843 3893 19855 3896
rect 19797 3887 19855 3893
rect 20162 3884 20168 3936
rect 20220 3884 20226 3936
rect 24394 3884 24400 3936
rect 24452 3884 24458 3936
rect 24946 3884 24952 3936
rect 25004 3884 25010 3936
rect 1104 3834 29440 3856
rect 1104 3782 4491 3834
rect 4543 3782 4555 3834
rect 4607 3782 4619 3834
rect 4671 3782 4683 3834
rect 4735 3782 4747 3834
rect 4799 3782 11574 3834
rect 11626 3782 11638 3834
rect 11690 3782 11702 3834
rect 11754 3782 11766 3834
rect 11818 3782 11830 3834
rect 11882 3782 18657 3834
rect 18709 3782 18721 3834
rect 18773 3782 18785 3834
rect 18837 3782 18849 3834
rect 18901 3782 18913 3834
rect 18965 3782 25740 3834
rect 25792 3782 25804 3834
rect 25856 3782 25868 3834
rect 25920 3782 25932 3834
rect 25984 3782 25996 3834
rect 26048 3782 29440 3834
rect 1104 3760 29440 3782
rect 2222 3680 2228 3732
rect 2280 3680 2286 3732
rect 12618 3680 12624 3732
rect 12676 3680 12682 3732
rect 14553 3723 14611 3729
rect 13188 3692 13952 3720
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 2240 3516 2268 3680
rect 12894 3584 12900 3596
rect 2746 3556 12900 3584
rect 1535 3488 2268 3516
rect 2409 3519 2467 3525
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 2746 3516 2774 3556
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 2455 3488 2774 3516
rect 12529 3519 12587 3525
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 12989 3519 13047 3525
rect 12575 3488 12940 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 934 3340 940 3392
rect 992 3380 998 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 992 3352 1593 3380
rect 992 3340 998 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 2222 3340 2228 3392
rect 2280 3340 2286 3392
rect 12802 3340 12808 3392
rect 12860 3340 12866 3392
rect 12912 3380 12940 3488
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13188 3516 13216 3692
rect 13924 3664 13952 3692
rect 14553 3689 14565 3723
rect 14599 3720 14611 3723
rect 14642 3720 14648 3732
rect 14599 3692 14648 3720
rect 14599 3689 14611 3692
rect 14553 3683 14611 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 24394 3720 24400 3732
rect 15488 3692 18184 3720
rect 13906 3612 13912 3664
rect 13964 3612 13970 3664
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14737 3655 14795 3661
rect 14737 3652 14749 3655
rect 14056 3624 14749 3652
rect 14056 3612 14062 3624
rect 14737 3621 14749 3624
rect 14783 3621 14795 3655
rect 14737 3615 14795 3621
rect 15102 3612 15108 3664
rect 15160 3612 15166 3664
rect 15488 3661 15516 3692
rect 15473 3655 15531 3661
rect 15473 3621 15485 3655
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 15654 3612 15660 3664
rect 15712 3652 15718 3664
rect 15712 3624 17448 3652
rect 15712 3612 15718 3624
rect 13630 3544 13636 3596
rect 13688 3584 13694 3596
rect 14090 3584 14096 3596
rect 13688 3556 14096 3584
rect 13688 3544 13694 3556
rect 13035 3488 13216 3516
rect 13265 3519 13323 3525
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13265 3485 13277 3519
rect 13311 3516 13323 3519
rect 13354 3516 13360 3528
rect 13311 3488 13360 3516
rect 13311 3485 13323 3488
rect 13265 3479 13323 3485
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13449 3519 13507 3525
rect 13449 3485 13461 3519
rect 13495 3516 13507 3519
rect 13538 3516 13544 3528
rect 13495 3488 13544 3516
rect 13495 3485 13507 3488
rect 13449 3479 13507 3485
rect 13538 3476 13544 3488
rect 13596 3516 13602 3528
rect 13740 3525 13768 3556
rect 14090 3544 14096 3556
rect 14148 3584 14154 3596
rect 16393 3587 16451 3593
rect 14148 3556 15608 3584
rect 14148 3544 14154 3556
rect 13725 3519 13783 3525
rect 13596 3488 13682 3516
rect 13596 3476 13602 3488
rect 13654 3448 13682 3488
rect 13725 3485 13737 3519
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 13872 3488 14228 3516
rect 13872 3476 13878 3488
rect 13654 3420 13860 3448
rect 13722 3380 13728 3392
rect 12912 3352 13728 3380
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13832 3389 13860 3420
rect 13906 3408 13912 3460
rect 13964 3448 13970 3460
rect 14093 3451 14151 3457
rect 14093 3448 14105 3451
rect 13964 3420 14105 3448
rect 13964 3408 13970 3420
rect 14093 3417 14105 3420
rect 14139 3417 14151 3451
rect 14200 3448 14228 3488
rect 14458 3476 14464 3528
rect 14516 3476 14522 3528
rect 14568 3525 14596 3556
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 14826 3476 14832 3528
rect 14884 3476 14890 3528
rect 15286 3476 15292 3528
rect 15344 3516 15350 3528
rect 15580 3525 15608 3556
rect 16393 3553 16405 3587
rect 16439 3553 16451 3587
rect 16393 3547 16451 3553
rect 15381 3519 15439 3525
rect 15381 3516 15393 3519
rect 15344 3488 15393 3516
rect 15344 3476 15350 3488
rect 15381 3485 15393 3488
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3516 15623 3519
rect 16408 3516 16436 3547
rect 16574 3544 16580 3596
rect 16632 3544 16638 3596
rect 15611 3488 16436 3516
rect 16592 3516 16620 3544
rect 16776 3525 16804 3624
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16592 3488 16681 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 17310 3516 17316 3528
rect 17083 3488 17316 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 14844 3448 14872 3476
rect 14200 3420 14872 3448
rect 16868 3448 16896 3479
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17420 3516 17448 3624
rect 18046 3544 18052 3596
rect 18104 3544 18110 3596
rect 17770 3516 17776 3528
rect 17420 3488 17776 3516
rect 17770 3476 17776 3488
rect 17828 3516 17834 3528
rect 17828 3488 17908 3516
rect 17828 3476 17834 3488
rect 17880 3457 17908 3488
rect 17865 3451 17923 3457
rect 16868 3420 17632 3448
rect 14093 3411 14151 3417
rect 17604 3392 17632 3420
rect 17865 3417 17877 3451
rect 17911 3417 17923 3451
rect 18156 3448 18184 3692
rect 22066 3692 24400 3720
rect 18874 3612 18880 3664
rect 18932 3652 18938 3664
rect 22066 3652 22094 3692
rect 24394 3680 24400 3692
rect 24452 3680 24458 3732
rect 24946 3680 24952 3732
rect 25004 3680 25010 3732
rect 18932 3624 22094 3652
rect 18932 3612 18938 3624
rect 18969 3587 19027 3593
rect 18969 3553 18981 3587
rect 19015 3584 19027 3587
rect 20162 3584 20168 3596
rect 19015 3556 20168 3584
rect 19015 3553 19027 3556
rect 18969 3547 19027 3553
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 18506 3476 18512 3528
rect 18564 3516 18570 3528
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 18564 3488 18705 3516
rect 18564 3476 18570 3488
rect 18693 3485 18705 3488
rect 18739 3485 18751 3519
rect 24964 3516 24992 3680
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 24964 3488 25421 3516
rect 18693 3479 18751 3485
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 25409 3479 25467 3485
rect 22094 3448 22100 3460
rect 18156 3420 22100 3448
rect 17865 3411 17923 3417
rect 22094 3408 22100 3420
rect 22152 3408 22158 3460
rect 13817 3383 13875 3389
rect 13817 3349 13829 3383
rect 13863 3380 13875 3383
rect 14274 3380 14280 3392
rect 13863 3352 14280 3380
rect 13863 3349 13875 3352
rect 13817 3343 13875 3349
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 15286 3340 15292 3392
rect 15344 3340 15350 3392
rect 17494 3340 17500 3392
rect 17552 3340 17558 3392
rect 17586 3340 17592 3392
rect 17644 3340 17650 3392
rect 17957 3383 18015 3389
rect 17957 3349 17969 3383
rect 18003 3380 18015 3383
rect 18325 3383 18383 3389
rect 18325 3380 18337 3383
rect 18003 3352 18337 3380
rect 18003 3349 18015 3352
rect 17957 3343 18015 3349
rect 18325 3349 18337 3352
rect 18371 3349 18383 3383
rect 18325 3343 18383 3349
rect 18782 3340 18788 3392
rect 18840 3340 18846 3392
rect 25222 3340 25228 3392
rect 25280 3340 25286 3392
rect 1104 3290 29440 3312
rect 1104 3238 5151 3290
rect 5203 3238 5215 3290
rect 5267 3238 5279 3290
rect 5331 3238 5343 3290
rect 5395 3238 5407 3290
rect 5459 3238 12234 3290
rect 12286 3238 12298 3290
rect 12350 3238 12362 3290
rect 12414 3238 12426 3290
rect 12478 3238 12490 3290
rect 12542 3238 19317 3290
rect 19369 3238 19381 3290
rect 19433 3238 19445 3290
rect 19497 3238 19509 3290
rect 19561 3238 19573 3290
rect 19625 3238 26400 3290
rect 26452 3238 26464 3290
rect 26516 3238 26528 3290
rect 26580 3238 26592 3290
rect 26644 3238 26656 3290
rect 26708 3238 29440 3290
rect 1104 3216 29440 3238
rect 12986 3136 12992 3188
rect 13044 3136 13050 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 13136 3148 14565 3176
rect 13136 3136 13142 3148
rect 13372 3049 13400 3148
rect 14553 3145 14565 3148
rect 14599 3176 14611 3179
rect 15102 3176 15108 3188
rect 14599 3148 15108 3176
rect 14599 3145 14611 3148
rect 14553 3139 14611 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 17494 3136 17500 3188
rect 17552 3136 17558 3188
rect 17586 3136 17592 3188
rect 17644 3136 17650 3188
rect 17678 3136 17684 3188
rect 17736 3136 17742 3188
rect 17957 3179 18015 3185
rect 17957 3145 17969 3179
rect 18003 3176 18015 3179
rect 18782 3176 18788 3188
rect 18003 3148 18788 3176
rect 18003 3145 18015 3148
rect 17957 3139 18015 3145
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 14090 3108 14096 3120
rect 13740 3080 14096 3108
rect 13740 3052 13768 3080
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 15286 3108 15292 3120
rect 14200 3080 15292 3108
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3009 13139 3043
rect 13081 3003 13139 3009
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 13538 3040 13544 3052
rect 13495 3012 13544 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 12912 2904 12940 3003
rect 13096 2972 13124 3003
rect 13464 2972 13492 3003
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 13096 2944 13492 2972
rect 13648 2972 13676 3003
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 13814 3000 13820 3052
rect 13872 3000 13878 3052
rect 13906 3000 13912 3052
rect 13964 3000 13970 3052
rect 13998 3000 14004 3052
rect 14056 3000 14062 3052
rect 14200 3049 14228 3080
rect 15286 3068 15292 3080
rect 15344 3068 15350 3120
rect 16868 3080 17172 3108
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 14642 3040 14648 3052
rect 14599 3012 14648 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 13832 2972 13860 3000
rect 13648 2944 13860 2972
rect 13924 2972 13952 3000
rect 14384 2972 14412 3003
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 16868 3049 16896 3080
rect 17144 3052 17172 3080
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17126 3000 17132 3052
rect 17184 3000 17190 3052
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3040 17279 3043
rect 17512 3040 17540 3136
rect 17696 3108 17724 3136
rect 17696 3080 18276 3108
rect 17267 3012 17540 3040
rect 17681 3043 17739 3049
rect 17267 3009 17279 3012
rect 17221 3003 17279 3009
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 13924 2944 14412 2972
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2972 17003 2975
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 16991 2944 17417 2972
rect 16991 2941 17003 2944
rect 16945 2935 17003 2941
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 17494 2932 17500 2984
rect 17552 2932 17558 2984
rect 17696 2972 17724 3003
rect 17770 3000 17776 3052
rect 17828 3000 17834 3052
rect 18248 3049 18276 3080
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17880 3012 18061 3040
rect 17880 2972 17908 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18233 3043 18291 3049
rect 18233 3009 18245 3043
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 17696 2944 17908 2972
rect 17954 2932 17960 2984
rect 18012 2932 18018 2984
rect 18064 2972 18092 3003
rect 19058 3000 19064 3052
rect 19116 3000 19122 3052
rect 28813 3043 28871 3049
rect 28813 3040 28825 3043
rect 22066 3012 28825 3040
rect 19076 2972 19104 3000
rect 18064 2944 19104 2972
rect 13354 2904 13360 2916
rect 12912 2876 13360 2904
rect 13354 2864 13360 2876
rect 13412 2864 13418 2916
rect 13817 2907 13875 2913
rect 13817 2873 13829 2907
rect 13863 2904 13875 2907
rect 22066 2904 22094 3012
rect 28813 3009 28825 3012
rect 28859 3009 28871 3043
rect 28813 3003 28871 3009
rect 13863 2876 22094 2904
rect 13863 2873 13875 2876
rect 13817 2867 13875 2873
rect 13170 2796 13176 2848
rect 13228 2796 13234 2848
rect 17126 2796 17132 2848
rect 17184 2836 17190 2848
rect 18049 2839 18107 2845
rect 18049 2836 18061 2839
rect 17184 2808 18061 2836
rect 17184 2796 17190 2808
rect 18049 2805 18061 2808
rect 18095 2836 18107 2839
rect 19886 2836 19892 2848
rect 18095 2808 19892 2836
rect 18095 2805 18107 2808
rect 18049 2799 18107 2805
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 28994 2796 29000 2848
rect 29052 2796 29058 2848
rect 1104 2746 29440 2768
rect 1104 2694 4491 2746
rect 4543 2694 4555 2746
rect 4607 2694 4619 2746
rect 4671 2694 4683 2746
rect 4735 2694 4747 2746
rect 4799 2694 11574 2746
rect 11626 2694 11638 2746
rect 11690 2694 11702 2746
rect 11754 2694 11766 2746
rect 11818 2694 11830 2746
rect 11882 2694 18657 2746
rect 18709 2694 18721 2746
rect 18773 2694 18785 2746
rect 18837 2694 18849 2746
rect 18901 2694 18913 2746
rect 18965 2694 25740 2746
rect 25792 2694 25804 2746
rect 25856 2694 25868 2746
rect 25920 2694 25932 2746
rect 25984 2694 25996 2746
rect 26048 2694 29440 2746
rect 1104 2672 29440 2694
rect 12802 2632 12808 2644
rect 6886 2604 12808 2632
rect 1489 2431 1547 2437
rect 1489 2397 1501 2431
rect 1535 2428 1547 2431
rect 2222 2428 2228 2440
rect 1535 2400 2228 2428
rect 1535 2397 1547 2400
rect 1489 2391 1547 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 6886 2428 6914 2604
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 13320 2604 13461 2632
rect 13320 2592 13326 2604
rect 13449 2601 13461 2604
rect 13495 2601 13507 2635
rect 13449 2595 13507 2601
rect 3927 2400 6914 2428
rect 7300 2468 13216 2496
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 7300 2369 7328 2468
rect 13188 2440 13216 2468
rect 13464 2468 13860 2496
rect 13170 2388 13176 2440
rect 13228 2388 13234 2440
rect 13464 2437 13492 2468
rect 13832 2440 13860 2468
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2428 13691 2431
rect 13722 2428 13728 2440
rect 13679 2400 13728 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 15059 2400 22232 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 7285 2363 7343 2369
rect 7285 2329 7297 2363
rect 7331 2329 7343 2363
rect 7285 2323 7343 2329
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 17494 2360 17500 2372
rect 11655 2332 17500 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 17494 2320 17500 2332
rect 17552 2320 17558 2372
rect 19337 2363 19395 2369
rect 19337 2329 19349 2363
rect 19383 2360 19395 2363
rect 20070 2360 20076 2372
rect 19383 2332 20076 2360
rect 19383 2329 19395 2332
rect 19337 2323 19395 2329
rect 20070 2320 20076 2332
rect 20128 2320 20134 2372
rect 22094 2320 22100 2372
rect 22152 2320 22158 2372
rect 22204 2360 22232 2400
rect 25222 2388 25228 2440
rect 25280 2428 25286 2440
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25280 2400 25973 2428
rect 25280 2388 25286 2400
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 28534 2388 28540 2440
rect 28592 2428 28598 2440
rect 28721 2431 28779 2437
rect 28721 2428 28733 2431
rect 28592 2400 28733 2428
rect 28592 2388 28598 2400
rect 28721 2397 28733 2400
rect 28767 2397 28779 2431
rect 28721 2391 28779 2397
rect 27062 2360 27068 2372
rect 22204 2332 27068 2360
rect 27062 2320 27068 2332
rect 27120 2320 27126 2372
rect 29089 2363 29147 2369
rect 29089 2329 29101 2363
rect 29135 2360 29147 2363
rect 29638 2360 29644 2372
rect 29135 2332 29644 2360
rect 29135 2329 29147 2332
rect 29089 2323 29147 2329
rect 29638 2320 29644 2332
rect 29696 2320 29702 2372
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 72 2264 1593 2292
rect 72 2252 78 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3476 2264 4169 2292
rect 3476 2252 3482 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11204 2264 11713 2292
rect 11204 2252 11210 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 14918 2252 14924 2304
rect 14976 2292 14982 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 14976 2264 15301 2292
rect 14976 2252 14982 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 18874 2252 18880 2304
rect 18932 2292 18938 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 18932 2264 19441 2292
rect 18932 2252 18938 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 22060 2264 22201 2292
rect 22060 2252 22066 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 26237 2295 26295 2301
rect 26237 2292 26249 2295
rect 26200 2264 26249 2292
rect 26200 2252 26206 2264
rect 26237 2261 26249 2264
rect 26283 2261 26295 2295
rect 26237 2255 26295 2261
rect 1104 2202 29440 2224
rect 1104 2150 5151 2202
rect 5203 2150 5215 2202
rect 5267 2150 5279 2202
rect 5331 2150 5343 2202
rect 5395 2150 5407 2202
rect 5459 2150 12234 2202
rect 12286 2150 12298 2202
rect 12350 2150 12362 2202
rect 12414 2150 12426 2202
rect 12478 2150 12490 2202
rect 12542 2150 19317 2202
rect 19369 2150 19381 2202
rect 19433 2150 19445 2202
rect 19497 2150 19509 2202
rect 19561 2150 19573 2202
rect 19625 2150 26400 2202
rect 26452 2150 26464 2202
rect 26516 2150 26528 2202
rect 26580 2150 26592 2202
rect 26644 2150 26656 2202
rect 26708 2150 29440 2202
rect 1104 2128 29440 2150
<< via1 >>
rect 5151 30438 5203 30490
rect 5215 30438 5267 30490
rect 5279 30438 5331 30490
rect 5343 30438 5395 30490
rect 5407 30438 5459 30490
rect 12234 30438 12286 30490
rect 12298 30438 12350 30490
rect 12362 30438 12414 30490
rect 12426 30438 12478 30490
rect 12490 30438 12542 30490
rect 19317 30438 19369 30490
rect 19381 30438 19433 30490
rect 19445 30438 19497 30490
rect 19509 30438 19561 30490
rect 19573 30438 19625 30490
rect 26400 30438 26452 30490
rect 26464 30438 26516 30490
rect 26528 30438 26580 30490
rect 26592 30438 26644 30490
rect 26656 30438 26708 30490
rect 6736 30379 6788 30388
rect 6736 30345 6745 30379
rect 6745 30345 6779 30379
rect 6779 30345 6788 30379
rect 6736 30336 6788 30345
rect 9680 30268 9732 30320
rect 21272 30268 21324 30320
rect 25412 30268 25464 30320
rect 1584 30243 1636 30252
rect 1584 30209 1593 30243
rect 1593 30209 1627 30243
rect 1627 30209 1636 30243
rect 1584 30200 1636 30209
rect 3332 30200 3384 30252
rect 6092 30200 6144 30252
rect 9864 30243 9916 30252
rect 9864 30209 9873 30243
rect 9873 30209 9907 30243
rect 9907 30209 9916 30243
rect 9864 30200 9916 30209
rect 14188 30243 14240 30252
rect 14188 30209 14197 30243
rect 14197 30209 14231 30243
rect 14231 30209 14240 30243
rect 14188 30200 14240 30209
rect 17592 30243 17644 30252
rect 17592 30209 17601 30243
rect 17601 30209 17635 30243
rect 17635 30209 17644 30243
rect 17592 30200 17644 30209
rect 21916 30243 21968 30252
rect 21916 30209 21925 30243
rect 21925 30209 21959 30243
rect 21959 30209 21968 30243
rect 21916 30200 21968 30209
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 29000 30268 29052 30320
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 28908 30132 28960 30184
rect 13820 30064 13872 30116
rect 17408 30064 17460 30116
rect 1584 29996 1636 30048
rect 2872 30039 2924 30048
rect 2872 30005 2881 30039
rect 2881 30005 2915 30039
rect 2915 30005 2924 30039
rect 2872 29996 2924 30005
rect 28540 30039 28592 30048
rect 28540 30005 28549 30039
rect 28549 30005 28583 30039
rect 28583 30005 28592 30039
rect 28540 29996 28592 30005
rect 4491 29894 4543 29946
rect 4555 29894 4607 29946
rect 4619 29894 4671 29946
rect 4683 29894 4735 29946
rect 4747 29894 4799 29946
rect 11574 29894 11626 29946
rect 11638 29894 11690 29946
rect 11702 29894 11754 29946
rect 11766 29894 11818 29946
rect 11830 29894 11882 29946
rect 18657 29894 18709 29946
rect 18721 29894 18773 29946
rect 18785 29894 18837 29946
rect 18849 29894 18901 29946
rect 18913 29894 18965 29946
rect 25740 29894 25792 29946
rect 25804 29894 25856 29946
rect 25868 29894 25920 29946
rect 25932 29894 25984 29946
rect 25996 29894 26048 29946
rect 21916 29792 21968 29844
rect 14096 29656 14148 29708
rect 23940 29724 23992 29776
rect 4988 29588 5040 29640
rect 5172 29588 5224 29640
rect 5632 29631 5684 29640
rect 5632 29597 5641 29631
rect 5641 29597 5675 29631
rect 5675 29597 5684 29631
rect 5632 29588 5684 29597
rect 5724 29631 5776 29640
rect 5724 29597 5733 29631
rect 5733 29597 5767 29631
rect 5767 29597 5776 29631
rect 5724 29588 5776 29597
rect 6000 29520 6052 29572
rect 8484 29588 8536 29640
rect 9036 29631 9088 29640
rect 9036 29597 9045 29631
rect 9045 29597 9079 29631
rect 9079 29597 9088 29631
rect 9036 29588 9088 29597
rect 11336 29588 11388 29640
rect 13268 29588 13320 29640
rect 16212 29656 16264 29708
rect 19156 29656 19208 29708
rect 4896 29495 4948 29504
rect 4896 29461 4905 29495
rect 4905 29461 4939 29495
rect 4939 29461 4948 29495
rect 4896 29452 4948 29461
rect 5816 29452 5868 29504
rect 5908 29452 5960 29504
rect 7288 29452 7340 29504
rect 7564 29563 7616 29572
rect 7564 29529 7573 29563
rect 7573 29529 7607 29563
rect 7607 29529 7616 29563
rect 7564 29520 7616 29529
rect 14280 29520 14332 29572
rect 16488 29520 16540 29572
rect 20812 29631 20864 29640
rect 20812 29597 20821 29631
rect 20821 29597 20855 29631
rect 20855 29597 20864 29631
rect 20812 29588 20864 29597
rect 25228 29588 25280 29640
rect 7472 29452 7524 29504
rect 7748 29495 7800 29504
rect 7748 29461 7757 29495
rect 7757 29461 7791 29495
rect 7791 29461 7800 29495
rect 7748 29452 7800 29461
rect 11244 29452 11296 29504
rect 17132 29452 17184 29504
rect 17316 29495 17368 29504
rect 17316 29461 17325 29495
rect 17325 29461 17359 29495
rect 17359 29461 17368 29495
rect 17316 29452 17368 29461
rect 20444 29452 20496 29504
rect 5151 29350 5203 29402
rect 5215 29350 5267 29402
rect 5279 29350 5331 29402
rect 5343 29350 5395 29402
rect 5407 29350 5459 29402
rect 12234 29350 12286 29402
rect 12298 29350 12350 29402
rect 12362 29350 12414 29402
rect 12426 29350 12478 29402
rect 12490 29350 12542 29402
rect 19317 29350 19369 29402
rect 19381 29350 19433 29402
rect 19445 29350 19497 29402
rect 19509 29350 19561 29402
rect 19573 29350 19625 29402
rect 26400 29350 26452 29402
rect 26464 29350 26516 29402
rect 26528 29350 26580 29402
rect 26592 29350 26644 29402
rect 26656 29350 26708 29402
rect 1584 29180 1636 29232
rect 3056 29180 3108 29232
rect 3240 29180 3292 29232
rect 5908 29248 5960 29300
rect 7104 29180 7156 29232
rect 7472 29248 7524 29300
rect 7288 29180 7340 29232
rect 3148 29019 3200 29028
rect 3148 28985 3157 29019
rect 3157 28985 3191 29019
rect 3191 28985 3200 29019
rect 3148 28976 3200 28985
rect 3516 29087 3568 29096
rect 3516 29053 3525 29087
rect 3525 29053 3559 29087
rect 3559 29053 3568 29087
rect 3516 29044 3568 29053
rect 5632 29044 5684 29096
rect 6184 29044 6236 29096
rect 5172 28976 5224 29028
rect 4160 28908 4212 28960
rect 4988 28951 5040 28960
rect 4988 28917 4997 28951
rect 4997 28917 5031 28951
rect 5031 28917 5040 28951
rect 4988 28908 5040 28917
rect 7656 29044 7708 29096
rect 11244 29248 11296 29300
rect 12624 29248 12676 29300
rect 13268 29291 13320 29300
rect 13268 29257 13277 29291
rect 13277 29257 13311 29291
rect 13311 29257 13320 29291
rect 13268 29248 13320 29257
rect 16488 29291 16540 29300
rect 16488 29257 16497 29291
rect 16497 29257 16531 29291
rect 16531 29257 16540 29291
rect 16488 29248 16540 29257
rect 9772 29044 9824 29096
rect 11244 29044 11296 29096
rect 12256 29180 12308 29232
rect 14280 29180 14332 29232
rect 16212 29155 16264 29164
rect 16212 29121 16221 29155
rect 16221 29121 16255 29155
rect 16255 29121 16264 29155
rect 16212 29112 16264 29121
rect 16672 29180 16724 29232
rect 17316 29248 17368 29300
rect 19156 29291 19208 29300
rect 19156 29257 19165 29291
rect 19165 29257 19199 29291
rect 19199 29257 19208 29291
rect 19156 29248 19208 29257
rect 28540 29248 28592 29300
rect 20444 29180 20496 29232
rect 18236 29112 18288 29164
rect 13452 29087 13504 29096
rect 13452 29053 13461 29087
rect 13461 29053 13495 29087
rect 13495 29053 13504 29087
rect 13452 29044 13504 29053
rect 13728 29087 13780 29096
rect 13728 29053 13737 29087
rect 13737 29053 13771 29087
rect 13771 29053 13780 29087
rect 13728 29044 13780 29053
rect 7840 28908 7892 28960
rect 8760 28951 8812 28960
rect 8760 28917 8769 28951
rect 8769 28917 8803 28951
rect 8803 28917 8812 28951
rect 8760 28908 8812 28917
rect 11152 28951 11204 28960
rect 11152 28917 11161 28951
rect 11161 28917 11195 28951
rect 11195 28917 11204 28951
rect 11152 28908 11204 28917
rect 16580 29044 16632 29096
rect 18420 29044 18472 29096
rect 21180 29112 21232 29164
rect 22836 29112 22888 29164
rect 22100 29044 22152 29096
rect 22192 29044 22244 29096
rect 23388 29087 23440 29096
rect 23388 29053 23397 29087
rect 23397 29053 23431 29087
rect 23431 29053 23440 29087
rect 23388 29044 23440 29053
rect 24492 29044 24544 29096
rect 15476 28908 15528 28960
rect 15936 28951 15988 28960
rect 15936 28917 15945 28951
rect 15945 28917 15979 28951
rect 15979 28917 15988 28951
rect 15936 28908 15988 28917
rect 18328 28908 18380 28960
rect 19892 28908 19944 28960
rect 21272 28908 21324 28960
rect 21364 28908 21416 28960
rect 21916 28976 21968 29028
rect 21732 28908 21784 28960
rect 22376 28976 22428 29028
rect 23020 28951 23072 28960
rect 23020 28917 23029 28951
rect 23029 28917 23063 28951
rect 23063 28917 23072 28951
rect 23020 28908 23072 28917
rect 23112 28951 23164 28960
rect 23112 28917 23121 28951
rect 23121 28917 23155 28951
rect 23155 28917 23164 28951
rect 23112 28908 23164 28917
rect 4491 28806 4543 28858
rect 4555 28806 4607 28858
rect 4619 28806 4671 28858
rect 4683 28806 4735 28858
rect 4747 28806 4799 28858
rect 11574 28806 11626 28858
rect 11638 28806 11690 28858
rect 11702 28806 11754 28858
rect 11766 28806 11818 28858
rect 11830 28806 11882 28858
rect 18657 28806 18709 28858
rect 18721 28806 18773 28858
rect 18785 28806 18837 28858
rect 18849 28806 18901 28858
rect 18913 28806 18965 28858
rect 25740 28806 25792 28858
rect 25804 28806 25856 28858
rect 25868 28806 25920 28858
rect 25932 28806 25984 28858
rect 25996 28806 26048 28858
rect 5172 28704 5224 28756
rect 5724 28704 5776 28756
rect 6460 28704 6512 28756
rect 7104 28704 7156 28756
rect 7748 28704 7800 28756
rect 3608 28407 3660 28416
rect 3608 28373 3617 28407
rect 3617 28373 3651 28407
rect 3651 28373 3660 28407
rect 3608 28364 3660 28373
rect 4252 28568 4304 28620
rect 6276 28636 6328 28688
rect 9772 28747 9824 28756
rect 9772 28713 9781 28747
rect 9781 28713 9815 28747
rect 9815 28713 9824 28747
rect 9772 28704 9824 28713
rect 12624 28747 12676 28756
rect 12624 28713 12633 28747
rect 12633 28713 12667 28747
rect 12667 28713 12676 28747
rect 12624 28704 12676 28713
rect 12900 28704 12952 28756
rect 13728 28704 13780 28756
rect 16212 28704 16264 28756
rect 16672 28747 16724 28756
rect 16672 28713 16681 28747
rect 16681 28713 16715 28747
rect 16715 28713 16724 28747
rect 16672 28704 16724 28713
rect 5080 28568 5132 28620
rect 4160 28500 4212 28552
rect 5908 28500 5960 28552
rect 6460 28543 6512 28552
rect 6460 28509 6469 28543
rect 6469 28509 6503 28543
rect 6503 28509 6512 28543
rect 6460 28500 6512 28509
rect 8760 28568 8812 28620
rect 9404 28568 9456 28620
rect 11152 28568 11204 28620
rect 11244 28568 11296 28620
rect 7012 28500 7064 28552
rect 4344 28364 4396 28416
rect 4896 28432 4948 28484
rect 6184 28475 6236 28484
rect 6184 28441 6193 28475
rect 6193 28441 6227 28475
rect 6227 28441 6236 28475
rect 6184 28432 6236 28441
rect 6828 28432 6880 28484
rect 4988 28364 5040 28416
rect 6368 28407 6420 28416
rect 6368 28373 6377 28407
rect 6377 28373 6411 28407
rect 6411 28373 6420 28407
rect 6368 28364 6420 28373
rect 7012 28407 7064 28416
rect 7012 28373 7021 28407
rect 7021 28373 7055 28407
rect 7055 28373 7064 28407
rect 7012 28364 7064 28373
rect 7196 28475 7248 28484
rect 7196 28441 7205 28475
rect 7205 28441 7239 28475
rect 7239 28441 7248 28475
rect 7196 28432 7248 28441
rect 7564 28432 7616 28484
rect 7656 28475 7708 28484
rect 7656 28441 7665 28475
rect 7665 28441 7699 28475
rect 7699 28441 7708 28475
rect 7656 28432 7708 28441
rect 7748 28432 7800 28484
rect 8760 28475 8812 28484
rect 8760 28441 8769 28475
rect 8769 28441 8803 28475
rect 8803 28441 8812 28475
rect 8760 28432 8812 28441
rect 9956 28475 10008 28484
rect 9956 28441 9965 28475
rect 9965 28441 9999 28475
rect 9999 28441 10008 28475
rect 9956 28432 10008 28441
rect 12164 28500 12216 28552
rect 13636 28611 13688 28620
rect 13636 28577 13645 28611
rect 13645 28577 13679 28611
rect 13679 28577 13688 28611
rect 13636 28568 13688 28577
rect 15936 28568 15988 28620
rect 12072 28432 12124 28484
rect 13544 28500 13596 28552
rect 14004 28500 14056 28552
rect 14464 28500 14516 28552
rect 13636 28432 13688 28484
rect 15476 28543 15528 28552
rect 15476 28509 15485 28543
rect 15485 28509 15519 28543
rect 15519 28509 15528 28543
rect 15476 28500 15528 28509
rect 17132 28568 17184 28620
rect 17776 28568 17828 28620
rect 18420 28636 18472 28688
rect 20812 28704 20864 28756
rect 21732 28747 21784 28756
rect 21732 28713 21741 28747
rect 21741 28713 21775 28747
rect 21775 28713 21784 28747
rect 21732 28704 21784 28713
rect 22008 28747 22060 28756
rect 22008 28713 22017 28747
rect 22017 28713 22051 28747
rect 22051 28713 22060 28747
rect 22008 28704 22060 28713
rect 22100 28704 22152 28756
rect 18236 28568 18288 28620
rect 16488 28543 16540 28552
rect 16488 28509 16497 28543
rect 16497 28509 16531 28543
rect 16531 28509 16540 28543
rect 16488 28500 16540 28509
rect 16580 28500 16632 28552
rect 21272 28568 21324 28620
rect 16304 28475 16356 28484
rect 8576 28364 8628 28416
rect 10324 28364 10376 28416
rect 10784 28364 10836 28416
rect 11704 28364 11756 28416
rect 16304 28441 16313 28475
rect 16313 28441 16347 28475
rect 16347 28441 16356 28475
rect 16304 28432 16356 28441
rect 19340 28543 19392 28552
rect 19340 28509 19349 28543
rect 19349 28509 19383 28543
rect 19383 28509 19392 28543
rect 19340 28500 19392 28509
rect 19800 28500 19852 28552
rect 20812 28543 20864 28552
rect 20812 28509 20821 28543
rect 20821 28509 20855 28543
rect 20855 28509 20864 28543
rect 20812 28500 20864 28509
rect 21364 28543 21416 28552
rect 13912 28407 13964 28416
rect 13912 28373 13921 28407
rect 13921 28373 13955 28407
rect 13955 28373 13964 28407
rect 13912 28364 13964 28373
rect 14740 28407 14792 28416
rect 14740 28373 14749 28407
rect 14749 28373 14783 28407
rect 14783 28373 14792 28407
rect 14740 28364 14792 28373
rect 15292 28364 15344 28416
rect 18052 28364 18104 28416
rect 19708 28364 19760 28416
rect 20260 28364 20312 28416
rect 21364 28509 21373 28543
rect 21373 28509 21407 28543
rect 21407 28509 21416 28543
rect 21364 28500 21416 28509
rect 21640 28500 21692 28552
rect 21916 28500 21968 28552
rect 22376 28543 22428 28552
rect 22376 28509 22385 28543
rect 22385 28509 22419 28543
rect 22419 28509 22428 28543
rect 22376 28500 22428 28509
rect 23112 28568 23164 28620
rect 24216 28679 24268 28688
rect 24216 28645 24225 28679
rect 24225 28645 24259 28679
rect 24259 28645 24268 28679
rect 24216 28636 24268 28645
rect 22008 28432 22060 28484
rect 22192 28432 22244 28484
rect 24308 28500 24360 28552
rect 21732 28364 21784 28416
rect 22744 28432 22796 28484
rect 22928 28364 22980 28416
rect 24216 28364 24268 28416
rect 24400 28364 24452 28416
rect 5151 28262 5203 28314
rect 5215 28262 5267 28314
rect 5279 28262 5331 28314
rect 5343 28262 5395 28314
rect 5407 28262 5459 28314
rect 12234 28262 12286 28314
rect 12298 28262 12350 28314
rect 12362 28262 12414 28314
rect 12426 28262 12478 28314
rect 12490 28262 12542 28314
rect 19317 28262 19369 28314
rect 19381 28262 19433 28314
rect 19445 28262 19497 28314
rect 19509 28262 19561 28314
rect 19573 28262 19625 28314
rect 26400 28262 26452 28314
rect 26464 28262 26516 28314
rect 26528 28262 26580 28314
rect 26592 28262 26644 28314
rect 26656 28262 26708 28314
rect 3516 28160 3568 28212
rect 3608 28160 3660 28212
rect 6000 28203 6052 28212
rect 6000 28169 6009 28203
rect 6009 28169 6043 28203
rect 6043 28169 6052 28203
rect 6000 28160 6052 28169
rect 6184 28160 6236 28212
rect 7564 28160 7616 28212
rect 8576 28160 8628 28212
rect 3608 28067 3660 28076
rect 3608 28033 3617 28067
rect 3617 28033 3651 28067
rect 3651 28033 3660 28067
rect 3608 28024 3660 28033
rect 5632 28024 5684 28076
rect 5908 28024 5960 28076
rect 6276 27956 6328 28008
rect 5816 27931 5868 27940
rect 5816 27897 5825 27931
rect 5825 27897 5859 27931
rect 5859 27897 5868 27931
rect 5816 27888 5868 27897
rect 6460 28024 6512 28076
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 7012 28024 7064 28076
rect 7472 28092 7524 28144
rect 7196 28024 7248 28076
rect 7564 28024 7616 28076
rect 7840 28092 7892 28144
rect 9036 28024 9088 28076
rect 9404 28203 9456 28212
rect 9404 28169 9413 28203
rect 9413 28169 9447 28203
rect 9447 28169 9456 28203
rect 9404 28160 9456 28169
rect 9956 28160 10008 28212
rect 9312 28024 9364 28076
rect 12900 28160 12952 28212
rect 15292 28160 15344 28212
rect 16304 28160 16356 28212
rect 11336 28092 11388 28144
rect 11704 28135 11756 28144
rect 11704 28101 11713 28135
rect 11713 28101 11747 28135
rect 11747 28101 11756 28135
rect 11704 28092 11756 28101
rect 9772 27956 9824 28008
rect 10324 27999 10376 28008
rect 10324 27965 10333 27999
rect 10333 27965 10367 27999
rect 10367 27965 10376 27999
rect 10324 27956 10376 27965
rect 11428 28024 11480 28076
rect 13084 28092 13136 28144
rect 12256 28024 12308 28076
rect 12716 28024 12768 28076
rect 14280 28092 14332 28144
rect 13452 28067 13504 28076
rect 13452 28033 13461 28067
rect 13461 28033 13495 28067
rect 13495 28033 13504 28067
rect 13452 28024 13504 28033
rect 17776 28160 17828 28212
rect 17868 28160 17920 28212
rect 22100 28160 22152 28212
rect 22744 28160 22796 28212
rect 23020 28160 23072 28212
rect 23388 28160 23440 28212
rect 16488 28024 16540 28076
rect 7196 27888 7248 27940
rect 11428 27888 11480 27940
rect 15292 27999 15344 28008
rect 15292 27965 15301 27999
rect 15301 27965 15335 27999
rect 15335 27965 15344 27999
rect 15292 27956 15344 27965
rect 4160 27820 4212 27872
rect 6368 27820 6420 27872
rect 6552 27820 6604 27872
rect 11060 27820 11112 27872
rect 11244 27820 11296 27872
rect 12072 27863 12124 27872
rect 12072 27829 12081 27863
rect 12081 27829 12115 27863
rect 12115 27829 12124 27863
rect 12072 27820 12124 27829
rect 17684 28024 17736 28076
rect 17776 28067 17828 28076
rect 17776 28033 17785 28067
rect 17785 28033 17819 28067
rect 17819 28033 17828 28067
rect 17776 28024 17828 28033
rect 18144 28024 18196 28076
rect 18052 27956 18104 28008
rect 18328 27999 18380 28008
rect 18328 27965 18337 27999
rect 18337 27965 18371 27999
rect 18371 27965 18380 27999
rect 18328 27956 18380 27965
rect 18420 27999 18472 28008
rect 18420 27965 18429 27999
rect 18429 27965 18463 27999
rect 18463 27965 18472 27999
rect 18420 27956 18472 27965
rect 14464 27820 14516 27872
rect 17132 27820 17184 27872
rect 17960 27863 18012 27872
rect 17960 27829 17969 27863
rect 17969 27829 18003 27863
rect 18003 27829 18012 27863
rect 17960 27820 18012 27829
rect 18052 27863 18104 27872
rect 18052 27829 18061 27863
rect 18061 27829 18095 27863
rect 18095 27829 18104 27863
rect 18052 27820 18104 27829
rect 19340 27956 19392 28008
rect 20720 28024 20772 28076
rect 21180 28024 21232 28076
rect 22284 28024 22336 28076
rect 22928 28067 22980 28076
rect 22928 28033 22937 28067
rect 22937 28033 22971 28067
rect 22971 28033 22980 28067
rect 22928 28024 22980 28033
rect 24308 28024 24360 28076
rect 21640 27956 21692 28008
rect 21916 27956 21968 28008
rect 20260 27888 20312 27940
rect 22652 27931 22704 27940
rect 22652 27897 22661 27931
rect 22661 27897 22695 27931
rect 22695 27897 22704 27931
rect 22652 27888 22704 27897
rect 19892 27820 19944 27872
rect 22468 27863 22520 27872
rect 22468 27829 22477 27863
rect 22477 27829 22511 27863
rect 22511 27829 22520 27863
rect 22468 27820 22520 27829
rect 22560 27863 22612 27872
rect 22560 27829 22569 27863
rect 22569 27829 22603 27863
rect 22603 27829 22612 27863
rect 22560 27820 22612 27829
rect 4491 27718 4543 27770
rect 4555 27718 4607 27770
rect 4619 27718 4671 27770
rect 4683 27718 4735 27770
rect 4747 27718 4799 27770
rect 11574 27718 11626 27770
rect 11638 27718 11690 27770
rect 11702 27718 11754 27770
rect 11766 27718 11818 27770
rect 11830 27718 11882 27770
rect 18657 27718 18709 27770
rect 18721 27718 18773 27770
rect 18785 27718 18837 27770
rect 18849 27718 18901 27770
rect 18913 27718 18965 27770
rect 25740 27718 25792 27770
rect 25804 27718 25856 27770
rect 25868 27718 25920 27770
rect 25932 27718 25984 27770
rect 25996 27718 26048 27770
rect 3608 27616 3660 27668
rect 3148 27480 3200 27532
rect 4252 27523 4304 27532
rect 4252 27489 4261 27523
rect 4261 27489 4295 27523
rect 4295 27489 4304 27523
rect 4252 27480 4304 27489
rect 4344 27412 4396 27464
rect 4988 27616 5040 27668
rect 6368 27616 6420 27668
rect 11060 27616 11112 27668
rect 11336 27616 11388 27668
rect 11888 27616 11940 27668
rect 12072 27616 12124 27668
rect 14004 27616 14056 27668
rect 14464 27616 14516 27668
rect 18144 27616 18196 27668
rect 19340 27616 19392 27668
rect 22560 27616 22612 27668
rect 7380 27548 7432 27600
rect 11152 27548 11204 27600
rect 9312 27523 9364 27532
rect 9312 27489 9321 27523
rect 9321 27489 9355 27523
rect 9355 27489 9364 27523
rect 9312 27480 9364 27489
rect 1492 27387 1544 27396
rect 1492 27353 1501 27387
rect 1501 27353 1535 27387
rect 1535 27353 1544 27387
rect 1492 27344 1544 27353
rect 5080 27344 5132 27396
rect 940 27276 992 27328
rect 3056 27276 3108 27328
rect 7932 27387 7984 27396
rect 7932 27353 7941 27387
rect 7941 27353 7975 27387
rect 7975 27353 7984 27387
rect 7932 27344 7984 27353
rect 9036 27344 9088 27396
rect 9772 27412 9824 27464
rect 9956 27412 10008 27464
rect 11428 27412 11480 27464
rect 11888 27412 11940 27464
rect 12256 27412 12308 27464
rect 22652 27548 22704 27600
rect 12716 27523 12768 27532
rect 12716 27489 12725 27523
rect 12725 27489 12759 27523
rect 12759 27489 12768 27523
rect 12716 27480 12768 27489
rect 13084 27480 13136 27532
rect 14004 27480 14056 27532
rect 15476 27480 15528 27532
rect 17132 27480 17184 27532
rect 19432 27480 19484 27532
rect 12992 27344 13044 27396
rect 8576 27319 8628 27328
rect 8576 27285 8585 27319
rect 8585 27285 8619 27319
rect 8619 27285 8628 27319
rect 8576 27276 8628 27285
rect 8944 27319 8996 27328
rect 8944 27285 8953 27319
rect 8953 27285 8987 27319
rect 8987 27285 8996 27319
rect 8944 27276 8996 27285
rect 11888 27276 11940 27328
rect 11980 27276 12032 27328
rect 12256 27276 12308 27328
rect 14004 27276 14056 27328
rect 14556 27276 14608 27328
rect 16396 27455 16448 27464
rect 16396 27421 16405 27455
rect 16405 27421 16439 27455
rect 16439 27421 16448 27455
rect 16396 27412 16448 27421
rect 16488 27455 16540 27464
rect 16488 27421 16497 27455
rect 16497 27421 16531 27455
rect 16531 27421 16540 27455
rect 16488 27412 16540 27421
rect 17776 27412 17828 27464
rect 18236 27412 18288 27464
rect 19800 27480 19852 27532
rect 19892 27523 19944 27532
rect 19892 27489 19901 27523
rect 19901 27489 19935 27523
rect 19935 27489 19944 27523
rect 19892 27480 19944 27489
rect 20720 27480 20772 27532
rect 19708 27412 19760 27464
rect 22100 27480 22152 27532
rect 22836 27548 22888 27600
rect 22008 27455 22060 27464
rect 22008 27421 22017 27455
rect 22017 27421 22051 27455
rect 22051 27421 22060 27455
rect 22008 27412 22060 27421
rect 22284 27412 22336 27464
rect 24400 27412 24452 27464
rect 20260 27344 20312 27396
rect 21180 27344 21232 27396
rect 22468 27344 22520 27396
rect 20996 27276 21048 27328
rect 21640 27319 21692 27328
rect 21640 27285 21649 27319
rect 21649 27285 21683 27319
rect 21683 27285 21692 27319
rect 21640 27276 21692 27285
rect 22192 27276 22244 27328
rect 5151 27174 5203 27226
rect 5215 27174 5267 27226
rect 5279 27174 5331 27226
rect 5343 27174 5395 27226
rect 5407 27174 5459 27226
rect 12234 27174 12286 27226
rect 12298 27174 12350 27226
rect 12362 27174 12414 27226
rect 12426 27174 12478 27226
rect 12490 27174 12542 27226
rect 19317 27174 19369 27226
rect 19381 27174 19433 27226
rect 19445 27174 19497 27226
rect 19509 27174 19561 27226
rect 19573 27174 19625 27226
rect 26400 27174 26452 27226
rect 26464 27174 26516 27226
rect 26528 27174 26580 27226
rect 26592 27174 26644 27226
rect 26656 27174 26708 27226
rect 8944 27072 8996 27124
rect 9036 27072 9088 27124
rect 9772 27072 9824 27124
rect 13636 27072 13688 27124
rect 14556 27115 14608 27124
rect 14556 27081 14565 27115
rect 14565 27081 14599 27115
rect 14599 27081 14608 27115
rect 14556 27072 14608 27081
rect 16396 27072 16448 27124
rect 19800 27072 19852 27124
rect 20904 27072 20956 27124
rect 22284 27072 22336 27124
rect 11336 27004 11388 27056
rect 12072 27004 12124 27056
rect 12900 27004 12952 27056
rect 14740 27004 14792 27056
rect 17132 27047 17184 27056
rect 17132 27013 17141 27047
rect 17141 27013 17175 27047
rect 17175 27013 17184 27047
rect 17132 27004 17184 27013
rect 9588 26936 9640 26988
rect 7840 26868 7892 26920
rect 8576 26868 8628 26920
rect 11888 26979 11940 26988
rect 11888 26945 11897 26979
rect 11897 26945 11931 26979
rect 11931 26945 11940 26979
rect 11888 26936 11940 26945
rect 12256 26936 12308 26988
rect 13912 26936 13964 26988
rect 14280 26936 14332 26988
rect 20720 27004 20772 27056
rect 22008 27004 22060 27056
rect 11980 26800 12032 26852
rect 12808 26868 12860 26920
rect 28264 26936 28316 26988
rect 15292 26868 15344 26920
rect 13912 26800 13964 26852
rect 14004 26800 14056 26852
rect 18052 26800 18104 26852
rect 11244 26732 11296 26784
rect 12808 26775 12860 26784
rect 12808 26741 12838 26775
rect 12838 26741 12860 26775
rect 12808 26732 12860 26741
rect 12900 26732 12952 26784
rect 20996 26775 21048 26784
rect 20996 26741 21005 26775
rect 21005 26741 21039 26775
rect 21039 26741 21048 26775
rect 20996 26732 21048 26741
rect 29000 26775 29052 26784
rect 29000 26741 29009 26775
rect 29009 26741 29043 26775
rect 29043 26741 29052 26775
rect 29000 26732 29052 26741
rect 4491 26630 4543 26682
rect 4555 26630 4607 26682
rect 4619 26630 4671 26682
rect 4683 26630 4735 26682
rect 4747 26630 4799 26682
rect 11574 26630 11626 26682
rect 11638 26630 11690 26682
rect 11702 26630 11754 26682
rect 11766 26630 11818 26682
rect 11830 26630 11882 26682
rect 18657 26630 18709 26682
rect 18721 26630 18773 26682
rect 18785 26630 18837 26682
rect 18849 26630 18901 26682
rect 18913 26630 18965 26682
rect 25740 26630 25792 26682
rect 25804 26630 25856 26682
rect 25868 26630 25920 26682
rect 25932 26630 25984 26682
rect 25996 26630 26048 26682
rect 1492 26528 1544 26580
rect 11244 26528 11296 26580
rect 12164 26528 12216 26580
rect 2412 26367 2464 26376
rect 2412 26333 2421 26367
rect 2421 26333 2455 26367
rect 2455 26333 2464 26367
rect 2412 26324 2464 26333
rect 10784 26435 10836 26444
rect 10784 26401 10793 26435
rect 10793 26401 10827 26435
rect 10827 26401 10836 26435
rect 10784 26392 10836 26401
rect 11428 26392 11480 26444
rect 12256 26392 12308 26444
rect 6460 26324 6512 26376
rect 9588 26324 9640 26376
rect 17960 26324 18012 26376
rect 7012 26256 7064 26308
rect 11336 26256 11388 26308
rect 5816 26231 5868 26240
rect 5816 26197 5825 26231
rect 5825 26197 5859 26231
rect 5859 26197 5868 26231
rect 5816 26188 5868 26197
rect 19800 26256 19852 26308
rect 19984 26256 20036 26308
rect 5151 26086 5203 26138
rect 5215 26086 5267 26138
rect 5279 26086 5331 26138
rect 5343 26086 5395 26138
rect 5407 26086 5459 26138
rect 12234 26086 12286 26138
rect 12298 26086 12350 26138
rect 12362 26086 12414 26138
rect 12426 26086 12478 26138
rect 12490 26086 12542 26138
rect 19317 26086 19369 26138
rect 19381 26086 19433 26138
rect 19445 26086 19497 26138
rect 19509 26086 19561 26138
rect 19573 26086 19625 26138
rect 26400 26086 26452 26138
rect 26464 26086 26516 26138
rect 26528 26086 26580 26138
rect 26592 26086 26644 26138
rect 26656 26086 26708 26138
rect 5816 25984 5868 26036
rect 7932 25984 7984 26036
rect 5080 25848 5132 25900
rect 4344 25712 4396 25764
rect 5448 25891 5500 25900
rect 5448 25857 5457 25891
rect 5457 25857 5491 25891
rect 5491 25857 5500 25891
rect 5448 25848 5500 25857
rect 5632 25848 5684 25900
rect 6460 25916 6512 25968
rect 6552 25848 6604 25900
rect 6920 25848 6972 25900
rect 7196 25848 7248 25900
rect 18236 25916 18288 25968
rect 6828 25780 6880 25832
rect 20076 25848 20128 25900
rect 4988 25687 5040 25696
rect 4988 25653 4997 25687
rect 4997 25653 5031 25687
rect 5031 25653 5040 25687
rect 4988 25644 5040 25653
rect 5632 25687 5684 25696
rect 5632 25653 5641 25687
rect 5641 25653 5675 25687
rect 5675 25653 5684 25687
rect 5632 25644 5684 25653
rect 5724 25687 5776 25696
rect 5724 25653 5733 25687
rect 5733 25653 5767 25687
rect 5767 25653 5776 25687
rect 5724 25644 5776 25653
rect 8576 25780 8628 25832
rect 17868 25780 17920 25832
rect 7748 25712 7800 25764
rect 6828 25644 6880 25696
rect 7288 25644 7340 25696
rect 7564 25644 7616 25696
rect 8760 25644 8812 25696
rect 20720 25644 20772 25696
rect 4491 25542 4543 25594
rect 4555 25542 4607 25594
rect 4619 25542 4671 25594
rect 4683 25542 4735 25594
rect 4747 25542 4799 25594
rect 11574 25542 11626 25594
rect 11638 25542 11690 25594
rect 11702 25542 11754 25594
rect 11766 25542 11818 25594
rect 11830 25542 11882 25594
rect 18657 25542 18709 25594
rect 18721 25542 18773 25594
rect 18785 25542 18837 25594
rect 18849 25542 18901 25594
rect 18913 25542 18965 25594
rect 25740 25542 25792 25594
rect 25804 25542 25856 25594
rect 25868 25542 25920 25594
rect 25932 25542 25984 25594
rect 25996 25542 26048 25594
rect 6368 25440 6420 25492
rect 6828 25440 6880 25492
rect 7012 25440 7064 25492
rect 7748 25440 7800 25492
rect 8760 25483 8812 25492
rect 8760 25449 8769 25483
rect 8769 25449 8803 25483
rect 8803 25449 8812 25483
rect 8760 25440 8812 25449
rect 18880 25440 18932 25492
rect 18144 25372 18196 25424
rect 4160 25304 4212 25356
rect 4344 25236 4396 25288
rect 4620 25279 4672 25288
rect 4620 25245 4629 25279
rect 4629 25245 4663 25279
rect 4663 25245 4672 25279
rect 4620 25236 4672 25245
rect 4988 25347 5040 25356
rect 4988 25313 4997 25347
rect 4997 25313 5031 25347
rect 5031 25313 5040 25347
rect 4988 25304 5040 25313
rect 5448 25304 5500 25356
rect 13452 25304 13504 25356
rect 15016 25347 15068 25356
rect 15016 25313 15025 25347
rect 15025 25313 15059 25347
rect 15059 25313 15068 25347
rect 15016 25304 15068 25313
rect 4896 25168 4948 25220
rect 5540 25168 5592 25220
rect 8392 25236 8444 25288
rect 9128 25236 9180 25288
rect 12992 25236 13044 25288
rect 17776 25304 17828 25356
rect 17868 25236 17920 25288
rect 19248 25304 19300 25356
rect 18788 25279 18840 25288
rect 18788 25245 18797 25279
rect 18797 25245 18831 25279
rect 18831 25245 18840 25279
rect 18788 25236 18840 25245
rect 18880 25279 18932 25288
rect 18880 25245 18915 25279
rect 18915 25245 18932 25279
rect 18880 25236 18932 25245
rect 19064 25279 19116 25288
rect 19064 25245 19073 25279
rect 19073 25245 19107 25279
rect 19107 25245 19116 25279
rect 19064 25236 19116 25245
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 19708 25304 19760 25356
rect 19892 25304 19944 25356
rect 21916 25304 21968 25356
rect 19800 25236 19852 25288
rect 7196 25168 7248 25220
rect 14924 25168 14976 25220
rect 16580 25168 16632 25220
rect 3056 25100 3108 25152
rect 4528 25100 4580 25152
rect 4804 25100 4856 25152
rect 5080 25100 5132 25152
rect 5356 25100 5408 25152
rect 6460 25143 6512 25152
rect 6460 25109 6469 25143
rect 6469 25109 6503 25143
rect 6503 25109 6512 25143
rect 6460 25100 6512 25109
rect 7380 25100 7432 25152
rect 11888 25143 11940 25152
rect 11888 25109 11897 25143
rect 11897 25109 11931 25143
rect 11931 25109 11940 25143
rect 11888 25100 11940 25109
rect 17408 25211 17460 25220
rect 17408 25177 17417 25211
rect 17417 25177 17451 25211
rect 17451 25177 17460 25211
rect 17408 25168 17460 25177
rect 17040 25143 17092 25152
rect 17040 25109 17049 25143
rect 17049 25109 17083 25143
rect 17083 25109 17092 25143
rect 17040 25100 17092 25109
rect 18420 25143 18472 25152
rect 18420 25109 18429 25143
rect 18429 25109 18463 25143
rect 18463 25109 18472 25143
rect 18420 25100 18472 25109
rect 20260 25236 20312 25288
rect 21180 25168 21232 25220
rect 22284 25168 22336 25220
rect 19156 25100 19208 25152
rect 19524 25100 19576 25152
rect 19984 25100 20036 25152
rect 20168 25100 20220 25152
rect 5151 24998 5203 25050
rect 5215 24998 5267 25050
rect 5279 24998 5331 25050
rect 5343 24998 5395 25050
rect 5407 24998 5459 25050
rect 12234 24998 12286 25050
rect 12298 24998 12350 25050
rect 12362 24998 12414 25050
rect 12426 24998 12478 25050
rect 12490 24998 12542 25050
rect 19317 24998 19369 25050
rect 19381 24998 19433 25050
rect 19445 24998 19497 25050
rect 19509 24998 19561 25050
rect 19573 24998 19625 25050
rect 26400 24998 26452 25050
rect 26464 24998 26516 25050
rect 26528 24998 26580 25050
rect 26592 24998 26644 25050
rect 26656 24998 26708 25050
rect 4896 24896 4948 24948
rect 5724 24896 5776 24948
rect 6460 24896 6512 24948
rect 7564 24896 7616 24948
rect 14924 24939 14976 24948
rect 14924 24905 14933 24939
rect 14933 24905 14967 24939
rect 14967 24905 14976 24939
rect 14924 24896 14976 24905
rect 15292 24896 15344 24948
rect 16120 24896 16172 24948
rect 4804 24828 4856 24880
rect 4528 24760 4580 24812
rect 3424 24735 3476 24744
rect 3424 24701 3433 24735
rect 3433 24701 3467 24735
rect 3467 24701 3476 24735
rect 3424 24692 3476 24701
rect 4620 24692 4672 24744
rect 5080 24760 5132 24812
rect 5632 24760 5684 24812
rect 7196 24828 7248 24880
rect 9588 24828 9640 24880
rect 11888 24828 11940 24880
rect 6368 24803 6420 24812
rect 6368 24769 6377 24803
rect 6377 24769 6411 24803
rect 6411 24769 6420 24803
rect 6368 24760 6420 24769
rect 7380 24760 7432 24812
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 6644 24692 6696 24744
rect 5080 24624 5132 24676
rect 6920 24624 6972 24676
rect 7840 24735 7892 24744
rect 7840 24701 7849 24735
rect 7849 24701 7883 24735
rect 7883 24701 7892 24735
rect 7840 24692 7892 24701
rect 5172 24556 5224 24608
rect 5540 24556 5592 24608
rect 6368 24556 6420 24608
rect 11428 24760 11480 24812
rect 10600 24692 10652 24744
rect 14096 24828 14148 24880
rect 15568 24828 15620 24880
rect 14280 24760 14332 24812
rect 13728 24692 13780 24744
rect 10416 24556 10468 24608
rect 14464 24735 14516 24744
rect 14464 24701 14473 24735
rect 14473 24701 14507 24735
rect 14507 24701 14516 24735
rect 14464 24692 14516 24701
rect 14556 24735 14608 24744
rect 14556 24701 14565 24735
rect 14565 24701 14599 24735
rect 14599 24701 14608 24735
rect 14556 24692 14608 24701
rect 14924 24624 14976 24676
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 15384 24803 15436 24812
rect 15384 24769 15419 24803
rect 15419 24769 15436 24803
rect 15384 24760 15436 24769
rect 15660 24803 15712 24812
rect 15660 24769 15669 24803
rect 15669 24769 15703 24803
rect 15703 24769 15712 24803
rect 15660 24760 15712 24769
rect 16028 24760 16080 24812
rect 17040 24828 17092 24880
rect 19064 24896 19116 24948
rect 18328 24828 18380 24880
rect 18420 24828 18472 24880
rect 20168 24828 20220 24880
rect 22284 24828 22336 24880
rect 15936 24692 15988 24744
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18144 24803 18196 24812
rect 18144 24769 18179 24803
rect 18179 24769 18196 24803
rect 18144 24760 18196 24769
rect 19800 24760 19852 24812
rect 20076 24760 20128 24812
rect 16948 24692 17000 24744
rect 15108 24556 15160 24608
rect 19892 24692 19944 24744
rect 19984 24692 20036 24744
rect 20720 24760 20772 24812
rect 18236 24624 18288 24676
rect 16304 24556 16356 24608
rect 17592 24556 17644 24608
rect 20076 24556 20128 24608
rect 4491 24454 4543 24506
rect 4555 24454 4607 24506
rect 4619 24454 4671 24506
rect 4683 24454 4735 24506
rect 4747 24454 4799 24506
rect 11574 24454 11626 24506
rect 11638 24454 11690 24506
rect 11702 24454 11754 24506
rect 11766 24454 11818 24506
rect 11830 24454 11882 24506
rect 18657 24454 18709 24506
rect 18721 24454 18773 24506
rect 18785 24454 18837 24506
rect 18849 24454 18901 24506
rect 18913 24454 18965 24506
rect 25740 24454 25792 24506
rect 25804 24454 25856 24506
rect 25868 24454 25920 24506
rect 25932 24454 25984 24506
rect 25996 24454 26048 24506
rect 3424 24352 3476 24404
rect 4988 24352 5040 24404
rect 5172 24284 5224 24336
rect 6644 24352 6696 24404
rect 7380 24352 7432 24404
rect 7656 24352 7708 24404
rect 14464 24352 14516 24404
rect 15292 24352 15344 24404
rect 15660 24352 15712 24404
rect 15844 24352 15896 24404
rect 19248 24395 19300 24404
rect 19248 24361 19257 24395
rect 19257 24361 19291 24395
rect 19291 24361 19300 24395
rect 19248 24352 19300 24361
rect 19708 24352 19760 24404
rect 13176 24284 13228 24336
rect 16212 24284 16264 24336
rect 4896 24216 4948 24268
rect 7840 24216 7892 24268
rect 15016 24216 15068 24268
rect 6552 24148 6604 24200
rect 7012 24148 7064 24200
rect 7288 24191 7340 24200
rect 7288 24157 7297 24191
rect 7297 24157 7331 24191
rect 7331 24157 7340 24191
rect 7288 24148 7340 24157
rect 10784 24148 10836 24200
rect 13912 24148 13964 24200
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 17224 24216 17276 24268
rect 16212 24148 16264 24200
rect 17776 24148 17828 24200
rect 19064 24148 19116 24200
rect 5632 24080 5684 24132
rect 11796 24080 11848 24132
rect 11888 24123 11940 24132
rect 11888 24089 11897 24123
rect 11897 24089 11931 24123
rect 11931 24089 11940 24123
rect 11888 24080 11940 24089
rect 13544 24080 13596 24132
rect 9680 24012 9732 24064
rect 15108 24080 15160 24132
rect 14280 24012 14332 24064
rect 15844 24012 15896 24064
rect 16028 24123 16080 24132
rect 16028 24089 16037 24123
rect 16037 24089 16071 24123
rect 16071 24089 16080 24123
rect 16028 24080 16080 24089
rect 18052 24080 18104 24132
rect 19708 24191 19760 24200
rect 19708 24157 19717 24191
rect 19717 24157 19751 24191
rect 19751 24157 19760 24191
rect 19708 24148 19760 24157
rect 19984 24123 20036 24132
rect 19984 24089 19993 24123
rect 19993 24089 20027 24123
rect 20027 24089 20036 24123
rect 19984 24080 20036 24089
rect 16764 24012 16816 24064
rect 17592 24012 17644 24064
rect 20168 24148 20220 24200
rect 20076 24012 20128 24064
rect 5151 23910 5203 23962
rect 5215 23910 5267 23962
rect 5279 23910 5331 23962
rect 5343 23910 5395 23962
rect 5407 23910 5459 23962
rect 12234 23910 12286 23962
rect 12298 23910 12350 23962
rect 12362 23910 12414 23962
rect 12426 23910 12478 23962
rect 12490 23910 12542 23962
rect 19317 23910 19369 23962
rect 19381 23910 19433 23962
rect 19445 23910 19497 23962
rect 19509 23910 19561 23962
rect 19573 23910 19625 23962
rect 26400 23910 26452 23962
rect 26464 23910 26516 23962
rect 26528 23910 26580 23962
rect 26592 23910 26644 23962
rect 26656 23910 26708 23962
rect 5816 23808 5868 23860
rect 11796 23808 11848 23860
rect 11888 23808 11940 23860
rect 12992 23851 13044 23860
rect 12992 23817 13001 23851
rect 13001 23817 13035 23851
rect 13035 23817 13044 23851
rect 12992 23808 13044 23817
rect 15568 23808 15620 23860
rect 16764 23808 16816 23860
rect 1492 23715 1544 23724
rect 1492 23681 1501 23715
rect 1501 23681 1535 23715
rect 1535 23681 1544 23715
rect 1492 23672 1544 23681
rect 10600 23672 10652 23724
rect 9128 23604 9180 23656
rect 12808 23672 12860 23724
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 10968 23511 11020 23520
rect 10968 23477 10977 23511
rect 10977 23477 11011 23511
rect 11011 23477 11020 23511
rect 10968 23468 11020 23477
rect 12164 23511 12216 23520
rect 12164 23477 12173 23511
rect 12173 23477 12207 23511
rect 12207 23477 12216 23511
rect 12164 23468 12216 23477
rect 16304 23740 16356 23792
rect 16948 23740 17000 23792
rect 13728 23604 13780 23656
rect 14280 23604 14332 23656
rect 14464 23647 14516 23656
rect 14464 23613 14473 23647
rect 14473 23613 14507 23647
rect 14507 23613 14516 23647
rect 14464 23604 14516 23613
rect 15016 23715 15068 23724
rect 15016 23681 15025 23715
rect 15025 23681 15059 23715
rect 15059 23681 15068 23715
rect 15016 23672 15068 23681
rect 15384 23672 15436 23724
rect 15200 23536 15252 23588
rect 15568 23715 15620 23724
rect 15568 23681 15577 23715
rect 15577 23681 15611 23715
rect 15611 23681 15620 23715
rect 15568 23672 15620 23681
rect 16028 23604 16080 23656
rect 17224 23715 17276 23724
rect 17224 23681 17233 23715
rect 17233 23681 17267 23715
rect 17267 23681 17276 23715
rect 17224 23672 17276 23681
rect 19708 23672 19760 23724
rect 17592 23604 17644 23656
rect 15844 23536 15896 23588
rect 16212 23536 16264 23588
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 19064 23604 19116 23656
rect 19708 23536 19760 23588
rect 19984 23536 20036 23588
rect 16120 23511 16172 23520
rect 16120 23477 16129 23511
rect 16129 23477 16163 23511
rect 16163 23477 16172 23511
rect 16120 23468 16172 23477
rect 4491 23366 4543 23418
rect 4555 23366 4607 23418
rect 4619 23366 4671 23418
rect 4683 23366 4735 23418
rect 4747 23366 4799 23418
rect 11574 23366 11626 23418
rect 11638 23366 11690 23418
rect 11702 23366 11754 23418
rect 11766 23366 11818 23418
rect 11830 23366 11882 23418
rect 18657 23366 18709 23418
rect 18721 23366 18773 23418
rect 18785 23366 18837 23418
rect 18849 23366 18901 23418
rect 18913 23366 18965 23418
rect 25740 23366 25792 23418
rect 25804 23366 25856 23418
rect 25868 23366 25920 23418
rect 25932 23366 25984 23418
rect 25996 23366 26048 23418
rect 6552 23128 6604 23180
rect 9128 23264 9180 23316
rect 11428 23264 11480 23316
rect 14556 23264 14608 23316
rect 15016 23307 15068 23316
rect 15016 23273 15025 23307
rect 15025 23273 15059 23307
rect 15059 23273 15068 23307
rect 15016 23264 15068 23273
rect 15108 23264 15160 23316
rect 15384 23264 15436 23316
rect 17408 23264 17460 23316
rect 25228 23307 25280 23316
rect 25228 23273 25237 23307
rect 25237 23273 25271 23307
rect 25271 23273 25280 23307
rect 25228 23264 25280 23273
rect 10600 23196 10652 23248
rect 10784 23239 10836 23248
rect 10784 23205 10793 23239
rect 10793 23205 10827 23239
rect 10827 23205 10836 23239
rect 10784 23196 10836 23205
rect 6184 23060 6236 23112
rect 15200 23239 15252 23248
rect 15200 23205 15209 23239
rect 15209 23205 15243 23239
rect 15243 23205 15252 23239
rect 15200 23196 15252 23205
rect 15568 23239 15620 23248
rect 15568 23205 15577 23239
rect 15577 23205 15611 23239
rect 15611 23205 15620 23239
rect 15568 23196 15620 23205
rect 15844 23196 15896 23248
rect 18144 23196 18196 23248
rect 11428 23128 11480 23180
rect 14556 23128 14608 23180
rect 14280 23060 14332 23112
rect 14464 23103 14516 23112
rect 14464 23069 14473 23103
rect 14473 23069 14507 23103
rect 14507 23069 14516 23103
rect 14464 23060 14516 23069
rect 14924 23060 14976 23112
rect 5080 22967 5132 22976
rect 5080 22933 5089 22967
rect 5089 22933 5123 22967
rect 5123 22933 5132 22967
rect 5080 22924 5132 22933
rect 5908 22924 5960 22976
rect 9312 23035 9364 23044
rect 9312 23001 9321 23035
rect 9321 23001 9355 23035
rect 9355 23001 9364 23035
rect 9312 22992 9364 23001
rect 10876 23035 10928 23044
rect 10876 23001 10885 23035
rect 10885 23001 10919 23035
rect 10919 23001 10928 23035
rect 10876 22992 10928 23001
rect 15292 23103 15344 23112
rect 15292 23069 15301 23103
rect 15301 23069 15335 23103
rect 15335 23069 15344 23103
rect 15292 23060 15344 23069
rect 16028 23171 16080 23180
rect 16028 23137 16037 23171
rect 16037 23137 16071 23171
rect 16071 23137 16080 23171
rect 16028 23128 16080 23137
rect 15200 22992 15252 23044
rect 15568 22992 15620 23044
rect 16120 23060 16172 23112
rect 21640 23128 21692 23180
rect 13728 22924 13780 22976
rect 14648 22924 14700 22976
rect 15016 22924 15068 22976
rect 17316 22992 17368 23044
rect 18328 23060 18380 23112
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 20812 23103 20864 23112
rect 20812 23069 20821 23103
rect 20821 23069 20855 23103
rect 20855 23069 20864 23103
rect 20812 23060 20864 23069
rect 21088 23103 21140 23112
rect 21088 23069 21097 23103
rect 21097 23069 21131 23103
rect 21131 23069 21140 23103
rect 21088 23060 21140 23069
rect 23756 23060 23808 23112
rect 24492 23103 24544 23112
rect 24492 23069 24501 23103
rect 24501 23069 24535 23103
rect 24535 23069 24544 23103
rect 24492 23060 24544 23069
rect 21180 23035 21232 23044
rect 21180 23001 21189 23035
rect 21189 23001 21223 23035
rect 21223 23001 21232 23035
rect 21180 22992 21232 23001
rect 22560 22992 22612 23044
rect 24676 23060 24728 23112
rect 17224 22924 17276 22976
rect 17592 22924 17644 22976
rect 18052 22924 18104 22976
rect 20996 22967 21048 22976
rect 20996 22933 21005 22967
rect 21005 22933 21039 22967
rect 21039 22933 21048 22967
rect 20996 22924 21048 22933
rect 23848 22924 23900 22976
rect 24400 22924 24452 22976
rect 24768 22924 24820 22976
rect 25504 22992 25556 23044
rect 25412 22924 25464 22976
rect 5151 22822 5203 22874
rect 5215 22822 5267 22874
rect 5279 22822 5331 22874
rect 5343 22822 5395 22874
rect 5407 22822 5459 22874
rect 12234 22822 12286 22874
rect 12298 22822 12350 22874
rect 12362 22822 12414 22874
rect 12426 22822 12478 22874
rect 12490 22822 12542 22874
rect 19317 22822 19369 22874
rect 19381 22822 19433 22874
rect 19445 22822 19497 22874
rect 19509 22822 19561 22874
rect 19573 22822 19625 22874
rect 26400 22822 26452 22874
rect 26464 22822 26516 22874
rect 26528 22822 26580 22874
rect 26592 22822 26644 22874
rect 26656 22822 26708 22874
rect 9312 22720 9364 22772
rect 9496 22720 9548 22772
rect 5908 22652 5960 22704
rect 9680 22652 9732 22704
rect 10968 22652 11020 22704
rect 12808 22763 12860 22772
rect 12808 22729 12817 22763
rect 12817 22729 12851 22763
rect 12851 22729 12860 22763
rect 12808 22720 12860 22729
rect 5724 22516 5776 22568
rect 6000 22559 6052 22568
rect 6000 22525 6009 22559
rect 6009 22525 6043 22559
rect 6043 22525 6052 22559
rect 6000 22516 6052 22525
rect 7104 22627 7156 22636
rect 7104 22593 7113 22627
rect 7113 22593 7147 22627
rect 7147 22593 7156 22627
rect 7104 22584 7156 22593
rect 8116 22584 8168 22636
rect 8668 22627 8720 22636
rect 8668 22593 8677 22627
rect 8677 22593 8711 22627
rect 8711 22593 8720 22627
rect 8668 22584 8720 22593
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 7656 22559 7708 22568
rect 7656 22525 7665 22559
rect 7665 22525 7699 22559
rect 7699 22525 7708 22559
rect 7656 22516 7708 22525
rect 9128 22584 9180 22636
rect 11336 22584 11388 22636
rect 12164 22584 12216 22636
rect 10140 22516 10192 22568
rect 10784 22516 10836 22568
rect 11428 22516 11480 22568
rect 8576 22448 8628 22500
rect 11244 22448 11296 22500
rect 12624 22627 12676 22636
rect 12624 22593 12633 22627
rect 12633 22593 12667 22627
rect 12667 22593 12676 22627
rect 12624 22584 12676 22593
rect 13176 22584 13228 22636
rect 14280 22584 14332 22636
rect 15844 22720 15896 22772
rect 20720 22720 20772 22772
rect 15384 22695 15436 22704
rect 15384 22661 15393 22695
rect 15393 22661 15427 22695
rect 15427 22661 15436 22695
rect 15384 22652 15436 22661
rect 15936 22652 15988 22704
rect 13728 22448 13780 22500
rect 15476 22516 15528 22568
rect 16488 22516 16540 22568
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 20536 22559 20588 22568
rect 20536 22525 20545 22559
rect 20545 22525 20579 22559
rect 20579 22525 20588 22559
rect 20536 22516 20588 22525
rect 4160 22380 4212 22432
rect 7288 22423 7340 22432
rect 7288 22389 7297 22423
rect 7297 22389 7331 22423
rect 7331 22389 7340 22423
rect 7288 22380 7340 22389
rect 7380 22380 7432 22432
rect 9404 22380 9456 22432
rect 10232 22380 10284 22432
rect 14832 22423 14884 22432
rect 14832 22389 14841 22423
rect 14841 22389 14875 22423
rect 14875 22389 14884 22423
rect 14832 22380 14884 22389
rect 15568 22448 15620 22500
rect 16396 22448 16448 22500
rect 20812 22584 20864 22636
rect 22836 22720 22888 22772
rect 21088 22652 21140 22704
rect 21732 22652 21784 22704
rect 21180 22516 21232 22568
rect 21640 22584 21692 22636
rect 21916 22584 21968 22636
rect 22652 22516 22704 22568
rect 23020 22584 23072 22636
rect 23112 22627 23164 22636
rect 23112 22593 23121 22627
rect 23121 22593 23155 22627
rect 23155 22593 23164 22627
rect 23112 22584 23164 22593
rect 23204 22584 23256 22636
rect 23296 22627 23348 22636
rect 23296 22593 23305 22627
rect 23305 22593 23339 22627
rect 23339 22593 23348 22627
rect 23296 22584 23348 22593
rect 25320 22720 25372 22772
rect 25412 22763 25464 22772
rect 25412 22729 25421 22763
rect 25421 22729 25455 22763
rect 25455 22729 25464 22763
rect 25412 22720 25464 22729
rect 21640 22448 21692 22500
rect 23848 22584 23900 22636
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 23480 22516 23532 22568
rect 24400 22584 24452 22636
rect 24032 22448 24084 22500
rect 24400 22448 24452 22500
rect 24768 22627 24820 22636
rect 24768 22593 24777 22627
rect 24777 22593 24811 22627
rect 24811 22593 24820 22627
rect 24768 22584 24820 22593
rect 25044 22627 25096 22636
rect 25044 22593 25053 22627
rect 25053 22593 25087 22627
rect 25087 22593 25096 22627
rect 25044 22584 25096 22593
rect 25228 22627 25280 22636
rect 25228 22593 25237 22627
rect 25237 22593 25271 22627
rect 25271 22593 25280 22627
rect 25228 22584 25280 22593
rect 28816 22627 28868 22636
rect 28816 22593 28825 22627
rect 28825 22593 28859 22627
rect 28859 22593 28868 22627
rect 28816 22584 28868 22593
rect 24952 22516 25004 22568
rect 24584 22448 24636 22500
rect 29000 22491 29052 22500
rect 29000 22457 29009 22491
rect 29009 22457 29043 22491
rect 29043 22457 29052 22491
rect 29000 22448 29052 22457
rect 20812 22380 20864 22432
rect 21088 22423 21140 22432
rect 21088 22389 21097 22423
rect 21097 22389 21131 22423
rect 21131 22389 21140 22423
rect 21088 22380 21140 22389
rect 22100 22380 22152 22432
rect 22744 22423 22796 22432
rect 22744 22389 22753 22423
rect 22753 22389 22787 22423
rect 22787 22389 22796 22423
rect 22744 22380 22796 22389
rect 23204 22423 23256 22432
rect 23204 22389 23213 22423
rect 23213 22389 23247 22423
rect 23247 22389 23256 22423
rect 23204 22380 23256 22389
rect 23388 22380 23440 22432
rect 24952 22380 25004 22432
rect 4491 22278 4543 22330
rect 4555 22278 4607 22330
rect 4619 22278 4671 22330
rect 4683 22278 4735 22330
rect 4747 22278 4799 22330
rect 11574 22278 11626 22330
rect 11638 22278 11690 22330
rect 11702 22278 11754 22330
rect 11766 22278 11818 22330
rect 11830 22278 11882 22330
rect 18657 22278 18709 22330
rect 18721 22278 18773 22330
rect 18785 22278 18837 22330
rect 18849 22278 18901 22330
rect 18913 22278 18965 22330
rect 25740 22278 25792 22330
rect 25804 22278 25856 22330
rect 25868 22278 25920 22330
rect 25932 22278 25984 22330
rect 25996 22278 26048 22330
rect 7288 22176 7340 22228
rect 7656 22176 7708 22228
rect 8668 22176 8720 22228
rect 11244 22176 11296 22228
rect 11336 22176 11388 22228
rect 12624 22176 12676 22228
rect 13728 22176 13780 22228
rect 14832 22176 14884 22228
rect 21640 22219 21692 22228
rect 21640 22185 21649 22219
rect 21649 22185 21683 22219
rect 21683 22185 21692 22219
rect 21640 22176 21692 22185
rect 21732 22176 21784 22228
rect 8116 22108 8168 22160
rect 9956 22108 10008 22160
rect 21272 22108 21324 22160
rect 3700 22040 3752 22092
rect 5448 22040 5500 22092
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 6368 22040 6420 22092
rect 4252 21972 4304 22024
rect 4988 21972 5040 22024
rect 5540 21972 5592 22024
rect 4896 21904 4948 21956
rect 3240 21836 3292 21888
rect 4712 21836 4764 21888
rect 5908 21879 5960 21888
rect 5908 21845 5917 21879
rect 5917 21845 5951 21879
rect 5951 21845 5960 21879
rect 5908 21836 5960 21845
rect 8576 21972 8628 22024
rect 7104 21836 7156 21888
rect 7840 21836 7892 21888
rect 8484 21879 8536 21888
rect 8484 21845 8493 21879
rect 8493 21845 8527 21879
rect 8527 21845 8536 21879
rect 8484 21836 8536 21845
rect 9128 21904 9180 21956
rect 10048 22040 10100 22092
rect 10140 22040 10192 22092
rect 10600 22040 10652 22092
rect 12900 22040 12952 22092
rect 14464 22083 14516 22092
rect 14464 22049 14473 22083
rect 14473 22049 14507 22083
rect 14507 22049 14516 22083
rect 14464 22040 14516 22049
rect 16488 22040 16540 22092
rect 9496 21836 9548 21888
rect 10232 21836 10284 21888
rect 10508 22015 10560 22024
rect 10508 21981 10518 22015
rect 10518 21981 10552 22015
rect 10552 21981 10560 22015
rect 10508 21972 10560 21981
rect 10784 22015 10836 22024
rect 10784 21981 10793 22015
rect 10793 21981 10827 22015
rect 10827 21981 10836 22015
rect 10784 21972 10836 21981
rect 18420 21972 18472 22024
rect 11980 21904 12032 21956
rect 12624 21904 12676 21956
rect 13452 21904 13504 21956
rect 17776 21904 17828 21956
rect 19800 21904 19852 21956
rect 20444 21972 20496 22024
rect 20720 21972 20772 22024
rect 20812 22015 20864 22024
rect 20812 21981 20821 22015
rect 20821 21981 20855 22015
rect 20855 21981 20864 22015
rect 20812 21972 20864 21981
rect 20996 21972 21048 22024
rect 21088 22015 21140 22024
rect 21088 21981 21097 22015
rect 21097 21981 21131 22015
rect 21131 21981 21140 22015
rect 21088 21972 21140 21981
rect 21548 22108 21600 22160
rect 22560 22176 22612 22228
rect 21456 22015 21508 22024
rect 21456 21981 21465 22015
rect 21465 21981 21499 22015
rect 21499 21981 21508 22015
rect 21456 21972 21508 21981
rect 21548 21972 21600 22024
rect 21824 21972 21876 22024
rect 23940 22108 23992 22160
rect 22560 22083 22612 22092
rect 22560 22049 22569 22083
rect 22569 22049 22603 22083
rect 22603 22049 22612 22083
rect 22560 22040 22612 22049
rect 22100 21972 22152 22024
rect 24584 22176 24636 22228
rect 22744 21972 22796 22024
rect 22836 22015 22888 22024
rect 22836 21981 22845 22015
rect 22845 21981 22879 22015
rect 22879 21981 22888 22015
rect 22836 21972 22888 21981
rect 23112 21972 23164 22024
rect 23204 22015 23256 22024
rect 23204 21981 23213 22015
rect 23213 21981 23247 22015
rect 23247 21981 23256 22015
rect 23204 21972 23256 21981
rect 23756 21972 23808 22024
rect 23940 22015 23992 22024
rect 23940 21981 23949 22015
rect 23949 21981 23983 22015
rect 23983 21981 23992 22015
rect 23940 21972 23992 21981
rect 24124 22015 24176 22024
rect 24124 21981 24133 22015
rect 24133 21981 24167 22015
rect 24167 21981 24176 22015
rect 24124 21972 24176 21981
rect 24400 22015 24452 22024
rect 24400 21981 24409 22015
rect 24409 21981 24443 22015
rect 24443 21981 24452 22015
rect 24400 21972 24452 21981
rect 24492 21972 24544 22024
rect 21180 21904 21232 21956
rect 10508 21836 10560 21888
rect 12072 21836 12124 21888
rect 12716 21836 12768 21888
rect 13544 21836 13596 21888
rect 16488 21836 16540 21888
rect 16672 21836 16724 21888
rect 17868 21879 17920 21888
rect 17868 21845 17877 21879
rect 17877 21845 17911 21879
rect 17911 21845 17920 21879
rect 17868 21836 17920 21845
rect 20352 21879 20404 21888
rect 20352 21845 20361 21879
rect 20361 21845 20395 21879
rect 20395 21845 20404 21879
rect 20352 21836 20404 21845
rect 20444 21836 20496 21888
rect 20996 21836 21048 21888
rect 22468 21836 22520 21888
rect 23480 21836 23532 21888
rect 24584 21836 24636 21888
rect 24768 21836 24820 21888
rect 24952 21972 25004 22024
rect 25044 21972 25096 22024
rect 25228 21972 25280 22024
rect 25504 21972 25556 22024
rect 28816 21972 28868 22024
rect 25596 21836 25648 21888
rect 5151 21734 5203 21786
rect 5215 21734 5267 21786
rect 5279 21734 5331 21786
rect 5343 21734 5395 21786
rect 5407 21734 5459 21786
rect 12234 21734 12286 21786
rect 12298 21734 12350 21786
rect 12362 21734 12414 21786
rect 12426 21734 12478 21786
rect 12490 21734 12542 21786
rect 19317 21734 19369 21786
rect 19381 21734 19433 21786
rect 19445 21734 19497 21786
rect 19509 21734 19561 21786
rect 19573 21734 19625 21786
rect 26400 21734 26452 21786
rect 26464 21734 26516 21786
rect 26528 21734 26580 21786
rect 26592 21734 26644 21786
rect 26656 21734 26708 21786
rect 4160 21632 4212 21684
rect 4068 21564 4120 21616
rect 4344 21564 4396 21616
rect 4896 21632 4948 21684
rect 5540 21675 5592 21684
rect 5540 21641 5549 21675
rect 5549 21641 5583 21675
rect 5583 21641 5592 21675
rect 5540 21632 5592 21641
rect 5632 21632 5684 21684
rect 3240 21496 3292 21548
rect 3700 21496 3752 21548
rect 5908 21632 5960 21684
rect 6184 21675 6236 21684
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 5080 21428 5132 21480
rect 6000 21539 6052 21548
rect 6000 21505 6009 21539
rect 6009 21505 6043 21539
rect 6043 21505 6052 21539
rect 6000 21496 6052 21505
rect 7932 21632 7984 21684
rect 7104 21564 7156 21616
rect 8392 21607 8444 21616
rect 8392 21573 8401 21607
rect 8401 21573 8435 21607
rect 8435 21573 8444 21607
rect 8392 21564 8444 21573
rect 8484 21607 8536 21616
rect 8484 21573 8493 21607
rect 8493 21573 8527 21607
rect 8527 21573 8536 21607
rect 8484 21564 8536 21573
rect 8116 21496 8168 21548
rect 5816 21360 5868 21412
rect 3700 21335 3752 21344
rect 3700 21301 3709 21335
rect 3709 21301 3743 21335
rect 3743 21301 3752 21335
rect 3700 21292 3752 21301
rect 3792 21292 3844 21344
rect 4068 21292 4120 21344
rect 8576 21539 8628 21548
rect 8576 21505 8585 21539
rect 8585 21505 8619 21539
rect 8619 21505 8628 21539
rect 8576 21496 8628 21505
rect 9956 21632 10008 21684
rect 10784 21632 10836 21684
rect 11060 21632 11112 21684
rect 10600 21564 10652 21616
rect 10968 21564 11020 21616
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 12164 21539 12216 21548
rect 12164 21505 12174 21539
rect 12174 21505 12208 21539
rect 12208 21505 12216 21539
rect 12164 21496 12216 21505
rect 6460 21292 6512 21344
rect 7380 21292 7432 21344
rect 7840 21292 7892 21344
rect 10048 21428 10100 21480
rect 12624 21496 12676 21548
rect 12716 21428 12768 21480
rect 9128 21292 9180 21344
rect 9496 21292 9548 21344
rect 10600 21292 10652 21344
rect 10784 21335 10836 21344
rect 10784 21301 10793 21335
rect 10793 21301 10827 21335
rect 10827 21301 10836 21335
rect 10784 21292 10836 21301
rect 12716 21335 12768 21344
rect 12716 21301 12725 21335
rect 12725 21301 12759 21335
rect 12759 21301 12768 21335
rect 12716 21292 12768 21301
rect 14464 21632 14516 21684
rect 17776 21632 17828 21684
rect 13084 21564 13136 21616
rect 13636 21564 13688 21616
rect 18420 21675 18472 21684
rect 18420 21641 18429 21675
rect 18429 21641 18463 21675
rect 18463 21641 18472 21675
rect 18420 21632 18472 21641
rect 19248 21564 19300 21616
rect 20812 21675 20864 21684
rect 20812 21641 20821 21675
rect 20821 21641 20855 21675
rect 20855 21641 20864 21675
rect 20812 21632 20864 21641
rect 20996 21632 21048 21684
rect 22652 21632 22704 21684
rect 23480 21632 23532 21684
rect 23572 21632 23624 21684
rect 24492 21632 24544 21684
rect 13268 21428 13320 21480
rect 16580 21428 16632 21480
rect 16948 21471 17000 21480
rect 16948 21437 16957 21471
rect 16957 21437 16991 21471
rect 16991 21437 17000 21471
rect 16948 21428 17000 21437
rect 18512 21496 18564 21548
rect 19156 21539 19208 21548
rect 19156 21505 19165 21539
rect 19165 21505 19199 21539
rect 19199 21505 19208 21539
rect 19156 21496 19208 21505
rect 19340 21539 19392 21548
rect 19340 21505 19349 21539
rect 19349 21505 19383 21539
rect 19383 21505 19392 21539
rect 19340 21496 19392 21505
rect 21180 21564 21232 21616
rect 21364 21564 21416 21616
rect 12992 21292 13044 21344
rect 14740 21292 14792 21344
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 20352 21428 20404 21480
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 21088 21539 21140 21548
rect 21088 21505 21097 21539
rect 21097 21505 21131 21539
rect 21131 21505 21140 21539
rect 21088 21496 21140 21505
rect 21272 21471 21324 21480
rect 19248 21292 19300 21344
rect 19524 21335 19576 21344
rect 19524 21301 19533 21335
rect 19533 21301 19567 21335
rect 19567 21301 19576 21335
rect 19524 21292 19576 21301
rect 21272 21437 21281 21471
rect 21281 21437 21315 21471
rect 21315 21437 21324 21471
rect 21272 21428 21324 21437
rect 21364 21471 21416 21480
rect 21364 21437 21373 21471
rect 21373 21437 21407 21471
rect 21407 21437 21416 21471
rect 21364 21428 21416 21437
rect 21916 21496 21968 21548
rect 23112 21564 23164 21616
rect 23756 21564 23808 21616
rect 22468 21539 22520 21548
rect 22468 21505 22477 21539
rect 22477 21505 22511 21539
rect 22511 21505 22520 21539
rect 22468 21496 22520 21505
rect 22744 21496 22796 21548
rect 23388 21496 23440 21548
rect 23572 21496 23624 21548
rect 24032 21496 24084 21548
rect 24400 21496 24452 21548
rect 24676 21539 24728 21548
rect 24676 21505 24685 21539
rect 24685 21505 24719 21539
rect 24719 21505 24728 21539
rect 24676 21496 24728 21505
rect 24952 21539 25004 21548
rect 24952 21505 24961 21539
rect 24961 21505 24995 21539
rect 24995 21505 25004 21539
rect 24952 21496 25004 21505
rect 25504 21539 25556 21548
rect 25504 21505 25513 21539
rect 25513 21505 25547 21539
rect 25547 21505 25556 21539
rect 25504 21496 25556 21505
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 27528 21539 27580 21548
rect 20720 21360 20772 21412
rect 20996 21292 21048 21344
rect 21456 21292 21508 21344
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 21824 21403 21876 21412
rect 21824 21369 21833 21403
rect 21833 21369 21867 21403
rect 21867 21369 21876 21403
rect 21824 21360 21876 21369
rect 22652 21292 22704 21344
rect 22928 21471 22980 21480
rect 22928 21437 22937 21471
rect 22937 21437 22971 21471
rect 22971 21437 22980 21471
rect 22928 21428 22980 21437
rect 23204 21403 23256 21412
rect 23204 21369 23213 21403
rect 23213 21369 23247 21403
rect 23247 21369 23256 21403
rect 23204 21360 23256 21369
rect 25596 21428 25648 21480
rect 27528 21505 27537 21539
rect 27537 21505 27571 21539
rect 27571 21505 27580 21539
rect 27528 21496 27580 21505
rect 27804 21496 27856 21548
rect 23664 21292 23716 21344
rect 23940 21335 23992 21344
rect 23940 21301 23949 21335
rect 23949 21301 23983 21335
rect 23983 21301 23992 21335
rect 23940 21292 23992 21301
rect 26240 21360 26292 21412
rect 27068 21403 27120 21412
rect 27068 21369 27077 21403
rect 27077 21369 27111 21403
rect 27111 21369 27120 21403
rect 27068 21360 27120 21369
rect 24952 21292 25004 21344
rect 27252 21292 27304 21344
rect 27620 21335 27672 21344
rect 27620 21301 27629 21335
rect 27629 21301 27663 21335
rect 27663 21301 27672 21335
rect 27620 21292 27672 21301
rect 4491 21190 4543 21242
rect 4555 21190 4607 21242
rect 4619 21190 4671 21242
rect 4683 21190 4735 21242
rect 4747 21190 4799 21242
rect 11574 21190 11626 21242
rect 11638 21190 11690 21242
rect 11702 21190 11754 21242
rect 11766 21190 11818 21242
rect 11830 21190 11882 21242
rect 18657 21190 18709 21242
rect 18721 21190 18773 21242
rect 18785 21190 18837 21242
rect 18849 21190 18901 21242
rect 18913 21190 18965 21242
rect 25740 21190 25792 21242
rect 25804 21190 25856 21242
rect 25868 21190 25920 21242
rect 25932 21190 25984 21242
rect 25996 21190 26048 21242
rect 3700 21088 3752 21140
rect 5724 21088 5776 21140
rect 3792 20995 3844 21004
rect 3792 20961 3801 20995
rect 3801 20961 3835 20995
rect 3835 20961 3844 20995
rect 6368 21088 6420 21140
rect 7472 21088 7524 21140
rect 10508 21088 10560 21140
rect 5908 21020 5960 21072
rect 8576 21020 8628 21072
rect 10232 21020 10284 21072
rect 3792 20952 3844 20961
rect 1860 20884 1912 20936
rect 5540 20884 5592 20936
rect 5908 20884 5960 20936
rect 6736 20884 6788 20936
rect 3424 20748 3476 20800
rect 4344 20748 4396 20800
rect 6184 20816 6236 20868
rect 5724 20748 5776 20800
rect 6920 20748 6972 20800
rect 7380 20927 7432 20936
rect 7380 20893 7390 20927
rect 7390 20893 7424 20927
rect 7424 20893 7432 20927
rect 7380 20884 7432 20893
rect 10784 20952 10836 21004
rect 7472 20816 7524 20868
rect 7656 20859 7708 20868
rect 7656 20825 7665 20859
rect 7665 20825 7699 20859
rect 7699 20825 7708 20859
rect 7656 20816 7708 20825
rect 10232 20884 10284 20936
rect 10876 20884 10928 20936
rect 11428 20927 11480 20936
rect 11428 20893 11437 20927
rect 11437 20893 11471 20927
rect 11471 20893 11480 20927
rect 11428 20884 11480 20893
rect 11520 20927 11572 20936
rect 11520 20893 11530 20927
rect 11530 20893 11564 20927
rect 11564 20893 11572 20927
rect 11520 20884 11572 20893
rect 14740 21131 14792 21140
rect 14740 21097 14749 21131
rect 14749 21097 14783 21131
rect 14783 21097 14792 21131
rect 14740 21088 14792 21097
rect 16948 21088 17000 21140
rect 17868 21088 17920 21140
rect 13452 21020 13504 21072
rect 11796 20952 11848 21004
rect 13912 20952 13964 21004
rect 9956 20816 10008 20868
rect 11152 20859 11204 20868
rect 11152 20825 11161 20859
rect 11161 20825 11195 20859
rect 11195 20825 11204 20859
rect 11152 20816 11204 20825
rect 8576 20748 8628 20800
rect 10140 20791 10192 20800
rect 10140 20757 10149 20791
rect 10149 20757 10183 20791
rect 10183 20757 10192 20791
rect 10140 20748 10192 20757
rect 10784 20748 10836 20800
rect 12900 20816 12952 20868
rect 11980 20748 12032 20800
rect 14188 20927 14240 20936
rect 14188 20893 14198 20927
rect 14198 20893 14232 20927
rect 14232 20893 14240 20927
rect 14188 20884 14240 20893
rect 19064 21088 19116 21140
rect 20996 21088 21048 21140
rect 18052 20952 18104 21004
rect 19156 20952 19208 21004
rect 16028 20884 16080 20936
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 17868 20884 17920 20936
rect 19524 20952 19576 21004
rect 20352 20995 20404 21004
rect 20352 20961 20361 20995
rect 20361 20961 20395 20995
rect 20395 20961 20404 20995
rect 20352 20952 20404 20961
rect 22192 21088 22244 21140
rect 23572 21088 23624 21140
rect 25596 21088 25648 21140
rect 26148 21088 26200 21140
rect 26976 21088 27028 21140
rect 21732 21020 21784 21072
rect 22836 21020 22888 21072
rect 13820 20748 13872 20800
rect 15752 20816 15804 20868
rect 16212 20859 16264 20868
rect 16212 20825 16221 20859
rect 16221 20825 16255 20859
rect 16255 20825 16264 20859
rect 16212 20816 16264 20825
rect 16948 20816 17000 20868
rect 18512 20816 18564 20868
rect 18604 20816 18656 20868
rect 14556 20748 14608 20800
rect 17500 20748 17552 20800
rect 19156 20748 19208 20800
rect 20536 20884 20588 20936
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 21364 20884 21416 20936
rect 21456 20927 21508 20936
rect 21456 20893 21465 20927
rect 21465 20893 21499 20927
rect 21499 20893 21508 20927
rect 21456 20884 21508 20893
rect 22192 20927 22244 20936
rect 21548 20816 21600 20868
rect 22192 20893 22201 20927
rect 22201 20893 22235 20927
rect 22235 20893 22244 20927
rect 22192 20884 22244 20893
rect 22652 20927 22704 20936
rect 22652 20893 22661 20927
rect 22661 20893 22695 20927
rect 22695 20893 22704 20927
rect 22652 20884 22704 20893
rect 22744 20884 22796 20936
rect 24860 20884 24912 20936
rect 24216 20816 24268 20868
rect 25320 20816 25372 20868
rect 25872 20859 25924 20868
rect 25872 20825 25881 20859
rect 25881 20825 25915 20859
rect 25915 20825 25924 20859
rect 25872 20816 25924 20825
rect 23296 20748 23348 20800
rect 23848 20748 23900 20800
rect 27068 20952 27120 21004
rect 27988 21020 28040 21072
rect 26240 20884 26292 20936
rect 26792 20927 26844 20936
rect 26792 20893 26801 20927
rect 26801 20893 26835 20927
rect 26835 20893 26844 20927
rect 26792 20884 26844 20893
rect 27528 20952 27580 21004
rect 27804 20952 27856 21004
rect 28908 20952 28960 21004
rect 27988 20816 28040 20868
rect 27436 20748 27488 20800
rect 28172 20791 28224 20800
rect 28172 20757 28181 20791
rect 28181 20757 28215 20791
rect 28215 20757 28224 20791
rect 28172 20748 28224 20757
rect 28540 20748 28592 20800
rect 5151 20646 5203 20698
rect 5215 20646 5267 20698
rect 5279 20646 5331 20698
rect 5343 20646 5395 20698
rect 5407 20646 5459 20698
rect 12234 20646 12286 20698
rect 12298 20646 12350 20698
rect 12362 20646 12414 20698
rect 12426 20646 12478 20698
rect 12490 20646 12542 20698
rect 19317 20646 19369 20698
rect 19381 20646 19433 20698
rect 19445 20646 19497 20698
rect 19509 20646 19561 20698
rect 19573 20646 19625 20698
rect 26400 20646 26452 20698
rect 26464 20646 26516 20698
rect 26528 20646 26580 20698
rect 26592 20646 26644 20698
rect 26656 20646 26708 20698
rect 4068 20476 4120 20528
rect 4344 20476 4396 20528
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 3976 20204 4028 20256
rect 6184 20544 6236 20596
rect 7472 20544 7524 20596
rect 9680 20544 9732 20596
rect 9864 20544 9916 20596
rect 7104 20476 7156 20528
rect 10048 20544 10100 20596
rect 13084 20544 13136 20596
rect 9680 20451 9732 20460
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 4896 20340 4948 20392
rect 6368 20383 6420 20392
rect 6368 20349 6377 20383
rect 6377 20349 6411 20383
rect 6411 20349 6420 20383
rect 6368 20340 6420 20349
rect 6644 20383 6696 20392
rect 6644 20349 6653 20383
rect 6653 20349 6687 20383
rect 6687 20349 6696 20383
rect 6644 20340 6696 20349
rect 4988 20204 5040 20256
rect 7012 20204 7064 20256
rect 7196 20204 7248 20256
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 12808 20476 12860 20528
rect 13912 20544 13964 20596
rect 15016 20544 15068 20596
rect 16212 20476 16264 20528
rect 10140 20408 10192 20460
rect 10600 20451 10652 20460
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 10968 20408 11020 20460
rect 11152 20408 11204 20460
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 8484 20272 8536 20324
rect 8208 20204 8260 20256
rect 10140 20204 10192 20256
rect 12072 20383 12124 20392
rect 12072 20349 12081 20383
rect 12081 20349 12115 20383
rect 12115 20349 12124 20383
rect 12072 20340 12124 20349
rect 14188 20408 14240 20460
rect 14464 20408 14516 20460
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 17408 20408 17460 20460
rect 17500 20451 17552 20460
rect 17500 20417 17509 20451
rect 17509 20417 17543 20451
rect 17543 20417 17552 20451
rect 17500 20408 17552 20417
rect 17592 20451 17644 20460
rect 17592 20417 17601 20451
rect 17601 20417 17635 20451
rect 17635 20417 17644 20451
rect 17592 20408 17644 20417
rect 17776 20408 17828 20460
rect 22560 20544 22612 20596
rect 22652 20544 22704 20596
rect 23112 20587 23164 20596
rect 23112 20553 23121 20587
rect 23121 20553 23155 20587
rect 23155 20553 23164 20587
rect 23112 20544 23164 20553
rect 24676 20544 24728 20596
rect 27068 20544 27120 20596
rect 18052 20408 18104 20460
rect 18328 20451 18380 20460
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 14648 20272 14700 20324
rect 18236 20340 18288 20392
rect 19064 20408 19116 20460
rect 21548 20476 21600 20528
rect 20904 20408 20956 20460
rect 21180 20451 21232 20460
rect 21180 20417 21189 20451
rect 21189 20417 21223 20451
rect 21223 20417 21232 20451
rect 21180 20408 21232 20417
rect 20536 20340 20588 20392
rect 21916 20408 21968 20460
rect 22744 20451 22796 20460
rect 22744 20417 22753 20451
rect 22753 20417 22787 20451
rect 22787 20417 22796 20451
rect 22744 20408 22796 20417
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 23664 20408 23716 20417
rect 23848 20451 23900 20460
rect 23848 20417 23857 20451
rect 23857 20417 23891 20451
rect 23891 20417 23900 20451
rect 23848 20408 23900 20417
rect 23940 20451 23992 20460
rect 23940 20417 23949 20451
rect 23949 20417 23983 20451
rect 23983 20417 23992 20451
rect 23940 20408 23992 20417
rect 25872 20476 25924 20528
rect 24216 20408 24268 20460
rect 26792 20476 26844 20528
rect 27344 20408 27396 20460
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 21732 20340 21784 20392
rect 28540 20476 28592 20528
rect 28080 20408 28132 20460
rect 28908 20451 28960 20460
rect 28908 20417 28917 20451
rect 28917 20417 28951 20451
rect 28951 20417 28960 20451
rect 28908 20408 28960 20417
rect 17040 20272 17092 20324
rect 19156 20272 19208 20324
rect 23664 20272 23716 20324
rect 27252 20272 27304 20324
rect 12532 20204 12584 20256
rect 14280 20247 14332 20256
rect 14280 20213 14289 20247
rect 14289 20213 14323 20247
rect 14323 20213 14332 20247
rect 14280 20204 14332 20213
rect 17868 20247 17920 20256
rect 17868 20213 17877 20247
rect 17877 20213 17911 20247
rect 17911 20213 17920 20247
rect 17868 20204 17920 20213
rect 24124 20204 24176 20256
rect 24492 20204 24544 20256
rect 27344 20247 27396 20256
rect 27344 20213 27353 20247
rect 27353 20213 27387 20247
rect 27387 20213 27396 20247
rect 27344 20204 27396 20213
rect 27528 20204 27580 20256
rect 27712 20247 27764 20256
rect 27712 20213 27721 20247
rect 27721 20213 27755 20247
rect 27755 20213 27764 20247
rect 27712 20204 27764 20213
rect 28356 20247 28408 20256
rect 28356 20213 28365 20247
rect 28365 20213 28399 20247
rect 28399 20213 28408 20247
rect 28356 20204 28408 20213
rect 4491 20102 4543 20154
rect 4555 20102 4607 20154
rect 4619 20102 4671 20154
rect 4683 20102 4735 20154
rect 4747 20102 4799 20154
rect 11574 20102 11626 20154
rect 11638 20102 11690 20154
rect 11702 20102 11754 20154
rect 11766 20102 11818 20154
rect 11830 20102 11882 20154
rect 18657 20102 18709 20154
rect 18721 20102 18773 20154
rect 18785 20102 18837 20154
rect 18849 20102 18901 20154
rect 18913 20102 18965 20154
rect 25740 20102 25792 20154
rect 25804 20102 25856 20154
rect 25868 20102 25920 20154
rect 25932 20102 25984 20154
rect 25996 20102 26048 20154
rect 3884 20000 3936 20052
rect 3976 20000 4028 20052
rect 6644 20000 6696 20052
rect 8208 20000 8260 20052
rect 9680 20000 9732 20052
rect 12072 20000 12124 20052
rect 14280 20000 14332 20052
rect 16856 20000 16908 20052
rect 16948 20000 17000 20052
rect 17040 20000 17092 20052
rect 21088 20000 21140 20052
rect 28080 20000 28132 20052
rect 7564 19932 7616 19984
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 3424 19728 3476 19780
rect 6460 19796 6512 19848
rect 6828 19796 6880 19848
rect 6920 19796 6972 19848
rect 7196 19839 7248 19848
rect 7196 19805 7203 19839
rect 7203 19805 7248 19839
rect 7196 19796 7248 19805
rect 9404 19864 9456 19916
rect 10508 19907 10560 19916
rect 10508 19873 10517 19907
rect 10517 19873 10551 19907
rect 10551 19873 10560 19907
rect 10508 19864 10560 19873
rect 8852 19796 8904 19848
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 10232 19839 10284 19848
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 11336 19864 11388 19916
rect 17868 19932 17920 19984
rect 6552 19771 6604 19780
rect 6552 19737 6561 19771
rect 6561 19737 6595 19771
rect 6595 19737 6604 19771
rect 6552 19728 6604 19737
rect 7288 19771 7340 19780
rect 7288 19737 7297 19771
rect 7297 19737 7331 19771
rect 7331 19737 7340 19771
rect 7288 19728 7340 19737
rect 10324 19728 10376 19780
rect 9588 19703 9640 19712
rect 9588 19669 9597 19703
rect 9597 19669 9631 19703
rect 9631 19669 9640 19703
rect 9588 19660 9640 19669
rect 10876 19771 10928 19780
rect 10876 19737 10885 19771
rect 10885 19737 10919 19771
rect 10919 19737 10928 19771
rect 10876 19728 10928 19737
rect 12716 19796 12768 19848
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 13176 19796 13228 19848
rect 14740 19796 14792 19848
rect 15108 19796 15160 19848
rect 18236 19864 18288 19916
rect 16856 19796 16908 19848
rect 19708 19796 19760 19848
rect 20168 19796 20220 19848
rect 27252 19839 27304 19848
rect 27252 19805 27261 19839
rect 27261 19805 27295 19839
rect 27295 19805 27304 19839
rect 27252 19796 27304 19805
rect 27344 19796 27396 19848
rect 27528 19839 27580 19848
rect 11060 19660 11112 19712
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 11336 19660 11388 19712
rect 12532 19728 12584 19780
rect 14648 19728 14700 19780
rect 15844 19728 15896 19780
rect 17592 19728 17644 19780
rect 19248 19728 19300 19780
rect 25044 19728 25096 19780
rect 27528 19805 27537 19839
rect 27537 19805 27571 19839
rect 27571 19805 27580 19839
rect 27528 19796 27580 19805
rect 27988 19796 28040 19848
rect 28172 19796 28224 19848
rect 12624 19660 12676 19712
rect 12900 19660 12952 19712
rect 19892 19660 19944 19712
rect 19984 19660 20036 19712
rect 26332 19660 26384 19712
rect 27068 19703 27120 19712
rect 27068 19669 27077 19703
rect 27077 19669 27111 19703
rect 27111 19669 27120 19703
rect 27068 19660 27120 19669
rect 27620 19660 27672 19712
rect 28724 19660 28776 19712
rect 5151 19558 5203 19610
rect 5215 19558 5267 19610
rect 5279 19558 5331 19610
rect 5343 19558 5395 19610
rect 5407 19558 5459 19610
rect 12234 19558 12286 19610
rect 12298 19558 12350 19610
rect 12362 19558 12414 19610
rect 12426 19558 12478 19610
rect 12490 19558 12542 19610
rect 19317 19558 19369 19610
rect 19381 19558 19433 19610
rect 19445 19558 19497 19610
rect 19509 19558 19561 19610
rect 19573 19558 19625 19610
rect 26400 19558 26452 19610
rect 26464 19558 26516 19610
rect 26528 19558 26580 19610
rect 26592 19558 26644 19610
rect 26656 19558 26708 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 1492 19363 1544 19372
rect 1492 19329 1501 19363
rect 1501 19329 1535 19363
rect 1535 19329 1544 19363
rect 1492 19320 1544 19329
rect 9588 19456 9640 19508
rect 11060 19456 11112 19508
rect 8116 19388 8168 19440
rect 8484 19388 8536 19440
rect 9772 19388 9824 19440
rect 10876 19388 10928 19440
rect 13084 19456 13136 19508
rect 13268 19456 13320 19508
rect 14556 19456 14608 19508
rect 14924 19456 14976 19508
rect 6552 19252 6604 19304
rect 7656 19363 7708 19372
rect 7656 19329 7665 19363
rect 7665 19329 7699 19363
rect 7699 19329 7708 19363
rect 7656 19320 7708 19329
rect 7932 19363 7984 19372
rect 7932 19329 7941 19363
rect 7941 19329 7975 19363
rect 7975 19329 7984 19363
rect 7932 19320 7984 19329
rect 9864 19320 9916 19372
rect 7564 19252 7616 19304
rect 8852 19252 8904 19304
rect 9220 19252 9272 19304
rect 12164 19252 12216 19304
rect 12900 19320 12952 19372
rect 13176 19363 13228 19372
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 15108 19431 15160 19440
rect 15108 19397 15117 19431
rect 15117 19397 15151 19431
rect 15151 19397 15160 19431
rect 15108 19388 15160 19397
rect 15476 19456 15528 19508
rect 4988 19184 5040 19236
rect 6460 19184 6512 19236
rect 7840 19159 7892 19168
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 9588 19184 9640 19236
rect 13820 19184 13872 19236
rect 16028 19320 16080 19372
rect 16856 19456 16908 19508
rect 17224 19499 17276 19508
rect 17224 19465 17233 19499
rect 17233 19465 17267 19499
rect 17267 19465 17276 19499
rect 17224 19456 17276 19465
rect 17960 19456 18012 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 19984 19456 20036 19508
rect 20536 19499 20588 19508
rect 20536 19465 20545 19499
rect 20545 19465 20579 19499
rect 20579 19465 20588 19499
rect 20536 19456 20588 19465
rect 28080 19456 28132 19508
rect 19432 19388 19484 19440
rect 19524 19431 19576 19440
rect 19524 19397 19533 19431
rect 19533 19397 19567 19431
rect 19567 19397 19576 19431
rect 19524 19388 19576 19397
rect 19892 19388 19944 19440
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 19340 19363 19392 19372
rect 19340 19329 19349 19363
rect 19349 19329 19383 19363
rect 19383 19329 19392 19363
rect 19340 19320 19392 19329
rect 20076 19388 20128 19440
rect 20168 19431 20220 19440
rect 20168 19397 20177 19431
rect 20177 19397 20211 19431
rect 20211 19397 20220 19431
rect 20168 19388 20220 19397
rect 22652 19388 22704 19440
rect 14188 19116 14240 19168
rect 15384 19116 15436 19168
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 19616 19184 19668 19236
rect 27436 19320 27488 19372
rect 20812 19252 20864 19304
rect 27804 19295 27856 19304
rect 27804 19261 27813 19295
rect 27813 19261 27847 19295
rect 27847 19261 27856 19295
rect 27804 19252 27856 19261
rect 20352 19184 20404 19236
rect 19340 19116 19392 19168
rect 4491 19014 4543 19066
rect 4555 19014 4607 19066
rect 4619 19014 4671 19066
rect 4683 19014 4735 19066
rect 4747 19014 4799 19066
rect 11574 19014 11626 19066
rect 11638 19014 11690 19066
rect 11702 19014 11754 19066
rect 11766 19014 11818 19066
rect 11830 19014 11882 19066
rect 18657 19014 18709 19066
rect 18721 19014 18773 19066
rect 18785 19014 18837 19066
rect 18849 19014 18901 19066
rect 18913 19014 18965 19066
rect 25740 19014 25792 19066
rect 25804 19014 25856 19066
rect 25868 19014 25920 19066
rect 25932 19014 25984 19066
rect 25996 19014 26048 19066
rect 7012 18912 7064 18964
rect 3608 18708 3660 18760
rect 6552 18844 6604 18896
rect 8944 18912 8996 18964
rect 9588 18955 9640 18964
rect 9588 18921 9597 18955
rect 9597 18921 9631 18955
rect 9631 18921 9640 18955
rect 9588 18912 9640 18921
rect 12164 18912 12216 18964
rect 15476 18912 15528 18964
rect 15844 18912 15896 18964
rect 16028 18912 16080 18964
rect 17776 18912 17828 18964
rect 19432 18912 19484 18964
rect 20260 18955 20312 18964
rect 20260 18921 20269 18955
rect 20269 18921 20303 18955
rect 20303 18921 20312 18955
rect 20260 18912 20312 18921
rect 21272 18912 21324 18964
rect 6368 18776 6420 18828
rect 7840 18776 7892 18828
rect 9220 18776 9272 18828
rect 6276 18640 6328 18692
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 6920 18708 6972 18760
rect 8576 18708 8628 18760
rect 9036 18751 9088 18760
rect 9036 18717 9046 18751
rect 9046 18717 9080 18751
rect 9080 18717 9088 18751
rect 9036 18708 9088 18717
rect 9404 18751 9456 18760
rect 9404 18717 9418 18751
rect 9418 18717 9452 18751
rect 9452 18717 9456 18751
rect 9404 18708 9456 18717
rect 7380 18640 7432 18692
rect 3976 18572 4028 18624
rect 5540 18572 5592 18624
rect 5816 18572 5868 18624
rect 7288 18572 7340 18624
rect 8208 18572 8260 18624
rect 9956 18776 10008 18828
rect 11152 18776 11204 18828
rect 12808 18844 12860 18896
rect 13084 18844 13136 18896
rect 11612 18776 11664 18828
rect 10416 18640 10468 18692
rect 10692 18640 10744 18692
rect 11152 18572 11204 18624
rect 12532 18776 12584 18828
rect 12900 18776 12952 18828
rect 13728 18776 13780 18828
rect 15568 18844 15620 18896
rect 18420 18844 18472 18896
rect 19340 18844 19392 18896
rect 12716 18708 12768 18760
rect 14096 18640 14148 18692
rect 14372 18640 14424 18692
rect 15476 18640 15528 18692
rect 12716 18572 12768 18624
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 12808 18572 12860 18581
rect 14648 18572 14700 18624
rect 16028 18751 16080 18760
rect 16028 18717 16037 18751
rect 16037 18717 16071 18751
rect 16071 18717 16080 18751
rect 16028 18708 16080 18717
rect 16396 18708 16448 18760
rect 17316 18708 17368 18760
rect 17776 18751 17828 18760
rect 17776 18717 17785 18751
rect 17785 18717 17819 18751
rect 17819 18717 17828 18751
rect 17776 18708 17828 18717
rect 18788 18708 18840 18760
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 15844 18572 15896 18624
rect 17500 18572 17552 18624
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 23296 18708 23348 18760
rect 27712 18708 27764 18760
rect 20076 18683 20128 18692
rect 20076 18649 20085 18683
rect 20085 18649 20119 18683
rect 20119 18649 20128 18683
rect 20076 18640 20128 18649
rect 19892 18572 19944 18624
rect 29000 18615 29052 18624
rect 29000 18581 29009 18615
rect 29009 18581 29043 18615
rect 29043 18581 29052 18615
rect 29000 18572 29052 18581
rect 5151 18470 5203 18522
rect 5215 18470 5267 18522
rect 5279 18470 5331 18522
rect 5343 18470 5395 18522
rect 5407 18470 5459 18522
rect 12234 18470 12286 18522
rect 12298 18470 12350 18522
rect 12362 18470 12414 18522
rect 12426 18470 12478 18522
rect 12490 18470 12542 18522
rect 19317 18470 19369 18522
rect 19381 18470 19433 18522
rect 19445 18470 19497 18522
rect 19509 18470 19561 18522
rect 19573 18470 19625 18522
rect 26400 18470 26452 18522
rect 26464 18470 26516 18522
rect 26528 18470 26580 18522
rect 26592 18470 26644 18522
rect 26656 18470 26708 18522
rect 1860 18368 1912 18420
rect 3700 18368 3752 18420
rect 3424 18300 3476 18352
rect 5540 18300 5592 18352
rect 6276 18368 6328 18420
rect 9864 18368 9916 18420
rect 12072 18368 12124 18420
rect 12624 18368 12676 18420
rect 12716 18368 12768 18420
rect 14372 18368 14424 18420
rect 7380 18300 7432 18352
rect 3608 18232 3660 18284
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 3424 18164 3476 18216
rect 5080 18096 5132 18148
rect 5172 18028 5224 18080
rect 6552 18232 6604 18284
rect 6644 18232 6696 18284
rect 6184 18164 6236 18216
rect 6920 18232 6972 18284
rect 7840 18232 7892 18284
rect 7012 18164 7064 18216
rect 7564 18164 7616 18216
rect 7932 18164 7984 18216
rect 6000 18096 6052 18148
rect 9128 18096 9180 18148
rect 9772 18275 9824 18284
rect 9772 18241 9781 18275
rect 9781 18241 9815 18275
rect 9815 18241 9824 18275
rect 9772 18232 9824 18241
rect 9864 18232 9916 18284
rect 13912 18300 13964 18352
rect 14648 18300 14700 18352
rect 10140 18232 10192 18284
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 11612 18232 11664 18284
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 11244 18164 11296 18216
rect 11336 18164 11388 18216
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 13360 18232 13412 18284
rect 13820 18164 13872 18216
rect 10324 18096 10376 18148
rect 16580 18368 16632 18420
rect 15476 18300 15528 18352
rect 17960 18368 18012 18420
rect 18052 18368 18104 18420
rect 18788 18411 18840 18420
rect 18788 18377 18797 18411
rect 18797 18377 18831 18411
rect 18831 18377 18840 18411
rect 18788 18368 18840 18377
rect 19616 18368 19668 18420
rect 19800 18368 19852 18420
rect 19892 18368 19944 18420
rect 25320 18368 25372 18420
rect 15476 18164 15528 18216
rect 15568 18164 15620 18216
rect 18052 18164 18104 18216
rect 19064 18232 19116 18284
rect 19432 18275 19484 18284
rect 19432 18241 19441 18275
rect 19441 18241 19475 18275
rect 19475 18241 19484 18275
rect 19432 18232 19484 18241
rect 19800 18275 19852 18284
rect 19800 18241 19809 18275
rect 19809 18241 19843 18275
rect 19843 18241 19852 18275
rect 19800 18232 19852 18241
rect 18512 18164 18564 18216
rect 19248 18207 19300 18216
rect 19248 18173 19257 18207
rect 19257 18173 19291 18207
rect 19291 18173 19300 18207
rect 19248 18164 19300 18173
rect 20720 18275 20772 18284
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 20812 18275 20864 18284
rect 20812 18241 20826 18275
rect 20826 18241 20860 18275
rect 20860 18241 20864 18275
rect 20812 18232 20864 18241
rect 21272 18232 21324 18284
rect 23480 18300 23532 18352
rect 24492 18300 24544 18352
rect 24952 18300 25004 18352
rect 27988 18300 28040 18352
rect 7656 18028 7708 18080
rect 9864 18028 9916 18080
rect 10140 18028 10192 18080
rect 11152 18028 11204 18080
rect 16764 18096 16816 18148
rect 18328 18096 18380 18148
rect 23204 18207 23256 18216
rect 23204 18173 23213 18207
rect 23213 18173 23247 18207
rect 23247 18173 23256 18207
rect 23204 18164 23256 18173
rect 20904 18096 20956 18148
rect 16120 18028 16172 18080
rect 22652 18028 22704 18080
rect 25504 18164 25556 18216
rect 26148 18164 26200 18216
rect 26884 18164 26936 18216
rect 27252 18207 27304 18216
rect 27252 18173 27261 18207
rect 27261 18173 27295 18207
rect 27295 18173 27304 18207
rect 27252 18164 27304 18173
rect 28448 18164 28500 18216
rect 24860 18028 24912 18080
rect 26608 18028 26660 18080
rect 26976 18028 27028 18080
rect 4491 17926 4543 17978
rect 4555 17926 4607 17978
rect 4619 17926 4671 17978
rect 4683 17926 4735 17978
rect 4747 17926 4799 17978
rect 11574 17926 11626 17978
rect 11638 17926 11690 17978
rect 11702 17926 11754 17978
rect 11766 17926 11818 17978
rect 11830 17926 11882 17978
rect 18657 17926 18709 17978
rect 18721 17926 18773 17978
rect 18785 17926 18837 17978
rect 18849 17926 18901 17978
rect 18913 17926 18965 17978
rect 25740 17926 25792 17978
rect 25804 17926 25856 17978
rect 25868 17926 25920 17978
rect 25932 17926 25984 17978
rect 25996 17926 26048 17978
rect 7380 17824 7432 17876
rect 10600 17824 10652 17876
rect 3700 17688 3752 17740
rect 5172 17620 5224 17672
rect 11336 17799 11388 17808
rect 11336 17765 11345 17799
rect 11345 17765 11379 17799
rect 11379 17765 11388 17799
rect 11336 17756 11388 17765
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 9956 17688 10008 17740
rect 3424 17552 3476 17604
rect 4528 17552 4580 17604
rect 5816 17552 5868 17604
rect 7104 17595 7156 17604
rect 7104 17561 7113 17595
rect 7113 17561 7147 17595
rect 7147 17561 7156 17595
rect 7104 17552 7156 17561
rect 4804 17484 4856 17536
rect 6368 17484 6420 17536
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 7932 17620 7984 17672
rect 10876 17620 10928 17672
rect 10140 17552 10192 17604
rect 10876 17484 10928 17536
rect 11244 17620 11296 17672
rect 11428 17663 11480 17672
rect 11428 17629 11437 17663
rect 11437 17629 11471 17663
rect 11471 17629 11480 17663
rect 11428 17620 11480 17629
rect 11980 17824 12032 17876
rect 12624 17824 12676 17876
rect 13912 17867 13964 17876
rect 13912 17833 13921 17867
rect 13921 17833 13955 17867
rect 13955 17833 13964 17867
rect 13912 17824 13964 17833
rect 15936 17824 15988 17876
rect 15108 17756 15160 17808
rect 19616 17824 19668 17876
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 23204 17824 23256 17876
rect 22744 17756 22796 17808
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 20076 17731 20128 17740
rect 20076 17697 20085 17731
rect 20085 17697 20119 17731
rect 20119 17697 20128 17731
rect 20076 17688 20128 17697
rect 20352 17731 20404 17740
rect 20352 17697 20361 17731
rect 20361 17697 20395 17731
rect 20395 17697 20404 17731
rect 20352 17688 20404 17697
rect 20720 17688 20772 17740
rect 22008 17688 22060 17740
rect 13084 17552 13136 17604
rect 14188 17595 14240 17604
rect 14188 17561 14197 17595
rect 14197 17561 14231 17595
rect 14231 17561 14240 17595
rect 14188 17552 14240 17561
rect 17592 17595 17644 17604
rect 17592 17561 17601 17595
rect 17601 17561 17635 17595
rect 17635 17561 17644 17595
rect 17592 17552 17644 17561
rect 18052 17552 18104 17604
rect 14648 17484 14700 17536
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 17132 17484 17184 17536
rect 17868 17484 17920 17536
rect 18420 17484 18472 17536
rect 19524 17663 19576 17672
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 19708 17620 19760 17672
rect 19800 17620 19852 17672
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 22652 17620 22704 17672
rect 23296 17620 23348 17672
rect 23756 17688 23808 17740
rect 24860 17688 24912 17740
rect 25964 17824 26016 17876
rect 26240 17756 26292 17808
rect 24400 17663 24452 17672
rect 24400 17629 24409 17663
rect 24409 17629 24443 17663
rect 24443 17629 24452 17663
rect 24400 17620 24452 17629
rect 26056 17731 26108 17740
rect 26056 17697 26065 17731
rect 26065 17697 26099 17731
rect 26099 17697 26108 17731
rect 26056 17688 26108 17697
rect 26148 17731 26200 17740
rect 26148 17697 26157 17731
rect 26157 17697 26191 17731
rect 26191 17697 26200 17731
rect 26148 17688 26200 17697
rect 26424 17688 26476 17740
rect 26516 17731 26568 17740
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 26516 17688 26568 17697
rect 18972 17552 19024 17604
rect 23572 17595 23624 17604
rect 23572 17561 23581 17595
rect 23581 17561 23615 17595
rect 23615 17561 23624 17595
rect 23572 17552 23624 17561
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 23112 17484 23164 17536
rect 24032 17552 24084 17604
rect 25320 17641 25372 17650
rect 25320 17607 25330 17641
rect 25330 17607 25364 17641
rect 25364 17607 25372 17641
rect 25320 17598 25372 17607
rect 25412 17595 25464 17604
rect 25412 17561 25421 17595
rect 25421 17561 25455 17595
rect 25455 17561 25464 17595
rect 25412 17552 25464 17561
rect 25964 17620 26016 17672
rect 26608 17663 26660 17672
rect 26608 17629 26617 17663
rect 26617 17629 26651 17663
rect 26651 17629 26660 17663
rect 26608 17620 26660 17629
rect 27252 17824 27304 17876
rect 27344 17756 27396 17808
rect 27528 17620 27580 17672
rect 27896 17663 27948 17672
rect 27896 17629 27905 17663
rect 27905 17629 27939 17663
rect 27939 17629 27948 17663
rect 27896 17620 27948 17629
rect 25136 17527 25188 17536
rect 25136 17493 25145 17527
rect 25145 17493 25179 17527
rect 25179 17493 25188 17527
rect 25136 17484 25188 17493
rect 25228 17484 25280 17536
rect 27160 17552 27212 17604
rect 25596 17484 25648 17536
rect 26148 17484 26200 17536
rect 26516 17484 26568 17536
rect 27620 17484 27672 17536
rect 28448 17552 28500 17604
rect 28080 17484 28132 17536
rect 28356 17484 28408 17536
rect 5151 17382 5203 17434
rect 5215 17382 5267 17434
rect 5279 17382 5331 17434
rect 5343 17382 5395 17434
rect 5407 17382 5459 17434
rect 12234 17382 12286 17434
rect 12298 17382 12350 17434
rect 12362 17382 12414 17434
rect 12426 17382 12478 17434
rect 12490 17382 12542 17434
rect 19317 17382 19369 17434
rect 19381 17382 19433 17434
rect 19445 17382 19497 17434
rect 19509 17382 19561 17434
rect 19573 17382 19625 17434
rect 26400 17382 26452 17434
rect 26464 17382 26516 17434
rect 26528 17382 26580 17434
rect 26592 17382 26644 17434
rect 26656 17382 26708 17434
rect 3240 17212 3292 17264
rect 3424 17076 3476 17128
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 4068 17280 4120 17332
rect 4528 17323 4580 17332
rect 4528 17289 4537 17323
rect 4537 17289 4571 17323
rect 4571 17289 4580 17323
rect 4528 17280 4580 17289
rect 4988 17280 5040 17332
rect 5080 17280 5132 17332
rect 5264 17280 5316 17332
rect 3976 17187 4028 17196
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 3976 17008 4028 17060
rect 5172 17144 5224 17196
rect 6000 17212 6052 17264
rect 9956 17280 10008 17332
rect 5540 17187 5592 17196
rect 5540 17153 5545 17187
rect 5545 17153 5579 17187
rect 5579 17153 5592 17187
rect 5540 17144 5592 17153
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 4804 17076 4856 17128
rect 7380 17144 7432 17196
rect 10876 17144 10928 17196
rect 12808 17280 12860 17332
rect 13820 17280 13872 17332
rect 9864 17119 9916 17128
rect 9864 17085 9873 17119
rect 9873 17085 9907 17119
rect 9907 17085 9916 17119
rect 9864 17076 9916 17085
rect 13084 17076 13136 17128
rect 13912 17144 13964 17196
rect 16672 17280 16724 17332
rect 16764 17280 16816 17332
rect 15108 17212 15160 17264
rect 15752 17212 15804 17264
rect 16120 17212 16172 17264
rect 14096 17076 14148 17128
rect 14372 17076 14424 17128
rect 11244 17008 11296 17060
rect 3332 16940 3384 16992
rect 4068 16940 4120 16992
rect 5816 16983 5868 16992
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 6000 16940 6052 16992
rect 6184 16940 6236 16992
rect 14096 16940 14148 16992
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 17592 17280 17644 17332
rect 19064 17280 19116 17332
rect 19248 17323 19300 17332
rect 19248 17289 19257 17323
rect 19257 17289 19291 17323
rect 19291 17289 19300 17323
rect 19248 17280 19300 17289
rect 20352 17280 20404 17332
rect 19156 17212 19208 17264
rect 23572 17280 23624 17332
rect 18328 17144 18380 17196
rect 15476 17076 15528 17128
rect 17500 17008 17552 17060
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 22008 17212 22060 17264
rect 25136 17280 25188 17332
rect 25412 17280 25464 17332
rect 26056 17280 26108 17332
rect 26148 17280 26200 17332
rect 26424 17280 26476 17332
rect 25044 17212 25096 17264
rect 16120 16940 16172 16992
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 22836 17187 22888 17196
rect 22836 17153 22845 17187
rect 22845 17153 22879 17187
rect 22879 17153 22888 17187
rect 22836 17144 22888 17153
rect 22376 17076 22428 17128
rect 22284 17008 22336 17060
rect 23204 17076 23256 17128
rect 23480 17119 23532 17128
rect 23480 17085 23489 17119
rect 23489 17085 23523 17119
rect 23523 17085 23532 17119
rect 23480 17076 23532 17085
rect 25412 17187 25464 17196
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 25504 17144 25556 17196
rect 24952 17076 25004 17128
rect 27896 17280 27948 17332
rect 27528 17212 27580 17264
rect 27712 17212 27764 17264
rect 26516 17144 26568 17196
rect 26700 17144 26752 17196
rect 27804 17144 27856 17196
rect 27896 17187 27948 17196
rect 27896 17153 27905 17187
rect 27905 17153 27939 17187
rect 27939 17153 27948 17187
rect 28448 17187 28500 17196
rect 27896 17144 27948 17153
rect 28448 17153 28457 17187
rect 28457 17153 28491 17187
rect 28491 17153 28500 17187
rect 28448 17144 28500 17153
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 23572 16940 23624 16992
rect 24400 16940 24452 16992
rect 27252 17119 27304 17128
rect 27252 17085 27261 17119
rect 27261 17085 27295 17119
rect 27295 17085 27304 17119
rect 27252 17076 27304 17085
rect 26516 17008 26568 17060
rect 26976 17051 27028 17060
rect 26976 17017 26985 17051
rect 26985 17017 27019 17051
rect 27019 17017 27028 17051
rect 26976 17008 27028 17017
rect 27436 17119 27488 17128
rect 27436 17085 27445 17119
rect 27445 17085 27479 17119
rect 27479 17085 27488 17119
rect 27436 17076 27488 17085
rect 27528 17076 27580 17128
rect 28356 17076 28408 17128
rect 26332 16940 26384 16992
rect 26608 16940 26660 16992
rect 27252 16940 27304 16992
rect 28632 16983 28684 16992
rect 28632 16949 28641 16983
rect 28641 16949 28675 16983
rect 28675 16949 28684 16983
rect 28632 16940 28684 16949
rect 4491 16838 4543 16890
rect 4555 16838 4607 16890
rect 4619 16838 4671 16890
rect 4683 16838 4735 16890
rect 4747 16838 4799 16890
rect 11574 16838 11626 16890
rect 11638 16838 11690 16890
rect 11702 16838 11754 16890
rect 11766 16838 11818 16890
rect 11830 16838 11882 16890
rect 18657 16838 18709 16890
rect 18721 16838 18773 16890
rect 18785 16838 18837 16890
rect 18849 16838 18901 16890
rect 18913 16838 18965 16890
rect 25740 16838 25792 16890
rect 25804 16838 25856 16890
rect 25868 16838 25920 16890
rect 25932 16838 25984 16890
rect 25996 16838 26048 16890
rect 3608 16736 3660 16788
rect 5172 16736 5224 16788
rect 5540 16736 5592 16788
rect 14648 16779 14700 16788
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 16948 16736 17000 16788
rect 19156 16736 19208 16788
rect 22192 16736 22244 16788
rect 22284 16736 22336 16788
rect 22652 16736 22704 16788
rect 3424 16668 3476 16720
rect 4988 16668 5040 16720
rect 7196 16668 7248 16720
rect 10508 16668 10560 16720
rect 16856 16668 16908 16720
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 4896 16532 4948 16584
rect 1676 16507 1728 16516
rect 1676 16473 1685 16507
rect 1685 16473 1719 16507
rect 1719 16473 1728 16507
rect 1676 16464 1728 16473
rect 3884 16464 3936 16516
rect 4436 16439 4488 16448
rect 4436 16405 4445 16439
rect 4445 16405 4479 16439
rect 4479 16405 4488 16439
rect 4436 16396 4488 16405
rect 5080 16532 5132 16584
rect 9772 16600 9824 16652
rect 10140 16600 10192 16652
rect 10968 16600 11020 16652
rect 22836 16736 22888 16788
rect 23388 16736 23440 16788
rect 23848 16736 23900 16788
rect 25320 16736 25372 16788
rect 26240 16736 26292 16788
rect 26516 16736 26568 16788
rect 27160 16736 27212 16788
rect 27804 16779 27856 16788
rect 27804 16745 27813 16779
rect 27813 16745 27847 16779
rect 27847 16745 27856 16779
rect 27804 16736 27856 16745
rect 23296 16711 23348 16720
rect 23296 16677 23305 16711
rect 23305 16677 23339 16711
rect 23339 16677 23348 16711
rect 23296 16668 23348 16677
rect 5724 16575 5776 16584
rect 5724 16541 5733 16575
rect 5733 16541 5767 16575
rect 5767 16541 5776 16575
rect 5724 16532 5776 16541
rect 7472 16532 7524 16584
rect 9956 16532 10008 16584
rect 14096 16575 14148 16584
rect 14096 16541 14105 16575
rect 14105 16541 14139 16575
rect 14139 16541 14148 16575
rect 14096 16532 14148 16541
rect 5080 16396 5132 16448
rect 5540 16439 5592 16448
rect 5540 16405 5549 16439
rect 5549 16405 5583 16439
rect 5583 16405 5592 16439
rect 5540 16396 5592 16405
rect 14372 16507 14424 16516
rect 14372 16473 14381 16507
rect 14381 16473 14415 16507
rect 14415 16473 14424 16507
rect 14372 16464 14424 16473
rect 10324 16396 10376 16448
rect 10416 16439 10468 16448
rect 10416 16405 10425 16439
rect 10425 16405 10459 16439
rect 10459 16405 10468 16439
rect 10416 16396 10468 16405
rect 12164 16396 12216 16448
rect 14740 16532 14792 16584
rect 14924 16532 14976 16584
rect 22008 16600 22060 16652
rect 15016 16464 15068 16516
rect 15476 16575 15528 16584
rect 15476 16541 15485 16575
rect 15485 16541 15519 16575
rect 15519 16541 15528 16575
rect 15476 16532 15528 16541
rect 22284 16532 22336 16584
rect 15660 16464 15712 16516
rect 17132 16464 17184 16516
rect 22744 16575 22796 16584
rect 22744 16541 22753 16575
rect 22753 16541 22787 16575
rect 22787 16541 22796 16575
rect 22744 16532 22796 16541
rect 15108 16396 15160 16448
rect 15292 16396 15344 16448
rect 23204 16439 23256 16448
rect 23204 16405 23213 16439
rect 23213 16405 23247 16439
rect 23247 16405 23256 16439
rect 23204 16396 23256 16405
rect 23388 16532 23440 16584
rect 23940 16532 23992 16584
rect 24676 16532 24728 16584
rect 25412 16600 25464 16652
rect 25596 16600 25648 16652
rect 26240 16600 26292 16652
rect 26792 16600 26844 16652
rect 23756 16464 23808 16516
rect 26424 16532 26476 16584
rect 26516 16575 26568 16584
rect 26516 16541 26525 16575
rect 26525 16541 26559 16575
rect 26559 16541 26568 16575
rect 26516 16532 26568 16541
rect 26792 16464 26844 16516
rect 27620 16575 27672 16584
rect 27620 16541 27629 16575
rect 27629 16541 27663 16575
rect 27663 16541 27672 16575
rect 27620 16532 27672 16541
rect 27160 16396 27212 16448
rect 27252 16439 27304 16448
rect 27252 16405 27261 16439
rect 27261 16405 27295 16439
rect 27295 16405 27304 16439
rect 27252 16396 27304 16405
rect 28080 16575 28132 16584
rect 28080 16541 28089 16575
rect 28089 16541 28123 16575
rect 28123 16541 28132 16575
rect 28080 16532 28132 16541
rect 28356 16575 28408 16584
rect 28356 16541 28373 16575
rect 28373 16541 28407 16575
rect 28407 16541 28408 16575
rect 28356 16532 28408 16541
rect 28632 16532 28684 16584
rect 5151 16294 5203 16346
rect 5215 16294 5267 16346
rect 5279 16294 5331 16346
rect 5343 16294 5395 16346
rect 5407 16294 5459 16346
rect 12234 16294 12286 16346
rect 12298 16294 12350 16346
rect 12362 16294 12414 16346
rect 12426 16294 12478 16346
rect 12490 16294 12542 16346
rect 19317 16294 19369 16346
rect 19381 16294 19433 16346
rect 19445 16294 19497 16346
rect 19509 16294 19561 16346
rect 19573 16294 19625 16346
rect 26400 16294 26452 16346
rect 26464 16294 26516 16346
rect 26528 16294 26580 16346
rect 26592 16294 26644 16346
rect 26656 16294 26708 16346
rect 1676 16192 1728 16244
rect 4436 16192 4488 16244
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 5080 16192 5132 16244
rect 7380 16192 7432 16244
rect 940 16056 992 16108
rect 3884 16056 3936 16108
rect 5172 16056 5224 16108
rect 5724 16056 5776 16108
rect 5908 16056 5960 16108
rect 6552 16124 6604 16176
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 1400 15988 1452 16040
rect 4344 15920 4396 15972
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 7012 16056 7064 16108
rect 9956 16192 10008 16244
rect 10048 16167 10100 16176
rect 10048 16133 10057 16167
rect 10057 16133 10091 16167
rect 10091 16133 10100 16167
rect 10048 16124 10100 16133
rect 11336 16192 11388 16244
rect 7196 16056 7248 16108
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 7932 16099 7984 16108
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 8116 16056 8168 16108
rect 9496 16056 9548 16108
rect 8300 15920 8352 15972
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 17960 16192 18012 16244
rect 22836 16192 22888 16244
rect 12900 16124 12952 16176
rect 14096 16124 14148 16176
rect 14924 16124 14976 16176
rect 23204 16124 23256 16176
rect 25412 16124 25464 16176
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 13176 16099 13228 16108
rect 13176 16065 13185 16099
rect 13185 16065 13219 16099
rect 13219 16065 13228 16099
rect 13176 16056 13228 16065
rect 13452 16056 13504 16108
rect 13912 16056 13964 16108
rect 15844 16056 15896 16108
rect 16120 16099 16172 16108
rect 16120 16065 16129 16099
rect 16129 16065 16163 16099
rect 16163 16065 16172 16099
rect 16120 16056 16172 16065
rect 17040 16056 17092 16108
rect 23940 16056 23992 16108
rect 10876 15988 10928 16040
rect 15292 15988 15344 16040
rect 26792 16192 26844 16244
rect 26332 16056 26384 16108
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 9956 15852 10008 15904
rect 23296 15920 23348 15972
rect 23664 15963 23716 15972
rect 23664 15929 23673 15963
rect 23673 15929 23707 15963
rect 23707 15929 23716 15963
rect 27528 15988 27580 16040
rect 23664 15920 23716 15929
rect 26240 15920 26292 15972
rect 26792 15920 26844 15972
rect 13820 15852 13872 15904
rect 15292 15852 15344 15904
rect 15660 15852 15712 15904
rect 16028 15852 16080 15904
rect 16120 15852 16172 15904
rect 16304 15895 16356 15904
rect 16304 15861 16313 15895
rect 16313 15861 16347 15895
rect 16347 15861 16356 15895
rect 16304 15852 16356 15861
rect 26148 15852 26200 15904
rect 4491 15750 4543 15802
rect 4555 15750 4607 15802
rect 4619 15750 4671 15802
rect 4683 15750 4735 15802
rect 4747 15750 4799 15802
rect 11574 15750 11626 15802
rect 11638 15750 11690 15802
rect 11702 15750 11754 15802
rect 11766 15750 11818 15802
rect 11830 15750 11882 15802
rect 18657 15750 18709 15802
rect 18721 15750 18773 15802
rect 18785 15750 18837 15802
rect 18849 15750 18901 15802
rect 18913 15750 18965 15802
rect 25740 15750 25792 15802
rect 25804 15750 25856 15802
rect 25868 15750 25920 15802
rect 25932 15750 25984 15802
rect 25996 15750 26048 15802
rect 4344 15648 4396 15700
rect 5724 15648 5776 15700
rect 5816 15580 5868 15632
rect 1400 15512 1452 15564
rect 3332 15512 3384 15564
rect 3240 15444 3292 15496
rect 3884 15444 3936 15496
rect 6092 15444 6144 15496
rect 7932 15648 7984 15700
rect 8668 15648 8720 15700
rect 9956 15648 10008 15700
rect 10876 15648 10928 15700
rect 15016 15648 15068 15700
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 16304 15648 16356 15700
rect 23572 15691 23624 15700
rect 23572 15657 23581 15691
rect 23581 15657 23615 15691
rect 23615 15657 23624 15691
rect 23572 15648 23624 15657
rect 24032 15648 24084 15700
rect 24952 15648 25004 15700
rect 26148 15648 26200 15700
rect 26700 15648 26752 15700
rect 27160 15648 27212 15700
rect 27620 15648 27672 15700
rect 7656 15512 7708 15564
rect 6552 15444 6604 15496
rect 8116 15512 8168 15564
rect 9496 15512 9548 15564
rect 10508 15512 10560 15564
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 10048 15376 10100 15428
rect 4160 15308 4212 15360
rect 5172 15308 5224 15360
rect 5816 15308 5868 15360
rect 7196 15308 7248 15360
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 12348 15512 12400 15564
rect 14372 15555 14424 15564
rect 14372 15521 14381 15555
rect 14381 15521 14415 15555
rect 14415 15521 14424 15555
rect 14372 15512 14424 15521
rect 19064 15580 19116 15632
rect 17408 15512 17460 15564
rect 17960 15512 18012 15564
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 11336 15376 11388 15428
rect 11796 15376 11848 15428
rect 11244 15308 11296 15360
rect 13912 15444 13964 15496
rect 18144 15444 18196 15496
rect 19800 15487 19852 15496
rect 19800 15453 19809 15487
rect 19809 15453 19843 15487
rect 19843 15453 19852 15487
rect 19800 15444 19852 15453
rect 23296 15580 23348 15632
rect 22284 15512 22336 15564
rect 12992 15376 13044 15428
rect 15660 15376 15712 15428
rect 16028 15376 16080 15428
rect 16856 15376 16908 15428
rect 17224 15376 17276 15428
rect 12624 15308 12676 15360
rect 13360 15308 13412 15360
rect 13544 15308 13596 15360
rect 18512 15376 18564 15428
rect 23204 15487 23256 15496
rect 23204 15453 23213 15487
rect 23213 15453 23247 15487
rect 23247 15453 23256 15487
rect 23204 15444 23256 15453
rect 24768 15580 24820 15632
rect 23756 15555 23808 15564
rect 23756 15521 23765 15555
rect 23765 15521 23799 15555
rect 23799 15521 23808 15555
rect 23756 15512 23808 15521
rect 24032 15555 24084 15564
rect 24032 15521 24041 15555
rect 24041 15521 24075 15555
rect 24075 15521 24084 15555
rect 24032 15512 24084 15521
rect 24676 15512 24728 15564
rect 27436 15580 27488 15632
rect 23940 15487 23992 15496
rect 23940 15453 23949 15487
rect 23949 15453 23983 15487
rect 23983 15453 23992 15487
rect 23940 15444 23992 15453
rect 18144 15308 18196 15360
rect 24216 15376 24268 15428
rect 19984 15308 20036 15360
rect 20076 15351 20128 15360
rect 20076 15317 20085 15351
rect 20085 15317 20119 15351
rect 20119 15317 20128 15351
rect 20076 15308 20128 15317
rect 24860 15376 24912 15428
rect 25228 15376 25280 15428
rect 27712 15512 27764 15564
rect 26700 15444 26752 15496
rect 26792 15487 26844 15496
rect 26792 15453 26801 15487
rect 26801 15453 26835 15487
rect 26835 15453 26844 15487
rect 26792 15444 26844 15453
rect 27252 15487 27304 15496
rect 27252 15453 27261 15487
rect 27261 15453 27295 15487
rect 27295 15453 27304 15487
rect 27252 15444 27304 15453
rect 27344 15444 27396 15496
rect 26332 15308 26384 15360
rect 27896 15376 27948 15428
rect 26608 15308 26660 15360
rect 26976 15308 27028 15360
rect 27252 15308 27304 15360
rect 5151 15206 5203 15258
rect 5215 15206 5267 15258
rect 5279 15206 5331 15258
rect 5343 15206 5395 15258
rect 5407 15206 5459 15258
rect 12234 15206 12286 15258
rect 12298 15206 12350 15258
rect 12362 15206 12414 15258
rect 12426 15206 12478 15258
rect 12490 15206 12542 15258
rect 19317 15206 19369 15258
rect 19381 15206 19433 15258
rect 19445 15206 19497 15258
rect 19509 15206 19561 15258
rect 19573 15206 19625 15258
rect 26400 15206 26452 15258
rect 26464 15206 26516 15258
rect 26528 15206 26580 15258
rect 26592 15206 26644 15258
rect 26656 15206 26708 15258
rect 1400 14900 1452 14952
rect 4160 15104 4212 15156
rect 5356 15104 5408 15156
rect 5632 15104 5684 15156
rect 8668 15104 8720 15156
rect 9404 15104 9456 15156
rect 8116 15036 8168 15088
rect 8208 15036 8260 15088
rect 5816 14968 5868 15020
rect 8300 14968 8352 15020
rect 10416 15104 10468 15156
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 11520 15104 11572 15156
rect 12164 15104 12216 15156
rect 10048 15036 10100 15088
rect 5540 14900 5592 14952
rect 6552 14943 6604 14952
rect 6552 14909 6561 14943
rect 6561 14909 6595 14943
rect 6595 14909 6604 14943
rect 6552 14900 6604 14909
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 8116 14764 8168 14816
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 12348 15036 12400 15088
rect 12624 15104 12676 15156
rect 12532 15036 12584 15088
rect 13912 15147 13964 15156
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 15476 15104 15528 15156
rect 15660 15104 15712 15156
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11520 14968 11572 14977
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 12072 14968 12124 15020
rect 13544 14968 13596 15020
rect 16028 15104 16080 15156
rect 16120 15104 16172 15156
rect 19984 15104 20036 15156
rect 16396 15036 16448 15088
rect 16028 14968 16080 15020
rect 16212 14968 16264 15020
rect 17408 15079 17460 15088
rect 17408 15045 17417 15079
rect 17417 15045 17451 15079
rect 17451 15045 17460 15079
rect 17408 15036 17460 15045
rect 18144 15036 18196 15088
rect 8576 14764 8628 14816
rect 12440 14900 12492 14952
rect 14372 14900 14424 14952
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 12624 14764 12676 14816
rect 15476 14900 15528 14952
rect 17224 14900 17276 14952
rect 14740 14764 14792 14816
rect 14832 14764 14884 14816
rect 17132 14832 17184 14884
rect 17960 14875 18012 14884
rect 17960 14841 17969 14875
rect 17969 14841 18003 14875
rect 18003 14841 18012 14875
rect 17960 14832 18012 14841
rect 19616 14968 19668 15020
rect 19800 14968 19852 15020
rect 20168 15036 20220 15088
rect 21180 14968 21232 15020
rect 25228 15104 25280 15156
rect 26240 15147 26292 15156
rect 26240 15113 26249 15147
rect 26249 15113 26283 15147
rect 26283 15113 26292 15147
rect 26240 15104 26292 15113
rect 24032 15079 24084 15088
rect 24032 15045 24041 15079
rect 24041 15045 24075 15079
rect 24075 15045 24084 15079
rect 24032 15036 24084 15045
rect 24676 15036 24728 15088
rect 24768 15079 24820 15088
rect 24768 15045 24777 15079
rect 24777 15045 24811 15079
rect 24811 15045 24820 15079
rect 24768 15036 24820 15045
rect 24860 15079 24912 15088
rect 24860 15045 24869 15079
rect 24869 15045 24903 15079
rect 24903 15045 24912 15079
rect 24860 15036 24912 15045
rect 24952 15079 25004 15088
rect 24952 15045 24987 15079
rect 24987 15045 25004 15079
rect 24952 15036 25004 15045
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 21548 14900 21600 14952
rect 22376 14968 22428 15020
rect 23204 14968 23256 15020
rect 23388 14968 23440 15020
rect 24860 14900 24912 14952
rect 25412 14943 25464 14952
rect 25412 14909 25421 14943
rect 25421 14909 25455 14943
rect 25455 14909 25464 14943
rect 25412 14900 25464 14909
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 16580 14764 16632 14816
rect 18144 14807 18196 14816
rect 18144 14773 18153 14807
rect 18153 14773 18187 14807
rect 18187 14773 18196 14807
rect 18144 14764 18196 14773
rect 19248 14807 19300 14816
rect 19248 14773 19257 14807
rect 19257 14773 19291 14807
rect 19291 14773 19300 14807
rect 19248 14764 19300 14773
rect 23848 14832 23900 14884
rect 26240 14968 26292 15020
rect 26976 15036 27028 15088
rect 27620 15104 27672 15156
rect 27252 14900 27304 14952
rect 27528 14900 27580 14952
rect 28356 15104 28408 15156
rect 28816 14968 28868 15020
rect 20720 14764 20772 14816
rect 24492 14807 24544 14816
rect 24492 14773 24501 14807
rect 24501 14773 24535 14807
rect 24535 14773 24544 14807
rect 24492 14764 24544 14773
rect 27068 14764 27120 14816
rect 27344 14764 27396 14816
rect 27712 14875 27764 14884
rect 27712 14841 27721 14875
rect 27721 14841 27755 14875
rect 27755 14841 27764 14875
rect 27712 14832 27764 14841
rect 4491 14662 4543 14714
rect 4555 14662 4607 14714
rect 4619 14662 4671 14714
rect 4683 14662 4735 14714
rect 4747 14662 4799 14714
rect 11574 14662 11626 14714
rect 11638 14662 11690 14714
rect 11702 14662 11754 14714
rect 11766 14662 11818 14714
rect 11830 14662 11882 14714
rect 18657 14662 18709 14714
rect 18721 14662 18773 14714
rect 18785 14662 18837 14714
rect 18849 14662 18901 14714
rect 18913 14662 18965 14714
rect 25740 14662 25792 14714
rect 25804 14662 25856 14714
rect 25868 14662 25920 14714
rect 25932 14662 25984 14714
rect 25996 14662 26048 14714
rect 6828 14560 6880 14612
rect 10416 14560 10468 14612
rect 11336 14560 11388 14612
rect 12072 14560 12124 14612
rect 13360 14603 13412 14612
rect 13360 14569 13369 14603
rect 13369 14569 13403 14603
rect 13403 14569 13412 14603
rect 13360 14560 13412 14569
rect 16120 14560 16172 14612
rect 16212 14560 16264 14612
rect 18144 14560 18196 14612
rect 19248 14560 19300 14612
rect 20168 14560 20220 14612
rect 20904 14560 20956 14612
rect 10508 14492 10560 14544
rect 10600 14492 10652 14544
rect 10876 14492 10928 14544
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 12440 14424 12492 14476
rect 14372 14424 14424 14476
rect 18512 14492 18564 14544
rect 18696 14492 18748 14544
rect 19064 14424 19116 14476
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 7840 14356 7892 14408
rect 9220 14356 9272 14408
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 7564 14288 7616 14340
rect 8576 14288 8628 14340
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 10876 14399 10928 14408
rect 10876 14365 10890 14399
rect 10890 14365 10924 14399
rect 10924 14365 10928 14399
rect 10876 14356 10928 14365
rect 14280 14356 14332 14408
rect 16028 14356 16080 14408
rect 16304 14356 16356 14408
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 20076 14424 20128 14476
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 19800 14356 19852 14408
rect 20168 14356 20220 14408
rect 20536 14356 20588 14408
rect 10692 14331 10744 14340
rect 10692 14297 10701 14331
rect 10701 14297 10735 14331
rect 10735 14297 10744 14331
rect 10692 14288 10744 14297
rect 13544 14288 13596 14340
rect 10968 14220 11020 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 11980 14220 12032 14272
rect 15568 14220 15620 14272
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 16764 14263 16816 14272
rect 16764 14229 16773 14263
rect 16773 14229 16807 14263
rect 16807 14229 16816 14263
rect 16764 14220 16816 14229
rect 18328 14263 18380 14272
rect 18328 14229 18337 14263
rect 18337 14229 18371 14263
rect 18371 14229 18380 14263
rect 18328 14220 18380 14229
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 19984 14331 20036 14340
rect 19984 14297 19993 14331
rect 19993 14297 20027 14331
rect 20027 14297 20036 14331
rect 19984 14288 20036 14297
rect 19616 14220 19668 14272
rect 19892 14220 19944 14272
rect 21088 14424 21140 14476
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 22284 14356 22336 14408
rect 22376 14399 22428 14408
rect 22376 14365 22385 14399
rect 22385 14365 22419 14399
rect 22419 14365 22428 14399
rect 22376 14356 22428 14365
rect 23388 14560 23440 14612
rect 23572 14603 23624 14612
rect 23572 14569 23581 14603
rect 23581 14569 23615 14603
rect 23615 14569 23624 14603
rect 23572 14560 23624 14569
rect 24492 14560 24544 14612
rect 26884 14560 26936 14612
rect 23848 14424 23900 14476
rect 24492 14467 24544 14476
rect 24492 14433 24501 14467
rect 24501 14433 24535 14467
rect 24535 14433 24544 14467
rect 24492 14424 24544 14433
rect 27068 14467 27120 14476
rect 27068 14433 27077 14467
rect 27077 14433 27111 14467
rect 27111 14433 27120 14467
rect 27068 14424 27120 14433
rect 28816 14467 28868 14476
rect 28816 14433 28825 14467
rect 28825 14433 28859 14467
rect 28859 14433 28868 14467
rect 28816 14424 28868 14433
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 22836 14356 22888 14408
rect 23664 14356 23716 14408
rect 25044 14288 25096 14340
rect 25320 14288 25372 14340
rect 22100 14220 22152 14272
rect 23940 14263 23992 14272
rect 23940 14229 23949 14263
rect 23949 14229 23983 14263
rect 23983 14229 23992 14263
rect 23940 14220 23992 14229
rect 25412 14220 25464 14272
rect 27528 14288 27580 14340
rect 5151 14118 5203 14170
rect 5215 14118 5267 14170
rect 5279 14118 5331 14170
rect 5343 14118 5395 14170
rect 5407 14118 5459 14170
rect 12234 14118 12286 14170
rect 12298 14118 12350 14170
rect 12362 14118 12414 14170
rect 12426 14118 12478 14170
rect 12490 14118 12542 14170
rect 19317 14118 19369 14170
rect 19381 14118 19433 14170
rect 19445 14118 19497 14170
rect 19509 14118 19561 14170
rect 19573 14118 19625 14170
rect 26400 14118 26452 14170
rect 26464 14118 26516 14170
rect 26528 14118 26580 14170
rect 26592 14118 26644 14170
rect 26656 14118 26708 14170
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 10324 14016 10376 14068
rect 10968 14016 11020 14068
rect 11060 14016 11112 14068
rect 13820 14016 13872 14068
rect 14372 14016 14424 14068
rect 3240 13948 3292 14000
rect 3608 13991 3660 14000
rect 3608 13957 3617 13991
rect 3617 13957 3651 13991
rect 3651 13957 3660 13991
rect 3608 13948 3660 13957
rect 1400 13880 1452 13932
rect 5632 13880 5684 13932
rect 9956 13880 10008 13932
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 5908 13812 5960 13864
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 6552 13744 6604 13796
rect 7288 13812 7340 13864
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 10508 13880 10560 13932
rect 7104 13744 7156 13796
rect 7196 13744 7248 13796
rect 10784 13855 10836 13864
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 14832 13880 14884 13932
rect 15660 14016 15712 14068
rect 18328 14016 18380 14068
rect 18420 14016 18472 14068
rect 19064 14016 19116 14068
rect 15568 13948 15620 14000
rect 6184 13676 6236 13728
rect 6368 13676 6420 13728
rect 10140 13676 10192 13728
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 11428 13744 11480 13796
rect 15108 13744 15160 13796
rect 11152 13676 11204 13728
rect 14096 13676 14148 13728
rect 17040 13880 17092 13932
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 19156 13948 19208 14000
rect 19708 13991 19760 14000
rect 19708 13957 19717 13991
rect 19717 13957 19751 13991
rect 19751 13957 19760 13991
rect 19708 13948 19760 13957
rect 19984 14016 20036 14068
rect 20628 14016 20680 14068
rect 22376 14016 22428 14068
rect 23388 14016 23440 14068
rect 27620 14016 27672 14068
rect 21456 13948 21508 14000
rect 21732 13948 21784 14000
rect 23572 13948 23624 14000
rect 24216 13948 24268 14000
rect 25044 13948 25096 14000
rect 25320 13948 25372 14000
rect 19524 13923 19576 13932
rect 19524 13889 19533 13923
rect 19533 13889 19567 13923
rect 19567 13889 19576 13923
rect 19524 13880 19576 13889
rect 20076 13880 20128 13932
rect 15476 13787 15528 13796
rect 15476 13753 15485 13787
rect 15485 13753 15519 13787
rect 15519 13753 15528 13787
rect 15476 13744 15528 13753
rect 16856 13744 16908 13796
rect 18144 13744 18196 13796
rect 20260 13855 20312 13864
rect 20260 13821 20269 13855
rect 20269 13821 20303 13855
rect 20303 13821 20312 13855
rect 20260 13812 20312 13821
rect 20720 13880 20772 13932
rect 23480 13923 23532 13932
rect 23480 13889 23489 13923
rect 23489 13889 23523 13923
rect 23523 13889 23532 13923
rect 24492 13923 24544 13932
rect 23480 13880 23532 13889
rect 24492 13889 24501 13923
rect 24501 13889 24535 13923
rect 24535 13889 24544 13923
rect 24492 13880 24544 13889
rect 27988 13923 28040 13932
rect 27988 13889 27997 13923
rect 27997 13889 28031 13923
rect 28031 13889 28040 13923
rect 27988 13880 28040 13889
rect 20996 13812 21048 13864
rect 22192 13812 22244 13864
rect 19800 13744 19852 13796
rect 21364 13787 21416 13796
rect 15752 13676 15804 13728
rect 18420 13719 18472 13728
rect 18420 13685 18429 13719
rect 18429 13685 18463 13719
rect 18463 13685 18472 13719
rect 18420 13676 18472 13685
rect 18880 13676 18932 13728
rect 21364 13753 21373 13787
rect 21373 13753 21407 13787
rect 21407 13753 21416 13787
rect 21364 13744 21416 13753
rect 24216 13812 24268 13864
rect 25320 13812 25372 13864
rect 27528 13812 27580 13864
rect 24952 13676 25004 13728
rect 4491 13574 4543 13626
rect 4555 13574 4607 13626
rect 4619 13574 4671 13626
rect 4683 13574 4735 13626
rect 4747 13574 4799 13626
rect 11574 13574 11626 13626
rect 11638 13574 11690 13626
rect 11702 13574 11754 13626
rect 11766 13574 11818 13626
rect 11830 13574 11882 13626
rect 18657 13574 18709 13626
rect 18721 13574 18773 13626
rect 18785 13574 18837 13626
rect 18849 13574 18901 13626
rect 18913 13574 18965 13626
rect 25740 13574 25792 13626
rect 25804 13574 25856 13626
rect 25868 13574 25920 13626
rect 25932 13574 25984 13626
rect 25996 13574 26048 13626
rect 1860 13472 1912 13524
rect 3608 13472 3660 13524
rect 6644 13472 6696 13524
rect 7196 13472 7248 13524
rect 13268 13472 13320 13524
rect 16948 13472 17000 13524
rect 18512 13472 18564 13524
rect 3056 13268 3108 13320
rect 9772 13404 9824 13456
rect 15292 13447 15344 13456
rect 15292 13413 15301 13447
rect 15301 13413 15335 13447
rect 15335 13413 15344 13447
rect 15292 13404 15344 13413
rect 17592 13404 17644 13456
rect 6920 13268 6972 13320
rect 7104 13268 7156 13320
rect 7196 13268 7248 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 8208 13268 8260 13320
rect 9404 13336 9456 13388
rect 13452 13336 13504 13388
rect 10324 13268 10376 13320
rect 10508 13311 10560 13320
rect 10508 13277 10518 13311
rect 10518 13277 10552 13311
rect 10552 13277 10560 13311
rect 10508 13268 10560 13277
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 10876 13311 10928 13320
rect 10876 13277 10890 13311
rect 10890 13277 10924 13311
rect 10924 13277 10928 13311
rect 10876 13268 10928 13277
rect 11428 13268 11480 13320
rect 11612 13268 11664 13320
rect 12164 13268 12216 13320
rect 12716 13268 12768 13320
rect 9864 13200 9916 13252
rect 10692 13243 10744 13252
rect 10692 13209 10701 13243
rect 10701 13209 10735 13243
rect 10735 13209 10744 13243
rect 10692 13200 10744 13209
rect 3240 13132 3292 13184
rect 7104 13175 7156 13184
rect 7104 13141 7113 13175
rect 7113 13141 7147 13175
rect 7147 13141 7156 13175
rect 7104 13132 7156 13141
rect 9404 13132 9456 13184
rect 10232 13132 10284 13184
rect 19524 13515 19576 13524
rect 19524 13481 19533 13515
rect 19533 13481 19567 13515
rect 19567 13481 19576 13515
rect 19524 13472 19576 13481
rect 20628 13472 20680 13524
rect 21364 13472 21416 13524
rect 24952 13472 25004 13524
rect 28908 13472 28960 13524
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 10968 13200 11020 13252
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 14464 13200 14516 13252
rect 15108 13200 15160 13252
rect 16488 13268 16540 13320
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17960 13268 18012 13320
rect 18144 13268 18196 13320
rect 16764 13200 16816 13252
rect 19248 13311 19300 13320
rect 19248 13277 19257 13311
rect 19257 13277 19291 13311
rect 19291 13277 19300 13311
rect 19248 13268 19300 13277
rect 19984 13268 20036 13320
rect 20260 13268 20312 13320
rect 22836 13404 22888 13456
rect 21456 13336 21508 13388
rect 22192 13336 22244 13388
rect 22652 13336 22704 13388
rect 25044 13336 25096 13388
rect 16580 13132 16632 13184
rect 19800 13132 19852 13184
rect 21824 13175 21876 13184
rect 21824 13141 21833 13175
rect 21833 13141 21867 13175
rect 21867 13141 21876 13175
rect 21824 13132 21876 13141
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 27620 13268 27672 13320
rect 23756 13132 23808 13184
rect 24032 13132 24084 13184
rect 5151 13030 5203 13082
rect 5215 13030 5267 13082
rect 5279 13030 5331 13082
rect 5343 13030 5395 13082
rect 5407 13030 5459 13082
rect 12234 13030 12286 13082
rect 12298 13030 12350 13082
rect 12362 13030 12414 13082
rect 12426 13030 12478 13082
rect 12490 13030 12542 13082
rect 19317 13030 19369 13082
rect 19381 13030 19433 13082
rect 19445 13030 19497 13082
rect 19509 13030 19561 13082
rect 19573 13030 19625 13082
rect 26400 13030 26452 13082
rect 26464 13030 26516 13082
rect 26528 13030 26580 13082
rect 26592 13030 26644 13082
rect 26656 13030 26708 13082
rect 1400 12792 1452 12844
rect 5172 12928 5224 12980
rect 3608 12860 3660 12912
rect 5540 12928 5592 12980
rect 7104 12928 7156 12980
rect 6736 12860 6788 12912
rect 10416 12928 10468 12980
rect 10784 12928 10836 12980
rect 11796 12928 11848 12980
rect 13268 12928 13320 12980
rect 3148 12792 3200 12844
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 4896 12792 4948 12844
rect 6368 12792 6420 12844
rect 6000 12656 6052 12708
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 10048 12860 10100 12912
rect 11428 12860 11480 12912
rect 15752 12928 15804 12980
rect 16488 12971 16540 12980
rect 16488 12937 16497 12971
rect 16497 12937 16531 12971
rect 16531 12937 16540 12971
rect 16488 12928 16540 12937
rect 17132 12928 17184 12980
rect 18420 12928 18472 12980
rect 21640 12928 21692 12980
rect 22284 12928 22336 12980
rect 10508 12792 10560 12844
rect 20720 12860 20772 12912
rect 22928 12860 22980 12912
rect 7288 12656 7340 12708
rect 7932 12724 7984 12776
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 10232 12724 10284 12776
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 12440 12792 12492 12801
rect 12716 12792 12768 12844
rect 13820 12792 13872 12844
rect 14372 12835 14424 12844
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14372 12792 14424 12801
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 16120 12792 16172 12844
rect 16580 12792 16632 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 17408 12792 17460 12844
rect 14556 12724 14608 12776
rect 14740 12767 14792 12776
rect 14740 12733 14749 12767
rect 14749 12733 14783 12767
rect 14783 12733 14792 12767
rect 14740 12724 14792 12733
rect 3884 12588 3936 12640
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 7012 12588 7064 12640
rect 10692 12656 10744 12708
rect 7932 12588 7984 12640
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 17132 12588 17184 12640
rect 19064 12588 19116 12640
rect 20536 12724 20588 12776
rect 21088 12792 21140 12844
rect 21824 12792 21876 12844
rect 21180 12724 21232 12776
rect 21732 12724 21784 12776
rect 22192 12724 22244 12776
rect 22744 12767 22796 12776
rect 22744 12733 22753 12767
rect 22753 12733 22787 12767
rect 22787 12733 22796 12767
rect 22744 12724 22796 12733
rect 22652 12656 22704 12708
rect 21640 12588 21692 12640
rect 23480 12588 23532 12640
rect 4491 12486 4543 12538
rect 4555 12486 4607 12538
rect 4619 12486 4671 12538
rect 4683 12486 4735 12538
rect 4747 12486 4799 12538
rect 11574 12486 11626 12538
rect 11638 12486 11690 12538
rect 11702 12486 11754 12538
rect 11766 12486 11818 12538
rect 11830 12486 11882 12538
rect 18657 12486 18709 12538
rect 18721 12486 18773 12538
rect 18785 12486 18837 12538
rect 18849 12486 18901 12538
rect 18913 12486 18965 12538
rect 25740 12486 25792 12538
rect 25804 12486 25856 12538
rect 25868 12486 25920 12538
rect 25932 12486 25984 12538
rect 25996 12486 26048 12538
rect 2044 12384 2096 12436
rect 4252 12316 4304 12368
rect 5908 12384 5960 12436
rect 6092 12384 6144 12436
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 3240 12180 3292 12232
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 6184 12248 6236 12300
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 5080 12180 5132 12232
rect 6920 12427 6972 12436
rect 6920 12393 6929 12427
rect 6929 12393 6963 12427
rect 6963 12393 6972 12427
rect 6920 12384 6972 12393
rect 7196 12384 7248 12436
rect 7564 12384 7616 12436
rect 10508 12384 10560 12436
rect 14740 12384 14792 12436
rect 16580 12384 16632 12436
rect 17408 12384 17460 12436
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7656 12223 7708 12232
rect 7288 12180 7340 12189
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 12072 12248 12124 12300
rect 17224 12316 17276 12368
rect 22928 12316 22980 12368
rect 3608 12044 3660 12096
rect 3884 12044 3936 12096
rect 5540 12044 5592 12096
rect 5632 12044 5684 12096
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 9772 12112 9824 12164
rect 9680 12044 9732 12096
rect 9956 12112 10008 12164
rect 10140 12044 10192 12096
rect 13452 12112 13504 12164
rect 16396 12248 16448 12300
rect 16764 12291 16816 12300
rect 16764 12257 16773 12291
rect 16773 12257 16807 12291
rect 16807 12257 16816 12291
rect 16764 12248 16816 12257
rect 14372 12180 14424 12232
rect 14556 12180 14608 12232
rect 15016 12223 15068 12232
rect 15016 12189 15025 12223
rect 15025 12189 15059 12223
rect 15059 12189 15068 12223
rect 15016 12180 15068 12189
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15200 12180 15252 12189
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 16948 12180 17000 12232
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 22192 12180 22244 12232
rect 22652 12180 22704 12232
rect 23112 12180 23164 12232
rect 23480 12180 23532 12232
rect 22284 12112 22336 12164
rect 23020 12112 23072 12164
rect 16212 12044 16264 12096
rect 19800 12087 19852 12096
rect 19800 12053 19809 12087
rect 19809 12053 19843 12087
rect 19843 12053 19852 12087
rect 19800 12044 19852 12053
rect 23756 12044 23808 12096
rect 23848 12087 23900 12096
rect 23848 12053 23857 12087
rect 23857 12053 23891 12087
rect 23891 12053 23900 12087
rect 23848 12044 23900 12053
rect 5151 11942 5203 11994
rect 5215 11942 5267 11994
rect 5279 11942 5331 11994
rect 5343 11942 5395 11994
rect 5407 11942 5459 11994
rect 12234 11942 12286 11994
rect 12298 11942 12350 11994
rect 12362 11942 12414 11994
rect 12426 11942 12478 11994
rect 12490 11942 12542 11994
rect 19317 11942 19369 11994
rect 19381 11942 19433 11994
rect 19445 11942 19497 11994
rect 19509 11942 19561 11994
rect 19573 11942 19625 11994
rect 26400 11942 26452 11994
rect 26464 11942 26516 11994
rect 26528 11942 26580 11994
rect 26592 11942 26644 11994
rect 26656 11942 26708 11994
rect 4436 11840 4488 11892
rect 5632 11840 5684 11892
rect 7196 11840 7248 11892
rect 7656 11840 7708 11892
rect 9864 11840 9916 11892
rect 3148 11772 3200 11824
rect 940 11704 992 11756
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 5080 11772 5132 11824
rect 5724 11772 5776 11824
rect 6552 11772 6604 11824
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 6368 11704 6420 11756
rect 7288 11704 7340 11756
rect 2228 11500 2280 11552
rect 4344 11636 4396 11688
rect 5448 11636 5500 11688
rect 6000 11568 6052 11620
rect 9772 11772 9824 11824
rect 12716 11840 12768 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 16120 11840 16172 11892
rect 19064 11840 19116 11892
rect 20168 11840 20220 11892
rect 20260 11840 20312 11892
rect 22284 11840 22336 11892
rect 14280 11772 14332 11824
rect 16212 11815 16264 11824
rect 16212 11781 16221 11815
rect 16221 11781 16255 11815
rect 16255 11781 16264 11815
rect 16212 11772 16264 11781
rect 23112 11840 23164 11892
rect 25504 11840 25556 11892
rect 8944 11636 8996 11688
rect 9772 11636 9824 11688
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 13452 11704 13504 11756
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14648 11704 14700 11756
rect 15660 11704 15712 11756
rect 13636 11636 13688 11688
rect 16488 11704 16540 11756
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 20076 11704 20128 11756
rect 20444 11704 20496 11756
rect 20536 11747 20588 11756
rect 20536 11713 20545 11747
rect 20545 11713 20579 11747
rect 20579 11713 20588 11747
rect 20536 11704 20588 11713
rect 16212 11636 16264 11688
rect 18052 11636 18104 11688
rect 19340 11636 19392 11688
rect 19984 11636 20036 11688
rect 16672 11568 16724 11620
rect 4252 11500 4304 11552
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 7380 11500 7432 11552
rect 14556 11500 14608 11552
rect 17592 11543 17644 11552
rect 17592 11509 17601 11543
rect 17601 11509 17635 11543
rect 17635 11509 17644 11543
rect 17592 11500 17644 11509
rect 22192 11704 22244 11756
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 22928 11704 22980 11756
rect 24032 11704 24084 11756
rect 26700 11704 26752 11756
rect 23296 11679 23348 11688
rect 23296 11645 23305 11679
rect 23305 11645 23339 11679
rect 23339 11645 23348 11679
rect 23296 11636 23348 11645
rect 22468 11568 22520 11620
rect 23756 11636 23808 11688
rect 22376 11500 22428 11552
rect 22652 11500 22704 11552
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 24584 11500 24636 11552
rect 26148 11500 26200 11552
rect 4491 11398 4543 11450
rect 4555 11398 4607 11450
rect 4619 11398 4671 11450
rect 4683 11398 4735 11450
rect 4747 11398 4799 11450
rect 11574 11398 11626 11450
rect 11638 11398 11690 11450
rect 11702 11398 11754 11450
rect 11766 11398 11818 11450
rect 11830 11398 11882 11450
rect 18657 11398 18709 11450
rect 18721 11398 18773 11450
rect 18785 11398 18837 11450
rect 18849 11398 18901 11450
rect 18913 11398 18965 11450
rect 25740 11398 25792 11450
rect 25804 11398 25856 11450
rect 25868 11398 25920 11450
rect 25932 11398 25984 11450
rect 25996 11398 26048 11450
rect 4344 11339 4396 11348
rect 4344 11305 4353 11339
rect 4353 11305 4387 11339
rect 4387 11305 4396 11339
rect 4344 11296 4396 11305
rect 11244 11296 11296 11348
rect 12164 11296 12216 11348
rect 15200 11296 15252 11348
rect 4068 11228 4120 11280
rect 2228 11160 2280 11212
rect 3884 11160 3936 11212
rect 3148 11092 3200 11144
rect 3700 11092 3752 11144
rect 2136 11067 2188 11076
rect 2136 11033 2145 11067
rect 2145 11033 2179 11067
rect 2179 11033 2188 11067
rect 2136 11024 2188 11033
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 7288 11228 7340 11280
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 6368 11160 6420 11212
rect 4620 11092 4672 11144
rect 7380 11092 7432 11144
rect 7840 11092 7892 11144
rect 8116 11092 8168 11144
rect 10140 11160 10192 11212
rect 17592 11296 17644 11348
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 19800 11296 19852 11348
rect 22100 11339 22152 11348
rect 22100 11305 22109 11339
rect 22109 11305 22143 11339
rect 22143 11305 22152 11339
rect 22100 11296 22152 11305
rect 22652 11296 22704 11348
rect 26700 11339 26752 11348
rect 26700 11305 26709 11339
rect 26709 11305 26743 11339
rect 26743 11305 26752 11339
rect 26700 11296 26752 11305
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 4712 10956 4764 11008
rect 5908 10956 5960 11008
rect 6184 11024 6236 11076
rect 7472 11067 7524 11076
rect 7472 11033 7481 11067
rect 7481 11033 7515 11067
rect 7515 11033 7524 11067
rect 7472 11024 7524 11033
rect 7564 11067 7616 11076
rect 7564 11033 7573 11067
rect 7573 11033 7607 11067
rect 7607 11033 7616 11067
rect 7564 11024 7616 11033
rect 8944 11024 8996 11076
rect 7104 10956 7156 11008
rect 13544 10956 13596 11008
rect 13820 10956 13872 11008
rect 14556 10956 14608 11008
rect 15936 11067 15988 11076
rect 15936 11033 15945 11067
rect 15945 11033 15979 11067
rect 15979 11033 15988 11067
rect 15936 11024 15988 11033
rect 18880 11271 18932 11280
rect 18880 11237 18889 11271
rect 18889 11237 18923 11271
rect 18923 11237 18932 11271
rect 18880 11228 18932 11237
rect 19340 11228 19392 11280
rect 22468 11271 22520 11280
rect 22468 11237 22477 11271
rect 22477 11237 22511 11271
rect 22511 11237 22520 11271
rect 22468 11228 22520 11237
rect 16580 11160 16632 11212
rect 19064 11160 19116 11212
rect 18144 11092 18196 11144
rect 18236 11092 18288 11144
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 22744 11160 22796 11212
rect 24952 11203 25004 11212
rect 24952 11169 24961 11203
rect 24961 11169 24995 11203
rect 24995 11169 25004 11203
rect 24952 11160 25004 11169
rect 28908 11160 28960 11212
rect 18696 11092 18748 11101
rect 19248 11092 19300 11144
rect 16856 11024 16908 11076
rect 16764 10956 16816 11008
rect 19708 11067 19760 11076
rect 19708 11033 19717 11067
rect 19717 11033 19751 11067
rect 19751 11033 19760 11067
rect 19708 11024 19760 11033
rect 22100 11135 22152 11144
rect 22100 11101 22109 11135
rect 22109 11101 22143 11135
rect 22143 11101 22152 11135
rect 22100 11092 22152 11101
rect 20352 11024 20404 11076
rect 21180 10956 21232 11008
rect 22376 11135 22428 11144
rect 22376 11101 22385 11135
rect 22385 11101 22419 11135
rect 22419 11101 22428 11135
rect 22376 11092 22428 11101
rect 22468 11024 22520 11076
rect 22928 11092 22980 11144
rect 23112 11067 23164 11076
rect 23112 11033 23121 11067
rect 23121 11033 23155 11067
rect 23155 11033 23164 11067
rect 23112 11024 23164 11033
rect 23572 11024 23624 11076
rect 23664 11024 23716 11076
rect 23940 10956 23992 11008
rect 24124 11024 24176 11076
rect 24308 10956 24360 11008
rect 28724 11135 28776 11144
rect 28724 11101 28733 11135
rect 28733 11101 28767 11135
rect 28767 11101 28776 11135
rect 28724 11092 28776 11101
rect 25228 11067 25280 11076
rect 25228 11033 25237 11067
rect 25237 11033 25271 11067
rect 25271 11033 25280 11067
rect 25228 11024 25280 11033
rect 25044 10956 25096 11008
rect 25320 10956 25372 11008
rect 27068 11024 27120 11076
rect 26792 10956 26844 11008
rect 5151 10854 5203 10906
rect 5215 10854 5267 10906
rect 5279 10854 5331 10906
rect 5343 10854 5395 10906
rect 5407 10854 5459 10906
rect 12234 10854 12286 10906
rect 12298 10854 12350 10906
rect 12362 10854 12414 10906
rect 12426 10854 12478 10906
rect 12490 10854 12542 10906
rect 19317 10854 19369 10906
rect 19381 10854 19433 10906
rect 19445 10854 19497 10906
rect 19509 10854 19561 10906
rect 19573 10854 19625 10906
rect 26400 10854 26452 10906
rect 26464 10854 26516 10906
rect 26528 10854 26580 10906
rect 26592 10854 26644 10906
rect 26656 10854 26708 10906
rect 4068 10752 4120 10804
rect 4160 10752 4212 10804
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 4712 10752 4764 10804
rect 4896 10727 4948 10736
rect 4896 10693 4905 10727
rect 4905 10693 4939 10727
rect 4939 10693 4948 10727
rect 4896 10684 4948 10693
rect 5264 10684 5316 10736
rect 5724 10752 5776 10804
rect 5908 10795 5960 10804
rect 5908 10761 5917 10795
rect 5917 10761 5951 10795
rect 5951 10761 5960 10795
rect 5908 10752 5960 10761
rect 6000 10795 6052 10804
rect 6000 10761 6009 10795
rect 6009 10761 6043 10795
rect 6043 10761 6052 10795
rect 6000 10752 6052 10761
rect 9772 10752 9824 10804
rect 14004 10752 14056 10804
rect 14556 10795 14608 10804
rect 14556 10761 14565 10795
rect 14565 10761 14599 10795
rect 14599 10761 14608 10795
rect 14556 10752 14608 10761
rect 18512 10752 18564 10804
rect 20352 10795 20404 10804
rect 20352 10761 20361 10795
rect 20361 10761 20395 10795
rect 20395 10761 20404 10795
rect 20352 10752 20404 10761
rect 23020 10752 23072 10804
rect 5540 10684 5592 10736
rect 4804 10548 4856 10600
rect 7196 10616 7248 10668
rect 4068 10412 4120 10464
rect 4160 10412 4212 10464
rect 5264 10480 5316 10532
rect 5632 10480 5684 10532
rect 5540 10412 5592 10464
rect 7012 10548 7064 10600
rect 19800 10684 19852 10736
rect 20076 10684 20128 10736
rect 23848 10752 23900 10804
rect 23940 10752 23992 10804
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 13544 10616 13596 10668
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 14924 10616 14976 10668
rect 15476 10616 15528 10668
rect 10416 10548 10468 10600
rect 11428 10548 11480 10600
rect 10600 10480 10652 10532
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 15292 10548 15344 10600
rect 16212 10616 16264 10668
rect 15936 10480 15988 10532
rect 16764 10548 16816 10600
rect 17316 10659 17368 10668
rect 17316 10625 17330 10659
rect 17330 10625 17364 10659
rect 17364 10625 17368 10659
rect 17316 10616 17368 10625
rect 17776 10616 17828 10668
rect 17868 10659 17920 10668
rect 17868 10625 17874 10659
rect 17874 10625 17908 10659
rect 17908 10625 17920 10659
rect 17868 10616 17920 10625
rect 18052 10616 18104 10668
rect 18420 10548 18472 10600
rect 9956 10412 10008 10464
rect 10048 10412 10100 10464
rect 10416 10412 10468 10464
rect 10508 10412 10560 10464
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 14740 10455 14792 10464
rect 14740 10421 14749 10455
rect 14749 10421 14783 10455
rect 14783 10421 14792 10455
rect 14740 10412 14792 10421
rect 17408 10412 17460 10464
rect 18972 10659 19024 10668
rect 18972 10625 18981 10659
rect 18981 10625 19015 10659
rect 19015 10625 19024 10659
rect 18972 10616 19024 10625
rect 19064 10616 19116 10668
rect 20536 10616 20588 10668
rect 20444 10548 20496 10600
rect 22008 10616 22060 10668
rect 22468 10616 22520 10668
rect 22744 10616 22796 10668
rect 25228 10752 25280 10804
rect 24584 10684 24636 10736
rect 25044 10684 25096 10736
rect 25780 10684 25832 10736
rect 26148 10616 26200 10668
rect 26424 10659 26476 10668
rect 26424 10625 26433 10659
rect 26433 10625 26467 10659
rect 26467 10625 26476 10659
rect 26424 10616 26476 10625
rect 26516 10659 26568 10668
rect 26516 10625 26525 10659
rect 26525 10625 26559 10659
rect 26559 10625 26568 10659
rect 26516 10616 26568 10625
rect 26608 10616 26660 10668
rect 20904 10548 20956 10600
rect 22192 10548 22244 10600
rect 25596 10591 25648 10600
rect 25596 10557 25605 10591
rect 25605 10557 25639 10591
rect 25639 10557 25648 10591
rect 25596 10548 25648 10557
rect 20536 10480 20588 10532
rect 24308 10480 24360 10532
rect 19892 10412 19944 10464
rect 22376 10455 22428 10464
rect 22376 10421 22385 10455
rect 22385 10421 22419 10455
rect 22419 10421 22428 10455
rect 22376 10412 22428 10421
rect 4491 10310 4543 10362
rect 4555 10310 4607 10362
rect 4619 10310 4671 10362
rect 4683 10310 4735 10362
rect 4747 10310 4799 10362
rect 11574 10310 11626 10362
rect 11638 10310 11690 10362
rect 11702 10310 11754 10362
rect 11766 10310 11818 10362
rect 11830 10310 11882 10362
rect 18657 10310 18709 10362
rect 18721 10310 18773 10362
rect 18785 10310 18837 10362
rect 18849 10310 18901 10362
rect 18913 10310 18965 10362
rect 25740 10310 25792 10362
rect 25804 10310 25856 10362
rect 25868 10310 25920 10362
rect 25932 10310 25984 10362
rect 25996 10310 26048 10362
rect 4068 10208 4120 10260
rect 9772 10208 9824 10260
rect 10048 10208 10100 10260
rect 10140 10208 10192 10260
rect 10968 10208 11020 10260
rect 12624 10208 12676 10260
rect 13544 10251 13596 10260
rect 13544 10217 13575 10251
rect 13575 10217 13596 10251
rect 13544 10208 13596 10217
rect 16488 10208 16540 10260
rect 17316 10208 17368 10260
rect 18144 10208 18196 10260
rect 19156 10208 19208 10260
rect 20260 10208 20312 10260
rect 22652 10208 22704 10260
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 10232 10115 10284 10124
rect 10232 10081 10241 10115
rect 10241 10081 10275 10115
rect 10275 10081 10284 10115
rect 10232 10072 10284 10081
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 10324 10004 10376 10056
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 13268 10183 13320 10192
rect 13268 10149 13277 10183
rect 13277 10149 13311 10183
rect 13311 10149 13320 10183
rect 13268 10140 13320 10149
rect 9956 9936 10008 9988
rect 10968 10004 11020 10056
rect 11060 10004 11112 10056
rect 11428 10049 11480 10056
rect 11428 10015 11437 10049
rect 11437 10015 11471 10049
rect 11471 10015 11480 10049
rect 11428 10004 11480 10015
rect 16580 10115 16632 10124
rect 16580 10081 16589 10115
rect 16589 10081 16623 10115
rect 16623 10081 16632 10115
rect 16580 10072 16632 10081
rect 17868 10140 17920 10192
rect 18236 10072 18288 10124
rect 19064 10072 19116 10124
rect 20904 10140 20956 10192
rect 20444 10115 20496 10124
rect 20444 10081 20453 10115
rect 20453 10081 20487 10115
rect 20487 10081 20496 10115
rect 20444 10072 20496 10081
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 10324 9868 10376 9920
rect 10876 9868 10928 9920
rect 11336 9936 11388 9988
rect 13360 9979 13412 9988
rect 13360 9945 13369 9979
rect 13369 9945 13403 9979
rect 13403 9945 13412 9979
rect 13360 9936 13412 9945
rect 12072 9868 12124 9920
rect 13084 9868 13136 9920
rect 15292 10004 15344 10056
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 15476 10047 15528 10056
rect 15476 10013 15486 10047
rect 15486 10013 15520 10047
rect 15520 10013 15528 10047
rect 15476 10004 15528 10013
rect 16488 10004 16540 10056
rect 18144 10004 18196 10056
rect 18328 10004 18380 10056
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 20076 10004 20128 10056
rect 22928 10208 22980 10260
rect 23388 10208 23440 10260
rect 25596 10208 25648 10260
rect 23204 10072 23256 10124
rect 13820 9868 13872 9920
rect 15200 9868 15252 9920
rect 16856 9979 16908 9988
rect 16856 9945 16865 9979
rect 16865 9945 16899 9979
rect 16899 9945 16908 9979
rect 16856 9936 16908 9945
rect 22192 9936 22244 9988
rect 22928 10004 22980 10056
rect 26516 10072 26568 10124
rect 26884 10072 26936 10124
rect 22836 9979 22888 9988
rect 22836 9945 22845 9979
rect 22845 9945 22879 9979
rect 22879 9945 22888 9979
rect 22836 9936 22888 9945
rect 18328 9911 18380 9920
rect 18328 9877 18337 9911
rect 18337 9877 18371 9911
rect 18371 9877 18380 9911
rect 18328 9868 18380 9877
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 22376 9911 22428 9920
rect 22376 9877 22385 9911
rect 22385 9877 22419 9911
rect 22419 9877 22428 9911
rect 22376 9868 22428 9877
rect 26424 10004 26476 10056
rect 26148 9868 26200 9920
rect 26240 9868 26292 9920
rect 5151 9766 5203 9818
rect 5215 9766 5267 9818
rect 5279 9766 5331 9818
rect 5343 9766 5395 9818
rect 5407 9766 5459 9818
rect 12234 9766 12286 9818
rect 12298 9766 12350 9818
rect 12362 9766 12414 9818
rect 12426 9766 12478 9818
rect 12490 9766 12542 9818
rect 19317 9766 19369 9818
rect 19381 9766 19433 9818
rect 19445 9766 19497 9818
rect 19509 9766 19561 9818
rect 19573 9766 19625 9818
rect 26400 9766 26452 9818
rect 26464 9766 26516 9818
rect 26528 9766 26580 9818
rect 26592 9766 26644 9818
rect 26656 9766 26708 9818
rect 6000 9664 6052 9716
rect 2228 9596 2280 9648
rect 4068 9596 4120 9648
rect 3332 9528 3384 9580
rect 4896 9528 4948 9580
rect 4160 9460 4212 9512
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 6276 9596 6328 9648
rect 9956 9664 10008 9716
rect 10508 9664 10560 9716
rect 10600 9707 10652 9716
rect 10600 9673 10609 9707
rect 10609 9673 10643 9707
rect 10643 9673 10652 9707
rect 10600 9664 10652 9673
rect 10692 9664 10744 9716
rect 10876 9664 10928 9716
rect 16856 9664 16908 9716
rect 18512 9707 18564 9716
rect 18512 9673 18521 9707
rect 18521 9673 18555 9707
rect 18555 9673 18564 9707
rect 18512 9664 18564 9673
rect 18972 9664 19024 9716
rect 21456 9664 21508 9716
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10232 9596 10284 9605
rect 9036 9528 9088 9580
rect 9864 9528 9916 9580
rect 9956 9528 10008 9580
rect 6184 9460 6236 9512
rect 4344 9324 4396 9376
rect 5080 9324 5132 9376
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 6552 9392 6604 9444
rect 6644 9324 6696 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9680 9460 9732 9512
rect 10324 9460 10376 9512
rect 10140 9392 10192 9444
rect 10692 9435 10744 9444
rect 10692 9401 10701 9435
rect 10701 9401 10735 9435
rect 10735 9401 10744 9435
rect 10692 9392 10744 9401
rect 10048 9324 10100 9376
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11336 9596 11388 9648
rect 13176 9639 13228 9648
rect 13176 9605 13185 9639
rect 13185 9605 13219 9639
rect 13219 9605 13228 9639
rect 13176 9596 13228 9605
rect 11980 9528 12032 9580
rect 13452 9596 13504 9648
rect 13820 9596 13872 9648
rect 14280 9596 14332 9648
rect 26884 9596 26936 9648
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 11060 9460 11112 9512
rect 14004 9460 14056 9512
rect 16580 9460 16632 9512
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 16028 9392 16080 9444
rect 18328 9528 18380 9580
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 17868 9392 17920 9444
rect 19064 9528 19116 9580
rect 22560 9528 22612 9580
rect 26332 9571 26384 9580
rect 26332 9537 26341 9571
rect 26341 9537 26375 9571
rect 26375 9537 26384 9571
rect 26332 9528 26384 9537
rect 13636 9324 13688 9376
rect 14280 9324 14332 9376
rect 17592 9367 17644 9376
rect 17592 9333 17601 9367
rect 17601 9333 17635 9367
rect 17635 9333 17644 9367
rect 17592 9324 17644 9333
rect 17960 9324 18012 9376
rect 18420 9324 18472 9376
rect 27804 9528 27856 9580
rect 28080 9596 28132 9648
rect 26884 9460 26936 9512
rect 28172 9571 28224 9580
rect 28172 9537 28181 9571
rect 28181 9537 28215 9571
rect 28215 9537 28224 9571
rect 28172 9528 28224 9537
rect 26148 9392 26200 9444
rect 19340 9324 19392 9376
rect 25596 9324 25648 9376
rect 28448 9324 28500 9376
rect 4491 9222 4543 9274
rect 4555 9222 4607 9274
rect 4619 9222 4671 9274
rect 4683 9222 4735 9274
rect 4747 9222 4799 9274
rect 11574 9222 11626 9274
rect 11638 9222 11690 9274
rect 11702 9222 11754 9274
rect 11766 9222 11818 9274
rect 11830 9222 11882 9274
rect 18657 9222 18709 9274
rect 18721 9222 18773 9274
rect 18785 9222 18837 9274
rect 18849 9222 18901 9274
rect 18913 9222 18965 9274
rect 25740 9222 25792 9274
rect 25804 9222 25856 9274
rect 25868 9222 25920 9274
rect 25932 9222 25984 9274
rect 25996 9222 26048 9274
rect 5632 9120 5684 9172
rect 3332 9052 3384 9104
rect 5080 9052 5132 9104
rect 5540 9052 5592 9104
rect 10416 9052 10468 9104
rect 13084 9163 13136 9172
rect 13084 9129 13093 9163
rect 13093 9129 13127 9163
rect 13127 9129 13136 9163
rect 13084 9120 13136 9129
rect 17500 9120 17552 9172
rect 2228 8984 2280 9036
rect 4344 8984 4396 9036
rect 6000 8984 6052 9036
rect 9128 8984 9180 9036
rect 9864 8984 9916 9036
rect 10140 8984 10192 9036
rect 17316 9052 17368 9104
rect 18328 9052 18380 9104
rect 22836 9120 22888 9172
rect 24952 9120 25004 9172
rect 24032 9052 24084 9104
rect 25596 9052 25648 9104
rect 25688 9052 25740 9104
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 11060 8984 11112 9036
rect 11244 8984 11296 9036
rect 12072 8984 12124 9036
rect 15660 8984 15712 9036
rect 6276 8848 6328 8900
rect 7104 8848 7156 8900
rect 9680 8848 9732 8900
rect 11336 8848 11388 8900
rect 4344 8780 4396 8832
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 5080 8780 5132 8832
rect 9956 8780 10008 8832
rect 12164 8916 12216 8968
rect 13728 8916 13780 8968
rect 13268 8848 13320 8900
rect 18144 8984 18196 9036
rect 18052 8916 18104 8968
rect 22192 9027 22244 9036
rect 22192 8993 22201 9027
rect 22201 8993 22235 9027
rect 22235 8993 22244 9027
rect 22192 8984 22244 8993
rect 22284 9027 22336 9036
rect 22284 8993 22293 9027
rect 22293 8993 22327 9027
rect 22327 8993 22336 9027
rect 22284 8984 22336 8993
rect 22468 8984 22520 9036
rect 19340 8959 19392 8968
rect 19340 8925 19349 8959
rect 19349 8925 19383 8959
rect 19383 8925 19392 8959
rect 19340 8916 19392 8925
rect 13912 8848 13964 8900
rect 16396 8848 16448 8900
rect 16856 8848 16908 8900
rect 18236 8891 18288 8900
rect 18236 8857 18245 8891
rect 18245 8857 18279 8891
rect 18279 8857 18288 8891
rect 18236 8848 18288 8857
rect 13636 8823 13688 8832
rect 13636 8789 13651 8823
rect 13651 8789 13685 8823
rect 13685 8789 13688 8823
rect 13636 8780 13688 8789
rect 18052 8780 18104 8832
rect 22376 8916 22428 8968
rect 22560 8891 22612 8900
rect 22560 8857 22569 8891
rect 22569 8857 22603 8891
rect 22603 8857 22612 8891
rect 22560 8848 22612 8857
rect 18512 8823 18564 8832
rect 18512 8789 18521 8823
rect 18521 8789 18555 8823
rect 18555 8789 18564 8823
rect 18512 8780 18564 8789
rect 20628 8780 20680 8832
rect 21732 8823 21784 8832
rect 21732 8789 21741 8823
rect 21741 8789 21775 8823
rect 21775 8789 21784 8823
rect 21732 8780 21784 8789
rect 22100 8780 22152 8832
rect 23388 8916 23440 8968
rect 27804 9120 27856 9172
rect 26148 8959 26200 8968
rect 26148 8925 26157 8959
rect 26157 8925 26191 8959
rect 26191 8925 26200 8959
rect 26148 8916 26200 8925
rect 25780 8891 25832 8900
rect 25780 8857 25789 8891
rect 25789 8857 25823 8891
rect 25823 8857 25832 8891
rect 25780 8848 25832 8857
rect 25872 8891 25924 8900
rect 25872 8857 25881 8891
rect 25881 8857 25915 8891
rect 25915 8857 25924 8891
rect 25872 8848 25924 8857
rect 22652 8780 22704 8832
rect 26792 8848 26844 8900
rect 27068 8848 27120 8900
rect 28448 8848 28500 8900
rect 5151 8678 5203 8730
rect 5215 8678 5267 8730
rect 5279 8678 5331 8730
rect 5343 8678 5395 8730
rect 5407 8678 5459 8730
rect 12234 8678 12286 8730
rect 12298 8678 12350 8730
rect 12362 8678 12414 8730
rect 12426 8678 12478 8730
rect 12490 8678 12542 8730
rect 19317 8678 19369 8730
rect 19381 8678 19433 8730
rect 19445 8678 19497 8730
rect 19509 8678 19561 8730
rect 19573 8678 19625 8730
rect 26400 8678 26452 8730
rect 26464 8678 26516 8730
rect 26528 8678 26580 8730
rect 26592 8678 26644 8730
rect 26656 8678 26708 8730
rect 2228 8576 2280 8628
rect 3332 8576 3384 8628
rect 1676 8440 1728 8492
rect 2688 8508 2740 8560
rect 4896 8576 4948 8628
rect 5540 8576 5592 8628
rect 6000 8576 6052 8628
rect 6736 8576 6788 8628
rect 5816 8508 5868 8560
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 4436 8440 4488 8492
rect 5448 8440 5500 8492
rect 4344 8304 4396 8356
rect 4988 8372 5040 8424
rect 5080 8415 5132 8424
rect 5080 8381 5089 8415
rect 5089 8381 5123 8415
rect 5123 8381 5132 8415
rect 5080 8372 5132 8381
rect 5724 8372 5776 8424
rect 6276 8440 6328 8492
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 9036 8551 9088 8560
rect 9036 8517 9045 8551
rect 9045 8517 9079 8551
rect 9079 8517 9088 8551
rect 9036 8508 9088 8517
rect 9956 8576 10008 8628
rect 13268 8576 13320 8628
rect 9772 8440 9824 8492
rect 13636 8508 13688 8560
rect 14280 8508 14332 8560
rect 16764 8576 16816 8628
rect 17592 8576 17644 8628
rect 18512 8576 18564 8628
rect 19156 8576 19208 8628
rect 15660 8508 15712 8560
rect 16580 8440 16632 8492
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 6736 8415 6788 8424
rect 6736 8381 6745 8415
rect 6745 8381 6779 8415
rect 6779 8381 6788 8415
rect 6736 8372 6788 8381
rect 8208 8372 8260 8424
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5080 8236 5132 8245
rect 5540 8236 5592 8288
rect 6184 8236 6236 8288
rect 9496 8372 9548 8424
rect 13360 8415 13412 8424
rect 13360 8381 13369 8415
rect 13369 8381 13403 8415
rect 13403 8381 13412 8415
rect 13360 8372 13412 8381
rect 13452 8415 13504 8424
rect 13452 8381 13461 8415
rect 13461 8381 13495 8415
rect 13495 8381 13504 8415
rect 13452 8372 13504 8381
rect 12164 8304 12216 8356
rect 16580 8304 16632 8356
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 17776 8440 17828 8492
rect 19248 8508 19300 8560
rect 20628 8619 20680 8628
rect 20628 8585 20637 8619
rect 20637 8585 20671 8619
rect 20671 8585 20680 8619
rect 20628 8576 20680 8585
rect 21732 8576 21784 8628
rect 23020 8576 23072 8628
rect 23664 8508 23716 8560
rect 22560 8440 22612 8492
rect 22928 8440 22980 8492
rect 23204 8440 23256 8492
rect 23480 8440 23532 8492
rect 24216 8508 24268 8560
rect 25780 8508 25832 8560
rect 26240 8508 26292 8560
rect 23388 8372 23440 8424
rect 23756 8415 23808 8424
rect 23756 8381 23765 8415
rect 23765 8381 23799 8415
rect 23799 8381 23808 8415
rect 23756 8372 23808 8381
rect 24032 8440 24084 8492
rect 26424 8440 26476 8492
rect 23020 8304 23072 8356
rect 23664 8347 23716 8356
rect 23664 8313 23673 8347
rect 23673 8313 23707 8347
rect 23707 8313 23716 8347
rect 23664 8304 23716 8313
rect 26332 8415 26384 8424
rect 26332 8381 26341 8415
rect 26341 8381 26375 8415
rect 26375 8381 26384 8415
rect 26332 8372 26384 8381
rect 26516 8304 26568 8356
rect 26608 8347 26660 8356
rect 26608 8313 26617 8347
rect 26617 8313 26651 8347
rect 26651 8313 26660 8347
rect 26608 8304 26660 8313
rect 26884 8440 26936 8492
rect 28448 8508 28500 8560
rect 27620 8440 27672 8492
rect 28080 8440 28132 8492
rect 28172 8440 28224 8492
rect 26884 8304 26936 8356
rect 27528 8304 27580 8356
rect 13912 8236 13964 8288
rect 17040 8236 17092 8288
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 22468 8236 22520 8288
rect 22928 8236 22980 8288
rect 24676 8236 24728 8288
rect 4491 8134 4543 8186
rect 4555 8134 4607 8186
rect 4619 8134 4671 8186
rect 4683 8134 4735 8186
rect 4747 8134 4799 8186
rect 11574 8134 11626 8186
rect 11638 8134 11690 8186
rect 11702 8134 11754 8186
rect 11766 8134 11818 8186
rect 11830 8134 11882 8186
rect 18657 8134 18709 8186
rect 18721 8134 18773 8186
rect 18785 8134 18837 8186
rect 18849 8134 18901 8186
rect 18913 8134 18965 8186
rect 25740 8134 25792 8186
rect 25804 8134 25856 8186
rect 25868 8134 25920 8186
rect 25932 8134 25984 8186
rect 25996 8134 26048 8186
rect 4068 7964 4120 8016
rect 6736 8007 6788 8016
rect 6736 7973 6745 8007
rect 6745 7973 6779 8007
rect 6779 7973 6788 8007
rect 6736 7964 6788 7973
rect 14096 8032 14148 8084
rect 14464 8032 14516 8084
rect 14740 8032 14792 8084
rect 14188 7964 14240 8016
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 3332 7828 3384 7880
rect 5448 7896 5500 7948
rect 5724 7939 5776 7948
rect 5724 7905 5733 7939
rect 5733 7905 5767 7939
rect 5767 7905 5776 7939
rect 5724 7896 5776 7905
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 7196 7896 7248 7948
rect 9956 7896 10008 7948
rect 14004 7896 14056 7948
rect 18052 8032 18104 8084
rect 22192 8032 22244 8084
rect 22284 8032 22336 8084
rect 17316 7964 17368 8016
rect 17776 7964 17828 8016
rect 23848 8032 23900 8084
rect 26608 8032 26660 8084
rect 27344 8032 27396 8084
rect 27528 8075 27580 8084
rect 27528 8041 27537 8075
rect 27537 8041 27571 8075
rect 27571 8041 27580 8075
rect 27528 8032 27580 8041
rect 4160 7760 4212 7812
rect 4896 7803 4948 7812
rect 4896 7769 4905 7803
rect 4905 7769 4939 7803
rect 4939 7769 4948 7803
rect 4896 7760 4948 7769
rect 6184 7760 6236 7812
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 6644 7760 6696 7812
rect 6828 7760 6880 7812
rect 4252 7692 4304 7744
rect 6276 7692 6328 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 9864 7760 9916 7812
rect 13636 7760 13688 7812
rect 13728 7803 13780 7812
rect 13728 7769 13769 7803
rect 13769 7769 13780 7803
rect 14464 7828 14516 7880
rect 14648 7828 14700 7880
rect 15108 7828 15160 7880
rect 15476 7828 15528 7880
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 16764 7828 16816 7880
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 17960 7871 18012 7880
rect 17960 7837 17967 7871
rect 17967 7837 18012 7871
rect 13728 7760 13780 7769
rect 7196 7735 7248 7744
rect 7196 7701 7205 7735
rect 7205 7701 7239 7735
rect 7239 7701 7248 7735
rect 7196 7692 7248 7701
rect 13360 7692 13412 7744
rect 13912 7735 13964 7744
rect 13912 7701 13921 7735
rect 13921 7701 13955 7735
rect 13955 7701 13964 7735
rect 13912 7692 13964 7701
rect 14004 7692 14056 7744
rect 17224 7803 17276 7812
rect 17224 7769 17233 7803
rect 17233 7769 17267 7803
rect 17267 7769 17276 7803
rect 17224 7760 17276 7769
rect 17960 7828 18012 7837
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 20904 7896 20956 7948
rect 20076 7871 20128 7880
rect 20076 7837 20085 7871
rect 20085 7837 20119 7871
rect 20119 7837 20128 7871
rect 20076 7828 20128 7837
rect 22008 7871 22060 7880
rect 22008 7837 22017 7871
rect 22017 7837 22051 7871
rect 22051 7837 22060 7871
rect 22008 7828 22060 7837
rect 22468 7896 22520 7948
rect 22284 7871 22336 7880
rect 22284 7837 22293 7871
rect 22293 7837 22327 7871
rect 22327 7837 22336 7871
rect 22284 7828 22336 7837
rect 22560 7871 22612 7880
rect 22560 7837 22569 7871
rect 22569 7837 22603 7871
rect 22603 7837 22612 7871
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 16764 7735 16816 7744
rect 16764 7701 16773 7735
rect 16773 7701 16807 7735
rect 16807 7701 16816 7735
rect 16764 7692 16816 7701
rect 17500 7692 17552 7744
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 21916 7760 21968 7812
rect 22560 7828 22612 7837
rect 23020 7964 23072 8016
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 22100 7692 22152 7744
rect 24032 7964 24084 8016
rect 26148 7964 26200 8016
rect 26332 7964 26384 8016
rect 23388 7828 23440 7880
rect 23480 7828 23532 7880
rect 23572 7828 23624 7880
rect 23664 7871 23716 7880
rect 23664 7837 23673 7871
rect 23673 7837 23707 7871
rect 23707 7837 23716 7871
rect 23664 7828 23716 7837
rect 23756 7871 23808 7880
rect 23756 7837 23765 7871
rect 23765 7837 23799 7871
rect 23799 7837 23808 7871
rect 23756 7828 23808 7837
rect 24216 7896 24268 7948
rect 24124 7828 24176 7880
rect 24676 7828 24728 7880
rect 22376 7735 22428 7744
rect 22376 7701 22385 7735
rect 22385 7701 22419 7735
rect 22419 7701 22428 7735
rect 22376 7692 22428 7701
rect 22468 7692 22520 7744
rect 24216 7760 24268 7812
rect 25504 7896 25556 7948
rect 27528 7939 27580 7948
rect 27528 7905 27537 7939
rect 27537 7905 27571 7939
rect 27571 7905 27580 7939
rect 27528 7896 27580 7905
rect 23296 7735 23348 7744
rect 23296 7701 23305 7735
rect 23305 7701 23339 7735
rect 23339 7701 23348 7735
rect 23296 7692 23348 7701
rect 23664 7692 23716 7744
rect 23756 7692 23808 7744
rect 25596 7735 25648 7744
rect 25596 7701 25605 7735
rect 25605 7701 25639 7735
rect 25639 7701 25648 7735
rect 25596 7692 25648 7701
rect 26516 7871 26568 7880
rect 26516 7837 26525 7871
rect 26525 7837 26559 7871
rect 26559 7837 26568 7871
rect 26516 7828 26568 7837
rect 26608 7828 26660 7880
rect 26976 7828 27028 7880
rect 25872 7803 25924 7812
rect 25872 7769 25881 7803
rect 25881 7769 25915 7803
rect 25915 7769 25924 7803
rect 25872 7760 25924 7769
rect 26240 7760 26292 7812
rect 26792 7760 26844 7812
rect 5151 7590 5203 7642
rect 5215 7590 5267 7642
rect 5279 7590 5331 7642
rect 5343 7590 5395 7642
rect 5407 7590 5459 7642
rect 12234 7590 12286 7642
rect 12298 7590 12350 7642
rect 12362 7590 12414 7642
rect 12426 7590 12478 7642
rect 12490 7590 12542 7642
rect 19317 7590 19369 7642
rect 19381 7590 19433 7642
rect 19445 7590 19497 7642
rect 19509 7590 19561 7642
rect 19573 7590 19625 7642
rect 26400 7590 26452 7642
rect 26464 7590 26516 7642
rect 26528 7590 26580 7642
rect 26592 7590 26644 7642
rect 26656 7590 26708 7642
rect 5080 7488 5132 7540
rect 5816 7488 5868 7540
rect 6552 7488 6604 7540
rect 12348 7488 12400 7540
rect 5724 7284 5776 7336
rect 5816 7327 5868 7336
rect 5816 7293 5825 7327
rect 5825 7293 5859 7327
rect 5859 7293 5868 7327
rect 5816 7284 5868 7293
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 11336 7352 11388 7404
rect 11428 7352 11480 7404
rect 12164 7352 12216 7404
rect 14648 7488 14700 7540
rect 16764 7488 16816 7540
rect 17132 7488 17184 7540
rect 14280 7420 14332 7472
rect 9680 7284 9732 7336
rect 10784 7284 10836 7336
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 14188 7284 14240 7336
rect 15108 7284 15160 7336
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 17408 7488 17460 7540
rect 17684 7488 17736 7540
rect 18052 7488 18104 7540
rect 22560 7531 22612 7540
rect 22560 7497 22569 7531
rect 22569 7497 22603 7531
rect 22603 7497 22612 7531
rect 22560 7488 22612 7497
rect 22928 7531 22980 7540
rect 22928 7497 22937 7531
rect 22937 7497 22971 7531
rect 22971 7497 22980 7531
rect 22928 7488 22980 7497
rect 23020 7488 23072 7540
rect 23664 7488 23716 7540
rect 17776 7420 17828 7472
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 17500 7395 17552 7404
rect 17500 7361 17509 7395
rect 17509 7361 17543 7395
rect 17543 7361 17552 7395
rect 17500 7352 17552 7361
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 18052 7395 18104 7404
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 24584 7420 24636 7472
rect 18420 7395 18472 7404
rect 18420 7361 18429 7395
rect 18429 7361 18463 7395
rect 18463 7361 18472 7395
rect 18420 7352 18472 7361
rect 18512 7352 18564 7404
rect 22284 7352 22336 7404
rect 22836 7352 22888 7404
rect 22192 7284 22244 7336
rect 22008 7216 22060 7268
rect 23296 7352 23348 7404
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 25596 7488 25648 7540
rect 25872 7488 25924 7540
rect 24952 7395 25004 7404
rect 24952 7361 24961 7395
rect 24961 7361 24995 7395
rect 24995 7361 25004 7395
rect 24952 7352 25004 7361
rect 25320 7284 25372 7336
rect 26884 7352 26936 7404
rect 26976 7395 27028 7404
rect 26976 7361 26985 7395
rect 26985 7361 27019 7395
rect 27019 7361 27028 7395
rect 26976 7352 27028 7361
rect 27068 7352 27120 7404
rect 27344 7352 27396 7404
rect 24124 7216 24176 7268
rect 26792 7216 26844 7268
rect 27528 7259 27580 7268
rect 27528 7225 27537 7259
rect 27537 7225 27571 7259
rect 27571 7225 27580 7259
rect 27528 7216 27580 7225
rect 6276 7148 6328 7200
rect 7748 7148 7800 7200
rect 11060 7148 11112 7200
rect 11152 7148 11204 7200
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 11980 7191 12032 7200
rect 11980 7157 11989 7191
rect 11989 7157 12023 7191
rect 12023 7157 12032 7191
rect 11980 7148 12032 7157
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 17408 7148 17460 7200
rect 17868 7191 17920 7200
rect 17868 7157 17877 7191
rect 17877 7157 17911 7191
rect 17911 7157 17920 7191
rect 17868 7148 17920 7157
rect 24400 7191 24452 7200
rect 24400 7157 24409 7191
rect 24409 7157 24443 7191
rect 24443 7157 24452 7191
rect 24400 7148 24452 7157
rect 28724 7395 28776 7404
rect 28724 7361 28733 7395
rect 28733 7361 28767 7395
rect 28767 7361 28776 7395
rect 28724 7352 28776 7361
rect 28908 7148 28960 7200
rect 4491 7046 4543 7098
rect 4555 7046 4607 7098
rect 4619 7046 4671 7098
rect 4683 7046 4735 7098
rect 4747 7046 4799 7098
rect 11574 7046 11626 7098
rect 11638 7046 11690 7098
rect 11702 7046 11754 7098
rect 11766 7046 11818 7098
rect 11830 7046 11882 7098
rect 18657 7046 18709 7098
rect 18721 7046 18773 7098
rect 18785 7046 18837 7098
rect 18849 7046 18901 7098
rect 18913 7046 18965 7098
rect 25740 7046 25792 7098
rect 25804 7046 25856 7098
rect 25868 7046 25920 7098
rect 25932 7046 25984 7098
rect 25996 7046 26048 7098
rect 4896 6944 4948 6996
rect 5080 6919 5132 6928
rect 5080 6885 5089 6919
rect 5089 6885 5123 6919
rect 5123 6885 5132 6919
rect 5080 6876 5132 6885
rect 5908 6808 5960 6860
rect 6276 6808 6328 6860
rect 6092 6740 6144 6792
rect 7288 6876 7340 6928
rect 7012 6808 7064 6860
rect 8116 6944 8168 6996
rect 10416 6944 10468 6996
rect 11244 6944 11296 6996
rect 11704 6944 11756 6996
rect 12348 6944 12400 6996
rect 10140 6876 10192 6928
rect 6736 6740 6788 6792
rect 6276 6715 6328 6724
rect 6276 6681 6285 6715
rect 6285 6681 6319 6715
rect 6319 6681 6328 6715
rect 6276 6672 6328 6681
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 8116 6740 8168 6792
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 6828 6604 6880 6656
rect 7748 6715 7800 6724
rect 7748 6681 7757 6715
rect 7757 6681 7791 6715
rect 7791 6681 7800 6715
rect 9864 6808 9916 6860
rect 8300 6740 8352 6792
rect 11152 6808 11204 6860
rect 11336 6919 11388 6928
rect 11336 6885 11345 6919
rect 11345 6885 11379 6919
rect 11379 6885 11388 6919
rect 11336 6876 11388 6885
rect 12072 6876 12124 6928
rect 11428 6851 11480 6860
rect 11428 6817 11437 6851
rect 11437 6817 11471 6851
rect 11471 6817 11480 6851
rect 11428 6808 11480 6817
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 11060 6740 11112 6792
rect 11336 6740 11388 6792
rect 11980 6740 12032 6792
rect 7748 6672 7800 6681
rect 9772 6672 9824 6724
rect 9864 6672 9916 6724
rect 10048 6715 10100 6724
rect 10048 6681 10057 6715
rect 10057 6681 10091 6715
rect 10091 6681 10100 6715
rect 10048 6672 10100 6681
rect 7656 6604 7708 6656
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 10600 6672 10652 6724
rect 11704 6715 11756 6724
rect 11704 6681 11713 6715
rect 11713 6681 11747 6715
rect 11747 6681 11756 6715
rect 11704 6672 11756 6681
rect 13636 6808 13688 6860
rect 13912 6876 13964 6928
rect 14464 6987 14516 6996
rect 14464 6953 14473 6987
rect 14473 6953 14507 6987
rect 14507 6953 14516 6987
rect 14464 6944 14516 6953
rect 16580 6944 16632 6996
rect 16764 6944 16816 6996
rect 17776 6944 17828 6996
rect 22376 6944 22428 6996
rect 24400 6944 24452 6996
rect 17592 6876 17644 6928
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 15476 6672 15528 6724
rect 17132 6740 17184 6792
rect 17224 6740 17276 6792
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 17592 6740 17644 6749
rect 17684 6740 17736 6792
rect 17776 6740 17828 6792
rect 22192 6876 22244 6928
rect 23848 6876 23900 6928
rect 24032 6876 24084 6928
rect 24124 6876 24176 6928
rect 20076 6808 20128 6860
rect 22744 6808 22796 6860
rect 21916 6740 21968 6792
rect 11152 6604 11204 6613
rect 12164 6604 12216 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 17132 6604 17184 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 17960 6647 18012 6656
rect 17960 6613 17969 6647
rect 17969 6613 18003 6647
rect 18003 6613 18012 6647
rect 17960 6604 18012 6613
rect 24216 6740 24268 6792
rect 24308 6672 24360 6724
rect 25320 6672 25372 6724
rect 5151 6502 5203 6554
rect 5215 6502 5267 6554
rect 5279 6502 5331 6554
rect 5343 6502 5395 6554
rect 5407 6502 5459 6554
rect 12234 6502 12286 6554
rect 12298 6502 12350 6554
rect 12362 6502 12414 6554
rect 12426 6502 12478 6554
rect 12490 6502 12542 6554
rect 19317 6502 19369 6554
rect 19381 6502 19433 6554
rect 19445 6502 19497 6554
rect 19509 6502 19561 6554
rect 19573 6502 19625 6554
rect 26400 6502 26452 6554
rect 26464 6502 26516 6554
rect 26528 6502 26580 6554
rect 26592 6502 26644 6554
rect 26656 6502 26708 6554
rect 5080 6400 5132 6452
rect 5908 6400 5960 6452
rect 6276 6400 6328 6452
rect 7472 6400 7524 6452
rect 10232 6400 10284 6452
rect 11428 6400 11480 6452
rect 12164 6400 12216 6452
rect 6828 6332 6880 6384
rect 9864 6332 9916 6384
rect 10600 6332 10652 6384
rect 2688 6264 2740 6316
rect 7104 6264 7156 6316
rect 7196 6264 7248 6316
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 5724 6196 5776 6248
rect 6736 6196 6788 6248
rect 9680 6196 9732 6248
rect 10140 6264 10192 6316
rect 10416 6264 10468 6316
rect 10508 6196 10560 6248
rect 6092 6128 6144 6180
rect 8116 6128 8168 6180
rect 10968 6307 11020 6316
rect 10968 6273 10983 6307
rect 10983 6273 11017 6307
rect 11017 6273 11020 6307
rect 10968 6264 11020 6273
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 14096 6400 14148 6452
rect 16580 6400 16632 6452
rect 17776 6400 17828 6452
rect 17960 6400 18012 6452
rect 20076 6443 20128 6452
rect 20076 6409 20085 6443
rect 20085 6409 20119 6443
rect 20119 6409 20128 6443
rect 20076 6400 20128 6409
rect 28724 6400 28776 6452
rect 14188 6332 14240 6384
rect 15476 6375 15528 6384
rect 15476 6341 15485 6375
rect 15485 6341 15519 6375
rect 15519 6341 15528 6375
rect 15476 6332 15528 6341
rect 16856 6332 16908 6384
rect 17868 6332 17920 6384
rect 20076 6264 20128 6316
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 9772 6060 9824 6112
rect 11152 6128 11204 6180
rect 12624 6196 12676 6248
rect 13452 6239 13504 6248
rect 13452 6205 13461 6239
rect 13461 6205 13495 6239
rect 13495 6205 13504 6239
rect 13452 6196 13504 6205
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 17592 6060 17644 6112
rect 20444 6060 20496 6112
rect 4491 5958 4543 6010
rect 4555 5958 4607 6010
rect 4619 5958 4671 6010
rect 4683 5958 4735 6010
rect 4747 5958 4799 6010
rect 11574 5958 11626 6010
rect 11638 5958 11690 6010
rect 11702 5958 11754 6010
rect 11766 5958 11818 6010
rect 11830 5958 11882 6010
rect 18657 5958 18709 6010
rect 18721 5958 18773 6010
rect 18785 5958 18837 6010
rect 18849 5958 18901 6010
rect 18913 5958 18965 6010
rect 25740 5958 25792 6010
rect 25804 5958 25856 6010
rect 25868 5958 25920 6010
rect 25932 5958 25984 6010
rect 25996 5958 26048 6010
rect 6552 5856 6604 5908
rect 7196 5856 7248 5908
rect 5724 5831 5776 5840
rect 5724 5797 5733 5831
rect 5733 5797 5767 5831
rect 5767 5797 5776 5831
rect 5724 5788 5776 5797
rect 2688 5720 2740 5772
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 7288 5720 7340 5772
rect 10048 5856 10100 5908
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 16948 5856 17000 5908
rect 9864 5720 9916 5772
rect 10140 5763 10192 5772
rect 10140 5729 10149 5763
rect 10149 5729 10183 5763
rect 10183 5729 10192 5763
rect 10140 5720 10192 5729
rect 17224 5788 17276 5840
rect 11428 5720 11480 5772
rect 7012 5584 7064 5636
rect 7104 5584 7156 5636
rect 10508 5652 10560 5704
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 17408 5720 17460 5772
rect 17500 5652 17552 5704
rect 18512 5720 18564 5772
rect 9312 5516 9364 5568
rect 11336 5584 11388 5636
rect 11428 5627 11480 5636
rect 11428 5593 11437 5627
rect 11437 5593 11471 5627
rect 11471 5593 11480 5627
rect 11428 5584 11480 5593
rect 16028 5584 16080 5636
rect 17776 5584 17828 5636
rect 18420 5697 18472 5704
rect 18420 5663 18429 5697
rect 18429 5663 18463 5697
rect 18463 5663 18472 5697
rect 18420 5652 18472 5663
rect 9680 5516 9732 5568
rect 9772 5559 9824 5568
rect 9772 5525 9781 5559
rect 9781 5525 9815 5559
rect 9815 5525 9824 5559
rect 9772 5516 9824 5525
rect 10140 5516 10192 5568
rect 11152 5516 11204 5568
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 17960 5516 18012 5568
rect 18236 5516 18288 5568
rect 5151 5414 5203 5466
rect 5215 5414 5267 5466
rect 5279 5414 5331 5466
rect 5343 5414 5395 5466
rect 5407 5414 5459 5466
rect 12234 5414 12286 5466
rect 12298 5414 12350 5466
rect 12362 5414 12414 5466
rect 12426 5414 12478 5466
rect 12490 5414 12542 5466
rect 19317 5414 19369 5466
rect 19381 5414 19433 5466
rect 19445 5414 19497 5466
rect 19509 5414 19561 5466
rect 19573 5414 19625 5466
rect 26400 5414 26452 5466
rect 26464 5414 26516 5466
rect 26528 5414 26580 5466
rect 26592 5414 26644 5466
rect 26656 5414 26708 5466
rect 8208 5312 8260 5364
rect 7104 5244 7156 5296
rect 8024 5244 8076 5296
rect 6276 5176 6328 5228
rect 8944 5312 8996 5364
rect 9772 5176 9824 5228
rect 10508 5244 10560 5296
rect 10232 5176 10284 5228
rect 12624 5312 12676 5364
rect 13820 5312 13872 5364
rect 16488 5312 16540 5364
rect 17224 5312 17276 5364
rect 17316 5355 17368 5364
rect 17316 5321 17325 5355
rect 17325 5321 17359 5355
rect 17359 5321 17368 5355
rect 17316 5312 17368 5321
rect 10140 5108 10192 5160
rect 10692 5108 10744 5160
rect 9680 5040 9732 5092
rect 11796 5176 11848 5228
rect 11336 5108 11388 5160
rect 12440 5108 12492 5160
rect 14188 5176 14240 5228
rect 16120 5176 16172 5228
rect 17040 5176 17092 5228
rect 17408 5176 17460 5228
rect 17684 5176 17736 5228
rect 17868 5176 17920 5228
rect 12716 5108 12768 5160
rect 18236 5219 18288 5228
rect 18236 5185 18245 5219
rect 18245 5185 18279 5219
rect 18279 5185 18288 5219
rect 18236 5176 18288 5185
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 20260 5312 20312 5364
rect 28264 5355 28316 5364
rect 28264 5321 28273 5355
rect 28273 5321 28307 5355
rect 28307 5321 28316 5355
rect 28264 5312 28316 5321
rect 18420 5108 18472 5160
rect 17408 5040 17460 5092
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 17132 4972 17184 5024
rect 18052 5040 18104 5092
rect 18236 5040 18288 5092
rect 28080 5219 28132 5228
rect 28080 5185 28089 5219
rect 28089 5185 28123 5219
rect 28123 5185 28132 5219
rect 28080 5176 28132 5185
rect 17868 5015 17920 5024
rect 17868 4981 17877 5015
rect 17877 4981 17911 5015
rect 17911 4981 17920 5015
rect 17868 4972 17920 4981
rect 17960 4972 18012 5024
rect 19064 4972 19116 5024
rect 19524 4972 19576 5024
rect 20720 4972 20772 5024
rect 4491 4870 4543 4922
rect 4555 4870 4607 4922
rect 4619 4870 4671 4922
rect 4683 4870 4735 4922
rect 4747 4870 4799 4922
rect 11574 4870 11626 4922
rect 11638 4870 11690 4922
rect 11702 4870 11754 4922
rect 11766 4870 11818 4922
rect 11830 4870 11882 4922
rect 18657 4870 18709 4922
rect 18721 4870 18773 4922
rect 18785 4870 18837 4922
rect 18849 4870 18901 4922
rect 18913 4870 18965 4922
rect 25740 4870 25792 4922
rect 25804 4870 25856 4922
rect 25868 4870 25920 4922
rect 25932 4870 25984 4922
rect 25996 4870 26048 4922
rect 10232 4768 10284 4820
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 11060 4768 11112 4820
rect 11428 4768 11480 4820
rect 16396 4768 16448 4820
rect 16488 4768 16540 4820
rect 16948 4811 17000 4820
rect 16948 4777 16957 4811
rect 16957 4777 16991 4811
rect 16991 4777 17000 4811
rect 16948 4768 17000 4777
rect 17592 4811 17644 4820
rect 17592 4777 17601 4811
rect 17601 4777 17635 4811
rect 17635 4777 17644 4811
rect 17592 4768 17644 4777
rect 17776 4811 17828 4820
rect 17776 4777 17785 4811
rect 17785 4777 17819 4811
rect 17819 4777 17828 4811
rect 17776 4768 17828 4777
rect 17868 4768 17920 4820
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 16120 4700 16172 4752
rect 19800 4768 19852 4820
rect 28080 4768 28132 4820
rect 16028 4632 16080 4684
rect 11336 4564 11388 4616
rect 12992 4564 13044 4616
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 17500 4632 17552 4684
rect 17776 4632 17828 4684
rect 17868 4632 17920 4684
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 20076 4700 20128 4752
rect 16488 4607 16540 4616
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 14004 4496 14056 4548
rect 16212 4539 16264 4548
rect 16212 4505 16221 4539
rect 16221 4505 16255 4539
rect 16255 4505 16264 4539
rect 16212 4496 16264 4505
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 16672 4496 16724 4548
rect 19340 4632 19392 4684
rect 19432 4675 19484 4684
rect 19432 4641 19442 4675
rect 19442 4641 19476 4675
rect 19476 4641 19484 4675
rect 19432 4632 19484 4641
rect 19524 4675 19576 4684
rect 19524 4641 19533 4675
rect 19533 4641 19567 4675
rect 19567 4641 19576 4675
rect 19524 4632 19576 4641
rect 19248 4564 19300 4616
rect 19800 4564 19852 4616
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 20444 4564 20496 4616
rect 20720 4607 20772 4616
rect 20720 4573 20729 4607
rect 20729 4573 20763 4607
rect 20763 4573 20772 4607
rect 20720 4564 20772 4573
rect 6460 4428 6512 4480
rect 16856 4428 16908 4480
rect 17132 4471 17184 4480
rect 17132 4437 17141 4471
rect 17141 4437 17175 4471
rect 17175 4437 17184 4471
rect 17132 4428 17184 4437
rect 17224 4471 17276 4480
rect 17224 4437 17233 4471
rect 17233 4437 17267 4471
rect 17267 4437 17276 4471
rect 17224 4428 17276 4437
rect 18052 4428 18104 4480
rect 18328 4428 18380 4480
rect 19432 4428 19484 4480
rect 19800 4428 19852 4480
rect 5151 4326 5203 4378
rect 5215 4326 5267 4378
rect 5279 4326 5331 4378
rect 5343 4326 5395 4378
rect 5407 4326 5459 4378
rect 12234 4326 12286 4378
rect 12298 4326 12350 4378
rect 12362 4326 12414 4378
rect 12426 4326 12478 4378
rect 12490 4326 12542 4378
rect 19317 4326 19369 4378
rect 19381 4326 19433 4378
rect 19445 4326 19497 4378
rect 19509 4326 19561 4378
rect 19573 4326 19625 4378
rect 26400 4326 26452 4378
rect 26464 4326 26516 4378
rect 26528 4326 26580 4378
rect 26592 4326 26644 4378
rect 26656 4326 26708 4378
rect 2412 4224 2464 4276
rect 12624 4224 12676 4276
rect 14832 4224 14884 4276
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 12992 4088 13044 4140
rect 3516 3952 3568 4004
rect 13360 4020 13412 4072
rect 14096 4063 14148 4072
rect 14096 4029 14105 4063
rect 14105 4029 14139 4063
rect 14139 4029 14148 4063
rect 14096 4020 14148 4029
rect 14648 4088 14700 4140
rect 15200 4088 15252 4140
rect 16396 4224 16448 4276
rect 16856 4224 16908 4276
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 13084 3884 13136 3936
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 13912 3884 13964 3936
rect 14464 3952 14516 4004
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16580 4088 16632 4140
rect 16948 4156 17000 4208
rect 17132 4088 17184 4140
rect 17224 4088 17276 4140
rect 19708 4224 19760 4276
rect 20444 4224 20496 4276
rect 18420 4088 18472 4140
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 19800 4156 19852 4208
rect 17316 3952 17368 4004
rect 17500 4020 17552 4072
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 24308 4156 24360 4208
rect 24492 4088 24544 4140
rect 19892 3952 19944 4004
rect 16488 3884 16540 3936
rect 17408 3884 17460 3936
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 24400 3927 24452 3936
rect 24400 3893 24409 3927
rect 24409 3893 24443 3927
rect 24443 3893 24452 3927
rect 24400 3884 24452 3893
rect 24952 3927 25004 3936
rect 24952 3893 24961 3927
rect 24961 3893 24995 3927
rect 24995 3893 25004 3927
rect 24952 3884 25004 3893
rect 4491 3782 4543 3834
rect 4555 3782 4607 3834
rect 4619 3782 4671 3834
rect 4683 3782 4735 3834
rect 4747 3782 4799 3834
rect 11574 3782 11626 3834
rect 11638 3782 11690 3834
rect 11702 3782 11754 3834
rect 11766 3782 11818 3834
rect 11830 3782 11882 3834
rect 18657 3782 18709 3834
rect 18721 3782 18773 3834
rect 18785 3782 18837 3834
rect 18849 3782 18901 3834
rect 18913 3782 18965 3834
rect 25740 3782 25792 3834
rect 25804 3782 25856 3834
rect 25868 3782 25920 3834
rect 25932 3782 25984 3834
rect 25996 3782 26048 3834
rect 2228 3680 2280 3732
rect 12624 3723 12676 3732
rect 12624 3689 12633 3723
rect 12633 3689 12667 3723
rect 12667 3689 12676 3723
rect 12624 3680 12676 3689
rect 12900 3544 12952 3596
rect 940 3340 992 3392
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 12808 3383 12860 3392
rect 12808 3349 12817 3383
rect 12817 3349 12851 3383
rect 12851 3349 12860 3383
rect 12808 3340 12860 3349
rect 14648 3680 14700 3732
rect 13912 3612 13964 3664
rect 14004 3612 14056 3664
rect 15108 3655 15160 3664
rect 15108 3621 15117 3655
rect 15117 3621 15151 3655
rect 15151 3621 15160 3655
rect 15108 3612 15160 3621
rect 15660 3612 15712 3664
rect 13636 3544 13688 3596
rect 13360 3476 13412 3528
rect 13544 3476 13596 3528
rect 14096 3544 14148 3596
rect 13820 3476 13872 3528
rect 13728 3340 13780 3392
rect 13912 3408 13964 3460
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 15292 3476 15344 3528
rect 16580 3544 16632 3596
rect 17316 3476 17368 3528
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 17776 3476 17828 3528
rect 18880 3612 18932 3664
rect 24400 3680 24452 3732
rect 24952 3680 25004 3732
rect 20168 3544 20220 3596
rect 18512 3476 18564 3528
rect 22100 3408 22152 3460
rect 14280 3340 14332 3392
rect 15292 3383 15344 3392
rect 15292 3349 15301 3383
rect 15301 3349 15335 3383
rect 15335 3349 15344 3383
rect 15292 3340 15344 3349
rect 17500 3383 17552 3392
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 17592 3340 17644 3392
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 5151 3238 5203 3290
rect 5215 3238 5267 3290
rect 5279 3238 5331 3290
rect 5343 3238 5395 3290
rect 5407 3238 5459 3290
rect 12234 3238 12286 3290
rect 12298 3238 12350 3290
rect 12362 3238 12414 3290
rect 12426 3238 12478 3290
rect 12490 3238 12542 3290
rect 19317 3238 19369 3290
rect 19381 3238 19433 3290
rect 19445 3238 19497 3290
rect 19509 3238 19561 3290
rect 19573 3238 19625 3290
rect 26400 3238 26452 3290
rect 26464 3238 26516 3290
rect 26528 3238 26580 3290
rect 26592 3238 26644 3290
rect 26656 3238 26708 3290
rect 12992 3179 13044 3188
rect 12992 3145 13001 3179
rect 13001 3145 13035 3179
rect 13035 3145 13044 3179
rect 12992 3136 13044 3145
rect 13084 3136 13136 3188
rect 15108 3136 15160 3188
rect 17500 3136 17552 3188
rect 17592 3179 17644 3188
rect 17592 3145 17601 3179
rect 17601 3145 17635 3179
rect 17635 3145 17644 3179
rect 17592 3136 17644 3145
rect 17684 3136 17736 3188
rect 18788 3136 18840 3188
rect 14096 3068 14148 3120
rect 13544 3000 13596 3052
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 13820 3000 13872 3052
rect 13912 3000 13964 3052
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 15292 3068 15344 3120
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14648 3000 14700 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 17500 2975 17552 2984
rect 17500 2941 17509 2975
rect 17509 2941 17543 2975
rect 17543 2941 17552 2975
rect 17500 2932 17552 2941
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 17960 2975 18012 2984
rect 17960 2941 17969 2975
rect 17969 2941 18003 2975
rect 18003 2941 18012 2975
rect 17960 2932 18012 2941
rect 19064 3000 19116 3052
rect 13360 2864 13412 2916
rect 13176 2839 13228 2848
rect 13176 2805 13185 2839
rect 13185 2805 13219 2839
rect 13219 2805 13228 2839
rect 13176 2796 13228 2805
rect 17132 2796 17184 2848
rect 19892 2796 19944 2848
rect 29000 2839 29052 2848
rect 29000 2805 29009 2839
rect 29009 2805 29043 2839
rect 29043 2805 29052 2839
rect 29000 2796 29052 2805
rect 4491 2694 4543 2746
rect 4555 2694 4607 2746
rect 4619 2694 4671 2746
rect 4683 2694 4735 2746
rect 4747 2694 4799 2746
rect 11574 2694 11626 2746
rect 11638 2694 11690 2746
rect 11702 2694 11754 2746
rect 11766 2694 11818 2746
rect 11830 2694 11882 2746
rect 18657 2694 18709 2746
rect 18721 2694 18773 2746
rect 18785 2694 18837 2746
rect 18849 2694 18901 2746
rect 18913 2694 18965 2746
rect 25740 2694 25792 2746
rect 25804 2694 25856 2746
rect 25868 2694 25920 2746
rect 25932 2694 25984 2746
rect 25996 2694 26048 2746
rect 2228 2388 2280 2440
rect 12808 2592 12860 2644
rect 13268 2592 13320 2644
rect 13176 2388 13228 2440
rect 13728 2388 13780 2440
rect 13820 2388 13872 2440
rect 17500 2320 17552 2372
rect 20076 2320 20128 2372
rect 22100 2363 22152 2372
rect 22100 2329 22109 2363
rect 22109 2329 22143 2363
rect 22143 2329 22152 2363
rect 22100 2320 22152 2329
rect 25228 2388 25280 2440
rect 28540 2388 28592 2440
rect 27068 2320 27120 2372
rect 29644 2320 29696 2372
rect 20 2252 72 2304
rect 3424 2252 3476 2304
rect 7104 2252 7156 2304
rect 11152 2252 11204 2304
rect 14924 2252 14976 2304
rect 18880 2252 18932 2304
rect 22008 2252 22060 2304
rect 26148 2252 26200 2304
rect 5151 2150 5203 2202
rect 5215 2150 5267 2202
rect 5279 2150 5331 2202
rect 5343 2150 5395 2202
rect 5407 2150 5459 2202
rect 12234 2150 12286 2202
rect 12298 2150 12350 2202
rect 12362 2150 12414 2202
rect 12426 2150 12478 2202
rect 12490 2150 12542 2202
rect 19317 2150 19369 2202
rect 19381 2150 19433 2202
rect 19445 2150 19497 2202
rect 19509 2150 19561 2202
rect 19573 2150 19625 2202
rect 26400 2150 26452 2202
rect 26464 2150 26516 2202
rect 26528 2150 26580 2202
rect 26592 2150 26644 2202
rect 26656 2150 26708 2202
<< metal2 >>
rect 2594 32042 2650 32725
rect 6458 32042 6514 32725
rect 2594 32014 2728 32042
rect 2594 31925 2650 32014
rect 1582 30968 1638 30977
rect 1582 30903 1638 30912
rect 1596 30258 1624 30903
rect 2700 30274 2728 32014
rect 6458 32014 6776 32042
rect 6458 31925 6514 32014
rect 5151 30492 5459 30501
rect 5151 30490 5157 30492
rect 5213 30490 5237 30492
rect 5293 30490 5317 30492
rect 5373 30490 5397 30492
rect 5453 30490 5459 30492
rect 5213 30438 5215 30490
rect 5395 30438 5397 30490
rect 5151 30436 5157 30438
rect 5213 30436 5237 30438
rect 5293 30436 5317 30438
rect 5373 30436 5397 30438
rect 5453 30436 5459 30438
rect 5151 30427 5459 30436
rect 6748 30394 6776 32014
rect 9678 31925 9734 32725
rect 13542 32042 13598 32725
rect 13542 32014 13768 32042
rect 13542 31925 13598 32014
rect 6736 30388 6788 30394
rect 6736 30330 6788 30336
rect 9692 30326 9720 31925
rect 12234 30492 12542 30501
rect 12234 30490 12240 30492
rect 12296 30490 12320 30492
rect 12376 30490 12400 30492
rect 12456 30490 12480 30492
rect 12536 30490 12542 30492
rect 12296 30438 12298 30490
rect 12478 30438 12480 30490
rect 12234 30436 12240 30438
rect 12296 30436 12320 30438
rect 12376 30436 12400 30438
rect 12456 30436 12480 30438
rect 12536 30436 12542 30438
rect 12234 30427 12542 30436
rect 9680 30320 9732 30326
rect 1584 30252 1636 30258
rect 2700 30246 2912 30274
rect 9680 30262 9732 30268
rect 13740 30274 13768 32014
rect 17406 31925 17462 32725
rect 21270 31925 21326 32725
rect 25134 32042 25190 32725
rect 25134 32014 25452 32042
rect 25134 31925 25190 32014
rect 1584 30194 1636 30200
rect 2884 30054 2912 30246
rect 3332 30252 3384 30258
rect 3332 30194 3384 30200
rect 6092 30252 6144 30258
rect 6092 30194 6144 30200
rect 9864 30252 9916 30258
rect 13740 30246 13860 30274
rect 9864 30194 9916 30200
rect 1584 30048 1636 30054
rect 1584 29990 1636 29996
rect 2872 30048 2924 30054
rect 2872 29990 2924 29996
rect 1596 29238 1624 29990
rect 1584 29232 1636 29238
rect 1584 29174 1636 29180
rect 3056 29232 3108 29238
rect 3240 29232 3292 29238
rect 3108 29192 3240 29220
rect 3056 29174 3108 29180
rect 3240 29174 3292 29180
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 3160 27538 3188 28970
rect 3148 27532 3200 27538
rect 3148 27474 3200 27480
rect 1492 27396 1544 27402
rect 1492 27338 1544 27344
rect 940 27328 992 27334
rect 938 27296 940 27305
rect 992 27296 994 27305
rect 938 27231 994 27240
rect 1504 26586 1532 27338
rect 3056 27328 3108 27334
rect 3056 27270 3108 27276
rect 1492 26580 1544 26586
rect 1492 26522 1544 26528
rect 2412 26376 2464 26382
rect 2412 26318 2464 26324
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1504 23089 1532 23666
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 1636 23488 1638 23497
rect 1582 23423 1638 23432
rect 1490 23080 1546 23089
rect 1490 23015 1546 23024
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1872 19854 1900 20878
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1582 19544 1638 19553
rect 1582 19479 1584 19488
rect 1636 19479 1638 19488
rect 1584 19450 1636 19456
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 940 16108 992 16114
rect 940 16050 992 16056
rect 952 15745 980 16050
rect 1412 16046 1440 16526
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 938 15736 994 15745
rect 938 15671 994 15680
rect 1412 15570 1440 15982
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 14958 1440 15506
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 13938 1440 14894
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 12850 1440 13874
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 1504 6361 1532 19314
rect 1872 18426 1900 19790
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 2424 16574 2452 26318
rect 3068 25158 3096 27270
rect 3056 25152 3108 25158
rect 3056 25094 3108 25100
rect 3344 22094 3372 30194
rect 4491 29948 4799 29957
rect 4491 29946 4497 29948
rect 4553 29946 4577 29948
rect 4633 29946 4657 29948
rect 4713 29946 4737 29948
rect 4793 29946 4799 29948
rect 4553 29894 4555 29946
rect 4735 29894 4737 29946
rect 4491 29892 4497 29894
rect 4553 29892 4577 29894
rect 4633 29892 4657 29894
rect 4713 29892 4737 29894
rect 4793 29892 4799 29894
rect 4491 29883 4799 29892
rect 4988 29640 5040 29646
rect 5172 29640 5224 29646
rect 4988 29582 5040 29588
rect 5092 29588 5172 29594
rect 5092 29582 5224 29588
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5724 29640 5776 29646
rect 5724 29582 5776 29588
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 3516 29096 3568 29102
rect 3516 29038 3568 29044
rect 3528 28218 3556 29038
rect 4160 28960 4212 28966
rect 4160 28902 4212 28908
rect 4172 28558 4200 28902
rect 4491 28860 4799 28869
rect 4491 28858 4497 28860
rect 4553 28858 4577 28860
rect 4633 28858 4657 28860
rect 4713 28858 4737 28860
rect 4793 28858 4799 28860
rect 4553 28806 4555 28858
rect 4735 28806 4737 28858
rect 4491 28804 4497 28806
rect 4553 28804 4577 28806
rect 4633 28804 4657 28806
rect 4713 28804 4737 28806
rect 4793 28804 4799 28806
rect 4491 28795 4799 28804
rect 4252 28620 4304 28626
rect 4252 28562 4304 28568
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 3608 28416 3660 28422
rect 3608 28358 3660 28364
rect 3620 28218 3648 28358
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3620 27674 3648 28018
rect 4172 27878 4200 28494
rect 4160 27872 4212 27878
rect 4160 27814 4212 27820
rect 3608 27668 3660 27674
rect 3608 27610 3660 27616
rect 4172 25362 4200 27814
rect 4264 27538 4292 28562
rect 4908 28490 4936 29446
rect 5000 28966 5028 29582
rect 5092 29566 5212 29582
rect 4988 28960 5040 28966
rect 4988 28902 5040 28908
rect 4896 28484 4948 28490
rect 4896 28426 4948 28432
rect 5000 28422 5028 28902
rect 5092 28626 5120 29566
rect 5151 29404 5459 29413
rect 5151 29402 5157 29404
rect 5213 29402 5237 29404
rect 5293 29402 5317 29404
rect 5373 29402 5397 29404
rect 5453 29402 5459 29404
rect 5213 29350 5215 29402
rect 5395 29350 5397 29402
rect 5151 29348 5157 29350
rect 5213 29348 5237 29350
rect 5293 29348 5317 29350
rect 5373 29348 5397 29350
rect 5453 29348 5459 29350
rect 5151 29339 5459 29348
rect 5644 29102 5672 29582
rect 5632 29096 5684 29102
rect 5632 29038 5684 29044
rect 5172 29028 5224 29034
rect 5172 28970 5224 28976
rect 5184 28762 5212 28970
rect 5736 28762 5764 29582
rect 6000 29572 6052 29578
rect 6000 29514 6052 29520
rect 5816 29504 5868 29510
rect 5816 29446 5868 29452
rect 5908 29504 5960 29510
rect 5908 29446 5960 29452
rect 5172 28756 5224 28762
rect 5172 28698 5224 28704
rect 5724 28756 5776 28762
rect 5724 28698 5776 28704
rect 5080 28620 5132 28626
rect 5080 28562 5132 28568
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 4252 27532 4304 27538
rect 4252 27474 4304 27480
rect 4356 27470 4384 28358
rect 4491 27772 4799 27781
rect 4491 27770 4497 27772
rect 4553 27770 4577 27772
rect 4633 27770 4657 27772
rect 4713 27770 4737 27772
rect 4793 27770 4799 27772
rect 4553 27718 4555 27770
rect 4735 27718 4737 27770
rect 4491 27716 4497 27718
rect 4553 27716 4577 27718
rect 4633 27716 4657 27718
rect 4713 27716 4737 27718
rect 4793 27716 4799 27718
rect 4491 27707 4799 27716
rect 5000 27674 5028 28358
rect 4988 27668 5040 27674
rect 4988 27610 5040 27616
rect 4344 27464 4396 27470
rect 4344 27406 4396 27412
rect 5092 27402 5120 28562
rect 5151 28316 5459 28325
rect 5151 28314 5157 28316
rect 5213 28314 5237 28316
rect 5293 28314 5317 28316
rect 5373 28314 5397 28316
rect 5453 28314 5459 28316
rect 5213 28262 5215 28314
rect 5395 28262 5397 28314
rect 5151 28260 5157 28262
rect 5213 28260 5237 28262
rect 5293 28260 5317 28262
rect 5373 28260 5397 28262
rect 5453 28260 5459 28262
rect 5151 28251 5459 28260
rect 5632 28076 5684 28082
rect 5552 28036 5632 28064
rect 5080 27396 5132 27402
rect 5080 27338 5132 27344
rect 4491 26684 4799 26693
rect 4491 26682 4497 26684
rect 4553 26682 4577 26684
rect 4633 26682 4657 26684
rect 4713 26682 4737 26684
rect 4793 26682 4799 26684
rect 4553 26630 4555 26682
rect 4735 26630 4737 26682
rect 4491 26628 4497 26630
rect 4553 26628 4577 26630
rect 4633 26628 4657 26630
rect 4713 26628 4737 26630
rect 4793 26628 4799 26630
rect 4491 26619 4799 26628
rect 5092 25906 5120 27338
rect 5151 27228 5459 27237
rect 5151 27226 5157 27228
rect 5213 27226 5237 27228
rect 5293 27226 5317 27228
rect 5373 27226 5397 27228
rect 5453 27226 5459 27228
rect 5213 27174 5215 27226
rect 5395 27174 5397 27226
rect 5151 27172 5157 27174
rect 5213 27172 5237 27174
rect 5293 27172 5317 27174
rect 5373 27172 5397 27174
rect 5453 27172 5459 27174
rect 5151 27163 5459 27172
rect 5151 26140 5459 26149
rect 5151 26138 5157 26140
rect 5213 26138 5237 26140
rect 5293 26138 5317 26140
rect 5373 26138 5397 26140
rect 5453 26138 5459 26140
rect 5213 26086 5215 26138
rect 5395 26086 5397 26138
rect 5151 26084 5157 26086
rect 5213 26084 5237 26086
rect 5293 26084 5317 26086
rect 5373 26084 5397 26086
rect 5453 26084 5459 26086
rect 5151 26075 5459 26084
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 4344 25764 4396 25770
rect 4344 25706 4396 25712
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 4356 25294 4384 25706
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 4491 25596 4799 25605
rect 4491 25594 4497 25596
rect 4553 25594 4577 25596
rect 4633 25594 4657 25596
rect 4713 25594 4737 25596
rect 4793 25594 4799 25596
rect 4553 25542 4555 25594
rect 4735 25542 4737 25594
rect 4491 25540 4497 25542
rect 4553 25540 4577 25542
rect 4633 25540 4657 25542
rect 4713 25540 4737 25542
rect 4793 25540 4799 25542
rect 4491 25531 4799 25540
rect 5000 25362 5028 25638
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4620 25288 4672 25294
rect 5092 25242 5120 25842
rect 5460 25362 5488 25842
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 5460 25242 5488 25298
rect 4620 25230 4672 25236
rect 4528 25152 4580 25158
rect 4528 25094 4580 25100
rect 4540 24818 4568 25094
rect 4528 24812 4580 24818
rect 4528 24754 4580 24760
rect 4632 24750 4660 25230
rect 4896 25220 4948 25226
rect 4896 25162 4948 25168
rect 5000 25214 5120 25242
rect 5368 25214 5488 25242
rect 5552 25226 5580 28036
rect 5632 28018 5684 28024
rect 5828 27946 5856 29446
rect 5920 29306 5948 29446
rect 5908 29300 5960 29306
rect 5908 29242 5960 29248
rect 5920 28558 5948 29242
rect 5908 28552 5960 28558
rect 5908 28494 5960 28500
rect 5920 28082 5948 28494
rect 6012 28218 6040 29514
rect 6000 28212 6052 28218
rect 6000 28154 6052 28160
rect 5908 28076 5960 28082
rect 5908 28018 5960 28024
rect 5816 27940 5868 27946
rect 5816 27882 5868 27888
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5828 26042 5856 26182
rect 5816 26036 5868 26042
rect 5816 25978 5868 25984
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 5644 25702 5672 25842
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 5724 25696 5776 25702
rect 5724 25638 5776 25644
rect 5540 25220 5592 25226
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4816 24886 4844 25094
rect 4908 24954 4936 25162
rect 4896 24948 4948 24954
rect 4896 24890 4948 24896
rect 4804 24880 4856 24886
rect 4804 24822 4856 24828
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 3436 24410 3464 24686
rect 4491 24508 4799 24517
rect 4491 24506 4497 24508
rect 4553 24506 4577 24508
rect 4633 24506 4657 24508
rect 4713 24506 4737 24508
rect 4793 24506 4799 24508
rect 4553 24454 4555 24506
rect 4735 24454 4737 24506
rect 4491 24452 4497 24454
rect 4553 24452 4577 24454
rect 4633 24452 4657 24454
rect 4713 24452 4737 24454
rect 4793 24452 4799 24454
rect 4491 24443 4799 24452
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 4908 24274 4936 24890
rect 5000 24410 5028 25214
rect 5368 25158 5396 25214
rect 5540 25162 5592 25168
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5092 24818 5120 25094
rect 5151 25052 5459 25061
rect 5151 25050 5157 25052
rect 5213 25050 5237 25052
rect 5293 25050 5317 25052
rect 5373 25050 5397 25052
rect 5453 25050 5459 25052
rect 5213 24998 5215 25050
rect 5395 24998 5397 25050
rect 5151 24996 5157 24998
rect 5213 24996 5237 24998
rect 5293 24996 5317 24998
rect 5373 24996 5397 24998
rect 5453 24996 5459 24998
rect 5151 24987 5459 24996
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 5080 24676 5132 24682
rect 5080 24618 5132 24624
rect 4988 24404 5040 24410
rect 4988 24346 5040 24352
rect 4896 24268 4948 24274
rect 4896 24210 4948 24216
rect 5092 24154 5120 24618
rect 5552 24614 5580 25162
rect 5644 24818 5672 25638
rect 5736 24954 5764 25638
rect 5724 24948 5776 24954
rect 5724 24890 5776 24896
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5184 24342 5212 24550
rect 5172 24336 5224 24342
rect 5172 24278 5224 24284
rect 4908 24126 5120 24154
rect 5552 24154 5580 24550
rect 5552 24138 5672 24154
rect 5552 24132 5684 24138
rect 5552 24126 5632 24132
rect 4491 23420 4799 23429
rect 4491 23418 4497 23420
rect 4553 23418 4577 23420
rect 4633 23418 4657 23420
rect 4713 23418 4737 23420
rect 4793 23418 4799 23420
rect 4553 23366 4555 23418
rect 4735 23366 4737 23418
rect 4491 23364 4497 23366
rect 4553 23364 4577 23366
rect 4633 23364 4657 23366
rect 4713 23364 4737 23366
rect 4793 23364 4799 23366
rect 4491 23355 4799 23364
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 3344 22066 3556 22094
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3252 21554 3280 21830
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3252 17270 3280 21490
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3436 19786 3464 20742
rect 3424 19780 3476 19786
rect 3424 19722 3476 19728
rect 3436 18358 3464 19722
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3436 17610 3464 18158
rect 3424 17604 3476 17610
rect 3424 17546 3476 17552
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 2332 16546 2452 16574
rect 1676 16516 1728 16522
rect 1676 16458 1728 16464
rect 1688 16250 1716 16458
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 13530 1900 13806
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 12442 2084 12718
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 2226 11792 2282 11801
rect 2226 11727 2228 11736
rect 2280 11727 2282 11736
rect 2228 11698 2280 11704
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11218 2268 11494
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2148 10713 2176 11018
rect 2134 10704 2190 10713
rect 2134 10639 2190 10648
rect 2240 9654 2268 11154
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2240 9042 2268 9590
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2240 8634 2268 8978
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1688 7886 1716 8434
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 2332 6914 2360 16546
rect 3344 15570 3372 16934
rect 3436 16726 3464 17070
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3252 14006 3280 15438
rect 3240 14000 3292 14006
rect 3160 13960 3240 13988
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3068 12345 3096 13262
rect 3160 12850 3188 13960
rect 3240 13942 3292 13948
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3054 12336 3110 12345
rect 3054 12271 3110 12280
rect 3068 12238 3096 12271
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3160 11830 3188 12786
rect 3252 12238 3280 13126
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3160 11150 3188 11766
rect 3148 11144 3200 11150
rect 3146 11112 3148 11121
rect 3200 11112 3202 11121
rect 3146 11047 3202 11056
rect 3160 9674 3188 11047
rect 3160 9646 3372 9674
rect 3344 9586 3372 9646
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3344 9110 3372 9522
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3344 8634 3372 9046
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2332 6886 2452 6914
rect 1490 6352 1546 6361
rect 1490 6287 1546 6296
rect 2424 4282 2452 6886
rect 2700 6322 2728 8502
rect 3344 7886 3372 8570
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 5778 2728 6258
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2424 4049 2452 4082
rect 2410 4040 2466 4049
rect 3528 4010 3556 22066
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3712 21554 3740 22034
rect 4172 21690 4200 22374
rect 4491 22332 4799 22341
rect 4491 22330 4497 22332
rect 4553 22330 4577 22332
rect 4633 22330 4657 22332
rect 4713 22330 4737 22332
rect 4793 22330 4799 22332
rect 4553 22278 4555 22330
rect 4735 22278 4737 22330
rect 4491 22276 4497 22278
rect 4553 22276 4577 22278
rect 4633 22276 4657 22278
rect 4713 22276 4737 22278
rect 4793 22276 4799 22278
rect 4491 22267 4799 22276
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 4068 21616 4120 21622
rect 4264 21570 4292 21966
rect 4908 21962 4936 24126
rect 5632 24074 5684 24080
rect 5151 23964 5459 23973
rect 5151 23962 5157 23964
rect 5213 23962 5237 23964
rect 5293 23962 5317 23964
rect 5373 23962 5397 23964
rect 5453 23962 5459 23964
rect 5213 23910 5215 23962
rect 5395 23910 5397 23962
rect 5151 23908 5157 23910
rect 5213 23908 5237 23910
rect 5293 23908 5317 23910
rect 5373 23908 5397 23910
rect 5453 23908 5459 23910
rect 5151 23899 5459 23908
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 5080 22976 5132 22982
rect 5080 22918 5132 22924
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4896 21956 4948 21962
rect 4896 21898 4948 21904
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4068 21558 4120 21564
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 4080 21350 4108 21558
rect 4172 21542 4292 21570
rect 4344 21616 4396 21622
rect 4724 21593 4752 21830
rect 4908 21690 4936 21898
rect 4896 21684 4948 21690
rect 4896 21626 4948 21632
rect 4344 21558 4396 21564
rect 4710 21584 4766 21593
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 3712 21146 3740 21286
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3804 21010 3832 21286
rect 3792 21004 3844 21010
rect 3792 20946 3844 20952
rect 4080 20534 4108 21286
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3896 20058 3924 20198
rect 3988 20058 4016 20198
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3620 18290 3648 18702
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3712 18290 3740 18362
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3712 17746 3740 18226
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 3988 17202 4016 18566
rect 4068 17332 4120 17338
rect 4172 17320 4200 21542
rect 4356 20806 4384 21558
rect 4710 21519 4766 21528
rect 4491 21244 4799 21253
rect 4491 21242 4497 21244
rect 4553 21242 4577 21244
rect 4633 21242 4657 21244
rect 4713 21242 4737 21244
rect 4793 21242 4799 21244
rect 4553 21190 4555 21242
rect 4735 21190 4737 21242
rect 4491 21188 4497 21190
rect 4553 21188 4577 21190
rect 4633 21188 4657 21190
rect 4713 21188 4737 21190
rect 4793 21188 4799 21190
rect 4491 21179 4799 21188
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 4344 20528 4396 20534
rect 4264 20488 4344 20516
rect 4264 17785 4292 20488
rect 4344 20470 4396 20476
rect 4896 20392 4948 20398
rect 4894 20360 4896 20369
rect 4948 20360 4950 20369
rect 4894 20295 4950 20304
rect 4491 20156 4799 20165
rect 4491 20154 4497 20156
rect 4553 20154 4577 20156
rect 4633 20154 4657 20156
rect 4713 20154 4737 20156
rect 4793 20154 4799 20156
rect 4553 20102 4555 20154
rect 4735 20102 4737 20154
rect 4491 20100 4497 20102
rect 4553 20100 4577 20102
rect 4633 20100 4657 20102
rect 4713 20100 4737 20102
rect 4793 20100 4799 20102
rect 4491 20091 4799 20100
rect 4491 19068 4799 19077
rect 4491 19066 4497 19068
rect 4553 19066 4577 19068
rect 4633 19066 4657 19068
rect 4713 19066 4737 19068
rect 4793 19066 4799 19068
rect 4553 19014 4555 19066
rect 4735 19014 4737 19066
rect 4491 19012 4497 19014
rect 4553 19012 4577 19014
rect 4633 19012 4657 19014
rect 4713 19012 4737 19014
rect 4793 19012 4799 19014
rect 4491 19003 4799 19012
rect 4491 17980 4799 17989
rect 4491 17978 4497 17980
rect 4553 17978 4577 17980
rect 4633 17978 4657 17980
rect 4713 17978 4737 17980
rect 4793 17978 4799 17980
rect 4553 17926 4555 17978
rect 4735 17926 4737 17978
rect 4491 17924 4497 17926
rect 4553 17924 4577 17926
rect 4633 17924 4657 17926
rect 4713 17924 4737 17926
rect 4793 17924 4799 17926
rect 4491 17915 4799 17924
rect 4250 17776 4306 17785
rect 4250 17711 4306 17720
rect 4120 17292 4200 17320
rect 4068 17274 4120 17280
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3620 16794 3648 17138
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3620 14006 3648 16730
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3896 16114 3924 16458
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3896 15502 3924 16050
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3620 13530 3648 13942
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3620 12918 3648 13466
rect 3608 12912 3660 12918
rect 3608 12854 3660 12860
rect 3620 12102 3648 12854
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3896 12102 3924 12582
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3698 11384 3754 11393
rect 3698 11319 3754 11328
rect 3712 11150 3740 11319
rect 3896 11257 3924 12038
rect 3882 11248 3938 11257
rect 3882 11183 3884 11192
rect 3936 11183 3938 11192
rect 3884 11154 3936 11160
rect 3988 11150 4016 17002
rect 4080 16998 4108 17274
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 11286 4108 16934
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 15162 4200 15302
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4264 13308 4292 17711
rect 4528 17604 4580 17610
rect 4528 17546 4580 17552
rect 4540 17338 4568 17546
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4816 17134 4844 17478
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4491 16892 4799 16901
rect 4491 16890 4497 16892
rect 4553 16890 4577 16892
rect 4633 16890 4657 16892
rect 4713 16890 4737 16892
rect 4793 16890 4799 16892
rect 4553 16838 4555 16890
rect 4735 16838 4737 16890
rect 4491 16836 4497 16838
rect 4553 16836 4577 16838
rect 4633 16836 4657 16838
rect 4713 16836 4737 16838
rect 4793 16836 4799 16838
rect 4491 16827 4799 16836
rect 4908 16590 4936 20295
rect 5000 20262 5028 21966
rect 5092 21486 5120 22918
rect 5151 22876 5459 22885
rect 5151 22874 5157 22876
rect 5213 22874 5237 22876
rect 5293 22874 5317 22876
rect 5373 22874 5397 22876
rect 5453 22874 5459 22876
rect 5213 22822 5215 22874
rect 5395 22822 5397 22874
rect 5151 22820 5157 22822
rect 5213 22820 5237 22822
rect 5293 22820 5317 22822
rect 5373 22820 5397 22822
rect 5453 22820 5459 22822
rect 5151 22811 5459 22820
rect 5724 22568 5776 22574
rect 5724 22510 5776 22516
rect 5448 22092 5500 22098
rect 5448 22034 5500 22040
rect 5460 22001 5488 22034
rect 5540 22024 5592 22030
rect 5446 21992 5502 22001
rect 5540 21966 5592 21972
rect 5446 21927 5502 21936
rect 5151 21788 5459 21797
rect 5151 21786 5157 21788
rect 5213 21786 5237 21788
rect 5293 21786 5317 21788
rect 5373 21786 5397 21788
rect 5453 21786 5459 21788
rect 5213 21734 5215 21786
rect 5395 21734 5397 21786
rect 5151 21732 5157 21734
rect 5213 21732 5237 21734
rect 5293 21732 5317 21734
rect 5373 21732 5397 21734
rect 5453 21732 5459 21734
rect 5151 21723 5459 21732
rect 5552 21690 5580 21966
rect 5630 21720 5686 21729
rect 5540 21684 5592 21690
rect 5630 21655 5632 21664
rect 5540 21626 5592 21632
rect 5684 21655 5686 21664
rect 5632 21626 5684 21632
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5552 20942 5580 21626
rect 5736 21146 5764 22510
rect 5828 21418 5856 23802
rect 5908 22976 5960 22982
rect 5908 22918 5960 22924
rect 5920 22710 5948 22918
rect 5908 22704 5960 22710
rect 5908 22646 5960 22652
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 6012 22098 6040 22510
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5920 21690 5948 21830
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 6000 21548 6052 21554
rect 5920 21508 6000 21536
rect 5816 21412 5868 21418
rect 5816 21354 5868 21360
rect 5920 21298 5948 21508
rect 6000 21490 6052 21496
rect 5828 21270 5948 21298
rect 5724 21140 5776 21146
rect 5724 21082 5776 21088
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5736 20806 5764 21082
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 5151 20700 5459 20709
rect 5151 20698 5157 20700
rect 5213 20698 5237 20700
rect 5293 20698 5317 20700
rect 5373 20698 5397 20700
rect 5453 20698 5459 20700
rect 5213 20646 5215 20698
rect 5395 20646 5397 20698
rect 5151 20644 5157 20646
rect 5213 20644 5237 20646
rect 5293 20644 5317 20646
rect 5373 20644 5397 20646
rect 5453 20644 5459 20646
rect 5151 20635 5459 20644
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 5151 19612 5459 19621
rect 5151 19610 5157 19612
rect 5213 19610 5237 19612
rect 5293 19610 5317 19612
rect 5373 19610 5397 19612
rect 5453 19610 5459 19612
rect 5213 19558 5215 19610
rect 5395 19558 5397 19610
rect 5151 19556 5157 19558
rect 5213 19556 5237 19558
rect 5293 19556 5317 19558
rect 5373 19556 5397 19558
rect 5453 19556 5459 19558
rect 5151 19547 5459 19556
rect 5828 19334 5856 21270
rect 5920 21078 5948 21270
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5644 19306 5856 19334
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 5000 17338 5028 19178
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5151 18524 5459 18533
rect 5151 18522 5157 18524
rect 5213 18522 5237 18524
rect 5293 18522 5317 18524
rect 5373 18522 5397 18524
rect 5453 18522 5459 18524
rect 5213 18470 5215 18522
rect 5395 18470 5397 18522
rect 5151 18468 5157 18470
rect 5213 18468 5237 18470
rect 5293 18468 5317 18470
rect 5373 18468 5397 18470
rect 5453 18468 5459 18470
rect 5151 18459 5459 18468
rect 5552 18358 5580 18566
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 5092 17338 5120 18090
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17678 5212 18022
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5151 17436 5459 17445
rect 5151 17434 5157 17436
rect 5213 17434 5237 17436
rect 5293 17434 5317 17436
rect 5373 17434 5397 17436
rect 5453 17434 5459 17436
rect 5213 17382 5215 17434
rect 5395 17382 5397 17434
rect 5151 17380 5157 17382
rect 5213 17380 5237 17382
rect 5293 17380 5317 17382
rect 5373 17380 5397 17382
rect 5453 17380 5459 17382
rect 5151 17371 5459 17380
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5264 17332 5316 17338
rect 5644 17320 5672 19306
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5828 17610 5856 18566
rect 5816 17604 5868 17610
rect 5816 17546 5868 17552
rect 5316 17292 5672 17320
rect 5264 17274 5316 17280
rect 5000 16810 5028 17274
rect 5644 17202 5672 17292
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5000 16782 5120 16810
rect 5184 16794 5212 17138
rect 5552 16794 5580 17138
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 4988 16720 5040 16726
rect 4988 16662 5040 16668
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 16250 4476 16390
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4356 15706 4384 15914
rect 4491 15804 4799 15813
rect 4491 15802 4497 15804
rect 4553 15802 4577 15804
rect 4633 15802 4657 15804
rect 4713 15802 4737 15804
rect 4793 15802 4799 15804
rect 4553 15750 4555 15802
rect 4735 15750 4737 15802
rect 4491 15748 4497 15750
rect 4553 15748 4577 15750
rect 4633 15748 4657 15750
rect 4713 15748 4737 15750
rect 4793 15748 4799 15750
rect 4491 15739 4799 15748
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4491 14716 4799 14725
rect 4491 14714 4497 14716
rect 4553 14714 4577 14716
rect 4633 14714 4657 14716
rect 4713 14714 4737 14716
rect 4793 14714 4799 14716
rect 4553 14662 4555 14714
rect 4735 14662 4737 14714
rect 4491 14660 4497 14662
rect 4553 14660 4577 14662
rect 4633 14660 4657 14662
rect 4713 14660 4737 14662
rect 4793 14660 4799 14662
rect 4491 14651 4799 14660
rect 4491 13628 4799 13637
rect 4491 13626 4497 13628
rect 4553 13626 4577 13628
rect 4633 13626 4657 13628
rect 4713 13626 4737 13628
rect 4793 13626 4799 13628
rect 4553 13574 4555 13626
rect 4735 13574 4737 13626
rect 4491 13572 4497 13574
rect 4553 13572 4577 13574
rect 4633 13572 4657 13574
rect 4713 13572 4737 13574
rect 4793 13572 4799 13574
rect 4491 13563 4799 13572
rect 4172 13280 4292 13308
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 9330 4016 11086
rect 4066 10840 4122 10849
rect 4172 10810 4200 13280
rect 4908 12968 4936 16526
rect 5000 16250 5028 16662
rect 5092 16590 5120 16782
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5092 16250 5120 16390
rect 5151 16348 5459 16357
rect 5151 16346 5157 16348
rect 5213 16346 5237 16348
rect 5293 16346 5317 16348
rect 5373 16346 5397 16348
rect 5453 16346 5459 16348
rect 5213 16294 5215 16346
rect 5395 16294 5397 16346
rect 5151 16292 5157 16294
rect 5213 16292 5237 16294
rect 5293 16292 5317 16294
rect 5373 16292 5397 16294
rect 5453 16292 5459 16294
rect 5151 16283 5459 16292
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5184 15366 5212 16050
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5151 15260 5459 15269
rect 5151 15258 5157 15260
rect 5213 15258 5237 15260
rect 5293 15258 5317 15260
rect 5373 15258 5397 15260
rect 5453 15258 5459 15260
rect 5213 15206 5215 15258
rect 5395 15206 5397 15258
rect 5151 15204 5157 15206
rect 5213 15204 5237 15206
rect 5293 15204 5317 15206
rect 5373 15204 5397 15206
rect 5453 15204 5459 15206
rect 5151 15195 5459 15204
rect 5356 15156 5408 15162
rect 5552 15144 5580 16390
rect 5736 16114 5764 16526
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5644 15162 5672 15982
rect 5736 15706 5764 16050
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5828 15638 5856 16934
rect 5920 16114 5948 20878
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 6012 17270 6040 18090
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 6104 17218 6132 30194
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 9036 29640 9088 29646
rect 9036 29582 9088 29588
rect 7564 29572 7616 29578
rect 7564 29514 7616 29520
rect 7288 29504 7340 29510
rect 7288 29446 7340 29452
rect 7472 29504 7524 29510
rect 7472 29446 7524 29452
rect 7300 29238 7328 29446
rect 7484 29306 7512 29446
rect 7472 29300 7524 29306
rect 7472 29242 7524 29248
rect 7104 29232 7156 29238
rect 7104 29174 7156 29180
rect 7288 29232 7340 29238
rect 7288 29174 7340 29180
rect 6184 29096 6236 29102
rect 6184 29038 6236 29044
rect 6196 28490 6224 29038
rect 7116 28762 7144 29174
rect 6460 28756 6512 28762
rect 6460 28698 6512 28704
rect 7104 28756 7156 28762
rect 7104 28698 7156 28704
rect 7208 28716 7420 28744
rect 6276 28688 6328 28694
rect 6276 28630 6328 28636
rect 6184 28484 6236 28490
rect 6184 28426 6236 28432
rect 6196 28218 6224 28426
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6288 28014 6316 28630
rect 6472 28558 6500 28698
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 7012 28552 7064 28558
rect 7064 28529 7144 28540
rect 7064 28520 7158 28529
rect 7064 28512 7102 28520
rect 7012 28494 7064 28500
rect 6368 28416 6420 28422
rect 6368 28358 6420 28364
rect 6276 28008 6328 28014
rect 6276 27950 6328 27956
rect 6380 27878 6408 28358
rect 6472 28082 6500 28494
rect 6828 28484 6880 28490
rect 7208 28490 7236 28716
rect 7102 28455 7158 28464
rect 7196 28484 7248 28490
rect 6828 28426 6880 28432
rect 7196 28426 7248 28432
rect 6840 28082 6868 28426
rect 7012 28416 7064 28422
rect 7012 28358 7064 28364
rect 7024 28082 7052 28358
rect 6460 28076 6512 28082
rect 6460 28018 6512 28024
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 7012 28076 7064 28082
rect 7012 28018 7064 28024
rect 7196 28076 7248 28082
rect 7196 28018 7248 28024
rect 7208 27946 7236 28018
rect 7196 27940 7248 27946
rect 7196 27882 7248 27888
rect 6368 27872 6420 27878
rect 6368 27814 6420 27820
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6380 27674 6408 27814
rect 6368 27668 6420 27674
rect 6368 27610 6420 27616
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6472 25974 6500 26318
rect 6460 25968 6512 25974
rect 6460 25910 6512 25916
rect 6368 25492 6420 25498
rect 6368 25434 6420 25440
rect 6380 24818 6408 25434
rect 6472 25158 6500 25910
rect 6564 25906 6592 27814
rect 7392 27606 7420 28716
rect 7484 28150 7512 29242
rect 7576 28994 7604 29514
rect 7748 29504 7800 29510
rect 7748 29446 7800 29452
rect 7656 29096 7708 29102
rect 7656 29038 7708 29044
rect 7668 28994 7696 29038
rect 7576 28966 7696 28994
rect 7668 28490 7696 28966
rect 7760 28762 7788 29446
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7748 28756 7800 28762
rect 7748 28698 7800 28704
rect 7564 28484 7616 28490
rect 7564 28426 7616 28432
rect 7656 28484 7708 28490
rect 7656 28426 7708 28432
rect 7748 28484 7800 28490
rect 7748 28426 7800 28432
rect 7576 28218 7604 28426
rect 7564 28212 7616 28218
rect 7564 28154 7616 28160
rect 7472 28144 7524 28150
rect 7472 28086 7524 28092
rect 7484 27962 7512 28086
rect 7564 28076 7616 28082
rect 7668 28064 7696 28426
rect 7616 28036 7696 28064
rect 7564 28018 7616 28024
rect 7760 27962 7788 28426
rect 7852 28150 7880 28902
rect 7840 28144 7892 28150
rect 7840 28086 7892 28092
rect 7484 27934 7788 27962
rect 7380 27600 7432 27606
rect 7380 27542 7432 27548
rect 7852 26926 7880 28086
rect 7932 27396 7984 27402
rect 7932 27338 7984 27344
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 7012 26308 7064 26314
rect 7012 26250 7064 26256
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 6828 25832 6880 25838
rect 6828 25774 6880 25780
rect 6840 25702 6868 25774
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6840 25498 6868 25638
rect 6828 25492 6880 25498
rect 6828 25434 6880 25440
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6472 24954 6500 25094
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 6380 24614 6408 24754
rect 6644 24744 6696 24750
rect 6644 24686 6696 24692
rect 6368 24608 6420 24614
rect 6368 24550 6420 24556
rect 6656 24410 6684 24686
rect 6932 24682 6960 25842
rect 7024 25498 7052 26250
rect 7196 25900 7248 25906
rect 7196 25842 7248 25848
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 6920 24676 6972 24682
rect 6920 24618 6972 24624
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 7024 24206 7052 25434
rect 7208 25226 7236 25842
rect 7748 25764 7800 25770
rect 7748 25706 7800 25712
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 7196 25220 7248 25226
rect 7196 25162 7248 25168
rect 7208 24886 7236 25162
rect 7196 24880 7248 24886
rect 7196 24822 7248 24828
rect 7300 24206 7328 25638
rect 7380 25152 7432 25158
rect 7380 25094 7432 25100
rect 7392 24818 7420 25094
rect 7576 24954 7604 25638
rect 7760 25498 7788 25706
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 7564 24948 7616 24954
rect 7564 24890 7616 24896
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7392 24410 7420 24754
rect 7668 24410 7696 24754
rect 7852 24750 7880 26862
rect 7944 26042 7972 27338
rect 8496 26738 8524 29582
rect 8760 28960 8812 28966
rect 8760 28902 8812 28908
rect 8772 28626 8800 28902
rect 8760 28620 8812 28626
rect 8760 28562 8812 28568
rect 8758 28520 8814 28529
rect 8758 28455 8760 28464
rect 8812 28455 8814 28464
rect 8760 28426 8812 28432
rect 8576 28416 8628 28422
rect 8576 28358 8628 28364
rect 8588 28218 8616 28358
rect 8576 28212 8628 28218
rect 8576 28154 8628 28160
rect 9048 28082 9076 29582
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 9784 28762 9812 29038
rect 9772 28756 9824 28762
rect 9772 28698 9824 28704
rect 9404 28620 9456 28626
rect 9404 28562 9456 28568
rect 9416 28218 9444 28562
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9312 28076 9364 28082
rect 9312 28018 9364 28024
rect 9324 27538 9352 28018
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9312 27532 9364 27538
rect 9312 27474 9364 27480
rect 9784 27470 9812 27950
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9036 27396 9088 27402
rect 9036 27338 9088 27344
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 8944 27328 8996 27334
rect 8944 27270 8996 27276
rect 8588 26926 8616 27270
rect 8956 27130 8984 27270
rect 9048 27130 9076 27338
rect 9784 27130 9812 27406
rect 8944 27124 8996 27130
rect 8944 27066 8996 27072
rect 9036 27124 9088 27130
rect 9036 27066 9088 27072
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 9588 26988 9640 26994
rect 9588 26930 9640 26936
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8404 26710 8524 26738
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 8404 25294 8432 26710
rect 8588 25838 8616 26862
rect 9600 26382 9628 26930
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8760 25696 8812 25702
rect 8760 25638 8812 25644
rect 8772 25498 8800 25638
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7656 24404 7708 24410
rect 7656 24346 7708 24352
rect 7852 24274 7880 24686
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 6564 23186 6592 24142
rect 9140 23662 9168 25230
rect 9600 24886 9628 26318
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9140 23322 9168 23598
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6196 21690 6224 23054
rect 9140 22642 9168 23258
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 9324 22778 9352 22986
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 7104 22636 7156 22642
rect 6932 22596 7104 22624
rect 6932 22137 6960 22596
rect 7104 22578 7156 22584
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 7300 22234 7328 22374
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 6918 22128 6974 22137
rect 6368 22092 6420 22098
rect 7392 22094 7420 22374
rect 7668 22234 7696 22510
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 6918 22063 6974 22072
rect 7208 22066 7420 22094
rect 6368 22034 6420 22040
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6380 21146 6408 22034
rect 6932 22001 6960 22063
rect 6918 21992 6974 22001
rect 6918 21927 6974 21936
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7116 21622 7144 21830
rect 7104 21616 7156 21622
rect 7208 21593 7236 22066
rect 7104 21558 7156 21564
rect 7194 21584 7250 21593
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6196 20602 6224 20810
rect 6184 20596 6236 20602
rect 6184 20538 6236 20544
rect 6196 18222 6224 20538
rect 6380 20398 6408 21082
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6380 18834 6408 20334
rect 6472 19854 6500 21286
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6656 20058 6684 20334
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6460 19848 6512 19854
rect 6460 19790 6512 19796
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6564 19310 6592 19722
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6460 19236 6512 19242
rect 6460 19178 6512 19184
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6472 18766 6500 19178
rect 6564 18902 6592 19246
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 6288 18426 6316 18634
rect 6748 18578 6776 20878
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 19854 6960 20742
rect 7116 20534 7144 21558
rect 7194 21519 7250 21528
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7392 20942 7420 21286
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 7484 20874 7512 21082
rect 7668 20874 7696 22170
rect 8128 22166 8156 22578
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 8116 22160 8168 22166
rect 8116 22102 8168 22108
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7852 21350 7880 21830
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7472 20868 7524 20874
rect 7472 20810 7524 20816
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 7484 20602 7512 20810
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6840 18748 6868 19790
rect 7024 18970 7052 20198
rect 7208 19854 7236 20198
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6920 18760 6972 18766
rect 6840 18720 6920 18748
rect 6920 18702 6972 18708
rect 6564 18550 6776 18578
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6564 18290 6592 18550
rect 6932 18290 6960 18702
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6012 16998 6040 17206
rect 6104 17190 6316 17218
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5408 15116 5580 15144
rect 5632 15156 5684 15162
rect 5356 15098 5408 15104
rect 5632 15098 5684 15104
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5151 14172 5459 14181
rect 5151 14170 5157 14172
rect 5213 14170 5237 14172
rect 5293 14170 5317 14172
rect 5373 14170 5397 14172
rect 5453 14170 5459 14172
rect 5213 14118 5215 14170
rect 5395 14118 5397 14170
rect 5151 14116 5157 14118
rect 5213 14116 5237 14118
rect 5293 14116 5317 14118
rect 5373 14116 5397 14118
rect 5453 14116 5459 14118
rect 5151 14107 5459 14116
rect 5151 13084 5459 13093
rect 5151 13082 5157 13084
rect 5213 13082 5237 13084
rect 5293 13082 5317 13084
rect 5373 13082 5397 13084
rect 5453 13082 5459 13084
rect 5213 13030 5215 13082
rect 5395 13030 5397 13082
rect 5151 13028 5157 13030
rect 5213 13028 5237 13030
rect 5293 13028 5317 13030
rect 5373 13028 5397 13030
rect 5453 13028 5459 13030
rect 5151 13019 5459 13028
rect 5552 12986 5580 14894
rect 5644 13938 5672 15098
rect 5828 15026 5856 15302
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5920 13870 5948 16050
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5172 12980 5224 12986
rect 4908 12940 5028 12968
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 12374 4292 12582
rect 4491 12540 4799 12549
rect 4491 12538 4497 12540
rect 4553 12538 4577 12540
rect 4633 12538 4657 12540
rect 4713 12538 4737 12540
rect 4793 12538 4799 12540
rect 4553 12486 4555 12538
rect 4735 12486 4737 12538
rect 4491 12484 4497 12486
rect 4553 12484 4577 12486
rect 4633 12484 4657 12486
rect 4713 12484 4737 12486
rect 4793 12484 4799 12486
rect 4491 12475 4799 12484
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4448 11898 4476 12174
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4908 11762 4936 12786
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11393 4292 11494
rect 4250 11384 4306 11393
rect 4356 11354 4384 11630
rect 4491 11452 4799 11461
rect 4491 11450 4497 11452
rect 4553 11450 4577 11452
rect 4633 11450 4657 11452
rect 4713 11450 4737 11452
rect 4793 11450 4799 11452
rect 4553 11398 4555 11450
rect 4735 11398 4737 11450
rect 4491 11396 4497 11398
rect 4553 11396 4577 11398
rect 4633 11396 4657 11398
rect 4713 11396 4737 11398
rect 4793 11396 4799 11398
rect 4491 11387 4799 11396
rect 4250 11319 4306 11328
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4894 11248 4950 11257
rect 4894 11183 4950 11192
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4066 10775 4068 10784
rect 4120 10775 4122 10784
rect 4160 10804 4212 10810
rect 4068 10746 4120 10752
rect 4160 10746 4212 10752
rect 4068 10668 4120 10674
rect 4120 10628 4384 10656
rect 4068 10610 4120 10616
rect 4250 10568 4306 10577
rect 4250 10503 4306 10512
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4080 10266 4108 10406
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9654 4108 9998
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4172 9518 4200 10406
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3988 9302 4200 9330
rect 4172 8498 4200 9302
rect 4264 8922 4292 10503
rect 4356 9674 4384 10628
rect 4632 10577 4660 11086
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4724 10810 4752 10950
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4908 10742 4936 11183
rect 5000 10849 5028 12940
rect 5172 12922 5224 12928
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5184 12306 5212 12922
rect 6012 12714 6040 16934
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5920 12186 5948 12378
rect 6012 12322 6040 12650
rect 6104 12442 6132 15438
rect 6196 13734 6224 16934
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6012 12294 6132 12322
rect 6196 12306 6224 12582
rect 6288 12434 6316 17190
rect 6380 14074 6408 17478
rect 6564 16182 6592 18226
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 6656 16114 6684 18226
rect 7024 18222 7052 18906
rect 7300 18630 7328 19722
rect 7576 19310 7604 19926
rect 7944 19378 7972 21626
rect 8128 21554 8156 22102
rect 8588 22030 8616 22442
rect 8680 22234 8708 22578
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8864 22094 8892 22578
rect 9404 22432 9456 22438
rect 9508 22386 9536 22714
rect 9456 22380 9536 22386
rect 9404 22374 9536 22380
rect 9416 22358 9536 22374
rect 9508 22114 9536 22358
rect 9600 22250 9628 24822
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9692 22710 9720 24006
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9600 22222 9812 22250
rect 8864 22066 9168 22094
rect 9508 22086 9720 22114
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8390 21720 8446 21729
rect 8390 21655 8446 21664
rect 8404 21622 8432 21655
rect 8496 21622 8524 21830
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8588 21554 8616 21966
rect 9140 21962 9168 22066
rect 9128 21956 9180 21962
rect 9128 21898 9180 21904
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8128 19446 8156 21490
rect 8588 21078 8616 21490
rect 9140 21350 9168 21898
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9508 21350 9536 21830
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 8576 21072 8628 21078
rect 8576 21014 8628 21020
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 20058 8248 20198
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8496 19446 8524 20266
rect 8116 19440 8168 19446
rect 8116 19382 8168 19388
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7380 18692 7432 18698
rect 7380 18634 7432 18640
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 7300 17678 7328 18566
rect 7392 18358 7420 18634
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7392 17882 7420 18294
rect 7576 18222 7604 19246
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7668 18170 7696 19314
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7852 18834 7880 19110
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 8588 18766 8616 20742
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8864 19310 8892 19790
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8956 18970 8984 19790
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8576 18760 8628 18766
rect 8956 18748 8984 18906
rect 9036 18760 9088 18766
rect 8956 18720 9036 18748
rect 8576 18702 8628 18708
rect 9036 18702 9088 18708
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7852 18170 7880 18226
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7378 17776 7434 17785
rect 7434 17734 7512 17762
rect 7378 17711 7434 17720
rect 7288 17672 7340 17678
rect 7102 17640 7158 17649
rect 7288 17614 7340 17620
rect 7102 17575 7104 17584
rect 7156 17575 7158 17584
rect 7104 17546 7156 17552
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7208 16114 7236 16662
rect 7392 16250 7420 17138
rect 7484 16590 7512 17734
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7392 16114 7420 16186
rect 7484 16114 7512 16526
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 6656 15858 6684 16050
rect 6656 15830 6776 15858
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6564 14958 6592 15438
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 12850 6408 13670
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6288 12406 6500 12434
rect 5092 11830 5120 12174
rect 5920 12158 6040 12186
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5151 11996 5459 12005
rect 5151 11994 5157 11996
rect 5213 11994 5237 11996
rect 5293 11994 5317 11996
rect 5373 11994 5397 11996
rect 5453 11994 5459 11996
rect 5213 11942 5215 11994
rect 5395 11942 5397 11994
rect 5151 11940 5157 11942
rect 5213 11940 5237 11942
rect 5293 11940 5317 11942
rect 5373 11940 5397 11942
rect 5453 11940 5459 11942
rect 5151 11931 5459 11940
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11218 5488 11630
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5151 10908 5459 10917
rect 5151 10906 5157 10908
rect 5213 10906 5237 10908
rect 5293 10906 5317 10908
rect 5373 10906 5397 10908
rect 5453 10906 5459 10908
rect 5213 10854 5215 10906
rect 5395 10854 5397 10906
rect 5151 10852 5157 10854
rect 5213 10852 5237 10854
rect 5293 10852 5317 10854
rect 5373 10852 5397 10854
rect 5453 10852 5459 10854
rect 4986 10840 5042 10849
rect 5151 10843 5459 10852
rect 4986 10775 5042 10784
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4804 10600 4856 10606
rect 4618 10568 4674 10577
rect 5000 10588 5028 10775
rect 5552 10742 5580 12038
rect 5644 11898 5672 12038
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5264 10736 5316 10742
rect 5262 10704 5264 10713
rect 5540 10736 5592 10742
rect 5316 10704 5318 10713
rect 5540 10678 5592 10684
rect 5262 10639 5318 10648
rect 4856 10560 5028 10588
rect 4804 10542 4856 10548
rect 4618 10503 4674 10512
rect 4491 10364 4799 10373
rect 4491 10362 4497 10364
rect 4553 10362 4577 10364
rect 4633 10362 4657 10364
rect 4713 10362 4737 10364
rect 4793 10362 4799 10364
rect 4553 10310 4555 10362
rect 4735 10310 4737 10362
rect 4491 10308 4497 10310
rect 4553 10308 4577 10310
rect 4633 10308 4657 10310
rect 4713 10308 4737 10310
rect 4793 10308 4799 10310
rect 4491 10299 4799 10308
rect 5000 9674 5028 10560
rect 5644 10538 5672 11834
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5736 10810 5764 11766
rect 6012 11626 6040 12158
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5920 10810 5948 10950
rect 6012 10810 6040 11562
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5264 10532 5316 10538
rect 4356 9646 4476 9674
rect 4448 9432 4476 9646
rect 4908 9646 5028 9674
rect 5092 10492 5264 10520
rect 4908 9586 4936 9646
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4448 9404 5028 9432
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 9042 4384 9318
rect 4491 9276 4799 9285
rect 4491 9274 4497 9276
rect 4553 9274 4577 9276
rect 4633 9274 4657 9276
rect 4713 9274 4737 9276
rect 4793 9274 4799 9276
rect 4553 9222 4555 9274
rect 4735 9222 4737 9274
rect 4491 9220 4497 9222
rect 4553 9220 4577 9222
rect 4633 9220 4657 9222
rect 4713 9220 4737 9222
rect 4793 9220 4799 9222
rect 4491 9211 4799 9220
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4264 8894 4476 8922
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 4080 7585 4108 7958
rect 4172 7818 4200 8434
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4264 7750 4292 8434
rect 4356 8362 4384 8774
rect 4448 8498 4476 8894
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8634 4936 8774
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5000 8514 5028 9404
rect 5092 9382 5120 10492
rect 5264 10474 5316 10480
rect 5632 10532 5684 10538
rect 5632 10474 5684 10480
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5151 9820 5459 9829
rect 5151 9818 5157 9820
rect 5213 9818 5237 9820
rect 5293 9818 5317 9820
rect 5373 9818 5397 9820
rect 5453 9818 5459 9820
rect 5213 9766 5215 9818
rect 5395 9766 5397 9818
rect 5151 9764 5157 9766
rect 5213 9764 5237 9766
rect 5293 9764 5317 9766
rect 5373 9764 5397 9766
rect 5453 9764 5459 9766
rect 5151 9755 5459 9764
rect 5552 9704 5580 10406
rect 6012 9722 6040 10746
rect 5460 9676 5580 9704
rect 6000 9716 6052 9722
rect 5460 9625 5488 9676
rect 6000 9658 6052 9664
rect 5446 9616 5502 9625
rect 5446 9551 5448 9560
rect 5500 9551 5502 9560
rect 5448 9522 5500 9528
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5092 9110 5120 9318
rect 5644 9178 5672 9318
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4908 8486 5028 8514
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4491 8188 4799 8197
rect 4491 8186 4497 8188
rect 4553 8186 4577 8188
rect 4633 8186 4657 8188
rect 4713 8186 4737 8188
rect 4793 8186 4799 8188
rect 4553 8134 4555 8186
rect 4735 8134 4737 8186
rect 4491 8132 4497 8134
rect 4553 8132 4577 8134
rect 4633 8132 4657 8134
rect 4713 8132 4737 8134
rect 4793 8132 4799 8134
rect 4491 8123 4799 8132
rect 4908 7818 4936 8486
rect 5092 8430 5120 8774
rect 5151 8732 5459 8741
rect 5151 8730 5157 8732
rect 5213 8730 5237 8732
rect 5293 8730 5317 8732
rect 5373 8730 5397 8732
rect 5453 8730 5459 8732
rect 5213 8678 5215 8730
rect 5395 8678 5397 8730
rect 5151 8676 5157 8678
rect 5213 8676 5237 8678
rect 5293 8676 5317 8678
rect 5373 8676 5397 8678
rect 5453 8676 5459 8678
rect 5151 8667 5459 8676
rect 5552 8634 5580 9046
rect 6012 9042 6040 9658
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6012 8634 6040 8978
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5816 8560 5868 8566
rect 5446 8528 5502 8537
rect 5816 8502 5868 8508
rect 5446 8463 5448 8472
rect 5500 8463 5502 8472
rect 5448 8434 5500 8440
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5000 7886 5028 8366
rect 5080 8288 5132 8294
rect 5540 8288 5592 8294
rect 5080 8230 5132 8236
rect 5460 8236 5540 8242
rect 5460 8230 5592 8236
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 4491 7100 4799 7109
rect 4491 7098 4497 7100
rect 4553 7098 4577 7100
rect 4633 7098 4657 7100
rect 4713 7098 4737 7100
rect 4793 7098 4799 7100
rect 4553 7046 4555 7098
rect 4735 7046 4737 7098
rect 4491 7044 4497 7046
rect 4553 7044 4577 7046
rect 4633 7044 4657 7046
rect 4713 7044 4737 7046
rect 4793 7044 4799 7046
rect 4491 7035 4799 7044
rect 4908 7002 4936 7754
rect 5092 7546 5120 8230
rect 5460 8214 5580 8230
rect 5460 7954 5488 8214
rect 5736 7954 5764 8366
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5151 7644 5459 7653
rect 5151 7642 5157 7644
rect 5213 7642 5237 7644
rect 5293 7642 5317 7644
rect 5373 7642 5397 7644
rect 5453 7642 5459 7644
rect 5213 7590 5215 7642
rect 5395 7590 5397 7642
rect 5151 7588 5157 7590
rect 5213 7588 5237 7590
rect 5293 7588 5317 7590
rect 5373 7588 5397 7590
rect 5453 7588 5459 7590
rect 5151 7579 5459 7588
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5736 7426 5764 7890
rect 5828 7886 5856 8502
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5828 7546 5856 7822
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5736 7398 5856 7426
rect 5828 7342 5856 7398
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 5092 6458 5120 6870
rect 5151 6556 5459 6565
rect 5151 6554 5157 6556
rect 5213 6554 5237 6556
rect 5293 6554 5317 6556
rect 5373 6554 5397 6556
rect 5453 6554 5459 6556
rect 5213 6502 5215 6554
rect 5395 6502 5397 6554
rect 5151 6500 5157 6502
rect 5213 6500 5237 6502
rect 5293 6500 5317 6502
rect 5373 6500 5397 6502
rect 5453 6500 5459 6502
rect 5151 6491 5459 6500
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5736 6254 5764 7278
rect 5920 6866 5948 7822
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5920 6458 5948 6802
rect 6104 6798 6132 12294
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 11218 6408 11698
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6182 11112 6238 11121
rect 6182 11047 6184 11056
rect 6236 11047 6238 11056
rect 6184 11018 6236 11024
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6196 8378 6224 9454
rect 6288 8906 6316 9590
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6288 8498 6316 8842
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6196 8350 6316 8378
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6196 7818 6224 8230
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6288 7750 6316 8350
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7206 6316 7686
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6866 6316 7142
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 4491 6012 4799 6021
rect 4491 6010 4497 6012
rect 4553 6010 4577 6012
rect 4633 6010 4657 6012
rect 4713 6010 4737 6012
rect 4793 6010 4799 6012
rect 4553 5958 4555 6010
rect 4735 5958 4737 6010
rect 4491 5956 4497 5958
rect 4553 5956 4577 5958
rect 4633 5956 4657 5958
rect 4713 5956 4737 5958
rect 4793 5956 4799 5958
rect 4491 5947 4799 5956
rect 5736 5846 5764 6190
rect 6104 6186 6132 6734
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6288 6458 6316 6666
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 5151 5468 5459 5477
rect 5151 5466 5157 5468
rect 5213 5466 5237 5468
rect 5293 5466 5317 5468
rect 5373 5466 5397 5468
rect 5453 5466 5459 5468
rect 5213 5414 5215 5466
rect 5395 5414 5397 5466
rect 5151 5412 5157 5414
rect 5213 5412 5237 5414
rect 5293 5412 5317 5414
rect 5373 5412 5397 5414
rect 5453 5412 5459 5414
rect 5151 5403 5459 5412
rect 6288 5234 6316 5714
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 4491 4924 4799 4933
rect 4491 4922 4497 4924
rect 4553 4922 4577 4924
rect 4633 4922 4657 4924
rect 4713 4922 4737 4924
rect 4793 4922 4799 4924
rect 4553 4870 4555 4922
rect 4735 4870 4737 4922
rect 4491 4868 4497 4870
rect 4553 4868 4577 4870
rect 4633 4868 4657 4870
rect 4713 4868 4737 4870
rect 4793 4868 4799 4870
rect 4491 4859 4799 4868
rect 6472 4486 6500 12406
rect 6564 11830 6592 13738
rect 6656 13530 6684 13806
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6748 12918 6776 15830
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14618 6868 14894
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6932 12442 6960 13262
rect 7024 12646 7052 16050
rect 7208 15366 7236 16050
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7392 14414 7420 16050
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7576 14346 7604 18158
rect 7668 18142 7880 18170
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7668 17678 7696 18022
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15570 7696 15846
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7852 14414 7880 18142
rect 7944 17678 7972 18158
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7944 15706 7972 16050
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 8128 15570 8156 16050
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 15094 8156 15506
rect 8220 15094 8248 18566
rect 9140 18154 9168 21286
rect 9692 20602 9720 22086
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9692 20058 9720 20402
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9232 18834 9260 19246
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9416 18766 9444 19858
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 19514 9628 19654
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9784 19446 9812 22222
rect 9876 22001 9904 30194
rect 13832 30122 13860 30246
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 13820 30116 13872 30122
rect 13820 30058 13872 30064
rect 11574 29948 11882 29957
rect 11574 29946 11580 29948
rect 11636 29946 11660 29948
rect 11716 29946 11740 29948
rect 11796 29946 11820 29948
rect 11876 29946 11882 29948
rect 11636 29894 11638 29946
rect 11818 29894 11820 29946
rect 11574 29892 11580 29894
rect 11636 29892 11660 29894
rect 11716 29892 11740 29894
rect 11796 29892 11820 29894
rect 11876 29892 11882 29894
rect 11574 29883 11882 29892
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 11244 29504 11296 29510
rect 11244 29446 11296 29452
rect 11256 29306 11284 29446
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11244 29096 11296 29102
rect 11244 29038 11296 29044
rect 11152 28960 11204 28966
rect 11152 28902 11204 28908
rect 11164 28626 11192 28902
rect 11256 28626 11284 29038
rect 11152 28620 11204 28626
rect 11152 28562 11204 28568
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 9956 28484 10008 28490
rect 9956 28426 10008 28432
rect 9968 28218 9996 28426
rect 10324 28416 10376 28422
rect 10324 28358 10376 28364
rect 10784 28416 10836 28422
rect 10784 28358 10836 28364
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 9968 27470 9996 28154
rect 10336 28014 10364 28358
rect 10324 28008 10376 28014
rect 10324 27950 10376 27956
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 10796 26450 10824 28358
rect 11058 28112 11114 28121
rect 11114 28070 11192 28098
rect 11058 28047 11114 28056
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 11072 27674 11100 27814
rect 11060 27668 11112 27674
rect 11060 27610 11112 27616
rect 11164 27606 11192 28070
rect 11256 27878 11284 28562
rect 11348 28150 11376 29582
rect 12234 29404 12542 29413
rect 12234 29402 12240 29404
rect 12296 29402 12320 29404
rect 12376 29402 12400 29404
rect 12456 29402 12480 29404
rect 12536 29402 12542 29404
rect 12296 29350 12298 29402
rect 12478 29350 12480 29402
rect 12234 29348 12240 29350
rect 12296 29348 12320 29350
rect 12376 29348 12400 29350
rect 12456 29348 12480 29350
rect 12536 29348 12542 29350
rect 12234 29339 12542 29348
rect 13280 29306 13308 29582
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 13268 29300 13320 29306
rect 13268 29242 13320 29248
rect 12256 29232 12308 29238
rect 12256 29174 12308 29180
rect 11574 28860 11882 28869
rect 11574 28858 11580 28860
rect 11636 28858 11660 28860
rect 11716 28858 11740 28860
rect 11796 28858 11820 28860
rect 11876 28858 11882 28860
rect 11636 28806 11638 28858
rect 11818 28806 11820 28858
rect 11574 28804 11580 28806
rect 11636 28804 11660 28806
rect 11716 28804 11740 28806
rect 11796 28804 11820 28806
rect 11876 28804 11882 28806
rect 11574 28795 11882 28804
rect 12268 28642 12296 29174
rect 12636 28762 12664 29242
rect 13452 29096 13504 29102
rect 13452 29038 13504 29044
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 12176 28614 12296 28642
rect 12176 28558 12204 28614
rect 12164 28552 12216 28558
rect 12164 28494 12216 28500
rect 12072 28484 12124 28490
rect 12072 28426 12124 28432
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11716 28150 11744 28358
rect 11336 28144 11388 28150
rect 11336 28086 11388 28092
rect 11704 28144 11756 28150
rect 12084 28121 12112 28426
rect 11704 28086 11756 28092
rect 12070 28112 12126 28121
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11348 27674 11376 28086
rect 11428 28076 11480 28082
rect 12070 28047 12126 28056
rect 11428 28018 11480 28024
rect 11440 27946 11468 28018
rect 12070 27976 12126 27985
rect 11428 27940 11480 27946
rect 11428 27882 11480 27888
rect 11992 27934 12070 27962
rect 11336 27668 11388 27674
rect 11336 27610 11388 27616
rect 11152 27600 11204 27606
rect 11152 27542 11204 27548
rect 11440 27470 11468 27882
rect 11574 27772 11882 27781
rect 11574 27770 11580 27772
rect 11636 27770 11660 27772
rect 11716 27770 11740 27772
rect 11796 27770 11820 27772
rect 11876 27770 11882 27772
rect 11636 27718 11638 27770
rect 11818 27718 11820 27770
rect 11574 27716 11580 27718
rect 11636 27716 11660 27718
rect 11716 27716 11740 27718
rect 11796 27716 11820 27718
rect 11876 27716 11882 27718
rect 11574 27707 11882 27716
rect 11888 27668 11940 27674
rect 11888 27610 11940 27616
rect 11900 27470 11928 27610
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 11992 27334 12020 27934
rect 12070 27911 12126 27920
rect 12072 27872 12124 27878
rect 12072 27814 12124 27820
rect 12084 27674 12112 27814
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 12176 27554 12204 28494
rect 12234 28316 12542 28325
rect 12234 28314 12240 28316
rect 12296 28314 12320 28316
rect 12376 28314 12400 28316
rect 12456 28314 12480 28316
rect 12536 28314 12542 28316
rect 12296 28262 12298 28314
rect 12478 28262 12480 28314
rect 12234 28260 12240 28262
rect 12296 28260 12320 28262
rect 12376 28260 12400 28262
rect 12456 28260 12480 28262
rect 12536 28260 12542 28262
rect 12234 28251 12542 28260
rect 12912 28218 12940 28698
rect 12900 28212 12952 28218
rect 12900 28154 12952 28160
rect 13084 28144 13136 28150
rect 13084 28086 13136 28092
rect 12256 28076 12308 28082
rect 12256 28018 12308 28024
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12084 27526 12204 27554
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11256 26586 11284 26726
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 11348 26314 11376 26998
rect 11900 26994 11928 27270
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 11992 26858 12020 27270
rect 12084 27062 12112 27526
rect 12268 27470 12296 28018
rect 12728 27538 12756 28018
rect 13096 27538 13124 28086
rect 13464 28082 13492 29038
rect 13740 28762 13768 29038
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13634 28656 13690 28665
rect 13634 28591 13636 28600
rect 13688 28591 13690 28600
rect 13636 28562 13688 28568
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 12268 27334 12296 27406
rect 12256 27328 12308 27334
rect 12176 27288 12256 27316
rect 12072 27056 12124 27062
rect 12072 26998 12124 27004
rect 11980 26852 12032 26858
rect 11980 26794 12032 26800
rect 11574 26684 11882 26693
rect 11574 26682 11580 26684
rect 11636 26682 11660 26684
rect 11716 26682 11740 26684
rect 11796 26682 11820 26684
rect 11876 26682 11882 26684
rect 11636 26630 11638 26682
rect 11818 26630 11820 26682
rect 11574 26628 11580 26630
rect 11636 26628 11660 26630
rect 11716 26628 11740 26630
rect 11796 26628 11820 26630
rect 11876 26628 11882 26630
rect 11574 26619 11882 26628
rect 12176 26586 12204 27288
rect 12256 27270 12308 27276
rect 12234 27228 12542 27237
rect 12234 27226 12240 27228
rect 12296 27226 12320 27228
rect 12376 27226 12400 27228
rect 12456 27226 12480 27228
rect 12536 27226 12542 27228
rect 12296 27174 12298 27226
rect 12478 27174 12480 27226
rect 12234 27172 12240 27174
rect 12296 27172 12320 27174
rect 12376 27172 12400 27174
rect 12456 27172 12480 27174
rect 12536 27172 12542 27174
rect 12234 27163 12542 27172
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 12164 26580 12216 26586
rect 12164 26522 12216 26528
rect 12268 26450 12296 26930
rect 12728 26874 12756 27474
rect 12992 27396 13044 27402
rect 12992 27338 13044 27344
rect 12900 27056 12952 27062
rect 12900 26998 12952 27004
rect 12808 26920 12860 26926
rect 12728 26868 12808 26874
rect 12728 26862 12860 26868
rect 12728 26846 12848 26862
rect 12912 26790 12940 26998
rect 12808 26784 12860 26790
rect 12808 26726 12860 26732
rect 12900 26784 12952 26790
rect 12900 26726 12952 26732
rect 12820 26602 12848 26726
rect 13004 26602 13032 27338
rect 12820 26574 13032 26602
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 11336 26308 11388 26314
rect 11336 26250 11388 26256
rect 11440 24818 11468 26386
rect 12234 26140 12542 26149
rect 12234 26138 12240 26140
rect 12296 26138 12320 26140
rect 12376 26138 12400 26140
rect 12456 26138 12480 26140
rect 12536 26138 12542 26140
rect 12296 26086 12298 26138
rect 12478 26086 12480 26138
rect 12234 26084 12240 26086
rect 12296 26084 12320 26086
rect 12376 26084 12400 26086
rect 12456 26084 12480 26086
rect 12536 26084 12542 26086
rect 12234 26075 12542 26084
rect 11574 25596 11882 25605
rect 11574 25594 11580 25596
rect 11636 25594 11660 25596
rect 11716 25594 11740 25596
rect 11796 25594 11820 25596
rect 11876 25594 11882 25596
rect 11636 25542 11638 25594
rect 11818 25542 11820 25594
rect 11574 25540 11580 25542
rect 11636 25540 11660 25542
rect 11716 25540 11740 25542
rect 11796 25540 11820 25542
rect 11876 25540 11882 25542
rect 11574 25531 11882 25540
rect 13464 25362 13492 28018
rect 13556 27985 13584 28494
rect 13636 28484 13688 28490
rect 13636 28426 13688 28432
rect 13648 28257 13676 28426
rect 13912 28416 13964 28422
rect 13832 28376 13912 28404
rect 13634 28248 13690 28257
rect 13634 28183 13690 28192
rect 13542 27976 13598 27985
rect 13542 27911 13598 27920
rect 13636 27124 13688 27130
rect 13636 27066 13688 27072
rect 13648 27010 13676 27066
rect 13832 27010 13860 28376
rect 13912 28358 13964 28364
rect 14016 27674 14044 28494
rect 14004 27668 14056 27674
rect 14004 27610 14056 27616
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 14016 27334 14044 27474
rect 14004 27328 14056 27334
rect 14004 27270 14056 27276
rect 13648 26982 13860 27010
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 13924 26858 13952 26930
rect 14016 26858 14044 27270
rect 13912 26852 13964 26858
rect 13912 26794 13964 26800
rect 14004 26852 14056 26858
rect 14004 26794 14056 26800
rect 13452 25356 13504 25362
rect 13452 25298 13504 25304
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 11888 25152 11940 25158
rect 11888 25094 11940 25100
rect 11900 24886 11928 25094
rect 12234 25052 12542 25061
rect 12234 25050 12240 25052
rect 12296 25050 12320 25052
rect 12376 25050 12400 25052
rect 12456 25050 12480 25052
rect 12536 25050 12542 25052
rect 12296 24998 12298 25050
rect 12478 24998 12480 25050
rect 12234 24996 12240 24998
rect 12296 24996 12320 24998
rect 12376 24996 12400 24998
rect 12456 24996 12480 24998
rect 12536 24996 12542 24998
rect 12234 24987 12542 24996
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 10600 24744 10652 24750
rect 10600 24686 10652 24692
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10140 22568 10192 22574
rect 10140 22510 10192 22516
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9862 21992 9918 22001
rect 9862 21927 9918 21936
rect 9968 21876 9996 22102
rect 10152 22098 10180 22510
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10060 21978 10088 22034
rect 10244 21978 10272 22374
rect 10060 21950 10272 21978
rect 9876 21848 9996 21876
rect 10232 21888 10284 21894
rect 9876 20602 9904 21848
rect 10232 21830 10284 21836
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9968 20874 9996 21626
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9876 20369 9904 20402
rect 9862 20360 9918 20369
rect 9862 20295 9918 20304
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9876 19378 9904 20295
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9600 18970 9628 19178
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9968 18834 9996 20810
rect 10060 20602 10088 21422
rect 10244 21078 10272 21830
rect 10232 21072 10284 21078
rect 10232 21014 10284 21020
rect 10244 20942 10272 21014
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 10152 20466 10180 20742
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14482 8156 14758
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7564 14340 7616 14346
rect 7484 14300 7564 14328
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7116 13326 7144 13738
rect 7208 13530 7236 13738
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7300 13326 7328 13806
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12986 7144 13126
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7208 12850 7236 13262
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7208 12442 7236 12786
rect 7300 12714 7328 13262
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7208 12238 7236 12378
rect 7300 12238 7328 12650
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 7024 10606 7052 12038
rect 7208 11898 7236 12174
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6564 8974 6592 9386
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6656 8430 6684 9318
rect 7116 8906 7144 10950
rect 7208 10674 7236 11494
rect 7300 11286 7328 11698
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 7392 11150 7420 11494
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7484 11082 7512 14300
rect 7564 14282 7616 14288
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7576 12442 7604 12786
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7668 11898 7696 12174
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7562 11248 7618 11257
rect 7562 11183 7618 11192
rect 7576 11082 7604 11183
rect 7852 11150 7880 14350
rect 8220 13326 8248 15030
rect 8312 15026 8340 15914
rect 8680 15706 8708 15982
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8680 15162 8708 15642
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 9232 14958 9260 15438
rect 9416 15162 9444 18702
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9876 18290 9904 18362
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9784 16658 9812 18226
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17134 9904 18022
rect 9968 17746 9996 18770
rect 10152 18290 10180 20198
rect 10244 19854 10272 20878
rect 10322 20360 10378 20369
rect 10322 20295 10378 20304
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10336 19786 10364 20295
rect 10324 19780 10376 19786
rect 10324 19722 10376 19728
rect 10428 19334 10456 24550
rect 10612 23730 10640 24686
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10612 23254 10640 23666
rect 10796 23254 10824 24142
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10600 23248 10652 23254
rect 10600 23190 10652 23196
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 10796 23066 10824 23190
rect 10520 23038 10824 23066
rect 10876 23044 10928 23050
rect 10520 22030 10548 23038
rect 10876 22986 10928 22992
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10690 22128 10746 22137
rect 10600 22092 10652 22098
rect 10796 22094 10824 22510
rect 10746 22072 10824 22094
rect 10690 22066 10824 22072
rect 10690 22063 10746 22066
rect 10600 22034 10652 22040
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10520 21146 10548 21830
rect 10612 21622 10640 22034
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10612 20466 10640 21286
rect 10704 20466 10732 22063
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10796 21690 10824 21966
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10796 21010 10824 21286
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10796 20806 10824 20946
rect 10888 20942 10916 22986
rect 10980 22794 11008 23462
rect 11440 23322 11468 24754
rect 11574 24508 11882 24517
rect 11574 24506 11580 24508
rect 11636 24506 11660 24508
rect 11716 24506 11740 24508
rect 11796 24506 11820 24508
rect 11876 24506 11882 24508
rect 11636 24454 11638 24506
rect 11818 24454 11820 24506
rect 11574 24452 11580 24454
rect 11636 24452 11660 24454
rect 11716 24452 11740 24454
rect 11796 24452 11820 24454
rect 11876 24452 11882 24454
rect 11574 24443 11882 24452
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11888 24132 11940 24138
rect 11888 24074 11940 24080
rect 11808 23866 11836 24074
rect 11900 23866 11928 24074
rect 12234 23964 12542 23973
rect 12234 23962 12240 23964
rect 12296 23962 12320 23964
rect 12376 23962 12400 23964
rect 12456 23962 12480 23964
rect 12536 23962 12542 23964
rect 12296 23910 12298 23962
rect 12478 23910 12480 23962
rect 12234 23908 12240 23910
rect 12296 23908 12320 23910
rect 12376 23908 12400 23910
rect 12456 23908 12480 23910
rect 12536 23908 12542 23910
rect 12234 23899 12542 23908
rect 13004 23866 13032 25230
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13176 24336 13228 24342
rect 13176 24278 13228 24284
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 11574 23420 11882 23429
rect 11574 23418 11580 23420
rect 11636 23418 11660 23420
rect 11716 23418 11740 23420
rect 11796 23418 11820 23420
rect 11876 23418 11882 23420
rect 11636 23366 11638 23418
rect 11818 23366 11820 23418
rect 11574 23364 11580 23366
rect 11636 23364 11660 23366
rect 11716 23364 11740 23366
rect 11796 23364 11820 23366
rect 11876 23364 11882 23366
rect 11574 23355 11882 23364
rect 11428 23316 11480 23322
rect 11428 23258 11480 23264
rect 11440 23186 11468 23258
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 10980 22766 11100 22794
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 10980 21622 11008 22646
rect 11072 21690 11100 22766
rect 12176 22642 12204 23462
rect 12234 22876 12542 22885
rect 12234 22874 12240 22876
rect 12296 22874 12320 22876
rect 12376 22874 12400 22876
rect 12456 22874 12480 22876
rect 12536 22874 12542 22876
rect 12296 22822 12298 22874
rect 12478 22822 12480 22874
rect 12234 22820 12240 22822
rect 12296 22820 12320 22822
rect 12376 22820 12400 22822
rect 12456 22820 12480 22822
rect 12536 22820 12542 22822
rect 12234 22811 12542 22820
rect 12820 22778 12848 23666
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 13188 22642 13216 24278
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 11244 22500 11296 22506
rect 11244 22442 11296 22448
rect 11256 22234 11284 22442
rect 11348 22234 11376 22578
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11244 22228 11296 22234
rect 11244 22170 11296 22176
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 11440 21128 11468 22510
rect 11574 22332 11882 22341
rect 11574 22330 11580 22332
rect 11636 22330 11660 22332
rect 11716 22330 11740 22332
rect 11796 22330 11820 22332
rect 11876 22330 11882 22332
rect 11636 22278 11638 22330
rect 11818 22278 11820 22330
rect 11574 22276 11580 22278
rect 11636 22276 11660 22278
rect 11716 22276 11740 22278
rect 11796 22276 11820 22278
rect 11876 22276 11882 22278
rect 11574 22267 11882 22276
rect 12636 22234 12664 22578
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 11574 21244 11882 21253
rect 11574 21242 11580 21244
rect 11636 21242 11660 21244
rect 11716 21242 11740 21244
rect 11796 21242 11820 21244
rect 11876 21242 11882 21244
rect 11636 21190 11638 21242
rect 11818 21190 11820 21242
rect 11574 21188 11580 21190
rect 11636 21188 11660 21190
rect 11716 21188 11740 21190
rect 11796 21188 11820 21190
rect 11876 21188 11882 21190
rect 11574 21179 11882 21188
rect 11440 21100 11560 21128
rect 11532 20942 11560 21100
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 11164 20466 11192 20810
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 10506 19952 10562 19961
rect 10506 19887 10508 19896
rect 10560 19887 10562 19896
rect 10508 19858 10560 19864
rect 10428 19306 10548 19334
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10428 18290 10456 18634
rect 10140 18284 10192 18290
rect 10060 18244 10140 18272
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9968 17338 9996 17682
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 16250 9996 16526
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 10060 16182 10088 18244
rect 10416 18284 10468 18290
rect 10140 18226 10192 18232
rect 10244 18244 10416 18272
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10152 17610 10180 18022
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9508 15570 9536 16050
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15706 9996 15846
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 10060 15586 10088 16118
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9968 15558 10088 15586
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8588 14346 8616 14758
rect 9232 14414 9260 14894
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 9232 12782 9260 14350
rect 9416 13394 9444 15098
rect 9968 13938 9996 15558
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 10060 15094 10088 15370
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9416 13190 9444 13330
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 7944 12646 7972 12718
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 9232 12306 9260 12718
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9784 12170 9812 13398
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11778 9720 12038
rect 9876 11898 9904 13194
rect 10060 12918 10088 15030
rect 10152 13734 10180 16594
rect 10244 16114 10272 18244
rect 10416 18226 10468 18232
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10336 16454 10364 18090
rect 10520 16726 10548 19306
rect 10704 18698 10732 20402
rect 10980 19825 11008 20402
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 10966 19816 11022 19825
rect 10876 19780 10928 19786
rect 10966 19751 11022 19760
rect 10876 19722 10928 19728
rect 10888 19446 10916 19722
rect 11348 19718 11376 19858
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11072 19514 11100 19654
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 11164 18834 11192 19654
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 18086 11192 18566
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10508 16720 10560 16726
rect 10508 16662 10560 16668
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10244 13938 10272 16050
rect 10336 14074 10364 16390
rect 10428 15162 10456 16390
rect 10506 15600 10562 15609
rect 10506 15535 10508 15544
rect 10560 15535 10562 15544
rect 10508 15506 10560 15512
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10428 14414 10456 14554
rect 10612 14550 10640 17818
rect 10876 17672 10928 17678
rect 10796 17620 10876 17626
rect 10796 17614 10928 17620
rect 10796 17598 10916 17614
rect 10796 17490 10824 17598
rect 10704 17462 10824 17490
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10508 14544 10560 14550
rect 10506 14512 10508 14521
rect 10600 14544 10652 14550
rect 10560 14512 10562 14521
rect 10600 14486 10652 14492
rect 10506 14447 10562 14456
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10428 13818 10456 14350
rect 10704 14346 10732 17462
rect 10888 17202 10916 17478
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15706 10916 15982
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10888 15178 10916 15642
rect 10796 15150 10916 15178
rect 10980 15162 11008 16594
rect 10968 15156 11020 15162
rect 10796 14414 10824 15150
rect 10968 15098 11020 15104
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10888 14414 10916 14486
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 13841 10548 13874
rect 10336 13790 10456 13818
rect 10506 13832 10562 13841
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13410 10180 13670
rect 10230 13424 10286 13433
rect 10152 13382 10230 13410
rect 10230 13359 10286 13368
rect 10336 13326 10364 13790
rect 10506 13767 10562 13776
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10324 13320 10376 13326
rect 10152 13268 10324 13274
rect 10152 13262 10376 13268
rect 10152 13246 10364 13262
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 10060 12434 10088 12854
rect 9968 12406 10088 12434
rect 9968 12170 9996 12406
rect 10152 12186 10180 13246
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10244 12782 10272 13126
rect 10428 12986 10456 13670
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10520 12850 10548 13262
rect 10704 13258 10732 14282
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10796 13326 10824 13806
rect 10888 13326 10916 14350
rect 10980 14278 11008 15098
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 14074 11100 14214
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10244 12434 10272 12718
rect 10520 12442 10548 12786
rect 10704 12714 10732 13194
rect 10796 12986 10824 13262
rect 10980 13258 11008 14010
rect 11164 13734 11192 18022
rect 11256 17678 11284 18158
rect 11348 17814 11376 18158
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11440 17678 11468 20878
rect 11808 20466 11836 20946
rect 11992 20806 12020 21898
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 12084 21554 12112 21830
rect 12234 21788 12542 21797
rect 12234 21786 12240 21788
rect 12296 21786 12320 21788
rect 12376 21786 12400 21788
rect 12456 21786 12480 21788
rect 12536 21786 12542 21788
rect 12296 21734 12298 21786
rect 12478 21734 12480 21786
rect 12234 21732 12240 21734
rect 12296 21732 12320 21734
rect 12376 21732 12400 21734
rect 12456 21732 12480 21734
rect 12536 21732 12542 21734
rect 12234 21723 12542 21732
rect 12636 21554 12664 21898
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11574 20156 11882 20165
rect 11574 20154 11580 20156
rect 11636 20154 11660 20156
rect 11716 20154 11740 20156
rect 11796 20154 11820 20156
rect 11876 20154 11882 20156
rect 11636 20102 11638 20154
rect 11818 20102 11820 20154
rect 11574 20100 11580 20102
rect 11636 20100 11660 20102
rect 11716 20100 11740 20102
rect 11796 20100 11820 20102
rect 11876 20100 11882 20102
rect 11574 20091 11882 20100
rect 11574 19068 11882 19077
rect 11574 19066 11580 19068
rect 11636 19066 11660 19068
rect 11716 19066 11740 19068
rect 11796 19066 11820 19068
rect 11876 19066 11882 19068
rect 11636 19014 11638 19066
rect 11818 19014 11820 19066
rect 11574 19012 11580 19014
rect 11636 19012 11660 19014
rect 11716 19012 11740 19014
rect 11796 19012 11820 19014
rect 11876 19012 11882 19014
rect 11574 19003 11882 19012
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11624 18290 11652 18770
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11574 17980 11882 17989
rect 11574 17978 11580 17980
rect 11636 17978 11660 17980
rect 11716 17978 11740 17980
rect 11796 17978 11820 17980
rect 11876 17978 11882 17980
rect 11636 17926 11638 17978
rect 11818 17926 11820 17978
rect 11574 17924 11580 17926
rect 11636 17924 11660 17926
rect 11716 17924 11740 17926
rect 11796 17924 11820 17926
rect 11876 17924 11882 17926
rect 11574 17915 11882 17924
rect 11992 17882 12020 20742
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 12084 20058 12112 20334
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12176 19310 12204 21490
rect 12728 21486 12756 21830
rect 12912 21570 12940 22034
rect 13084 21616 13136 21622
rect 12912 21564 13084 21570
rect 12912 21558 13136 21564
rect 12912 21542 13124 21558
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12234 20700 12542 20709
rect 12234 20698 12240 20700
rect 12296 20698 12320 20700
rect 12376 20698 12400 20700
rect 12456 20698 12480 20700
rect 12536 20698 12542 20700
rect 12296 20646 12298 20698
rect 12478 20646 12480 20698
rect 12234 20644 12240 20646
rect 12296 20644 12320 20646
rect 12376 20644 12400 20646
rect 12456 20644 12480 20646
rect 12536 20644 12542 20646
rect 12234 20635 12542 20644
rect 12728 20505 12756 21286
rect 12912 20874 12940 21542
rect 13188 21468 13216 22578
rect 13556 22094 13584 24074
rect 13740 23662 13768 24686
rect 13924 24206 13952 26794
rect 14108 24886 14136 29650
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13740 22982 13768 23598
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13740 22506 13768 22918
rect 13728 22500 13780 22506
rect 13728 22442 13780 22448
rect 13740 22234 13768 22442
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 14200 22094 14228 30194
rect 17420 30122 17448 31925
rect 19317 30492 19625 30501
rect 19317 30490 19323 30492
rect 19379 30490 19403 30492
rect 19459 30490 19483 30492
rect 19539 30490 19563 30492
rect 19619 30490 19625 30492
rect 19379 30438 19381 30490
rect 19561 30438 19563 30490
rect 19317 30436 19323 30438
rect 19379 30436 19403 30438
rect 19459 30436 19483 30438
rect 19539 30436 19563 30438
rect 19619 30436 19625 30438
rect 19317 30427 19625 30436
rect 21284 30326 21312 31925
rect 25424 30326 25452 32014
rect 28998 31925 29054 32725
rect 28906 30696 28962 30705
rect 28906 30631 28962 30640
rect 26400 30492 26708 30501
rect 26400 30490 26406 30492
rect 26462 30490 26486 30492
rect 26542 30490 26566 30492
rect 26622 30490 26646 30492
rect 26702 30490 26708 30492
rect 26462 30438 26464 30490
rect 26644 30438 26646 30490
rect 26400 30436 26406 30438
rect 26462 30436 26486 30438
rect 26542 30436 26566 30438
rect 26622 30436 26646 30438
rect 26702 30436 26708 30438
rect 26400 30427 26708 30436
rect 21272 30320 21324 30326
rect 21272 30262 21324 30268
rect 25412 30320 25464 30326
rect 25412 30262 25464 30268
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 17408 30116 17460 30122
rect 17408 30058 17460 30064
rect 16212 29708 16264 29714
rect 16212 29650 16264 29656
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 14292 29238 14320 29514
rect 14280 29232 14332 29238
rect 14280 29174 14332 29180
rect 14292 28150 14320 29174
rect 16224 29170 16252 29650
rect 16488 29572 16540 29578
rect 16488 29514 16540 29520
rect 16500 29306 16528 29514
rect 17132 29504 17184 29510
rect 17132 29446 17184 29452
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 16488 29300 16540 29306
rect 16488 29242 16540 29248
rect 16672 29232 16724 29238
rect 16672 29174 16724 29180
rect 16212 29164 16264 29170
rect 16212 29106 16264 29112
rect 15476 28960 15528 28966
rect 15476 28902 15528 28908
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15488 28558 15516 28902
rect 15948 28626 15976 28902
rect 16224 28762 16252 29106
rect 16580 29096 16632 29102
rect 16580 29038 16632 29044
rect 16212 28756 16264 28762
rect 16212 28698 16264 28704
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 16592 28558 16620 29038
rect 16684 28762 16712 29174
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 17144 28626 17172 29446
rect 17328 29306 17356 29446
rect 17316 29300 17368 29306
rect 17316 29242 17368 29248
rect 17132 28620 17184 28626
rect 17132 28562 17184 28568
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 14280 28144 14332 28150
rect 14280 28086 14332 28092
rect 14292 26994 14320 28086
rect 14476 27878 14504 28494
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14476 27674 14504 27814
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14568 27130 14596 27270
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14752 27062 14780 28358
rect 15304 28218 15332 28358
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 15292 28008 15344 28014
rect 15292 27950 15344 27956
rect 14740 27056 14792 27062
rect 14740 26998 14792 27004
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 15304 26926 15332 27950
rect 15488 27538 15516 28494
rect 16304 28484 16356 28490
rect 16304 28426 16356 28432
rect 16316 28218 16344 28426
rect 16304 28212 16356 28218
rect 16304 28154 16356 28160
rect 16500 28082 16528 28494
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 15476 27532 15528 27538
rect 15476 27474 15528 27480
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16488 27464 16540 27470
rect 16592 27452 16620 28494
rect 17132 27872 17184 27878
rect 17132 27814 17184 27820
rect 17144 27538 17172 27814
rect 17132 27532 17184 27538
rect 17132 27474 17184 27480
rect 16540 27424 16620 27452
rect 16488 27406 16540 27412
rect 16408 27130 16436 27406
rect 16396 27124 16448 27130
rect 16396 27066 16448 27072
rect 15292 26920 15344 26926
rect 15292 26862 15344 26868
rect 15016 25356 15068 25362
rect 15016 25298 15068 25304
rect 14924 25220 14976 25226
rect 14924 25162 14976 25168
rect 14936 24954 14964 25162
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14280 24812 14332 24818
rect 14332 24772 14412 24800
rect 14280 24754 14332 24760
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14292 23662 14320 24006
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14292 22642 14320 23054
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 13556 22066 13768 22094
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 13096 21440 13216 21468
rect 13268 21480 13320 21486
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12808 20528 12860 20534
rect 12714 20496 12770 20505
rect 12912 20516 12940 20810
rect 12860 20488 12940 20516
rect 12808 20470 12860 20476
rect 12714 20431 12770 20440
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12544 19786 12572 20198
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12532 19780 12584 19786
rect 12532 19722 12584 19728
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12234 19612 12542 19621
rect 12234 19610 12240 19612
rect 12296 19610 12320 19612
rect 12376 19610 12400 19612
rect 12456 19610 12480 19612
rect 12536 19610 12542 19612
rect 12296 19558 12298 19610
rect 12478 19558 12480 19610
rect 12234 19556 12240 19558
rect 12296 19556 12320 19558
rect 12376 19556 12400 19558
rect 12456 19556 12480 19558
rect 12536 19556 12542 19558
rect 12234 19547 12542 19556
rect 12636 19334 12664 19654
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12544 19306 12664 19334
rect 12176 18970 12204 19246
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12544 18834 12572 19306
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12728 18766 12756 19790
rect 12820 18902 12848 20470
rect 13004 19854 13032 21286
rect 13096 20602 13124 21440
rect 13268 21422 13320 21428
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12912 19378 12940 19654
rect 13096 19514 13124 20538
rect 13176 19848 13228 19854
rect 13174 19816 13176 19825
rect 13228 19816 13230 19825
rect 13174 19751 13230 19760
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13188 19378 13216 19751
rect 13280 19514 13308 21422
rect 13464 21078 13492 21898
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12716 18760 12768 18766
rect 12636 18720 12716 18748
rect 12234 18524 12542 18533
rect 12234 18522 12240 18524
rect 12296 18522 12320 18524
rect 12376 18522 12400 18524
rect 12456 18522 12480 18524
rect 12536 18522 12542 18524
rect 12296 18470 12298 18522
rect 12478 18470 12480 18522
rect 12234 18468 12240 18470
rect 12296 18468 12320 18470
rect 12376 18468 12400 18470
rect 12456 18468 12480 18470
rect 12536 18468 12542 18470
rect 12234 18459 12542 18468
rect 12636 18426 12664 18720
rect 12716 18702 12768 18708
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12728 18426 12756 18566
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11256 17066 11284 17614
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11348 15434 11376 16186
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10508 12436 10560 12442
rect 10244 12406 10364 12434
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 10060 12158 10180 12186
rect 9864 11892 9916 11898
rect 9916 11852 9996 11880
rect 9864 11834 9916 11840
rect 9772 11824 9824 11830
rect 9692 11772 9772 11778
rect 9692 11766 9824 11772
rect 9692 11750 9812 11766
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7484 9674 7512 11018
rect 7484 9646 7696 9674
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6748 8430 6776 8570
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6656 7818 6684 8366
rect 6748 8022 6776 8366
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6840 7818 6868 8434
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7546 6592 7686
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6736 6792 6788 6798
rect 7024 6769 7052 6802
rect 6736 6734 6788 6740
rect 7010 6760 7066 6769
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6564 5914 6592 6598
rect 6748 6254 6776 6734
rect 7010 6695 7066 6704
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 6390 6868 6598
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 7116 6322 7144 8842
rect 7208 7954 7236 9318
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 6322 7236 7686
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 7116 5658 7144 6258
rect 7208 5914 7236 6258
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7300 5778 7328 6870
rect 7668 6798 7696 9646
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7484 6458 7512 6734
rect 7668 6662 7696 6734
rect 7760 6730 7788 7142
rect 8128 7002 8156 11086
rect 8956 11082 8984 11630
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8852 9512 8904 9518
rect 8850 9480 8852 9489
rect 8904 9480 8906 9489
rect 8850 9415 8906 9424
rect 8956 8974 8984 11018
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9586 9076 9862
rect 9600 9674 9628 10066
rect 9508 9646 9628 9674
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9140 9042 9168 9454
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8128 6798 8156 6938
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7024 5642 7144 5658
rect 7012 5636 7156 5642
rect 7064 5630 7104 5636
rect 7012 5578 7064 5584
rect 7104 5578 7156 5584
rect 7116 5302 7144 5578
rect 8036 5302 8064 6598
rect 8128 6186 8156 6734
rect 8220 6322 8248 8366
rect 8300 6792 8352 6798
rect 8298 6760 8300 6769
rect 8352 6760 8354 6769
rect 8298 6695 8354 6704
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8220 5370 8248 6258
rect 8956 5370 8984 8910
rect 9036 8560 9088 8566
rect 9034 8528 9036 8537
rect 9088 8528 9090 8537
rect 9034 8463 9090 8472
rect 9508 8430 9536 9646
rect 9692 9602 9720 11750
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9784 10810 9812 11630
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9968 10674 9996 11852
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10060 10470 10088 12158
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11218 10180 12038
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10336 10674 10364 12406
rect 10704 12434 10732 12650
rect 10704 12406 10824 12434
rect 10508 12378 10560 12384
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9600 9574 9720 9602
rect 9600 9330 9628 9574
rect 9680 9512 9732 9518
rect 9784 9500 9812 10202
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9876 9874 9904 9998
rect 9968 9994 9996 10406
rect 10060 10266 10088 10406
rect 10152 10266 10180 10610
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10060 10146 10088 10202
rect 10060 10118 10180 10146
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9954 9888 10010 9897
rect 9876 9846 9954 9874
rect 9954 9823 10010 9832
rect 9968 9722 9996 9823
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9732 9472 9812 9500
rect 9680 9454 9732 9460
rect 9600 9302 9720 9330
rect 9692 8906 9720 9302
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9784 8498 9812 9472
rect 9876 9042 9904 9522
rect 9968 9081 9996 9522
rect 10060 9382 10088 9998
rect 10152 9450 10180 10118
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10244 9654 10272 10066
rect 10336 10062 10364 10610
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10428 10470 10456 10542
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10336 9926 10364 9998
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10336 9518 10364 9862
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10428 9110 10456 9998
rect 10520 9722 10548 10406
rect 10612 9722 10640 10474
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10704 9722 10732 10066
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10796 9602 10824 12406
rect 11256 11354 11284 15302
rect 11440 14906 11468 17614
rect 11574 16892 11882 16901
rect 11574 16890 11580 16892
rect 11636 16890 11660 16892
rect 11716 16890 11740 16892
rect 11796 16890 11820 16892
rect 11876 16890 11882 16892
rect 11636 16838 11638 16890
rect 11818 16838 11820 16890
rect 11574 16836 11580 16838
rect 11636 16836 11660 16838
rect 11716 16836 11740 16838
rect 11796 16836 11820 16838
rect 11876 16836 11882 16838
rect 11574 16827 11882 16836
rect 11574 15804 11882 15813
rect 11574 15802 11580 15804
rect 11636 15802 11660 15804
rect 11716 15802 11740 15804
rect 11796 15802 11820 15804
rect 11876 15802 11882 15804
rect 11636 15750 11638 15802
rect 11818 15750 11820 15802
rect 11574 15748 11580 15750
rect 11636 15748 11660 15750
rect 11716 15748 11740 15750
rect 11796 15748 11820 15750
rect 11876 15748 11882 15750
rect 11574 15739 11882 15748
rect 11888 15496 11940 15502
rect 11978 15464 12034 15473
rect 11940 15444 11978 15450
rect 11888 15438 11978 15444
rect 11796 15428 11848 15434
rect 11900 15422 11978 15438
rect 11978 15399 12034 15408
rect 11796 15370 11848 15376
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11532 15026 11560 15098
rect 11808 15026 11836 15370
rect 12084 15026 12112 18362
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12636 17882 12664 18226
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12234 17436 12542 17445
rect 12234 17434 12240 17436
rect 12296 17434 12320 17436
rect 12376 17434 12400 17436
rect 12456 17434 12480 17436
rect 12536 17434 12542 17436
rect 12296 17382 12298 17434
rect 12478 17382 12480 17434
rect 12234 17380 12240 17382
rect 12296 17380 12320 17382
rect 12376 17380 12400 17382
rect 12456 17380 12480 17382
rect 12536 17380 12542 17382
rect 12234 17371 12542 17380
rect 12820 17338 12848 18566
rect 12912 18290 12940 18770
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12176 16130 12204 16390
rect 12234 16348 12542 16357
rect 12234 16346 12240 16348
rect 12296 16346 12320 16348
rect 12376 16346 12400 16348
rect 12456 16346 12480 16348
rect 12536 16346 12542 16348
rect 12296 16294 12298 16346
rect 12478 16294 12480 16346
rect 12234 16292 12240 16294
rect 12296 16292 12320 16294
rect 12376 16292 12400 16294
rect 12456 16292 12480 16294
rect 12536 16292 12542 16294
rect 12234 16283 12542 16292
rect 12912 16182 12940 18226
rect 13096 17610 13124 18838
rect 13360 18284 13412 18290
rect 13464 18272 13492 21014
rect 13556 20482 13584 21830
rect 13740 21706 13768 22066
rect 13648 21678 13768 21706
rect 14016 22066 14228 22094
rect 13648 21622 13676 21678
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13832 20482 13860 20742
rect 13924 20602 13952 20946
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13556 20454 13860 20482
rect 13740 18834 13768 20454
rect 13818 19272 13874 19281
rect 13818 19207 13820 19216
rect 13872 19207 13874 19216
rect 13820 19178 13872 19184
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13412 18244 13492 18272
rect 13360 18226 13412 18232
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 13096 17134 13124 17546
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12900 16176 12952 16182
rect 12176 16102 12296 16130
rect 12900 16118 12952 16124
rect 13464 16114 13492 18244
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 17338 13860 18158
rect 13924 17882 13952 18294
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13924 17202 13952 17818
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 12268 15502 12296 16102
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12360 15348 12388 15506
rect 13004 15434 13032 16050
rect 13188 15994 13216 16050
rect 13188 15966 13308 15994
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 12176 15320 12388 15348
rect 12624 15360 12676 15366
rect 12176 15162 12204 15320
rect 12624 15302 12676 15308
rect 12234 15260 12542 15269
rect 12234 15258 12240 15260
rect 12296 15258 12320 15260
rect 12376 15258 12400 15260
rect 12456 15258 12480 15260
rect 12536 15258 12542 15260
rect 12296 15206 12298 15258
rect 12478 15206 12480 15258
rect 12234 15204 12240 15206
rect 12296 15204 12320 15206
rect 12376 15204 12400 15206
rect 12456 15204 12480 15206
rect 12536 15204 12542 15206
rect 12234 15195 12542 15204
rect 12636 15162 12664 15302
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12348 15088 12400 15094
rect 12532 15088 12584 15094
rect 12400 15036 12532 15042
rect 12348 15030 12584 15036
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 12072 15020 12124 15026
rect 12360 15014 12572 15030
rect 12124 14980 12204 15008
rect 12072 14962 12124 14968
rect 11348 14878 11468 14906
rect 11348 14618 11376 14878
rect 11808 14872 11836 14962
rect 11808 14844 12020 14872
rect 11574 14716 11882 14725
rect 11574 14714 11580 14716
rect 11636 14714 11660 14716
rect 11716 14714 11740 14716
rect 11796 14714 11820 14716
rect 11876 14714 11882 14716
rect 11636 14662 11638 14714
rect 11818 14662 11820 14714
rect 11574 14660 11580 14662
rect 11636 14660 11660 14662
rect 11716 14660 11740 14662
rect 11796 14660 11820 14662
rect 11876 14660 11882 14662
rect 11574 14651 11882 14660
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11992 14278 12020 14844
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12084 14618 12112 14758
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12176 14521 12204 14980
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12162 14512 12218 14521
rect 12452 14482 12480 14894
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12162 14447 12218 14456
rect 12440 14476 12492 14482
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11440 13326 11468 13738
rect 11574 13628 11882 13637
rect 11574 13626 11580 13628
rect 11636 13626 11660 13628
rect 11716 13626 11740 13628
rect 11796 13626 11820 13628
rect 11876 13626 11882 13628
rect 11636 13574 11638 13626
rect 11818 13574 11820 13626
rect 11574 13572 11580 13574
rect 11636 13572 11660 13574
rect 11716 13572 11740 13574
rect 11796 13572 11820 13574
rect 11876 13572 11882 13574
rect 11574 13563 11882 13572
rect 12176 13326 12204 14447
rect 12440 14418 12492 14424
rect 12234 14172 12542 14181
rect 12234 14170 12240 14172
rect 12296 14170 12320 14172
rect 12376 14170 12400 14172
rect 12456 14170 12480 14172
rect 12536 14170 12542 14172
rect 12296 14118 12298 14170
rect 12478 14118 12480 14170
rect 12234 14116 12240 14118
rect 12296 14116 12320 14118
rect 12376 14116 12400 14118
rect 12456 14116 12480 14118
rect 12536 14116 12542 14118
rect 12234 14107 12542 14116
rect 11428 13320 11480 13326
rect 11612 13320 11664 13326
rect 11428 13262 11480 13268
rect 11518 13288 11574 13297
rect 11440 12918 11468 13262
rect 11574 13268 11612 13274
rect 11574 13262 11664 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11574 13246 11652 13262
rect 11796 13252 11848 13258
rect 11518 13223 11574 13232
rect 11796 13194 11848 13200
rect 11808 12986 11836 13194
rect 12234 13084 12542 13093
rect 12234 13082 12240 13084
rect 12296 13082 12320 13084
rect 12376 13082 12400 13084
rect 12456 13082 12480 13084
rect 12536 13082 12542 13084
rect 12296 13030 12298 13082
rect 12478 13030 12480 13082
rect 12234 13028 12240 13030
rect 12296 13028 12320 13030
rect 12376 13028 12400 13030
rect 12456 13028 12480 13030
rect 12536 13028 12542 13030
rect 12234 13019 12542 13028
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 12440 12844 12492 12850
rect 12636 12832 12664 14758
rect 13280 13530 13308 15966
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13372 14618 13400 15302
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12728 12850 12756 13262
rect 13280 12986 13308 13466
rect 13464 13394 13492 16050
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13542 15464 13598 15473
rect 13542 15399 13598 15408
rect 13556 15366 13584 15399
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14346 13584 14962
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12492 12804 12664 12832
rect 12716 12844 12768 12850
rect 12440 12786 12492 12792
rect 12716 12786 12768 12792
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 11574 12540 11882 12549
rect 11574 12538 11580 12540
rect 11636 12538 11660 12540
rect 11716 12538 11740 12540
rect 11796 12538 11820 12540
rect 11876 12538 11882 12540
rect 11636 12486 11638 12538
rect 11818 12486 11820 12538
rect 11574 12484 11580 12486
rect 11636 12484 11660 12486
rect 11716 12484 11740 12486
rect 11796 12484 11820 12486
rect 11876 12484 11882 12486
rect 11574 12475 11882 12484
rect 12820 12434 12848 12582
rect 13556 12434 13584 14282
rect 13832 14074 13860 15846
rect 13924 15502 13952 16050
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13924 15162 13952 15438
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 12728 12406 12848 12434
rect 13464 12406 13584 12434
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12084 11762 12112 12242
rect 12234 11996 12542 12005
rect 12234 11994 12240 11996
rect 12296 11994 12320 11996
rect 12376 11994 12400 11996
rect 12456 11994 12480 11996
rect 12536 11994 12542 11996
rect 12296 11942 12298 11994
rect 12478 11942 12480 11994
rect 12234 11940 12240 11942
rect 12296 11940 12320 11942
rect 12376 11940 12400 11942
rect 12456 11940 12480 11942
rect 12536 11940 12542 11942
rect 12234 11931 12542 11940
rect 12728 11898 12756 12406
rect 13464 12170 13492 12406
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 13464 11762 13492 12106
rect 13832 11898 13860 12786
rect 14016 12434 14044 22066
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14200 20466 14228 20878
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14292 20346 14320 22578
rect 14200 20318 14320 20346
rect 14200 19174 14228 20318
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14292 20058 14320 20198
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14384 18850 14412 24772
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14476 24410 14504 24686
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14476 23118 14504 23598
rect 14568 23322 14596 24686
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14568 23186 14596 23258
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14936 23118 14964 24618
rect 15028 24274 15056 25298
rect 16500 25208 16528 27406
rect 17144 27062 17172 27474
rect 17132 27056 17184 27062
rect 17132 26998 17184 27004
rect 17604 26194 17632 30194
rect 18657 29948 18965 29957
rect 18657 29946 18663 29948
rect 18719 29946 18743 29948
rect 18799 29946 18823 29948
rect 18879 29946 18903 29948
rect 18959 29946 18965 29948
rect 18719 29894 18721 29946
rect 18901 29894 18903 29946
rect 18657 29892 18663 29894
rect 18719 29892 18743 29894
rect 18799 29892 18823 29894
rect 18879 29892 18903 29894
rect 18959 29892 18965 29894
rect 18657 29883 18965 29892
rect 21928 29850 21956 30194
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 23940 29776 23992 29782
rect 23940 29718 23992 29724
rect 19156 29708 19208 29714
rect 19156 29650 19208 29656
rect 19168 29306 19196 29650
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 19317 29404 19625 29413
rect 19317 29402 19323 29404
rect 19379 29402 19403 29404
rect 19459 29402 19483 29404
rect 19539 29402 19563 29404
rect 19619 29402 19625 29404
rect 19379 29350 19381 29402
rect 19561 29350 19563 29402
rect 19317 29348 19323 29350
rect 19379 29348 19403 29350
rect 19459 29348 19483 29350
rect 19539 29348 19563 29350
rect 19619 29348 19625 29350
rect 19317 29339 19625 29348
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 20456 29238 20484 29446
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 18236 29164 18288 29170
rect 18236 29106 18288 29112
rect 18248 28626 18276 29106
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 18236 28620 18288 28626
rect 18236 28562 18288 28568
rect 17788 28218 17816 28562
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 17958 28248 18014 28257
rect 17776 28212 17828 28218
rect 17776 28154 17828 28160
rect 17868 28212 17920 28218
rect 17958 28183 18014 28192
rect 17868 28154 17920 28160
rect 17788 28082 17816 28154
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17776 28076 17828 28082
rect 17776 28018 17828 28024
rect 17696 27962 17724 28018
rect 17880 27962 17908 28154
rect 17696 27934 17908 27962
rect 17972 27878 18000 28183
rect 18064 28014 18092 28358
rect 18144 28076 18196 28082
rect 18144 28018 18196 28024
rect 18052 28008 18104 28014
rect 18052 27950 18104 27956
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 17776 27464 17828 27470
rect 17776 27406 17828 27412
rect 17604 26166 17724 26194
rect 16580 25220 16632 25226
rect 16408 25180 16580 25208
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 16120 24948 16172 24954
rect 16120 24890 16172 24896
rect 15304 24818 15332 24890
rect 15568 24880 15620 24886
rect 15568 24822 15620 24828
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15120 24313 15148 24550
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15106 24304 15162 24313
rect 15016 24268 15068 24274
rect 15106 24239 15162 24248
rect 15016 24210 15068 24216
rect 15108 24132 15160 24138
rect 15108 24074 15160 24080
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 15028 23322 15056 23666
rect 15120 23322 15148 24074
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14924 23112 14976 23118
rect 14924 23054 14976 23060
rect 15028 22982 15056 23258
rect 15212 23254 15240 23530
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 15304 23118 15332 24346
rect 15396 23730 15424 24754
rect 15580 23882 15608 24822
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15672 24698 15700 24754
rect 15936 24744 15988 24750
rect 15672 24692 15936 24698
rect 15672 24686 15988 24692
rect 15672 24670 15976 24686
rect 15672 24410 15700 24670
rect 16040 24562 16068 24754
rect 15764 24534 16068 24562
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15488 23866 15608 23882
rect 15488 23860 15620 23866
rect 15488 23854 15568 23860
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15384 23316 15436 23322
rect 15384 23258 15436 23264
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14476 21690 14504 22034
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14556 20800 14608 20806
rect 14476 20760 14556 20788
rect 14476 20466 14504 20760
rect 14556 20742 14608 20748
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14568 19514 14596 20402
rect 14660 20330 14688 22918
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 22234 14872 22374
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14752 21146 14780 21286
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 14660 19786 14688 20266
rect 14752 19854 14780 20402
rect 15028 20369 15056 20538
rect 15014 20360 15070 20369
rect 15014 20295 15070 20304
rect 15212 20074 15240 22986
rect 15396 22710 15424 23258
rect 15384 22704 15436 22710
rect 15384 22646 15436 22652
rect 15488 22574 15516 23854
rect 15568 23802 15620 23808
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15580 23254 15608 23666
rect 15568 23248 15620 23254
rect 15568 23190 15620 23196
rect 15764 23066 15792 24534
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15856 24070 15884 24346
rect 16028 24132 16080 24138
rect 16132 24120 16160 24890
rect 16304 24608 16356 24614
rect 16224 24568 16304 24596
rect 16224 24342 16252 24568
rect 16304 24550 16356 24556
rect 16212 24336 16264 24342
rect 16212 24278 16264 24284
rect 16302 24304 16358 24313
rect 16408 24274 16436 25180
rect 16580 25162 16632 25168
rect 17408 25220 17460 25226
rect 17408 25162 17460 25168
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17052 24886 17080 25094
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 16302 24239 16358 24248
rect 16396 24268 16448 24274
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16080 24092 16160 24120
rect 16028 24074 16080 24080
rect 15844 24064 15896 24070
rect 15844 24006 15896 24012
rect 16040 23662 16068 24074
rect 16224 24052 16252 24142
rect 16132 24024 16252 24052
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 15844 23588 15896 23594
rect 15844 23530 15896 23536
rect 15856 23254 15884 23530
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 15580 23050 15792 23066
rect 15568 23044 15792 23050
rect 15620 23038 15792 23044
rect 15568 22986 15620 22992
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15580 22506 15608 22986
rect 15856 22778 15884 23190
rect 16040 23186 16068 23598
rect 16132 23526 16160 24024
rect 16316 23798 16344 24239
rect 16396 24210 16448 24216
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16776 23866 16804 24006
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16960 23798 16988 24686
rect 17224 24268 17276 24274
rect 17224 24210 17276 24216
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16948 23792 17000 23798
rect 16948 23734 17000 23740
rect 17236 23730 17264 24210
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 16212 23588 16264 23594
rect 16212 23530 16264 23536
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 16028 23180 16080 23186
rect 16028 23122 16080 23128
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15936 22704 15988 22710
rect 15936 22646 15988 22652
rect 15568 22500 15620 22506
rect 15568 22442 15620 22448
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 14936 20046 15516 20074
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14292 18822 14412 18850
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 14108 17134 14136 18634
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16590 14136 16934
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14108 15609 14136 16118
rect 14094 15600 14150 15609
rect 14094 15535 14150 15544
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 13924 12406 14044 12434
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 11574 11452 11882 11461
rect 11574 11450 11580 11452
rect 11636 11450 11660 11452
rect 11716 11450 11740 11452
rect 11796 11450 11820 11452
rect 11876 11450 11882 11452
rect 11636 11398 11638 11450
rect 11818 11398 11820 11450
rect 11574 11396 11580 11398
rect 11636 11396 11660 11398
rect 11716 11396 11740 11398
rect 11796 11396 11820 11398
rect 11876 11396 11882 11398
rect 11574 11387 11882 11396
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11428 10600 11480 10606
rect 11334 10568 11390 10577
rect 11428 10542 11480 10548
rect 11334 10503 11390 10512
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10980 10062 11008 10202
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9722 10916 9862
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10796 9586 11008 9602
rect 10796 9580 11020 9586
rect 10796 9574 10968 9580
rect 10796 9466 10824 9574
rect 10968 9522 11020 9528
rect 11072 9518 11100 9998
rect 11348 9994 11376 10503
rect 11440 10062 11468 10542
rect 11574 10364 11882 10373
rect 11574 10362 11580 10364
rect 11636 10362 11660 10364
rect 11716 10362 11740 10364
rect 11796 10362 11820 10364
rect 11876 10362 11882 10364
rect 11636 10310 11638 10362
rect 11818 10310 11820 10362
rect 11574 10308 11580 10310
rect 11636 10308 11660 10310
rect 11716 10308 11740 10310
rect 11796 10308 11820 10310
rect 11876 10308 11882 10310
rect 11574 10299 11882 10308
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11348 9897 11376 9930
rect 11334 9888 11390 9897
rect 11334 9823 11390 9832
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 10704 9450 10824 9466
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10692 9444 10824 9450
rect 10744 9438 10824 9444
rect 10692 9386 10744 9392
rect 10416 9104 10468 9110
rect 9954 9072 10010 9081
rect 9864 9036 9916 9042
rect 10416 9046 10468 9052
rect 11242 9072 11298 9081
rect 9954 9007 10010 9016
rect 10140 9036 10192 9042
rect 9864 8978 9916 8984
rect 10140 8978 10192 8984
rect 11060 9036 11112 9042
rect 11242 9007 11244 9016
rect 11060 8978 11112 8984
rect 11296 9007 11298 9016
rect 11244 8978 11296 8984
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9968 8634 9996 8774
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 6254 9720 7278
rect 9876 6866 9904 7754
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9864 6724 9916 6730
rect 9968 6712 9996 7890
rect 10152 6934 10180 8978
rect 10782 8256 10838 8265
rect 10782 8191 10838 8200
rect 10598 8120 10654 8129
rect 10598 8055 10654 8064
rect 10612 7410 10640 8055
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10796 7342 10824 8191
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 11072 7206 11100 8978
rect 11348 8906 11376 9590
rect 11992 9586 12020 10066
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11574 9276 11882 9285
rect 11574 9274 11580 9276
rect 11636 9274 11660 9276
rect 11716 9274 11740 9276
rect 11796 9274 11820 9276
rect 11876 9274 11882 9276
rect 11636 9222 11638 9274
rect 11818 9222 11820 9274
rect 11574 9220 11580 9222
rect 11636 9220 11660 9222
rect 11716 9220 11740 9222
rect 11796 9220 11820 9222
rect 11876 9220 11882 9222
rect 11574 9211 11882 9220
rect 11336 8900 11388 8906
rect 11256 8860 11336 8888
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 10152 6798 10180 6870
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9916 6684 9996 6712
rect 10048 6724 10100 6730
rect 9864 6666 9916 6672
rect 10048 6666 10100 6672
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9784 6118 9812 6666
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9876 5778 9904 6326
rect 10060 5914 10088 6666
rect 10152 6322 10180 6734
rect 10244 6458 10272 6734
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10428 6322 10456 6938
rect 11072 6882 11100 7142
rect 10520 6854 11100 6882
rect 11164 6866 11192 7142
rect 11256 7002 11284 8860
rect 11336 8842 11388 8848
rect 11574 8188 11882 8197
rect 11574 8186 11580 8188
rect 11636 8186 11660 8188
rect 11716 8186 11740 8188
rect 11796 8186 11820 8188
rect 11876 8186 11882 8188
rect 11636 8134 11638 8186
rect 11818 8134 11820 8186
rect 11574 8132 11580 8134
rect 11636 8132 11660 8134
rect 11716 8132 11740 8134
rect 11796 8132 11820 8134
rect 11876 8132 11882 8134
rect 11574 8123 11882 8132
rect 11992 8072 12020 9522
rect 12084 9042 12112 9862
rect 12176 9625 12204 11290
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 12234 10908 12542 10917
rect 12234 10906 12240 10908
rect 12296 10906 12320 10908
rect 12376 10906 12400 10908
rect 12456 10906 12480 10908
rect 12536 10906 12542 10908
rect 12296 10854 12298 10906
rect 12478 10854 12480 10906
rect 12234 10852 12240 10854
rect 12296 10852 12320 10854
rect 12376 10852 12400 10854
rect 12456 10852 12480 10854
rect 12536 10852 12542 10854
rect 12234 10843 12542 10852
rect 12622 10840 12678 10849
rect 12622 10775 12678 10784
rect 12636 10266 12664 10775
rect 13266 10704 13322 10713
rect 13556 10674 13584 10950
rect 13266 10639 13322 10648
rect 13544 10668 13596 10674
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 13280 10198 13308 10639
rect 13544 10610 13596 10616
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10266 13584 10406
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13358 10024 13414 10033
rect 13358 9959 13360 9968
rect 13412 9959 13414 9968
rect 13360 9930 13412 9936
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12234 9820 12542 9829
rect 12234 9818 12240 9820
rect 12296 9818 12320 9820
rect 12376 9818 12400 9820
rect 12456 9818 12480 9820
rect 12536 9818 12542 9820
rect 12296 9766 12298 9818
rect 12478 9766 12480 9818
rect 12234 9764 12240 9766
rect 12296 9764 12320 9766
rect 12376 9764 12400 9766
rect 12456 9764 12480 9766
rect 12536 9764 12542 9766
rect 12234 9755 12542 9764
rect 12162 9616 12218 9625
rect 12162 9551 12218 9560
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11900 8044 12020 8072
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11348 6934 11376 7346
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11440 6866 11468 7346
rect 11900 7206 11928 8044
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11574 7100 11882 7109
rect 11574 7098 11580 7100
rect 11636 7098 11660 7100
rect 11716 7098 11740 7100
rect 11796 7098 11820 7100
rect 11876 7098 11882 7100
rect 11636 7046 11638 7098
rect 11818 7046 11820 7098
rect 11574 7044 11580 7046
rect 11636 7044 11660 7046
rect 11716 7044 11740 7046
rect 11796 7044 11820 7046
rect 11876 7044 11882 7046
rect 11574 7035 11882 7044
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11152 6860 11204 6866
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10152 5778 10180 6258
rect 10520 6254 10548 6854
rect 11152 6802 11204 6808
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11060 6792 11112 6798
rect 10966 6760 11022 6769
rect 10600 6724 10652 6730
rect 11060 6734 11112 6740
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 10966 6695 11022 6704
rect 10600 6666 10652 6672
rect 10612 6390 10640 6666
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10980 6322 11008 6695
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10152 5574 10180 5714
rect 10520 5710 10548 6190
rect 11072 5914 11100 6734
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6322 11192 6598
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11164 6186 11192 6258
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 8956 4690 8984 5306
rect 9324 4690 9352 5510
rect 9692 5098 9720 5510
rect 9784 5234 9812 5510
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 10152 5166 10180 5510
rect 10520 5302 10548 5646
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 10244 4826 10272 5170
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10704 4826 10732 5102
rect 11072 4826 11100 5850
rect 11164 5794 11192 6122
rect 11164 5766 11284 5794
rect 11256 5710 11284 5766
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11164 5574 11192 5646
rect 11348 5642 11376 6734
rect 11716 6730 11744 6938
rect 11992 6798 12020 7142
rect 12084 6934 12112 8978
rect 12176 8974 12204 9551
rect 13096 9178 13124 9862
rect 13176 9648 13228 9654
rect 13174 9616 13176 9625
rect 13228 9616 13230 9625
rect 13174 9551 13230 9560
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 12234 8732 12542 8741
rect 12234 8730 12240 8732
rect 12296 8730 12320 8732
rect 12376 8730 12400 8732
rect 12456 8730 12480 8732
rect 12536 8730 12542 8732
rect 12296 8678 12298 8730
rect 12478 8678 12480 8730
rect 12234 8676 12240 8678
rect 12296 8676 12320 8678
rect 12376 8676 12400 8678
rect 12456 8676 12480 8678
rect 12536 8676 12542 8678
rect 12234 8667 12542 8676
rect 13280 8634 13308 8842
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8430 13400 9930
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13464 8430 13492 9590
rect 13648 9382 13676 11630
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10690 13860 10950
rect 13740 10674 13860 10690
rect 13728 10668 13860 10674
rect 13780 10662 13860 10668
rect 13728 10610 13780 10616
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9654 13860 9862
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13924 9024 13952 12406
rect 14108 12209 14136 13670
rect 14094 12200 14150 12209
rect 14094 12135 14150 12144
rect 14108 11762 14136 12135
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 14016 10606 14044 10746
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14016 9518 14044 10542
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 13832 8996 13952 9024
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 8566 13676 8774
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12176 7410 12204 8298
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 12234 7644 12542 7653
rect 12234 7642 12240 7644
rect 12296 7642 12320 7644
rect 12376 7642 12400 7644
rect 12456 7642 12480 7644
rect 12536 7642 12542 7644
rect 12296 7590 12298 7642
rect 12478 7590 12480 7642
rect 12234 7588 12240 7590
rect 12296 7588 12320 7590
rect 12376 7588 12400 7590
rect 12456 7588 12480 7590
rect 12536 7588 12542 7590
rect 12234 7579 12542 7588
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12360 7002 12388 7482
rect 13372 7410 13400 7686
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13464 7392 13492 8366
rect 13740 7818 13768 8910
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13544 7404 13596 7410
rect 13464 7364 13544 7392
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6458 12204 6598
rect 12234 6556 12542 6565
rect 12234 6554 12240 6556
rect 12296 6554 12320 6556
rect 12376 6554 12400 6556
rect 12456 6554 12480 6556
rect 12536 6554 12542 6556
rect 12296 6502 12298 6554
rect 12478 6502 12480 6554
rect 12234 6500 12240 6502
rect 12296 6500 12320 6502
rect 12376 6500 12400 6502
rect 12456 6500 12480 6502
rect 12536 6500 12542 6502
rect 12234 6491 12542 6500
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 11440 5778 11468 6394
rect 13464 6254 13492 7364
rect 13544 7346 13596 7352
rect 13648 6866 13676 7754
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 11574 6012 11882 6021
rect 11574 6010 11580 6012
rect 11636 6010 11660 6012
rect 11716 6010 11740 6012
rect 11796 6010 11820 6012
rect 11876 6010 11882 6012
rect 11636 5958 11638 6010
rect 11818 5958 11820 6010
rect 11574 5956 11580 5958
rect 11636 5956 11660 5958
rect 11716 5956 11740 5958
rect 11796 5956 11820 5958
rect 11876 5956 11882 5958
rect 11574 5947 11882 5956
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11348 5166 11376 5578
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 11348 4622 11376 5102
rect 11440 4826 11468 5578
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5234 11836 5510
rect 12234 5468 12542 5477
rect 12234 5466 12240 5468
rect 12296 5466 12320 5468
rect 12376 5466 12400 5468
rect 12456 5466 12480 5468
rect 12536 5466 12542 5468
rect 12296 5414 12298 5466
rect 12478 5414 12480 5466
rect 12234 5412 12240 5414
rect 12296 5412 12320 5414
rect 12376 5412 12400 5414
rect 12456 5412 12480 5414
rect 12536 5412 12542 5414
rect 12234 5403 12542 5412
rect 12636 5370 12664 6190
rect 13832 5370 13860 8996
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13924 8294 13952 8842
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7750 13952 8230
rect 14016 7954 14044 9454
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14108 7886 14136 8026
rect 14200 8022 14228 17546
rect 14292 14414 14320 18822
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14384 18426 14412 18634
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14660 18358 14688 18566
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14384 16522 14412 17070
rect 14660 16794 14688 17478
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14752 16590 14780 19790
rect 14936 19514 14964 20046
rect 15106 19952 15162 19961
rect 15106 19887 15162 19896
rect 15120 19854 15148 19887
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15488 19514 15516 20046
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15108 19440 15160 19446
rect 15160 19400 15424 19428
rect 15108 19382 15160 19388
rect 15396 19334 15424 19400
rect 15764 19334 15792 20810
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15396 19306 15792 19334
rect 15856 19310 15884 19722
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15396 18850 15424 19110
rect 15488 18970 15516 19110
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15568 18896 15620 18902
rect 15396 18844 15568 18850
rect 15396 18838 15620 18844
rect 15396 18822 15608 18838
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15488 18358 15516 18634
rect 15764 18612 15792 19306
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15856 18970 15884 19246
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15844 18624 15896 18630
rect 15764 18584 15844 18612
rect 15476 18352 15528 18358
rect 15528 18312 15608 18340
rect 15476 18294 15528 18300
rect 15580 18222 15608 18312
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 15120 17270 15148 17750
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 15488 17134 15516 18158
rect 15764 17270 15792 18584
rect 15844 18566 15896 18572
rect 15948 17882 15976 22646
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 16040 19378 16068 20878
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16040 18970 16068 19314
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 16040 18766 16068 18906
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 14740 16584 14792 16590
rect 14924 16584 14976 16590
rect 14740 16526 14792 16532
rect 14844 16544 14924 16572
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14384 14958 14412 15506
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14844 14822 14872 16544
rect 14924 16526 14976 16532
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14384 14074 14412 14418
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14476 12850 14504 13194
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14292 11830 14320 12271
rect 14384 12238 14412 12786
rect 14752 12782 14780 14758
rect 14844 13938 14872 14758
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14568 12238 14596 12718
rect 14752 12442 14780 12718
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14372 12232 14424 12238
rect 14556 12232 14608 12238
rect 14372 12174 14424 12180
rect 14476 12192 14556 12220
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14292 9382 14320 9590
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 8566 14320 9318
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14096 7880 14148 7886
rect 14148 7840 14228 7868
rect 14096 7822 14148 7828
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13924 6934 13952 7686
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 13912 6792 13964 6798
rect 13910 6760 13912 6769
rect 14016 6780 14044 7686
rect 14200 7342 14228 7840
rect 14292 7478 14320 8502
rect 14476 8090 14504 12192
rect 14556 12174 14608 12180
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14568 11014 14596 11494
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14568 10810 14596 10950
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14660 7886 14688 11698
rect 14936 10674 14964 16118
rect 15028 15706 15056 16458
rect 15108 16448 15160 16454
rect 15292 16448 15344 16454
rect 15160 16408 15240 16436
rect 15108 16390 15160 16396
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15028 12238 15056 15642
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15120 13258 15148 13738
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15212 12434 15240 16408
rect 15292 16390 15344 16396
rect 15304 16046 15332 16390
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15304 13462 15332 15846
rect 15488 15162 15516 16526
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 15910 15700 16458
rect 15764 16096 15792 17206
rect 15844 16108 15896 16114
rect 15764 16068 15844 16096
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15672 15162 15700 15370
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 13802 15516 14894
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15580 14006 15608 14214
rect 15672 14074 15700 14214
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15212 12406 15424 12434
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15212 11354 15240 12174
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 8090 14780 10406
rect 15304 10062 15332 10542
rect 15396 10062 15424 12406
rect 15580 11744 15608 13942
rect 15764 13734 15792 16068
rect 15844 16050 15896 16056
rect 15948 15144 15976 17818
rect 16040 16980 16068 18702
rect 16132 18442 16160 23054
rect 16224 20874 16252 23530
rect 17236 22982 17264 23666
rect 17420 23322 17448 25162
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17604 24070 17632 24550
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17604 23662 17632 24006
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16396 22500 16448 22506
rect 16396 22442 16448 22448
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16224 20534 16252 20810
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 16408 18766 16436 22442
rect 16500 22098 16528 22510
rect 16488 22094 16540 22098
rect 16488 22092 16620 22094
rect 16540 22066 16620 22092
rect 16488 22034 16540 22040
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16132 18414 16252 18442
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16132 17678 16160 18022
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16132 17270 16160 17614
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 16120 16992 16172 16998
rect 16040 16952 16120 16980
rect 16120 16934 16172 16940
rect 16132 16114 16160 16934
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16040 15434 16068 15846
rect 16132 15706 16160 15846
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16028 15428 16080 15434
rect 16028 15370 16080 15376
rect 16028 15156 16080 15162
rect 15948 15116 16028 15144
rect 16028 15098 16080 15104
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16040 14498 16068 14962
rect 16132 14618 16160 15098
rect 16224 15026 16252 18414
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16316 15706 16344 15846
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16224 14906 16252 14962
rect 16224 14878 16344 14906
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14618 16252 14758
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16040 14470 16160 14498
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15764 12986 15792 13262
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15660 11756 15712 11762
rect 15580 11716 15660 11744
rect 15660 11698 15712 11704
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15488 10062 15516 10610
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 14476 7750 14504 7822
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14292 7188 14320 7414
rect 13964 6760 14044 6780
rect 13966 6752 14044 6760
rect 14200 7160 14320 7188
rect 13910 6695 13966 6704
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6458 14136 6598
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14200 6390 14228 7160
rect 14476 7002 14504 7686
rect 14660 7546 14688 7686
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 15120 7342 15148 7822
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 14200 5234 14228 6326
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 12440 5160 12492 5166
rect 12716 5160 12768 5166
rect 12492 5120 12716 5148
rect 12440 5102 12492 5108
rect 12716 5102 12768 5108
rect 11574 4924 11882 4933
rect 11574 4922 11580 4924
rect 11636 4922 11660 4924
rect 11716 4922 11740 4924
rect 11796 4922 11820 4924
rect 11876 4922 11882 4924
rect 11636 4870 11638 4922
rect 11818 4870 11820 4922
rect 11574 4868 11580 4870
rect 11636 4868 11660 4870
rect 11716 4868 11740 4870
rect 11796 4868 11820 4870
rect 11876 4868 11882 4870
rect 11574 4859 11882 4868
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 5151 4380 5459 4389
rect 5151 4378 5157 4380
rect 5213 4378 5237 4380
rect 5293 4378 5317 4380
rect 5373 4378 5397 4380
rect 5453 4378 5459 4380
rect 5213 4326 5215 4378
rect 5395 4326 5397 4378
rect 5151 4324 5157 4326
rect 5213 4324 5237 4326
rect 5293 4324 5317 4326
rect 5373 4324 5397 4326
rect 5453 4324 5459 4326
rect 5151 4315 5459 4324
rect 12234 4380 12542 4389
rect 12234 4378 12240 4380
rect 12296 4378 12320 4380
rect 12376 4378 12400 4380
rect 12456 4378 12480 4380
rect 12536 4378 12542 4380
rect 12296 4326 12298 4378
rect 12478 4326 12480 4378
rect 12234 4324 12240 4326
rect 12296 4324 12320 4326
rect 12376 4324 12400 4326
rect 12456 4324 12480 4326
rect 12536 4324 12542 4326
rect 12234 4315 12542 4324
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 2410 3975 2466 3984
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3738 2268 3878
rect 4491 3836 4799 3845
rect 4491 3834 4497 3836
rect 4553 3834 4577 3836
rect 4633 3834 4657 3836
rect 4713 3834 4737 3836
rect 4793 3834 4799 3836
rect 4553 3782 4555 3834
rect 4735 3782 4737 3834
rect 4491 3780 4497 3782
rect 4553 3780 4577 3782
rect 4633 3780 4657 3782
rect 4713 3780 4737 3782
rect 4793 3780 4799 3782
rect 4491 3771 4799 3780
rect 11574 3836 11882 3845
rect 11574 3834 11580 3836
rect 11636 3834 11660 3836
rect 11716 3834 11740 3836
rect 11796 3834 11820 3836
rect 11876 3834 11882 3836
rect 11636 3782 11638 3834
rect 11818 3782 11820 3834
rect 11574 3780 11580 3782
rect 11636 3780 11660 3782
rect 11716 3780 11740 3782
rect 11796 3780 11820 3782
rect 11876 3780 11882 3782
rect 11574 3771 11882 3780
rect 12636 3738 12664 4218
rect 13004 4146 13032 4558
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12898 3632 12954 3641
rect 12898 3567 12900 3576
rect 12952 3567 12954 3576
rect 12900 3538 12952 3544
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 952 3398 980 3431
rect 940 3392 992 3398
rect 940 3334 992 3340
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 2240 2446 2268 3334
rect 5151 3292 5459 3301
rect 5151 3290 5157 3292
rect 5213 3290 5237 3292
rect 5293 3290 5317 3292
rect 5373 3290 5397 3292
rect 5453 3290 5459 3292
rect 5213 3238 5215 3290
rect 5395 3238 5397 3290
rect 5151 3236 5157 3238
rect 5213 3236 5237 3238
rect 5293 3236 5317 3238
rect 5373 3236 5397 3238
rect 5453 3236 5459 3238
rect 5151 3227 5459 3236
rect 12234 3292 12542 3301
rect 12234 3290 12240 3292
rect 12296 3290 12320 3292
rect 12376 3290 12400 3292
rect 12456 3290 12480 3292
rect 12536 3290 12542 3292
rect 12296 3238 12298 3290
rect 12478 3238 12480 3290
rect 12234 3236 12240 3238
rect 12296 3236 12320 3238
rect 12376 3236 12400 3238
rect 12456 3236 12480 3238
rect 12536 3236 12542 3238
rect 12234 3227 12542 3236
rect 4491 2748 4799 2757
rect 4491 2746 4497 2748
rect 4553 2746 4577 2748
rect 4633 2746 4657 2748
rect 4713 2746 4737 2748
rect 4793 2746 4799 2748
rect 4553 2694 4555 2746
rect 4735 2694 4737 2746
rect 4491 2692 4497 2694
rect 4553 2692 4577 2694
rect 4633 2692 4657 2694
rect 4713 2692 4737 2694
rect 4793 2692 4799 2694
rect 4491 2683 4799 2692
rect 11574 2748 11882 2757
rect 11574 2746 11580 2748
rect 11636 2746 11660 2748
rect 11716 2746 11740 2748
rect 11796 2746 11820 2748
rect 11876 2746 11882 2748
rect 11636 2694 11638 2746
rect 11818 2694 11820 2746
rect 11574 2692 11580 2694
rect 11636 2692 11660 2694
rect 11716 2692 11740 2694
rect 11796 2692 11820 2694
rect 11876 2692 11882 2694
rect 11574 2683 11882 2692
rect 12820 2650 12848 3334
rect 13004 3194 13032 4082
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13096 3194 13124 3878
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13188 2446 13216 2790
rect 13280 2650 13308 4558
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13372 3534 13400 4014
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13556 3534 13584 3878
rect 13924 3670 13952 3878
rect 14016 3670 14044 4490
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14646 4176 14702 4185
rect 14646 4111 14648 4120
rect 14700 4111 14702 4120
rect 14648 4082 14700 4088
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13372 2922 13400 3470
rect 13544 3052 13596 3058
rect 13648 3040 13676 3538
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3058 13768 3334
rect 13832 3058 13860 3470
rect 13924 3466 13952 3606
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13924 3058 13952 3402
rect 14016 3058 14044 3606
rect 14108 3602 14136 4014
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14476 3534 14504 3946
rect 14660 3738 14688 4082
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14464 3528 14516 3534
rect 14108 3476 14464 3482
rect 14108 3470 14516 3476
rect 14108 3454 14504 3470
rect 14108 3126 14136 3454
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14292 3058 14320 3334
rect 14660 3058 14688 3674
rect 14844 3534 14872 4218
rect 15212 4146 15240 9862
rect 15672 9042 15700 11698
rect 16040 11642 16068 14350
rect 16132 12850 16160 14470
rect 16316 14414 16344 14878
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16132 12753 16160 12786
rect 16118 12744 16174 12753
rect 16118 12679 16174 12688
rect 16408 12306 16436 15030
rect 16500 14414 16528 21830
rect 16592 21486 16620 22066
rect 16684 21894 16712 22510
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16592 20942 16620 21422
rect 16960 21146 16988 21422
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16592 18426 16620 20878
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16868 20058 16896 20402
rect 16960 20058 16988 20810
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 17052 20058 17080 20266
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 16868 19514 16896 19790
rect 17236 19514 17264 20402
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17328 18766 17356 22986
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 17500 20800 17552 20806
rect 17420 20760 17500 20788
rect 17420 20466 17448 20760
rect 17500 20742 17552 20748
rect 17604 20466 17632 22918
rect 17696 22001 17724 26166
rect 17788 25362 17816 27406
rect 18064 26858 18092 27814
rect 18156 27674 18184 28018
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 18248 27470 18276 28562
rect 18340 28014 18368 28902
rect 18432 28694 18460 29038
rect 19892 28960 19944 28966
rect 19892 28902 19944 28908
rect 18657 28860 18965 28869
rect 18657 28858 18663 28860
rect 18719 28858 18743 28860
rect 18799 28858 18823 28860
rect 18879 28858 18903 28860
rect 18959 28858 18965 28860
rect 18719 28806 18721 28858
rect 18901 28806 18903 28858
rect 18657 28804 18663 28806
rect 18719 28804 18743 28806
rect 18799 28804 18823 28806
rect 18879 28804 18903 28806
rect 18959 28804 18965 28806
rect 18657 28795 18965 28804
rect 18420 28688 18472 28694
rect 18420 28630 18472 28636
rect 18432 28014 18460 28630
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19352 28404 19380 28494
rect 19260 28376 19380 28404
rect 19708 28416 19760 28422
rect 19260 28200 19288 28376
rect 19708 28358 19760 28364
rect 19317 28316 19625 28325
rect 19317 28314 19323 28316
rect 19379 28314 19403 28316
rect 19459 28314 19483 28316
rect 19539 28314 19563 28316
rect 19619 28314 19625 28316
rect 19379 28262 19381 28314
rect 19561 28262 19563 28314
rect 19317 28260 19323 28262
rect 19379 28260 19403 28262
rect 19459 28260 19483 28262
rect 19539 28260 19563 28262
rect 19619 28260 19625 28262
rect 19317 28251 19625 28260
rect 19260 28172 19472 28200
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 18420 28008 18472 28014
rect 18420 27950 18472 27956
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 18657 27772 18965 27781
rect 18657 27770 18663 27772
rect 18719 27770 18743 27772
rect 18799 27770 18823 27772
rect 18879 27770 18903 27772
rect 18959 27770 18965 27772
rect 18719 27718 18721 27770
rect 18901 27718 18903 27770
rect 18657 27716 18663 27718
rect 18719 27716 18743 27718
rect 18799 27716 18823 27718
rect 18879 27716 18903 27718
rect 18959 27716 18965 27718
rect 18657 27707 18965 27716
rect 19352 27674 19380 27950
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19444 27538 19472 28172
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19720 27470 19748 28358
rect 19812 28121 19840 28494
rect 19798 28112 19854 28121
rect 19798 28047 19854 28056
rect 19904 27878 19932 28902
rect 20824 28762 20852 29582
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 20812 28756 20864 28762
rect 20812 28698 20864 28704
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 20260 28416 20312 28422
rect 20260 28358 20312 28364
rect 20272 27946 20300 28358
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20260 27940 20312 27946
rect 20260 27882 20312 27888
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 19904 27538 19932 27814
rect 19800 27532 19852 27538
rect 19800 27474 19852 27480
rect 19892 27532 19944 27538
rect 19892 27474 19944 27480
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 19708 27464 19760 27470
rect 19708 27406 19760 27412
rect 19317 27228 19625 27237
rect 19317 27226 19323 27228
rect 19379 27226 19403 27228
rect 19459 27226 19483 27228
rect 19539 27226 19563 27228
rect 19619 27226 19625 27228
rect 19379 27174 19381 27226
rect 19561 27174 19563 27226
rect 19317 27172 19323 27174
rect 19379 27172 19403 27174
rect 19459 27172 19483 27174
rect 19539 27172 19563 27174
rect 19619 27172 19625 27174
rect 19317 27163 19625 27172
rect 19812 27130 19840 27474
rect 19800 27124 19852 27130
rect 19800 27066 19852 27072
rect 18052 26852 18104 26858
rect 18052 26794 18104 26800
rect 18657 26684 18965 26693
rect 18657 26682 18663 26684
rect 18719 26682 18743 26684
rect 18799 26682 18823 26684
rect 18879 26682 18903 26684
rect 18959 26682 18965 26684
rect 18719 26630 18721 26682
rect 18901 26630 18903 26682
rect 18657 26628 18663 26630
rect 18719 26628 18743 26630
rect 18799 26628 18823 26630
rect 18879 26628 18903 26630
rect 18959 26628 18965 26630
rect 18657 26619 18965 26628
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17776 25356 17828 25362
rect 17776 25298 17828 25304
rect 17788 24206 17816 25298
rect 17880 25294 17908 25774
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 17972 24818 18000 26318
rect 19800 26308 19852 26314
rect 19800 26250 19852 26256
rect 19317 26140 19625 26149
rect 19317 26138 19323 26140
rect 19379 26138 19403 26140
rect 19459 26138 19483 26140
rect 19539 26138 19563 26140
rect 19619 26138 19625 26140
rect 19379 26086 19381 26138
rect 19561 26086 19563 26138
rect 19317 26084 19323 26086
rect 19379 26084 19403 26086
rect 19459 26084 19483 26086
rect 19539 26084 19563 26086
rect 19619 26084 19625 26086
rect 19317 26075 19625 26084
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 18144 25424 18196 25430
rect 18144 25366 18196 25372
rect 18156 24818 18184 25366
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17682 21992 17738 22001
rect 17788 21962 17816 24142
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 18064 23662 18092 24074
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18064 22982 18092 23598
rect 18156 23254 18184 24754
rect 18248 24682 18276 25910
rect 18657 25596 18965 25605
rect 18657 25594 18663 25596
rect 18719 25594 18743 25596
rect 18799 25594 18823 25596
rect 18879 25594 18903 25596
rect 18959 25594 18965 25596
rect 18719 25542 18721 25594
rect 18901 25542 18903 25594
rect 18657 25540 18663 25542
rect 18719 25540 18743 25542
rect 18799 25540 18823 25542
rect 18879 25540 18903 25542
rect 18959 25540 18965 25542
rect 18657 25531 18965 25540
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18892 25294 18920 25434
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19708 25356 19760 25362
rect 19708 25298 19760 25304
rect 18788 25288 18840 25294
rect 18340 25248 18788 25276
rect 18340 24886 18368 25248
rect 18788 25230 18840 25236
rect 18880 25288 18932 25294
rect 19064 25288 19116 25294
rect 18880 25230 18932 25236
rect 18984 25248 19064 25276
rect 18420 25152 18472 25158
rect 18420 25094 18472 25100
rect 18432 24886 18460 25094
rect 18328 24880 18380 24886
rect 18328 24822 18380 24828
rect 18420 24880 18472 24886
rect 18420 24822 18472 24828
rect 18984 24834 19012 25248
rect 19064 25230 19116 25236
rect 19156 25152 19208 25158
rect 19156 25094 19208 25100
rect 19168 24970 19196 25094
rect 19076 24954 19196 24970
rect 19064 24948 19196 24954
rect 19116 24942 19196 24948
rect 19064 24890 19116 24896
rect 18236 24676 18288 24682
rect 18236 24618 18288 24624
rect 18144 23248 18196 23254
rect 18144 23190 18196 23196
rect 18340 23118 18368 24822
rect 18984 24806 19104 24834
rect 18657 24508 18965 24517
rect 18657 24506 18663 24508
rect 18719 24506 18743 24508
rect 18799 24506 18823 24508
rect 18879 24506 18903 24508
rect 18959 24506 18965 24508
rect 18719 24454 18721 24506
rect 18901 24454 18903 24506
rect 18657 24452 18663 24454
rect 18719 24452 18743 24454
rect 18799 24452 18823 24454
rect 18879 24452 18903 24454
rect 18959 24452 18965 24454
rect 18657 24443 18965 24452
rect 19076 24206 19104 24806
rect 19260 24410 19288 25298
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19536 25158 19564 25230
rect 19524 25152 19576 25158
rect 19524 25094 19576 25100
rect 19317 25052 19625 25061
rect 19317 25050 19323 25052
rect 19379 25050 19403 25052
rect 19459 25050 19483 25052
rect 19539 25050 19563 25052
rect 19619 25050 19625 25052
rect 19379 24998 19381 25050
rect 19561 24998 19563 25050
rect 19317 24996 19323 24998
rect 19379 24996 19403 24998
rect 19459 24996 19483 24998
rect 19539 24996 19563 24998
rect 19619 24996 19625 24998
rect 19317 24987 19625 24996
rect 19720 24410 19748 25298
rect 19812 25294 19840 26250
rect 19904 25362 19932 27474
rect 20272 27402 20300 27882
rect 20732 27538 20760 28018
rect 20720 27532 20772 27538
rect 20720 27474 20772 27480
rect 20260 27396 20312 27402
rect 20260 27338 20312 27344
rect 20732 27062 20760 27474
rect 20824 27112 20852 28494
rect 21192 28082 21220 29106
rect 22100 29096 22152 29102
rect 22100 29038 22152 29044
rect 22192 29096 22244 29102
rect 22192 29038 22244 29044
rect 21916 29028 21968 29034
rect 21916 28970 21968 28976
rect 21272 28960 21324 28966
rect 21272 28902 21324 28908
rect 21364 28960 21416 28966
rect 21364 28902 21416 28908
rect 21732 28960 21784 28966
rect 21732 28902 21784 28908
rect 21284 28626 21312 28902
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 21376 28558 21404 28902
rect 21744 28762 21772 28902
rect 21732 28756 21784 28762
rect 21732 28698 21784 28704
rect 21364 28552 21416 28558
rect 21364 28494 21416 28500
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 21192 27402 21220 28018
rect 21652 28014 21680 28494
rect 21744 28422 21772 28698
rect 21928 28558 21956 28970
rect 22112 28762 22140 29038
rect 22008 28756 22060 28762
rect 22008 28698 22060 28704
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 22020 28665 22048 28698
rect 22006 28656 22062 28665
rect 22006 28591 22062 28600
rect 21916 28552 21968 28558
rect 21916 28494 21968 28500
rect 22204 28490 22232 29038
rect 22376 29028 22428 29034
rect 22376 28970 22428 28976
rect 22388 28558 22416 28970
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22008 28484 22060 28490
rect 22192 28484 22244 28490
rect 22060 28444 22140 28472
rect 22008 28426 22060 28432
rect 21732 28416 21784 28422
rect 21732 28358 21784 28364
rect 22112 28218 22140 28444
rect 22192 28426 22244 28432
rect 22744 28484 22796 28490
rect 22744 28426 22796 28432
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 21640 28008 21692 28014
rect 21916 28008 21968 28014
rect 21640 27950 21692 27956
rect 21914 27976 21916 27985
rect 21968 27976 21970 27985
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 20904 27124 20956 27130
rect 20824 27084 20904 27112
rect 20904 27066 20956 27072
rect 20720 27056 20772 27062
rect 20720 26998 20772 27004
rect 21008 26790 21036 27270
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 19892 25356 19944 25362
rect 19892 25298 19944 25304
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19800 24812 19852 24818
rect 19800 24754 19852 24760
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19076 23662 19104 24142
rect 19317 23964 19625 23973
rect 19317 23962 19323 23964
rect 19379 23962 19403 23964
rect 19459 23962 19483 23964
rect 19539 23962 19563 23964
rect 19619 23962 19625 23964
rect 19379 23910 19381 23962
rect 19561 23910 19563 23962
rect 19317 23908 19323 23910
rect 19379 23908 19403 23910
rect 19459 23908 19483 23910
rect 19539 23908 19563 23910
rect 19619 23908 19625 23910
rect 19317 23899 19625 23908
rect 19720 23730 19748 24142
rect 19708 23724 19760 23730
rect 19708 23666 19760 23672
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 18657 23420 18965 23429
rect 18657 23418 18663 23420
rect 18719 23418 18743 23420
rect 18799 23418 18823 23420
rect 18879 23418 18903 23420
rect 18959 23418 18965 23420
rect 18719 23366 18721 23418
rect 18901 23366 18903 23418
rect 18657 23364 18663 23366
rect 18719 23364 18743 23366
rect 18799 23364 18823 23366
rect 18879 23364 18903 23366
rect 18959 23364 18965 23366
rect 18657 23355 18965 23364
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 19317 22876 19625 22885
rect 19317 22874 19323 22876
rect 19379 22874 19403 22876
rect 19459 22874 19483 22876
rect 19539 22874 19563 22876
rect 19619 22874 19625 22876
rect 19379 22822 19381 22874
rect 19561 22822 19563 22874
rect 19317 22820 19323 22822
rect 19379 22820 19403 22822
rect 19459 22820 19483 22822
rect 19539 22820 19563 22822
rect 19619 22820 19625 22822
rect 19317 22811 19625 22820
rect 18657 22332 18965 22341
rect 18657 22330 18663 22332
rect 18719 22330 18743 22332
rect 18799 22330 18823 22332
rect 18879 22330 18903 22332
rect 18959 22330 18965 22332
rect 18719 22278 18721 22330
rect 18901 22278 18903 22330
rect 18657 22276 18663 22278
rect 18719 22276 18743 22278
rect 18799 22276 18823 22278
rect 18879 22276 18903 22278
rect 18959 22276 18965 22278
rect 18657 22267 18965 22276
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 17682 21927 17738 21936
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17788 21690 17816 21898
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17788 20924 17816 21626
rect 17880 21146 17908 21830
rect 18432 21690 18460 21966
rect 19317 21788 19625 21797
rect 19317 21786 19323 21788
rect 19379 21786 19403 21788
rect 19459 21786 19483 21788
rect 19539 21786 19563 21788
rect 19619 21786 19625 21788
rect 19379 21734 19381 21786
rect 19561 21734 19563 21786
rect 19317 21732 19323 21734
rect 19379 21732 19403 21734
rect 19459 21732 19483 21734
rect 19539 21732 19563 21734
rect 19619 21732 19625 21734
rect 19317 21723 19625 21732
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 17868 20936 17920 20942
rect 17788 20896 17868 20924
rect 17868 20878 17920 20884
rect 18064 20466 18092 20946
rect 18432 20890 18460 21626
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19720 21570 19748 23530
rect 19812 21962 19840 24754
rect 19904 24750 19932 25298
rect 19996 25158 20024 26250
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 25242 20116 25842
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20260 25288 20312 25294
rect 20088 25236 20260 25242
rect 20088 25230 20312 25236
rect 20088 25214 20300 25230
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19996 24750 20024 25094
rect 20088 24818 20116 25214
rect 20168 25152 20220 25158
rect 20168 25094 20220 25100
rect 20180 24886 20208 25094
rect 20168 24880 20220 24886
rect 20168 24822 20220 24828
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19996 24138 20024 24686
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 19984 24132 20036 24138
rect 19984 24074 20036 24080
rect 19996 23594 20024 24074
rect 20088 24070 20116 24550
rect 20180 24206 20208 24822
rect 20732 24818 20760 25638
rect 21192 25226 21220 27338
rect 21652 27334 21680 27950
rect 21914 27911 21970 27920
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21928 25362 21956 27911
rect 22112 27538 22140 28154
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22008 27464 22060 27470
rect 22008 27406 22060 27412
rect 22020 27062 22048 27406
rect 22204 27334 22232 28426
rect 22756 28218 22784 28426
rect 22744 28212 22796 28218
rect 22744 28154 22796 28160
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22296 27470 22324 28018
rect 22652 27940 22704 27946
rect 22652 27882 22704 27888
rect 22468 27872 22520 27878
rect 22468 27814 22520 27820
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22296 27130 22324 27406
rect 22480 27402 22508 27814
rect 22572 27674 22600 27814
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 22664 27606 22692 27882
rect 22848 27606 22876 29106
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23020 28960 23072 28966
rect 23020 28902 23072 28908
rect 23112 28960 23164 28966
rect 23112 28902 23164 28908
rect 22928 28416 22980 28422
rect 22928 28358 22980 28364
rect 22940 28082 22968 28358
rect 23032 28218 23060 28902
rect 23124 28626 23152 28902
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 23400 28218 23428 29038
rect 23952 28994 23980 29718
rect 25228 29640 25280 29646
rect 25228 29582 25280 29588
rect 24492 29096 24544 29102
rect 24492 29038 24544 29044
rect 24504 28994 24532 29038
rect 23952 28966 24532 28994
rect 24216 28688 24268 28694
rect 24216 28630 24268 28636
rect 24228 28422 24256 28630
rect 24320 28558 24348 28966
rect 24308 28552 24360 28558
rect 24308 28494 24360 28500
rect 24216 28416 24268 28422
rect 24216 28358 24268 28364
rect 23020 28212 23072 28218
rect 23020 28154 23072 28160
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 24320 28082 24348 28494
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 24308 28076 24360 28082
rect 24308 28018 24360 28024
rect 22652 27600 22704 27606
rect 22652 27542 22704 27548
rect 22836 27600 22888 27606
rect 22836 27542 22888 27548
rect 22468 27396 22520 27402
rect 22468 27338 22520 27344
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 22008 27056 22060 27062
rect 22008 26998 22060 27004
rect 21916 25356 21968 25362
rect 21916 25298 21968 25304
rect 21180 25220 21232 25226
rect 21180 25162 21232 25168
rect 22284 25220 22336 25226
rect 22284 25162 22336 25168
rect 22296 24886 22324 25162
rect 22284 24880 22336 24886
rect 22284 24822 22336 24828
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19984 23588 20036 23594
rect 19984 23530 20036 23536
rect 19800 21956 19852 21962
rect 19800 21898 19852 21904
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 18524 20992 18552 21490
rect 18880 21480 18932 21486
rect 18932 21440 19104 21468
rect 18880 21422 18932 21428
rect 18657 21244 18965 21253
rect 18657 21242 18663 21244
rect 18719 21242 18743 21244
rect 18799 21242 18823 21244
rect 18879 21242 18903 21244
rect 18959 21242 18965 21244
rect 18719 21190 18721 21242
rect 18901 21190 18903 21242
rect 18657 21188 18663 21190
rect 18719 21188 18743 21190
rect 18799 21188 18823 21190
rect 18879 21188 18903 21190
rect 18959 21188 18965 21190
rect 18657 21179 18965 21188
rect 19076 21146 19104 21440
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19168 21010 19196 21490
rect 19260 21350 19288 21558
rect 19340 21548 19392 21554
rect 19720 21542 19840 21570
rect 19340 21490 19392 21496
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19156 21004 19208 21010
rect 18524 20964 18644 20992
rect 18340 20862 18460 20890
rect 18616 20874 18644 20964
rect 19156 20946 19208 20952
rect 19352 20913 19380 21490
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 21010 19564 21286
rect 19524 21004 19576 21010
rect 19524 20946 19576 20952
rect 19338 20904 19394 20913
rect 18512 20868 18564 20874
rect 18234 20632 18290 20641
rect 18234 20567 18290 20576
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17512 18630 17540 20402
rect 17604 19786 17632 20402
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17788 18970 17816 20402
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 19990 17908 20198
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17972 19281 18000 19450
rect 17958 19272 18014 19281
rect 17958 19207 18014 19216
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17788 18766 17816 18906
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 17338 16712 17478
rect 16776 17338 16804 18090
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 17144 17202 17172 17478
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 16960 16794 16988 17138
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16868 15434 16896 16662
rect 17144 16522 17172 17138
rect 17512 17066 17540 18566
rect 17972 18426 18000 18566
rect 18064 18426 18092 20402
rect 18248 20398 18276 20567
rect 18340 20466 18368 20862
rect 18512 20810 18564 20816
rect 18604 20868 18656 20874
rect 19338 20839 19394 20848
rect 18604 20810 18656 20816
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18248 19922 18276 20334
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18248 19417 18276 19858
rect 18234 19408 18290 19417
rect 18234 19343 18290 19352
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18064 18306 18092 18362
rect 17880 18278 18092 18306
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17604 17338 17632 17546
rect 17880 17542 17908 18278
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18064 17610 18092 18158
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 18340 17202 18368 18090
rect 18432 17542 18460 18838
rect 18524 18222 18552 20810
rect 19156 20800 19208 20806
rect 19156 20742 19208 20748
rect 19062 20496 19118 20505
rect 19062 20431 19064 20440
rect 19116 20431 19118 20440
rect 19064 20402 19116 20408
rect 19168 20330 19196 20742
rect 19317 20700 19625 20709
rect 19317 20698 19323 20700
rect 19379 20698 19403 20700
rect 19459 20698 19483 20700
rect 19539 20698 19563 20700
rect 19619 20698 19625 20700
rect 19379 20646 19381 20698
rect 19561 20646 19563 20698
rect 19317 20644 19323 20646
rect 19379 20644 19403 20646
rect 19459 20644 19483 20646
rect 19539 20644 19563 20646
rect 19619 20644 19625 20646
rect 19317 20635 19625 20644
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 18657 20156 18965 20165
rect 18657 20154 18663 20156
rect 18719 20154 18743 20156
rect 18799 20154 18823 20156
rect 18879 20154 18903 20156
rect 18959 20154 18965 20156
rect 18719 20102 18721 20154
rect 18901 20102 18903 20154
rect 18657 20100 18663 20102
rect 18719 20100 18743 20102
rect 18799 20100 18823 20102
rect 18879 20100 18903 20102
rect 18959 20100 18965 20102
rect 18657 20091 18965 20100
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18892 19281 18920 19314
rect 18878 19272 18934 19281
rect 18878 19207 18934 19216
rect 18657 19068 18965 19077
rect 18657 19066 18663 19068
rect 18719 19066 18743 19068
rect 18799 19066 18823 19068
rect 18879 19066 18903 19068
rect 18959 19066 18965 19068
rect 18719 19014 18721 19066
rect 18901 19014 18903 19066
rect 18657 19012 18663 19014
rect 18719 19012 18743 19014
rect 18799 19012 18823 19014
rect 18879 19012 18903 19014
rect 18959 19012 18965 19014
rect 18657 19003 18965 19012
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 18426 18828 18702
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 19076 18290 19104 19450
rect 19154 19408 19210 19417
rect 19260 19394 19288 19722
rect 19317 19612 19625 19621
rect 19317 19610 19323 19612
rect 19379 19610 19403 19612
rect 19459 19610 19483 19612
rect 19539 19610 19563 19612
rect 19619 19610 19625 19612
rect 19379 19558 19381 19610
rect 19561 19558 19563 19610
rect 19317 19556 19323 19558
rect 19379 19556 19403 19558
rect 19459 19556 19483 19558
rect 19539 19556 19563 19558
rect 19619 19556 19625 19558
rect 19317 19547 19625 19556
rect 19432 19440 19484 19446
rect 19260 19378 19380 19394
rect 19432 19382 19484 19388
rect 19524 19440 19576 19446
rect 19720 19428 19748 19790
rect 19576 19400 19748 19428
rect 19524 19382 19576 19388
rect 19260 19372 19392 19378
rect 19260 19366 19340 19372
rect 19154 19343 19210 19352
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18524 17592 18552 18158
rect 18657 17980 18965 17989
rect 18657 17978 18663 17980
rect 18719 17978 18743 17980
rect 18799 17978 18823 17980
rect 18879 17978 18903 17980
rect 18959 17978 18965 17980
rect 18719 17926 18721 17978
rect 18901 17926 18903 17978
rect 18657 17924 18663 17926
rect 18719 17924 18743 17926
rect 18799 17924 18823 17926
rect 18879 17924 18903 17926
rect 18959 17924 18965 17926
rect 18657 17915 18965 17924
rect 18972 17604 19024 17610
rect 18524 17564 18972 17592
rect 18972 17546 19024 17552
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18328 17196 18380 17202
rect 18432 17184 18460 17478
rect 19076 17338 19104 17478
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19168 17270 19196 19343
rect 19340 19314 19392 19320
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19352 18902 19380 19110
rect 19444 18970 19472 19382
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19432 18760 19484 18766
rect 19536 18748 19564 19382
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19628 18766 19656 19178
rect 19484 18720 19564 18748
rect 19616 18760 19668 18766
rect 19432 18702 19484 18708
rect 19668 18720 19748 18748
rect 19616 18702 19668 18708
rect 19317 18524 19625 18533
rect 19317 18522 19323 18524
rect 19379 18522 19403 18524
rect 19459 18522 19483 18524
rect 19539 18522 19563 18524
rect 19619 18522 19625 18524
rect 19379 18470 19381 18522
rect 19561 18470 19563 18522
rect 19317 18468 19323 18470
rect 19379 18468 19403 18470
rect 19459 18468 19483 18470
rect 19539 18468 19563 18470
rect 19619 18468 19625 18470
rect 19317 18459 19625 18468
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19260 17338 19288 18158
rect 19444 17649 19472 18226
rect 19628 17882 19656 18362
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19522 17776 19578 17785
rect 19522 17711 19578 17720
rect 19536 17678 19564 17711
rect 19720 17678 19748 18720
rect 19812 18426 19840 21542
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19904 19446 19932 19654
rect 19996 19514 20024 19654
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 20088 19446 20116 24006
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 21178 23080 21234 23089
rect 20732 22778 20760 23054
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20824 22642 20852 23054
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20548 22094 20576 22510
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20456 22066 20576 22094
rect 20456 22030 20484 22066
rect 20824 22030 20852 22374
rect 21008 22030 21036 22918
rect 21100 22710 21128 23054
rect 21178 23015 21180 23024
rect 21232 23015 21234 23024
rect 21180 22986 21232 22992
rect 21192 22760 21220 22986
rect 21192 22732 21496 22760
rect 21088 22704 21140 22710
rect 21088 22646 21140 22652
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 21100 22030 21128 22374
rect 21192 22250 21220 22510
rect 21192 22222 21404 22250
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 20456 21894 20484 21966
rect 20352 21888 20404 21894
rect 20350 21856 20352 21865
rect 20444 21888 20496 21894
rect 20404 21856 20406 21865
rect 20444 21830 20496 21836
rect 20350 21791 20406 21800
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20364 21010 20392 21422
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20180 19446 20208 19790
rect 19892 19440 19944 19446
rect 20076 19440 20128 19446
rect 19892 19382 19944 19388
rect 19982 19408 20038 19417
rect 20076 19382 20128 19388
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 19982 19343 20038 19352
rect 19996 19292 20024 19343
rect 19996 19264 20029 19292
rect 20001 19258 20029 19264
rect 20258 19272 20314 19281
rect 20001 19230 20116 19258
rect 20088 18698 20116 19230
rect 20364 19242 20392 20946
rect 20548 20942 20576 21422
rect 20732 21418 20760 21966
rect 20824 21690 20852 21966
rect 21192 21962 21220 22222
rect 21272 22160 21324 22166
rect 21272 22102 21324 22108
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21008 21690 21036 21830
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21008 21146 21036 21286
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20548 19514 20576 20334
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20258 19207 20314 19216
rect 20352 19236 20404 19242
rect 20272 18970 20300 19207
rect 20352 19178 20404 19184
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19904 18426 19932 18566
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19812 17882 19840 18226
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19524 17672 19576 17678
rect 19430 17640 19486 17649
rect 19524 17614 19576 17620
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 19800 17672 19852 17678
rect 19904 17660 19932 18362
rect 20824 18290 20852 19246
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20732 17746 20760 18226
rect 20916 18154 20944 20402
rect 21100 20058 21128 21490
rect 21192 21162 21220 21558
rect 21284 21486 21312 22102
rect 21376 21622 21404 22222
rect 21468 22030 21496 22732
rect 21652 22642 21680 23122
rect 21732 22704 21784 22710
rect 21732 22646 21784 22652
rect 21640 22636 21692 22642
rect 21560 22596 21640 22624
rect 21560 22166 21588 22596
rect 21640 22578 21692 22584
rect 21640 22500 21692 22506
rect 21640 22442 21692 22448
rect 21652 22234 21680 22442
rect 21744 22234 21772 22646
rect 21916 22636 21968 22642
rect 21836 22596 21916 22624
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21732 22228 21784 22234
rect 21732 22170 21784 22176
rect 21548 22160 21600 22166
rect 21548 22102 21600 22108
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21364 21616 21416 21622
rect 21364 21558 21416 21564
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21364 21480 21416 21486
rect 21560 21468 21588 21966
rect 21416 21440 21588 21468
rect 21364 21422 21416 21428
rect 21376 21162 21404 21422
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21192 21134 21404 21162
rect 21192 20466 21220 21134
rect 21376 20942 21404 21134
rect 21468 20942 21496 21286
rect 21744 21078 21772 22170
rect 21836 22030 21864 22596
rect 21916 22578 21968 22584
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22112 22030 22140 22374
rect 22190 22264 22246 22273
rect 22190 22199 22246 22208
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 21822 21584 21878 21593
rect 21822 21519 21878 21528
rect 21916 21548 21968 21554
rect 21836 21418 21864 21519
rect 21916 21490 21968 21496
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21732 21072 21784 21078
rect 21732 21014 21784 21020
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21284 20380 21312 20878
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21560 20534 21588 20810
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 21928 20466 21956 21490
rect 22204 21146 22232 22199
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22190 21040 22246 21049
rect 22190 20975 22246 20984
rect 22204 20942 22232 20975
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21732 20392 21784 20398
rect 21284 20352 21732 20380
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21284 18970 21312 20352
rect 21732 20334 21784 20340
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20076 17740 20128 17746
rect 20352 17740 20404 17746
rect 20128 17700 20208 17728
rect 20076 17682 20128 17688
rect 19852 17632 19932 17660
rect 19800 17614 19852 17620
rect 19430 17575 19486 17584
rect 19812 17490 19840 17614
rect 19720 17462 19840 17490
rect 19317 17436 19625 17445
rect 19317 17434 19323 17436
rect 19379 17434 19403 17436
rect 19459 17434 19483 17436
rect 19539 17434 19563 17436
rect 19619 17434 19625 17436
rect 19379 17382 19381 17434
rect 19561 17382 19563 17434
rect 19317 17380 19323 17382
rect 19379 17380 19403 17382
rect 19459 17380 19483 17382
rect 19539 17380 19563 17382
rect 19619 17380 19625 17382
rect 19317 17371 19625 17380
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 18512 17196 18564 17202
rect 18432 17156 18512 17184
rect 18328 17138 18380 17144
rect 18512 17138 18564 17144
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 18657 16892 18965 16901
rect 18657 16890 18663 16892
rect 18719 16890 18743 16892
rect 18799 16890 18823 16892
rect 18879 16890 18903 16892
rect 18959 16890 18965 16892
rect 18719 16838 18721 16890
rect 18901 16838 18903 16890
rect 18657 16836 18663 16838
rect 18719 16836 18743 16838
rect 18799 16836 18823 16838
rect 18879 16836 18903 16838
rect 18959 16836 18965 16838
rect 18657 16827 18965 16836
rect 19168 16794 19196 17206
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 19317 16348 19625 16357
rect 19317 16346 19323 16348
rect 19379 16346 19403 16348
rect 19459 16346 19483 16348
rect 19539 16346 19563 16348
rect 19619 16346 19625 16348
rect 19379 16294 19381 16346
rect 19561 16294 19563 16346
rect 19317 16292 19323 16294
rect 19379 16292 19403 16294
rect 19459 16292 19483 16294
rect 19539 16292 19563 16294
rect 19619 16292 19625 16294
rect 19317 16283 19625 16292
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 14414 16620 14758
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16764 14272 16816 14278
rect 16684 14232 16764 14260
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16500 12986 16528 13262
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16592 12850 16620 13126
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 11898 16160 12174
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16224 11830 16252 12038
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16212 11688 16264 11694
rect 16040 11636 16212 11642
rect 16040 11630 16264 11636
rect 16040 11614 16252 11630
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15948 10538 15976 11018
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 16040 9625 16068 11086
rect 16224 10674 16252 11614
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16500 10266 16528 11698
rect 16592 11218 16620 12378
rect 16684 12345 16712 14232
rect 16764 14214 16816 14220
rect 17052 13938 17080 16050
rect 17972 15570 18000 16186
rect 18657 15804 18965 15813
rect 18657 15802 18663 15804
rect 18719 15802 18743 15804
rect 18799 15802 18823 15804
rect 18879 15802 18903 15804
rect 18959 15802 18965 15804
rect 18719 15750 18721 15802
rect 18901 15750 18903 15802
rect 18657 15748 18663 15750
rect 18719 15748 18743 15750
rect 18799 15748 18823 15750
rect 18879 15748 18903 15750
rect 18959 15748 18965 15750
rect 18657 15739 18965 15748
rect 19064 15632 19116 15638
rect 19064 15574 19116 15580
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17236 14958 17264 15370
rect 17420 15094 17448 15506
rect 17408 15088 17460 15094
rect 17408 15030 17460 15036
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16670 12336 16726 12345
rect 16776 12306 16804 13194
rect 16868 12850 16896 13738
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16670 12271 16726 12280
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16684 11626 16712 12174
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16500 10062 16528 10202
rect 16592 10130 16620 11154
rect 16868 11082 16896 12786
rect 16960 12238 16988 13466
rect 17052 12850 17080 13874
rect 17144 13326 17172 14826
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16856 11076 16908 11082
rect 16908 11036 16988 11064
rect 16856 11018 16908 11024
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16776 10606 16804 10950
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16026 9616 16082 9625
rect 16026 9551 16082 9560
rect 16040 9450 16068 9551
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8566 15700 8978
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 16408 7886 16436 8842
rect 16592 8498 16620 9454
rect 16776 8634 16804 10542
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16868 9722 16896 9930
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16856 9580 16908 9586
rect 16960 9568 16988 11036
rect 17052 9586 17080 12786
rect 17144 12646 17172 12922
rect 17420 12850 17448 15030
rect 17972 14890 18000 15506
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18156 15366 18184 15438
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18156 15094 18184 15302
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18156 14618 18184 14758
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18156 13802 18184 14554
rect 18524 14550 18552 15370
rect 18657 14716 18965 14725
rect 18657 14714 18663 14716
rect 18719 14714 18743 14716
rect 18799 14714 18823 14716
rect 18879 14714 18903 14716
rect 18959 14714 18965 14716
rect 18719 14662 18721 14714
rect 18901 14662 18903 14714
rect 18657 14660 18663 14662
rect 18719 14660 18743 14662
rect 18799 14660 18823 14662
rect 18879 14660 18903 14662
rect 18959 14660 18965 14662
rect 18657 14651 18965 14660
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18604 14408 18656 14414
rect 18524 14368 18604 14396
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 14074 18368 14214
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18432 13818 18460 14010
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 18248 13790 18460 13818
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17420 12442 17448 12786
rect 17408 12436 17460 12442
rect 17604 12434 17632 13398
rect 18156 13326 18184 13738
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 17604 12406 17724 12434
rect 17408 12378 17460 12384
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17236 9674 17264 12310
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17604 11354 17632 11494
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17328 10266 17356 10610
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17144 9646 17264 9674
rect 16908 9540 16988 9568
rect 17040 9580 17092 9586
rect 16856 9522 16908 9528
rect 17040 9522 17092 9528
rect 16868 8906 16896 9522
rect 17052 9353 17080 9522
rect 17038 9344 17094 9353
rect 17038 9279 17094 9288
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 15488 6730 15516 7822
rect 16592 7002 16620 8298
rect 16776 7886 16804 8570
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7546 16804 7686
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 17052 7410 17080 8230
rect 17144 7546 17172 9646
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17328 8022 17356 9046
rect 17420 8072 17448 10406
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17512 8498 17540 9114
rect 17604 8634 17632 9318
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17420 8044 17632 8072
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17406 7984 17462 7993
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 7002 16804 7142
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15488 6390 15516 6666
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 16040 4690 16068 5578
rect 16486 5400 16542 5409
rect 16486 5335 16488 5344
rect 16540 5335 16542 5344
rect 16488 5306 16540 5312
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16132 4758 16160 5170
rect 16210 5128 16266 5137
rect 16210 5063 16266 5072
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16224 4554 16252 5063
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16408 4729 16436 4762
rect 16394 4720 16450 4729
rect 16394 4655 16450 4664
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16408 4282 16436 4655
rect 16500 4622 16528 4762
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 16500 3942 16528 4558
rect 16592 4536 16620 6394
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16868 5030 16896 6326
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16672 4548 16724 4554
rect 16592 4508 16672 4536
rect 16592 4146 16620 4508
rect 16672 4490 16724 4496
rect 16868 4486 16896 4966
rect 16960 4826 16988 5850
rect 17052 5234 17080 7346
rect 17144 6798 17172 7482
rect 17236 7449 17264 7754
rect 17222 7440 17278 7449
rect 17222 7375 17278 7384
rect 17328 7392 17356 7958
rect 17406 7919 17462 7928
rect 17420 7886 17448 7919
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17500 7744 17552 7750
rect 17406 7712 17462 7721
rect 17500 7686 17552 7692
rect 17406 7647 17462 7656
rect 17420 7546 17448 7647
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17512 7410 17540 7686
rect 17408 7404 17460 7410
rect 17236 6798 17264 7375
rect 17328 7364 17408 7392
rect 17408 7346 17460 7352
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 6798 17448 7142
rect 17604 6934 17632 8044
rect 17696 7546 17724 12406
rect 17972 11778 18000 13262
rect 18248 12209 18276 13790
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18432 12986 18460 13670
rect 18524 13530 18552 14368
rect 18604 14350 18656 14356
rect 18708 13938 18736 14486
rect 19076 14482 19104 15574
rect 19317 15260 19625 15269
rect 19317 15258 19323 15260
rect 19379 15258 19403 15260
rect 19459 15258 19483 15260
rect 19539 15258 19563 15260
rect 19619 15258 19625 15260
rect 19379 15206 19381 15258
rect 19561 15206 19563 15258
rect 19317 15204 19323 15206
rect 19379 15204 19403 15206
rect 19459 15204 19483 15206
rect 19539 15204 19563 15206
rect 19619 15204 19625 15206
rect 19317 15195 19625 15204
rect 19616 15020 19668 15026
rect 19720 15008 19748 17462
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19812 15026 19840 15438
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19996 15162 20024 15302
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19668 14980 19748 15008
rect 19800 15020 19852 15026
rect 19616 14962 19668 14968
rect 19800 14962 19852 14968
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19260 14618 19288 14758
rect 19248 14612 19300 14618
rect 19168 14572 19248 14600
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 19062 14376 19118 14385
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18892 13734 18920 14350
rect 19062 14311 19118 14320
rect 19076 14074 19104 14311
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19168 14006 19196 14572
rect 19248 14554 19300 14560
rect 19628 14414 19656 14962
rect 19812 14414 19840 14962
rect 20088 14482 20116 15302
rect 20180 15094 20208 17700
rect 20352 17682 20404 17688
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20364 17338 20392 17682
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20180 14618 20208 14894
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20536 14408 20588 14414
rect 20588 14356 20668 14362
rect 20536 14350 20668 14356
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19616 14272 19668 14278
rect 19892 14272 19944 14278
rect 19668 14232 19840 14260
rect 19616 14214 19668 14220
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18657 13628 18965 13637
rect 18657 13626 18663 13628
rect 18719 13626 18743 13628
rect 18799 13626 18823 13628
rect 18879 13626 18903 13628
rect 18959 13626 18965 13628
rect 18719 13574 18721 13626
rect 18901 13574 18903 13626
rect 18657 13572 18663 13574
rect 18719 13572 18743 13574
rect 18799 13572 18823 13574
rect 18879 13572 18903 13574
rect 18959 13572 18965 13574
rect 18657 13563 18965 13572
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 19260 13326 19288 14214
rect 19317 14172 19625 14181
rect 19317 14170 19323 14172
rect 19379 14170 19403 14172
rect 19459 14170 19483 14172
rect 19539 14170 19563 14172
rect 19619 14170 19625 14172
rect 19379 14118 19381 14170
rect 19561 14118 19563 14170
rect 19317 14116 19323 14118
rect 19379 14116 19403 14118
rect 19459 14116 19483 14118
rect 19539 14116 19563 14118
rect 19619 14116 19625 14118
rect 19317 14107 19625 14116
rect 19706 14104 19762 14113
rect 19706 14039 19762 14048
rect 19720 14006 19748 14039
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19536 13530 19564 13874
rect 19812 13802 19840 14232
rect 19892 14214 19944 14220
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19904 13682 19932 14214
rect 19996 14074 20024 14282
rect 20180 14113 20208 14350
rect 20548 14334 20668 14350
rect 20166 14104 20222 14113
rect 19984 14068 20036 14074
rect 20640 14074 20668 14334
rect 20166 14039 20222 14048
rect 20628 14068 20680 14074
rect 19984 14010 20036 14016
rect 20628 14010 20680 14016
rect 20076 13932 20128 13938
rect 20128 13892 20208 13920
rect 20076 13874 20128 13880
rect 19720 13654 19932 13682
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19317 13084 19625 13093
rect 19317 13082 19323 13084
rect 19379 13082 19403 13084
rect 19459 13082 19483 13084
rect 19539 13082 19563 13084
rect 19619 13082 19625 13084
rect 19379 13030 19381 13082
rect 19561 13030 19563 13082
rect 19317 13028 19323 13030
rect 19379 13028 19403 13030
rect 19459 13028 19483 13030
rect 19539 13028 19563 13030
rect 19619 13028 19625 13030
rect 19317 13019 19625 13028
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 19062 12744 19118 12753
rect 19062 12679 19118 12688
rect 19076 12646 19104 12679
rect 19064 12640 19116 12646
rect 19116 12600 19196 12628
rect 19064 12582 19116 12588
rect 18657 12540 18965 12549
rect 18657 12538 18663 12540
rect 18719 12538 18743 12540
rect 18799 12538 18823 12540
rect 18879 12538 18903 12540
rect 18959 12538 18965 12540
rect 18719 12486 18721 12538
rect 18901 12486 18903 12538
rect 18657 12484 18663 12486
rect 18719 12484 18743 12486
rect 18799 12484 18823 12486
rect 18879 12484 18903 12486
rect 18959 12484 18965 12486
rect 18657 12475 18965 12484
rect 18234 12200 18290 12209
rect 18234 12135 18290 12144
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 17972 11750 18460 11778
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18064 11354 18092 11630
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18064 10674 18092 11290
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17788 9625 17816 10610
rect 17880 10198 17908 10610
rect 18156 10266 18184 11086
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 17774 9616 17830 9625
rect 17774 9551 17830 9560
rect 17788 8498 17816 9551
rect 17880 9450 17908 10134
rect 18156 10062 18184 10202
rect 18248 10130 18276 11086
rect 18432 10606 18460 11750
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18524 10810 18552 11698
rect 18657 11452 18965 11461
rect 18657 11450 18663 11452
rect 18719 11450 18743 11452
rect 18799 11450 18823 11452
rect 18879 11450 18903 11452
rect 18959 11450 18965 11452
rect 18719 11398 18721 11450
rect 18901 11398 18903 11450
rect 18657 11396 18663 11398
rect 18719 11396 18743 11398
rect 18799 11396 18823 11398
rect 18879 11396 18903 11398
rect 18959 11396 18965 11398
rect 18657 11387 18965 11396
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18340 9926 18368 9998
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18340 9586 18368 9862
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18236 9512 18288 9518
rect 18432 9489 18460 10542
rect 18524 9722 18552 10746
rect 18708 10713 18736 11086
rect 18694 10704 18750 10713
rect 18694 10639 18750 10648
rect 18892 10577 18920 11222
rect 19076 11218 19104 11834
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 18970 10840 19026 10849
rect 18970 10775 19026 10784
rect 18984 10674 19012 10775
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 18878 10568 18934 10577
rect 18878 10503 18934 10512
rect 18657 10364 18965 10373
rect 18657 10362 18663 10364
rect 18719 10362 18743 10364
rect 18799 10362 18823 10364
rect 18879 10362 18903 10364
rect 18959 10362 18965 10364
rect 18719 10310 18721 10362
rect 18901 10310 18903 10362
rect 18657 10308 18663 10310
rect 18719 10308 18743 10310
rect 18799 10308 18823 10310
rect 18879 10308 18903 10310
rect 18959 10308 18965 10310
rect 18657 10299 18965 10308
rect 19076 10130 19104 10610
rect 19168 10266 19196 12600
rect 19317 11996 19625 12005
rect 19317 11994 19323 11996
rect 19379 11994 19403 11996
rect 19459 11994 19483 11996
rect 19539 11994 19563 11996
rect 19619 11994 19625 11996
rect 19379 11942 19381 11994
rect 19561 11942 19563 11994
rect 19317 11940 19323 11942
rect 19379 11940 19403 11942
rect 19459 11940 19483 11942
rect 19539 11940 19563 11942
rect 19619 11940 19625 11942
rect 19317 11931 19625 11940
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19352 11286 19380 11630
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18984 9625 19012 9658
rect 18970 9616 19026 9625
rect 19076 9586 19104 9862
rect 18970 9551 19026 9560
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 18418 9480 18474 9489
rect 18288 9460 18418 9466
rect 18236 9454 18418 9460
rect 17868 9444 17920 9450
rect 18248 9438 18418 9454
rect 18418 9415 18474 9424
rect 17868 9386 17920 9392
rect 18432 9382 18460 9415
rect 17960 9376 18012 9382
rect 18420 9376 18472 9382
rect 17960 9318 18012 9324
rect 18326 9344 18382 9353
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17788 8022 17816 8434
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17592 6928 17644 6934
rect 17512 6888 17592 6916
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16868 4282 16896 4422
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16960 4214 16988 4762
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 15672 3670 15700 3878
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15120 3194 15148 3606
rect 16592 3602 16620 4082
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15304 3398 15332 3470
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15304 3126 15332 3334
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 17052 3058 17080 5170
rect 17144 5030 17172 6598
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17236 5370 17264 5782
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17144 4146 17172 4422
rect 17236 4146 17264 4422
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17328 4010 17356 5306
rect 17420 5234 17448 5714
rect 17512 5710 17540 6888
rect 17592 6870 17644 6876
rect 17696 6798 17724 7482
rect 17788 7478 17816 7958
rect 17972 7886 18000 9318
rect 18420 9318 18472 9324
rect 18326 9279 18382 9288
rect 18340 9110 18368 9279
rect 18657 9276 18965 9285
rect 18657 9274 18663 9276
rect 18719 9274 18743 9276
rect 18799 9274 18823 9276
rect 18879 9274 18903 9276
rect 18959 9274 18965 9276
rect 18719 9222 18721 9274
rect 18901 9222 18903 9274
rect 18657 9220 18663 9222
rect 18719 9220 18743 9222
rect 18799 9220 18823 9222
rect 18879 9220 18903 9222
rect 18959 9220 18965 9222
rect 18657 9211 18965 9220
rect 18328 9104 18380 9110
rect 18328 9046 18380 9052
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18064 8838 18092 8910
rect 18156 8888 18184 8978
rect 18236 8900 18288 8906
rect 18156 8860 18236 8888
rect 18236 8842 18288 8848
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18524 8634 18552 8774
rect 19168 8634 19196 10202
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19260 8566 19288 11086
rect 19720 11082 19748 13654
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19812 12220 19840 13126
rect 19996 12434 20024 13262
rect 19996 12406 20116 12434
rect 19984 12232 20036 12238
rect 19812 12192 19984 12220
rect 19984 12174 20036 12180
rect 19800 12096 19852 12102
rect 20088 12050 20116 12406
rect 19800 12038 19852 12044
rect 19812 11354 19840 12038
rect 19996 12022 20116 12050
rect 19996 11694 20024 12022
rect 20180 11898 20208 13892
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20272 13326 20300 13806
rect 20640 13530 20668 14010
rect 20732 13938 20760 14758
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20916 14385 20944 14554
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 20902 14376 20958 14385
rect 20902 14311 20958 14320
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 11898 20300 13262
rect 20732 12918 20760 13874
rect 20996 13864 21048 13870
rect 21100 13852 21128 14418
rect 21048 13824 21128 13852
rect 20996 13806 21048 13812
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 21100 12850 21128 13824
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21192 12782 21220 14962
rect 21284 13376 21312 18226
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 22020 17270 22048 17682
rect 22296 17678 22324 24822
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22572 22234 22600 22986
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22572 22098 22600 22170
rect 22560 22092 22612 22098
rect 22560 22034 22612 22040
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22480 21554 22508 21830
rect 22664 21690 22692 22510
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22756 22030 22784 22374
rect 22848 22030 22876 22714
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 23112 22636 23164 22642
rect 23112 22578 23164 22584
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22836 22024 22888 22030
rect 23032 22012 23060 22578
rect 23124 22273 23152 22578
rect 23216 22438 23244 22578
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 23110 22264 23166 22273
rect 23110 22199 23166 22208
rect 23216 22030 23244 22374
rect 23112 22024 23164 22030
rect 23032 21984 23112 22012
rect 22836 21966 22888 21972
rect 23112 21966 23164 21972
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22756 21554 22784 21966
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22572 20602 22600 21422
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 22664 20942 22692 21286
rect 22848 21078 22876 21966
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 22836 21072 22888 21078
rect 22940 21049 22968 21422
rect 22836 21014 22888 21020
rect 22926 21040 22982 21049
rect 22926 20975 22982 20984
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22664 20602 22692 20878
rect 22560 20596 22612 20602
rect 22560 20538 22612 20544
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22756 20466 22784 20878
rect 23124 20602 23152 21558
rect 23216 21418 23244 21966
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23308 20806 23336 22578
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23400 21554 23428 22374
rect 23492 21894 23520 22510
rect 23768 22030 23796 23054
rect 23848 22976 23900 22982
rect 23848 22918 23900 22924
rect 23860 22642 23888 22918
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 24044 22506 24072 22578
rect 24032 22500 24084 22506
rect 24032 22442 24084 22448
rect 23938 22400 23994 22409
rect 23938 22335 23994 22344
rect 23952 22166 23980 22335
rect 23940 22160 23992 22166
rect 23940 22102 23992 22108
rect 23756 22024 23808 22030
rect 23676 21984 23756 22012
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21690 23520 21830
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23572 21684 23624 21690
rect 23676 21672 23704 21984
rect 23756 21966 23808 21972
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23624 21644 23704 21672
rect 23572 21626 23624 21632
rect 23756 21616 23808 21622
rect 23754 21584 23756 21593
rect 23808 21584 23810 21593
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23572 21548 23624 21554
rect 23754 21519 23810 21528
rect 23572 21490 23624 21496
rect 23584 21146 23612 21490
rect 23952 21350 23980 21966
rect 24044 21554 24072 22442
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23676 20466 23704 21286
rect 23848 20800 23900 20806
rect 23848 20742 23900 20748
rect 23860 20466 23888 20742
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23940 20460 23992 20466
rect 24136 20448 24164 21966
rect 24216 20868 24268 20874
rect 24216 20810 24268 20816
rect 24228 20466 24256 20810
rect 23992 20420 24164 20448
rect 24216 20460 24268 20466
rect 23940 20402 23992 20408
rect 24216 20402 24268 20408
rect 23676 20330 23704 20402
rect 23664 20324 23716 20330
rect 23664 20266 23716 20272
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22664 18086 22692 19382
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22664 17678 22692 18022
rect 23216 17882 23244 18158
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 22744 17808 22796 17814
rect 22744 17750 22796 17756
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22008 17264 22060 17270
rect 22008 17206 22060 17212
rect 22296 17218 22324 17614
rect 22020 16658 22048 17206
rect 22192 17196 22244 17202
rect 22296 17190 22416 17218
rect 22192 17138 22244 17144
rect 22204 16794 22232 17138
rect 22388 17134 22416 17190
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22296 16794 22324 17002
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22296 15570 22324 16526
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21560 14414 21588 14894
rect 22296 14414 22324 15506
rect 22388 15026 22416 17070
rect 22664 16794 22692 17614
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22756 16590 22784 17750
rect 23308 17678 23336 18702
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22848 16794 22876 17138
rect 23124 16998 23152 17478
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 22848 16250 22876 16730
rect 23216 16538 23244 17070
rect 23308 16726 23336 17614
rect 23492 17134 23520 18294
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 23584 17338 23612 17546
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23400 16590 23428 16730
rect 23388 16584 23440 16590
rect 23216 16510 23336 16538
rect 23388 16526 23440 16532
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 23216 16182 23244 16390
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23216 15502 23244 16118
rect 23308 15978 23336 16510
rect 23296 15972 23348 15978
rect 23296 15914 23348 15920
rect 23296 15632 23348 15638
rect 23296 15574 23348 15580
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 23204 15020 23256 15026
rect 23308 15008 23336 15574
rect 23256 14980 23336 15008
rect 23388 15020 23440 15026
rect 23204 14962 23256 14968
rect 23388 14962 23440 14968
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 21456 14000 21508 14006
rect 21560 13988 21588 14350
rect 21508 13960 21588 13988
rect 21456 13942 21508 13948
rect 21364 13796 21416 13802
rect 21364 13738 21416 13744
rect 21376 13530 21404 13738
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21456 13388 21508 13394
rect 21284 13348 21456 13376
rect 21456 13330 21508 13336
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19317 10908 19625 10917
rect 19317 10906 19323 10908
rect 19379 10906 19403 10908
rect 19459 10906 19483 10908
rect 19539 10906 19563 10908
rect 19619 10906 19625 10908
rect 19379 10854 19381 10906
rect 19561 10854 19563 10906
rect 19317 10852 19323 10854
rect 19379 10852 19403 10854
rect 19459 10852 19483 10854
rect 19539 10852 19563 10854
rect 19619 10852 19625 10854
rect 19317 10843 19625 10852
rect 20088 10742 20116 11698
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 19812 10305 19840 10678
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19798 10296 19854 10305
rect 19798 10231 19854 10240
rect 19904 10062 19932 10406
rect 20088 10062 20116 10678
rect 20272 10266 20300 11834
rect 20548 11762 20576 12718
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20364 10810 20392 11018
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20456 10606 20484 11698
rect 20548 10674 20576 11698
rect 21192 11014 21220 12718
rect 21180 11008 21232 11014
rect 21180 10950 21232 10956
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20456 10130 20484 10542
rect 20548 10538 20576 10610
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20536 10532 20588 10538
rect 20536 10474 20588 10480
rect 20916 10198 20944 10542
rect 20904 10192 20956 10198
rect 20904 10134 20956 10140
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19317 9820 19625 9829
rect 19317 9818 19323 9820
rect 19379 9818 19403 9820
rect 19459 9818 19483 9820
rect 19539 9818 19563 9820
rect 19619 9818 19625 9820
rect 19379 9766 19381 9818
rect 19561 9766 19563 9818
rect 19317 9764 19323 9766
rect 19379 9764 19403 9766
rect 19459 9764 19483 9766
rect 19539 9764 19563 9766
rect 19619 9764 19625 9766
rect 19317 9755 19625 9764
rect 21468 9722 21496 13330
rect 21652 12986 21680 14350
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 21732 14000 21784 14006
rect 21732 13942 21784 13948
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21652 12646 21680 12922
rect 21744 12782 21772 13942
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21836 12850 21864 13126
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 22112 11354 22140 14214
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22204 13394 22232 13806
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22296 12986 22324 14350
rect 22388 14074 22416 14350
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22664 13394 22692 14350
rect 22848 13462 22876 14350
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22204 12238 22232 12718
rect 22652 12708 22704 12714
rect 22652 12650 22704 12656
rect 22664 12238 22692 12650
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22204 11762 22232 12174
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 22296 11898 22324 12106
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22100 11144 22152 11150
rect 22020 11104 22100 11132
rect 22020 10674 22048 11104
rect 22100 11086 22152 11092
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22204 10606 22232 11698
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22296 10282 22324 11834
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22468 11620 22520 11626
rect 22468 11562 22520 11568
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22388 11150 22416 11494
rect 22480 11286 22508 11562
rect 22664 11558 22692 11698
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22468 11280 22520 11286
rect 22468 11222 22520 11228
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22388 10470 22416 11086
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22480 10674 22508 11018
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22296 10254 22508 10282
rect 22664 10266 22692 11290
rect 22756 11218 22784 12718
rect 22940 12374 22968 12854
rect 22928 12368 22980 12374
rect 22848 12328 22928 12356
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22756 10674 22784 11154
rect 22848 10690 22876 12328
rect 22928 12310 22980 12316
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22940 11150 22968 11698
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 23032 10810 23060 12106
rect 23124 11898 23152 12174
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23112 11076 23164 11082
rect 23112 11018 23164 11024
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 22744 10668 22796 10674
rect 22848 10662 23060 10690
rect 22744 10610 22796 10616
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 8974 19380 9318
rect 22204 9042 22232 9930
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22284 9036 22336 9042
rect 22284 8978 22336 8984
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 19317 8732 19625 8741
rect 19317 8730 19323 8732
rect 19379 8730 19403 8732
rect 19459 8730 19483 8732
rect 19539 8730 19563 8732
rect 19619 8730 19625 8732
rect 19379 8678 19381 8730
rect 19561 8678 19563 8730
rect 19317 8676 19323 8678
rect 19379 8676 19403 8678
rect 19459 8676 19483 8678
rect 19539 8676 19563 8678
rect 19619 8676 19625 8678
rect 19317 8667 19625 8676
rect 20640 8634 20668 8774
rect 21744 8634 21772 8774
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 18657 8188 18965 8197
rect 18657 8186 18663 8188
rect 18719 8186 18743 8188
rect 18799 8186 18823 8188
rect 18879 8186 18903 8188
rect 18959 8186 18965 8188
rect 18719 8134 18721 8186
rect 18901 8134 18903 8186
rect 18657 8132 18663 8134
rect 18719 8132 18743 8134
rect 18799 8132 18823 8134
rect 18879 8132 18903 8134
rect 18959 8132 18965 8134
rect 18657 8123 18965 8132
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18064 7886 18092 8026
rect 20916 7954 20944 8230
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 17972 7721 18000 7822
rect 18420 7744 18472 7750
rect 17958 7712 18014 7721
rect 18420 7686 18472 7692
rect 17958 7647 18014 7656
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17866 7440 17922 7449
rect 18064 7410 18092 7482
rect 18432 7410 18460 7686
rect 19317 7644 19625 7653
rect 19317 7642 19323 7644
rect 19379 7642 19403 7644
rect 19459 7642 19483 7644
rect 19539 7642 19563 7644
rect 19619 7642 19625 7644
rect 19379 7590 19381 7642
rect 19561 7590 19563 7642
rect 19317 7588 19323 7590
rect 19379 7588 19403 7590
rect 19459 7588 19483 7590
rect 19539 7588 19563 7590
rect 19619 7588 19625 7590
rect 19317 7579 19625 7588
rect 17866 7375 17868 7384
rect 17920 7375 17922 7384
rect 18052 7404 18104 7410
rect 17868 7346 17920 7352
rect 18052 7346 18104 7352
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17788 6798 17816 6938
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17604 6202 17632 6734
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6458 17816 6598
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17880 6390 17908 7142
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6458 18000 6598
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17604 6174 17724 6202
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17408 5092 17460 5098
rect 17460 5052 17540 5080
rect 17408 5034 17460 5040
rect 17512 4690 17540 5052
rect 17604 4826 17632 6054
rect 17696 5234 17724 6174
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17696 4672 17724 5170
rect 17788 5001 17816 5578
rect 17880 5234 17908 6326
rect 18432 5710 18460 7346
rect 18524 5778 18552 7346
rect 18657 7100 18965 7109
rect 18657 7098 18663 7100
rect 18719 7098 18743 7100
rect 18799 7098 18823 7100
rect 18879 7098 18903 7100
rect 18959 7098 18965 7100
rect 18719 7046 18721 7098
rect 18901 7046 18903 7098
rect 18657 7044 18663 7046
rect 18719 7044 18743 7046
rect 18799 7044 18823 7046
rect 18879 7044 18903 7046
rect 18959 7044 18965 7046
rect 18657 7035 18965 7044
rect 20088 6866 20116 7822
rect 21916 7812 21968 7818
rect 21916 7754 21968 7760
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 21928 6798 21956 7754
rect 22020 7274 22048 7822
rect 22112 7750 22140 8774
rect 22204 8090 22232 8978
rect 22296 8090 22324 8978
rect 22388 8974 22416 9862
rect 22480 9042 22508 10254
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22572 8906 22600 9522
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22204 7970 22232 8026
rect 22204 7942 22324 7970
rect 22480 7954 22508 8230
rect 22296 7886 22324 7942
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22572 7886 22600 8434
rect 22664 7993 22692 8774
rect 22650 7984 22706 7993
rect 22650 7919 22706 7928
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22296 7410 22324 7822
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 22204 6934 22232 7278
rect 22388 7002 22416 7686
rect 22480 7528 22508 7686
rect 22560 7540 22612 7546
rect 22480 7500 22560 7528
rect 22560 7482 22612 7488
rect 22376 6996 22428 7002
rect 22376 6938 22428 6944
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 22756 6866 22784 10610
rect 22926 10296 22982 10305
rect 22926 10231 22928 10240
rect 22980 10231 22982 10240
rect 22928 10202 22980 10208
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 22836 9988 22888 9994
rect 22836 9930 22888 9936
rect 22848 9178 22876 9930
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22940 8498 22968 9998
rect 23032 8634 23060 10662
rect 23124 10033 23152 11018
rect 23216 10130 23244 14962
rect 23400 14618 23428 14962
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23308 11694 23336 13262
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 23400 10266 23428 14010
rect 23492 13938 23520 17070
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23584 15706 23612 16934
rect 23768 16810 23796 17682
rect 24032 17604 24084 17610
rect 24032 17546 24084 17552
rect 23768 16794 23888 16810
rect 23768 16788 23900 16794
rect 23768 16782 23848 16788
rect 23848 16730 23900 16736
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23584 14618 23612 15642
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23676 14414 23704 15914
rect 23768 15570 23796 16458
rect 23952 16114 23980 16526
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23952 15502 23980 16050
rect 24044 15706 24072 17546
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 24044 15570 24072 15642
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23848 14884 23900 14890
rect 23848 14826 23900 14832
rect 23860 14482 23888 14826
rect 23952 14532 23980 15438
rect 24044 15094 24072 15506
rect 24032 15088 24084 15094
rect 24032 15030 24084 15036
rect 23952 14504 24072 14532
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23860 14090 23888 14418
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23676 14062 23888 14090
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23492 12238 23520 12582
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23584 11082 23612 13942
rect 23676 11082 23704 14062
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 12102 23796 13126
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23768 11694 23796 12038
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 23860 10810 23888 12038
rect 23952 11642 23980 14214
rect 24044 13190 24072 14504
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24136 12434 24164 20198
rect 24320 19334 24348 28018
rect 24412 27470 24440 28358
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 25240 23322 25268 29582
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24400 22976 24452 22982
rect 24400 22918 24452 22924
rect 24412 22642 24440 22918
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24400 22500 24452 22506
rect 24400 22442 24452 22448
rect 24412 22409 24440 22442
rect 24398 22400 24454 22409
rect 24398 22335 24454 22344
rect 24504 22030 24532 23054
rect 24688 22522 24716 23054
rect 24768 22976 24820 22982
rect 24768 22918 24820 22924
rect 24780 22681 24808 22918
rect 25332 22778 25360 30194
rect 28540 30048 28592 30054
rect 28540 29990 28592 29996
rect 25740 29948 26048 29957
rect 25740 29946 25746 29948
rect 25802 29946 25826 29948
rect 25882 29946 25906 29948
rect 25962 29946 25986 29948
rect 26042 29946 26048 29948
rect 25802 29894 25804 29946
rect 25984 29894 25986 29946
rect 25740 29892 25746 29894
rect 25802 29892 25826 29894
rect 25882 29892 25906 29894
rect 25962 29892 25986 29894
rect 26042 29892 26048 29894
rect 25740 29883 26048 29892
rect 26400 29404 26708 29413
rect 26400 29402 26406 29404
rect 26462 29402 26486 29404
rect 26542 29402 26566 29404
rect 26622 29402 26646 29404
rect 26702 29402 26708 29404
rect 26462 29350 26464 29402
rect 26644 29350 26646 29402
rect 26400 29348 26406 29350
rect 26462 29348 26486 29350
rect 26542 29348 26566 29350
rect 26622 29348 26646 29350
rect 26702 29348 26708 29350
rect 26400 29339 26708 29348
rect 28552 29306 28580 29990
rect 28540 29300 28592 29306
rect 28540 29242 28592 29248
rect 28736 29073 28764 30194
rect 28920 30190 28948 30631
rect 29012 30326 29040 31925
rect 29000 30320 29052 30326
rect 29000 30262 29052 30268
rect 28908 30184 28960 30190
rect 28908 30126 28960 30132
rect 28722 29064 28778 29073
rect 28722 28999 28778 29008
rect 25740 28860 26048 28869
rect 25740 28858 25746 28860
rect 25802 28858 25826 28860
rect 25882 28858 25906 28860
rect 25962 28858 25986 28860
rect 26042 28858 26048 28860
rect 25802 28806 25804 28858
rect 25984 28806 25986 28858
rect 25740 28804 25746 28806
rect 25802 28804 25826 28806
rect 25882 28804 25906 28806
rect 25962 28804 25986 28806
rect 26042 28804 26048 28806
rect 25740 28795 26048 28804
rect 26400 28316 26708 28325
rect 26400 28314 26406 28316
rect 26462 28314 26486 28316
rect 26542 28314 26566 28316
rect 26622 28314 26646 28316
rect 26702 28314 26708 28316
rect 26462 28262 26464 28314
rect 26644 28262 26646 28314
rect 26400 28260 26406 28262
rect 26462 28260 26486 28262
rect 26542 28260 26566 28262
rect 26622 28260 26646 28262
rect 26702 28260 26708 28262
rect 26400 28251 26708 28260
rect 25740 27772 26048 27781
rect 25740 27770 25746 27772
rect 25802 27770 25826 27772
rect 25882 27770 25906 27772
rect 25962 27770 25986 27772
rect 26042 27770 26048 27772
rect 25802 27718 25804 27770
rect 25984 27718 25986 27770
rect 25740 27716 25746 27718
rect 25802 27716 25826 27718
rect 25882 27716 25906 27718
rect 25962 27716 25986 27718
rect 26042 27716 26048 27718
rect 25740 27707 26048 27716
rect 26400 27228 26708 27237
rect 26400 27226 26406 27228
rect 26462 27226 26486 27228
rect 26542 27226 26566 27228
rect 26622 27226 26646 27228
rect 26702 27226 26708 27228
rect 26462 27174 26464 27226
rect 26644 27174 26646 27226
rect 26400 27172 26406 27174
rect 26462 27172 26486 27174
rect 26542 27172 26566 27174
rect 26622 27172 26646 27174
rect 26702 27172 26708 27174
rect 26400 27163 26708 27172
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 25740 26684 26048 26693
rect 25740 26682 25746 26684
rect 25802 26682 25826 26684
rect 25882 26682 25906 26684
rect 25962 26682 25986 26684
rect 26042 26682 26048 26684
rect 25802 26630 25804 26682
rect 25984 26630 25986 26682
rect 25740 26628 25746 26630
rect 25802 26628 25826 26630
rect 25882 26628 25906 26630
rect 25962 26628 25986 26630
rect 26042 26628 26048 26630
rect 25740 26619 26048 26628
rect 26400 26140 26708 26149
rect 26400 26138 26406 26140
rect 26462 26138 26486 26140
rect 26542 26138 26566 26140
rect 26622 26138 26646 26140
rect 26702 26138 26708 26140
rect 26462 26086 26464 26138
rect 26644 26086 26646 26138
rect 26400 26084 26406 26086
rect 26462 26084 26486 26086
rect 26542 26084 26566 26086
rect 26622 26084 26646 26086
rect 26702 26084 26708 26086
rect 26400 26075 26708 26084
rect 25740 25596 26048 25605
rect 25740 25594 25746 25596
rect 25802 25594 25826 25596
rect 25882 25594 25906 25596
rect 25962 25594 25986 25596
rect 26042 25594 26048 25596
rect 25802 25542 25804 25594
rect 25984 25542 25986 25594
rect 25740 25540 25746 25542
rect 25802 25540 25826 25542
rect 25882 25540 25906 25542
rect 25962 25540 25986 25542
rect 26042 25540 26048 25542
rect 25740 25531 26048 25540
rect 26400 25052 26708 25061
rect 26400 25050 26406 25052
rect 26462 25050 26486 25052
rect 26542 25050 26566 25052
rect 26622 25050 26646 25052
rect 26702 25050 26708 25052
rect 26462 24998 26464 25050
rect 26644 24998 26646 25050
rect 26400 24996 26406 24998
rect 26462 24996 26486 24998
rect 26542 24996 26566 24998
rect 26622 24996 26646 24998
rect 26702 24996 26708 24998
rect 26400 24987 26708 24996
rect 25740 24508 26048 24517
rect 25740 24506 25746 24508
rect 25802 24506 25826 24508
rect 25882 24506 25906 24508
rect 25962 24506 25986 24508
rect 26042 24506 26048 24508
rect 25802 24454 25804 24506
rect 25984 24454 25986 24506
rect 25740 24452 25746 24454
rect 25802 24452 25826 24454
rect 25882 24452 25906 24454
rect 25962 24452 25986 24454
rect 26042 24452 26048 24454
rect 25740 24443 26048 24452
rect 26400 23964 26708 23973
rect 26400 23962 26406 23964
rect 26462 23962 26486 23964
rect 26542 23962 26566 23964
rect 26622 23962 26646 23964
rect 26702 23962 26708 23964
rect 26462 23910 26464 23962
rect 26644 23910 26646 23962
rect 26400 23908 26406 23910
rect 26462 23908 26486 23910
rect 26542 23908 26566 23910
rect 26622 23908 26646 23910
rect 26702 23908 26708 23910
rect 26400 23899 26708 23908
rect 25740 23420 26048 23429
rect 25740 23418 25746 23420
rect 25802 23418 25826 23420
rect 25882 23418 25906 23420
rect 25962 23418 25986 23420
rect 26042 23418 26048 23420
rect 25802 23366 25804 23418
rect 25984 23366 25986 23418
rect 25740 23364 25746 23366
rect 25802 23364 25826 23366
rect 25882 23364 25906 23366
rect 25962 23364 25986 23366
rect 26042 23364 26048 23366
rect 25740 23355 26048 23364
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25412 22976 25464 22982
rect 25412 22918 25464 22924
rect 25424 22778 25452 22918
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 24766 22672 24822 22681
rect 24766 22607 24768 22616
rect 24820 22607 24822 22616
rect 25044 22636 25096 22642
rect 24768 22578 24820 22584
rect 25044 22578 25096 22584
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 24952 22568 25004 22574
rect 24584 22500 24636 22506
rect 24688 22494 24808 22522
rect 24952 22510 25004 22516
rect 24584 22442 24636 22448
rect 24596 22234 24624 22442
rect 24584 22228 24636 22234
rect 24584 22170 24636 22176
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24412 21554 24440 21966
rect 24780 21894 24808 22494
rect 24964 22438 24992 22510
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 24858 22264 24914 22273
rect 24858 22199 24914 22208
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24504 20262 24532 21626
rect 24492 20256 24544 20262
rect 24492 20198 24544 20204
rect 24320 19306 24532 19334
rect 24504 18358 24532 19306
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24412 16998 24440 17614
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24228 14006 24256 15370
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24504 14618 24532 14758
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24216 14000 24268 14006
rect 24216 13942 24268 13948
rect 24228 13870 24256 13942
rect 24504 13938 24532 14418
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 24596 12434 24624 21830
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24688 20602 24716 21490
rect 24872 20942 24900 22199
rect 24964 22030 24992 22374
rect 25056 22030 25084 22578
rect 25240 22030 25268 22578
rect 25516 22030 25544 22986
rect 26400 22876 26708 22885
rect 26400 22874 26406 22876
rect 26462 22874 26486 22876
rect 26542 22874 26566 22876
rect 26622 22874 26646 22876
rect 26702 22874 26708 22876
rect 26462 22822 26464 22874
rect 26644 22822 26646 22874
rect 26400 22820 26406 22822
rect 26462 22820 26486 22822
rect 26542 22820 26566 22822
rect 26622 22820 26646 22822
rect 26702 22820 26708 22822
rect 26400 22811 26708 22820
rect 25740 22332 26048 22341
rect 25740 22330 25746 22332
rect 25802 22330 25826 22332
rect 25882 22330 25906 22332
rect 25962 22330 25986 22332
rect 26042 22330 26048 22332
rect 25802 22278 25804 22330
rect 25984 22278 25986 22330
rect 25740 22276 25746 22278
rect 25802 22276 25826 22278
rect 25882 22276 25906 22278
rect 25962 22276 25986 22278
rect 26042 22276 26048 22278
rect 25740 22267 26048 22276
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 26146 21992 26202 22001
rect 25042 21856 25098 21865
rect 25240 21842 25268 21966
rect 25098 21814 25268 21842
rect 25042 21791 25098 21800
rect 25516 21554 25544 21966
rect 26146 21927 26202 21936
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 24952 21548 25004 21554
rect 24952 21490 25004 21496
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 24964 21350 24992 21490
rect 25608 21486 25636 21830
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 25608 21146 25636 21422
rect 25740 21244 26048 21253
rect 25740 21242 25746 21244
rect 25802 21242 25826 21244
rect 25882 21242 25906 21244
rect 25962 21242 25986 21244
rect 26042 21242 26048 21244
rect 25802 21190 25804 21242
rect 25984 21190 25986 21242
rect 25740 21188 25746 21190
rect 25802 21188 25826 21190
rect 25882 21188 25906 21190
rect 25962 21188 25986 21190
rect 26042 21188 26048 21190
rect 25740 21179 26048 21188
rect 26160 21146 26188 21927
rect 26400 21788 26708 21797
rect 26400 21786 26406 21788
rect 26462 21786 26486 21788
rect 26542 21786 26566 21788
rect 26622 21786 26646 21788
rect 26702 21786 26708 21788
rect 26462 21734 26464 21786
rect 26644 21734 26646 21786
rect 26400 21732 26406 21734
rect 26462 21732 26486 21734
rect 26542 21732 26566 21734
rect 26622 21732 26646 21734
rect 26702 21732 26708 21734
rect 26400 21723 26708 21732
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 25596 21140 25648 21146
rect 25596 21082 25648 21088
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 26252 20942 26280 21354
rect 26988 21146 27016 21490
rect 27066 21448 27122 21457
rect 27066 21383 27068 21392
rect 27120 21383 27122 21392
rect 27068 21354 27120 21360
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 25872 20868 25924 20874
rect 25872 20810 25924 20816
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24872 17746 24900 18022
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24964 17241 24992 18294
rect 25056 17270 25084 19722
rect 25332 18426 25360 20810
rect 25884 20534 25912 20810
rect 26400 20700 26708 20709
rect 26400 20698 26406 20700
rect 26462 20698 26486 20700
rect 26542 20698 26566 20700
rect 26622 20698 26646 20700
rect 26702 20698 26708 20700
rect 26462 20646 26464 20698
rect 26644 20646 26646 20698
rect 26400 20644 26406 20646
rect 26462 20644 26486 20646
rect 26542 20644 26566 20646
rect 26622 20644 26646 20646
rect 26702 20644 26708 20646
rect 26400 20635 26708 20644
rect 26804 20534 26832 20878
rect 27080 20602 27108 20946
rect 27068 20596 27120 20602
rect 27068 20538 27120 20544
rect 25872 20528 25924 20534
rect 25872 20470 25924 20476
rect 26792 20528 26844 20534
rect 26792 20470 26844 20476
rect 27264 20330 27292 21286
rect 27540 21010 27568 21490
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27528 21004 27580 21010
rect 27356 20964 27528 20992
rect 27356 20466 27384 20964
rect 27528 20946 27580 20952
rect 27436 20800 27488 20806
rect 27436 20742 27488 20748
rect 27448 20466 27476 20742
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 25740 20156 26048 20165
rect 25740 20154 25746 20156
rect 25802 20154 25826 20156
rect 25882 20154 25906 20156
rect 25962 20154 25986 20156
rect 26042 20154 26048 20156
rect 25802 20102 25804 20154
rect 25984 20102 25986 20154
rect 25740 20100 25746 20102
rect 25802 20100 25826 20102
rect 25882 20100 25906 20102
rect 25962 20100 25986 20102
rect 26042 20100 26048 20102
rect 25740 20091 26048 20100
rect 27264 19854 27292 20266
rect 27356 20262 27384 20402
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27356 19854 27384 20198
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 25740 19068 26048 19077
rect 25740 19066 25746 19068
rect 25802 19066 25826 19068
rect 25882 19066 25906 19068
rect 25962 19066 25986 19068
rect 26042 19066 26048 19068
rect 25802 19014 25804 19066
rect 25984 19014 25986 19066
rect 25740 19012 25746 19014
rect 25802 19012 25826 19014
rect 25882 19012 25906 19014
rect 25962 19012 25986 19014
rect 26042 19012 26048 19014
rect 25740 19003 26048 19012
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 25320 17650 25372 17656
rect 25320 17592 25372 17598
rect 25412 17604 25464 17610
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25148 17338 25176 17478
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25044 17264 25096 17270
rect 24950 17232 25006 17241
rect 25044 17206 25096 17212
rect 24950 17167 25006 17176
rect 24964 17134 24992 17167
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24688 15570 24716 16526
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24780 15314 24808 15574
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24688 15286 24808 15314
rect 24688 15094 24716 15286
rect 24872 15178 24900 15370
rect 24780 15150 24900 15178
rect 24780 15094 24808 15150
rect 24964 15094 24992 15642
rect 25240 15434 25268 17478
rect 25332 16794 25360 17592
rect 25412 17546 25464 17552
rect 25424 17338 25452 17546
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25516 17202 25544 18158
rect 25740 17980 26048 17989
rect 25740 17978 25746 17980
rect 25802 17978 25826 17980
rect 25882 17978 25906 17980
rect 25962 17978 25986 17980
rect 26042 17978 26048 17980
rect 25802 17926 25804 17978
rect 25984 17926 25986 17978
rect 25740 17924 25746 17926
rect 25802 17924 25826 17926
rect 25882 17924 25906 17926
rect 25962 17924 25986 17926
rect 26042 17924 26048 17926
rect 25740 17915 26048 17924
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 25594 17776 25650 17785
rect 25594 17711 25650 17720
rect 25608 17542 25636 17711
rect 25976 17678 26004 17818
rect 26160 17746 26188 18158
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 26056 17740 26108 17746
rect 26056 17682 26108 17688
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 26068 17338 26096 17682
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17338 26188 17478
rect 26056 17332 26108 17338
rect 26056 17274 26108 17280
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25504 17196 25556 17202
rect 25556 17156 25636 17184
rect 25504 17138 25556 17144
rect 25320 16788 25372 16794
rect 25320 16730 25372 16736
rect 25424 16658 25452 17138
rect 25608 16658 25636 17156
rect 25740 16892 26048 16901
rect 25740 16890 25746 16892
rect 25802 16890 25826 16892
rect 25882 16890 25906 16892
rect 25962 16890 25986 16892
rect 26042 16890 26048 16892
rect 25802 16838 25804 16890
rect 25984 16838 25986 16890
rect 25740 16836 25746 16838
rect 25802 16836 25826 16838
rect 25882 16836 25906 16838
rect 25962 16836 25986 16838
rect 26042 16836 26048 16838
rect 25740 16827 26048 16836
rect 26252 16794 26280 17750
rect 26344 17728 26372 19654
rect 26400 19612 26708 19621
rect 26400 19610 26406 19612
rect 26462 19610 26486 19612
rect 26542 19610 26566 19612
rect 26622 19610 26646 19612
rect 26702 19610 26708 19612
rect 26462 19558 26464 19610
rect 26644 19558 26646 19610
rect 26400 19556 26406 19558
rect 26462 19556 26486 19558
rect 26542 19556 26566 19558
rect 26622 19556 26646 19558
rect 26702 19556 26708 19558
rect 26400 19547 26708 19556
rect 26400 18524 26708 18533
rect 26400 18522 26406 18524
rect 26462 18522 26486 18524
rect 26542 18522 26566 18524
rect 26622 18522 26646 18524
rect 26702 18522 26708 18524
rect 26462 18470 26464 18522
rect 26644 18470 26646 18522
rect 26400 18468 26406 18470
rect 26462 18468 26486 18470
rect 26542 18468 26566 18470
rect 26622 18468 26646 18470
rect 26702 18468 26708 18470
rect 26400 18459 26708 18468
rect 26884 18216 26936 18222
rect 26884 18158 26936 18164
rect 26608 18080 26660 18086
rect 26608 18022 26660 18028
rect 26424 17740 26476 17746
rect 26344 17700 26424 17728
rect 26344 17105 26372 17700
rect 26516 17740 26568 17746
rect 26476 17700 26516 17728
rect 26424 17682 26476 17688
rect 26516 17682 26568 17688
rect 26620 17678 26648 18022
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26516 17536 26568 17542
rect 26568 17496 26832 17524
rect 26516 17478 26568 17484
rect 26400 17436 26708 17445
rect 26400 17434 26406 17436
rect 26462 17434 26486 17436
rect 26542 17434 26566 17436
rect 26622 17434 26646 17436
rect 26702 17434 26708 17436
rect 26462 17382 26464 17434
rect 26644 17382 26646 17434
rect 26400 17380 26406 17382
rect 26462 17380 26486 17382
rect 26542 17380 26566 17382
rect 26622 17380 26646 17382
rect 26702 17380 26708 17382
rect 26400 17371 26708 17380
rect 26424 17332 26476 17338
rect 26476 17292 26740 17320
rect 26424 17274 26476 17280
rect 26712 17202 26740 17292
rect 26516 17196 26568 17202
rect 26700 17196 26752 17202
rect 26568 17156 26648 17184
rect 26516 17138 26568 17144
rect 26330 17096 26386 17105
rect 26330 17031 26386 17040
rect 26516 17060 26568 17066
rect 26344 16998 26372 17031
rect 26516 17002 26568 17008
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26528 16794 26556 17002
rect 26620 16998 26648 17156
rect 26700 17138 26752 17144
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26516 16788 26568 16794
rect 26516 16730 26568 16736
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 25424 16182 25452 16594
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 25240 15162 25268 15370
rect 25228 15156 25280 15162
rect 25228 15098 25280 15104
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 24872 14958 24900 15030
rect 25424 14958 25452 16118
rect 26252 15978 26280 16594
rect 26528 16590 26556 16730
rect 26804 16658 26832 17496
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 26424 16584 26476 16590
rect 26344 16544 26424 16572
rect 26344 16114 26372 16544
rect 26424 16526 26476 16532
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26792 16516 26844 16522
rect 26792 16458 26844 16464
rect 26400 16348 26708 16357
rect 26400 16346 26406 16348
rect 26462 16346 26486 16348
rect 26542 16346 26566 16348
rect 26622 16346 26646 16348
rect 26702 16346 26708 16348
rect 26462 16294 26464 16346
rect 26644 16294 26646 16346
rect 26400 16292 26406 16294
rect 26462 16292 26486 16294
rect 26542 16292 26566 16294
rect 26622 16292 26646 16294
rect 26702 16292 26708 16294
rect 26400 16283 26708 16292
rect 26804 16250 26832 16458
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26240 15972 26292 15978
rect 26240 15914 26292 15920
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 25740 15804 26048 15813
rect 25740 15802 25746 15804
rect 25802 15802 25826 15804
rect 25882 15802 25906 15804
rect 25962 15802 25986 15804
rect 26042 15802 26048 15804
rect 25802 15750 25804 15802
rect 25984 15750 25986 15802
rect 25740 15748 25746 15750
rect 25802 15748 25826 15750
rect 25882 15748 25906 15750
rect 25962 15748 25986 15750
rect 26042 15748 26048 15750
rect 25740 15739 26048 15748
rect 26160 15706 26188 15846
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26700 15700 26752 15706
rect 26700 15642 26752 15648
rect 26712 15502 26740 15642
rect 26804 15502 26832 15914
rect 26700 15496 26752 15502
rect 26606 15464 26662 15473
rect 26700 15438 26752 15444
rect 26792 15496 26844 15502
rect 26792 15438 26844 15444
rect 26606 15399 26662 15408
rect 26620 15366 26648 15399
rect 26332 15360 26384 15366
rect 26608 15360 26660 15366
rect 26384 15320 26608 15348
rect 26332 15302 26384 15308
rect 26608 15302 26660 15308
rect 26400 15260 26708 15269
rect 26400 15258 26406 15260
rect 26462 15258 26486 15260
rect 26542 15258 26566 15260
rect 26622 15258 26646 15260
rect 26702 15258 26708 15260
rect 26462 15206 26464 15258
rect 26644 15206 26646 15258
rect 26400 15204 26406 15206
rect 26462 15204 26486 15206
rect 26542 15204 26566 15206
rect 26622 15204 26646 15206
rect 26702 15204 26708 15206
rect 26400 15195 26708 15204
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26252 15026 26280 15098
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25044 14340 25096 14346
rect 25044 14282 25096 14288
rect 25320 14340 25372 14346
rect 25320 14282 25372 14288
rect 25056 14006 25084 14282
rect 25332 14006 25360 14282
rect 25424 14278 25452 14894
rect 25740 14716 26048 14725
rect 25740 14714 25746 14716
rect 25802 14714 25826 14716
rect 25882 14714 25906 14716
rect 25962 14714 25986 14716
rect 26042 14714 26048 14716
rect 25802 14662 25804 14714
rect 25984 14662 25986 14714
rect 25740 14660 25746 14662
rect 25802 14660 25826 14662
rect 25882 14660 25906 14662
rect 25962 14660 25986 14662
rect 26042 14660 26048 14662
rect 25740 14651 26048 14660
rect 26896 14618 26924 18158
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 26988 17066 27016 18022
rect 26976 17060 27028 17066
rect 26976 17002 27028 17008
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26988 15094 27016 15302
rect 26976 15088 27028 15094
rect 26976 15030 27028 15036
rect 27080 15042 27108 19654
rect 27448 19378 27476 20402
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27540 19854 27568 20198
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27632 19718 27660 21286
rect 27816 21010 27844 21490
rect 27988 21072 28040 21078
rect 27988 21014 28040 21020
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 28000 20874 28028 21014
rect 27988 20868 28040 20874
rect 27988 20810 28040 20816
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27724 18766 27752 20198
rect 28000 19854 28028 20810
rect 28172 20800 28224 20806
rect 28172 20742 28224 20748
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 28092 20058 28120 20402
rect 28080 20052 28132 20058
rect 28080 19994 28132 20000
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28092 19514 28120 19994
rect 28184 19854 28212 20742
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 27804 19304 27856 19310
rect 27804 19246 27856 19252
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27252 18216 27304 18222
rect 27252 18158 27304 18164
rect 27264 17882 27292 18158
rect 27816 18057 27844 19246
rect 27988 18352 28040 18358
rect 27988 18294 28040 18300
rect 27802 18048 27858 18057
rect 27802 17983 27858 17992
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 27344 17808 27396 17814
rect 27344 17750 27396 17756
rect 27160 17604 27212 17610
rect 27160 17546 27212 17552
rect 27172 16794 27200 17546
rect 27356 17252 27384 17750
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 27540 17270 27568 17614
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27264 17224 27384 17252
rect 27528 17264 27580 17270
rect 27264 17134 27292 17224
rect 27528 17206 27580 17212
rect 27632 17252 27660 17478
rect 27908 17338 27936 17614
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 27712 17264 27764 17270
rect 27632 17224 27712 17252
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27436 17128 27488 17134
rect 27436 17070 27488 17076
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 27160 16788 27212 16794
rect 27160 16730 27212 16736
rect 27264 16538 27292 16934
rect 27172 16510 27292 16538
rect 27172 16454 27200 16510
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27172 15706 27200 16390
rect 27160 15700 27212 15706
rect 27160 15642 27212 15648
rect 27264 15502 27292 16390
rect 27448 15638 27476 17070
rect 27540 16046 27568 17070
rect 27632 16590 27660 17224
rect 28000 17241 28028 18294
rect 28080 17536 28132 17542
rect 28080 17478 28132 17484
rect 27712 17206 27764 17212
rect 27986 17232 28042 17241
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27896 17196 27948 17202
rect 27986 17167 28042 17176
rect 27896 17138 27948 17144
rect 27816 16794 27844 17138
rect 27908 17105 27936 17138
rect 27894 17096 27950 17105
rect 27894 17031 27950 17040
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27436 15632 27488 15638
rect 27436 15574 27488 15580
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27344 15496 27396 15502
rect 27344 15438 27396 15444
rect 27252 15360 27304 15366
rect 27252 15302 27304 15308
rect 27080 15014 27200 15042
rect 27068 14816 27120 14822
rect 27068 14758 27120 14764
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 27080 14482 27108 14758
rect 27068 14476 27120 14482
rect 27068 14418 27120 14424
rect 25412 14272 25464 14278
rect 25412 14214 25464 14220
rect 26400 14172 26708 14181
rect 26400 14170 26406 14172
rect 26462 14170 26486 14172
rect 26542 14170 26566 14172
rect 26622 14170 26646 14172
rect 26702 14170 26708 14172
rect 26462 14118 26464 14170
rect 26644 14118 26646 14170
rect 26400 14116 26406 14118
rect 26462 14116 26486 14118
rect 26542 14116 26566 14118
rect 26622 14116 26646 14118
rect 26702 14116 26708 14118
rect 26400 14107 26708 14116
rect 25044 14000 25096 14006
rect 25044 13942 25096 13948
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24964 13530 24992 13670
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 25056 13394 25084 13942
rect 25332 13870 25360 13942
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24136 12406 24256 12434
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 24044 11642 24072 11698
rect 23952 11614 24072 11642
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24136 11082 24164 11494
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 23952 10810 23980 10950
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23110 10024 23166 10033
rect 23110 9959 23166 9968
rect 24228 9194 24256 12406
rect 24504 12406 24624 12434
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24320 10538 24348 10950
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 23952 9166 24256 9194
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 22928 8492 22980 8498
rect 22848 8452 22928 8480
rect 22848 7410 22876 8452
rect 22928 8434 22980 8440
rect 23032 8362 23060 8570
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23020 8356 23072 8362
rect 23020 8298 23072 8304
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22940 7546 22968 8230
rect 23032 8022 23060 8298
rect 23216 8294 23244 8434
rect 23400 8430 23428 8910
rect 23664 8560 23716 8566
rect 23584 8520 23664 8548
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23216 8266 23428 8294
rect 23020 8016 23072 8022
rect 23020 7958 23072 7964
rect 23400 7886 23428 8266
rect 23492 7886 23520 8434
rect 23584 7886 23612 8520
rect 23664 8502 23716 8508
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23676 7886 23704 8298
rect 23768 7886 23796 8366
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23032 7546 23060 7822
rect 23296 7744 23348 7750
rect 23492 7732 23520 7822
rect 23768 7750 23796 7822
rect 23348 7704 23520 7732
rect 23664 7744 23716 7750
rect 23296 7686 23348 7692
rect 23664 7686 23716 7692
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23308 7410 23336 7686
rect 23676 7546 23704 7686
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23860 6934 23888 8026
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 21916 6792 21968 6798
rect 20074 6760 20130 6769
rect 21916 6734 21968 6740
rect 20074 6695 20130 6704
rect 19317 6556 19625 6565
rect 19317 6554 19323 6556
rect 19379 6554 19403 6556
rect 19459 6554 19483 6556
rect 19539 6554 19563 6556
rect 19619 6554 19625 6556
rect 19379 6502 19381 6554
rect 19561 6502 19563 6554
rect 19317 6500 19323 6502
rect 19379 6500 19403 6502
rect 19459 6500 19483 6502
rect 19539 6500 19563 6502
rect 19619 6500 19625 6502
rect 19317 6491 19625 6500
rect 20088 6458 20116 6695
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20258 6352 20314 6361
rect 20076 6316 20128 6322
rect 20258 6287 20260 6296
rect 20076 6258 20128 6264
rect 20312 6287 20314 6296
rect 20536 6316 20588 6322
rect 20260 6258 20312 6264
rect 20536 6258 20588 6264
rect 18657 6012 18965 6021
rect 18657 6010 18663 6012
rect 18719 6010 18743 6012
rect 18799 6010 18823 6012
rect 18879 6010 18903 6012
rect 18959 6010 18965 6012
rect 18719 5958 18721 6010
rect 18901 5958 18903 6010
rect 18657 5956 18663 5958
rect 18719 5956 18743 5958
rect 18799 5956 18823 5958
rect 18879 5956 18903 5958
rect 18959 5956 18965 5958
rect 18657 5947 18965 5956
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17972 5030 18000 5510
rect 18248 5234 18276 5510
rect 18326 5400 18382 5409
rect 18326 5335 18382 5344
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18234 5128 18290 5137
rect 18052 5092 18104 5098
rect 18234 5063 18236 5072
rect 18052 5034 18104 5040
rect 18288 5063 18290 5072
rect 18236 5034 18288 5040
rect 17868 5024 17920 5030
rect 17774 4992 17830 5001
rect 17868 4966 17920 4972
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17774 4927 17830 4936
rect 17774 4856 17830 4865
rect 17880 4826 17908 4966
rect 17774 4791 17776 4800
rect 17828 4791 17830 4800
rect 17868 4820 17920 4826
rect 17776 4762 17828 4768
rect 17868 4762 17920 4768
rect 17866 4720 17922 4729
rect 17776 4684 17828 4690
rect 17696 4644 17776 4672
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17328 3534 17356 3946
rect 17420 3942 17448 4558
rect 17498 4176 17554 4185
rect 17498 4111 17554 4120
rect 17512 4078 17540 4111
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 13596 3012 13676 3040
rect 13728 3052 13780 3058
rect 13544 2994 13596 3000
rect 13728 2994 13780 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13740 2446 13768 2994
rect 13832 2446 13860 2994
rect 17144 2854 17172 2994
rect 17420 2972 17448 3878
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17512 3194 17540 3334
rect 17604 3194 17632 3334
rect 17696 3194 17724 4644
rect 17866 4655 17868 4664
rect 17776 4626 17828 4632
rect 17920 4655 17922 4664
rect 17868 4626 17920 4632
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17788 3058 17816 3470
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17972 2990 18000 4966
rect 18064 4672 18092 5034
rect 18236 4684 18288 4690
rect 18064 4644 18236 4672
rect 18236 4626 18288 4632
rect 18340 4486 18368 5335
rect 18432 5166 18460 5646
rect 18524 5234 18552 5714
rect 19317 5468 19625 5477
rect 19317 5466 19323 5468
rect 19379 5466 19403 5468
rect 19459 5466 19483 5468
rect 19539 5466 19563 5468
rect 19619 5466 19625 5468
rect 19379 5414 19381 5466
rect 19561 5414 19563 5466
rect 19317 5412 19323 5414
rect 19379 5412 19403 5414
rect 19459 5412 19483 5414
rect 19539 5412 19563 5414
rect 19619 5412 19625 5414
rect 19317 5403 19625 5412
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18418 4992 18474 5001
rect 18418 4927 18474 4936
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18064 3602 18092 4422
rect 18432 4146 18460 4927
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18524 3534 18552 5170
rect 19064 5024 19116 5030
rect 19524 5024 19576 5030
rect 19064 4966 19116 4972
rect 19352 4972 19524 4978
rect 19352 4966 19576 4972
rect 18657 4924 18965 4933
rect 18657 4922 18663 4924
rect 18719 4922 18743 4924
rect 18799 4922 18823 4924
rect 18879 4922 18903 4924
rect 18959 4922 18965 4924
rect 18719 4870 18721 4922
rect 18901 4870 18903 4922
rect 18657 4868 18663 4870
rect 18719 4868 18743 4870
rect 18799 4868 18823 4870
rect 18879 4868 18903 4870
rect 18959 4868 18965 4870
rect 18657 4859 18965 4868
rect 18602 4720 18658 4729
rect 18602 4655 18658 4664
rect 18616 4622 18644 4655
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18657 3836 18965 3845
rect 18657 3834 18663 3836
rect 18719 3834 18743 3836
rect 18799 3834 18823 3836
rect 18879 3834 18903 3836
rect 18959 3834 18965 3836
rect 18719 3782 18721 3834
rect 18901 3782 18903 3834
rect 18657 3780 18663 3782
rect 18719 3780 18743 3782
rect 18799 3780 18823 3782
rect 18879 3780 18903 3782
rect 18959 3780 18965 3782
rect 18657 3771 18965 3780
rect 18880 3664 18932 3670
rect 18878 3632 18880 3641
rect 18932 3632 18934 3641
rect 18878 3567 18934 3576
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 3194 18828 3334
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 19076 3058 19104 4966
rect 19352 4950 19564 4966
rect 19352 4690 19380 4950
rect 19536 4690 19564 4950
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19524 4684 19576 4690
rect 19576 4644 19748 4672
rect 19524 4626 19576 4632
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19260 4146 19288 4558
rect 19444 4486 19472 4626
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19317 4380 19625 4389
rect 19317 4378 19323 4380
rect 19379 4378 19403 4380
rect 19459 4378 19483 4380
rect 19539 4378 19563 4380
rect 19619 4378 19625 4380
rect 19379 4326 19381 4378
rect 19561 4326 19563 4378
rect 19317 4324 19323 4326
rect 19379 4324 19403 4326
rect 19459 4324 19483 4326
rect 19539 4324 19563 4326
rect 19619 4324 19625 4326
rect 19317 4315 19625 4324
rect 19720 4282 19748 4644
rect 19812 4622 19840 4762
rect 20088 4758 20116 6258
rect 20272 5370 20300 6258
rect 20548 6202 20576 6258
rect 20456 6174 20576 6202
rect 20456 6118 20484 6174
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 19800 4616 19852 4622
rect 19852 4564 19932 4570
rect 19800 4558 19932 4564
rect 19812 4542 19932 4558
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19812 4214 19840 4422
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19904 4010 19932 4542
rect 20088 4146 20116 4694
rect 20456 4622 20484 6054
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20732 4622 20760 4966
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19892 4004 19944 4010
rect 19892 3946 19944 3952
rect 19317 3292 19625 3301
rect 19317 3290 19323 3292
rect 19379 3290 19403 3292
rect 19459 3290 19483 3292
rect 19539 3290 19563 3292
rect 19619 3290 19625 3292
rect 19379 3238 19381 3290
rect 19561 3238 19563 3290
rect 19317 3236 19323 3238
rect 19379 3236 19403 3238
rect 19459 3236 19483 3238
rect 19539 3236 19563 3238
rect 19619 3236 19625 3238
rect 19317 3227 19625 3236
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 17500 2984 17552 2990
rect 17420 2944 17500 2972
rect 17500 2926 17552 2932
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 17512 2378 17540 2926
rect 19904 2854 19932 3946
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 18657 2748 18965 2757
rect 18657 2746 18663 2748
rect 18719 2746 18743 2748
rect 18799 2746 18823 2748
rect 18879 2746 18903 2748
rect 18959 2746 18965 2748
rect 18719 2694 18721 2746
rect 18901 2694 18903 2746
rect 18657 2692 18663 2694
rect 18719 2692 18743 2694
rect 18799 2692 18823 2694
rect 18879 2692 18903 2694
rect 18959 2692 18965 2694
rect 18657 2683 18965 2692
rect 20088 2378 20116 4082
rect 20180 3942 20208 4558
rect 20456 4282 20484 4558
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 23952 4049 23980 9166
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 24044 8498 24072 9046
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24044 8106 24072 8434
rect 24044 8078 24164 8106
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 24044 7410 24072 7958
rect 24136 7886 24164 8078
rect 24228 7954 24256 8502
rect 24216 7948 24268 7954
rect 24216 7890 24268 7896
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24044 6934 24072 7346
rect 24136 7274 24164 7822
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24228 7410 24256 7754
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 24136 6934 24164 7210
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 24124 6928 24176 6934
rect 24124 6870 24176 6876
rect 24228 6798 24256 7346
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 24320 6730 24348 10474
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24412 7002 24440 7142
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24308 6724 24360 6730
rect 24308 6666 24360 6672
rect 24306 5536 24362 5545
rect 24306 5471 24362 5480
rect 24320 4214 24348 5471
rect 24308 4208 24360 4214
rect 24308 4150 24360 4156
rect 24504 4146 24532 12406
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 10742 24624 11494
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 24584 10736 24636 10742
rect 24584 10678 24636 10684
rect 24964 9178 24992 11154
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 25056 10742 25084 10950
rect 25240 10810 25268 11018
rect 25332 11014 25360 13806
rect 25740 13628 26048 13637
rect 25740 13626 25746 13628
rect 25802 13626 25826 13628
rect 25882 13626 25906 13628
rect 25962 13626 25986 13628
rect 26042 13626 26048 13628
rect 25802 13574 25804 13626
rect 25984 13574 25986 13626
rect 25740 13572 25746 13574
rect 25802 13572 25826 13574
rect 25882 13572 25906 13574
rect 25962 13572 25986 13574
rect 26042 13572 26048 13574
rect 25740 13563 26048 13572
rect 26400 13084 26708 13093
rect 26400 13082 26406 13084
rect 26462 13082 26486 13084
rect 26542 13082 26566 13084
rect 26622 13082 26646 13084
rect 26702 13082 26708 13084
rect 26462 13030 26464 13082
rect 26644 13030 26646 13082
rect 26400 13028 26406 13030
rect 26462 13028 26486 13030
rect 26542 13028 26566 13030
rect 26622 13028 26646 13030
rect 26702 13028 26708 13030
rect 26400 13019 26708 13028
rect 25740 12540 26048 12549
rect 25740 12538 25746 12540
rect 25802 12538 25826 12540
rect 25882 12538 25906 12540
rect 25962 12538 25986 12540
rect 26042 12538 26048 12540
rect 25802 12486 25804 12538
rect 25984 12486 25986 12538
rect 25740 12484 25746 12486
rect 25802 12484 25826 12486
rect 25882 12484 25906 12486
rect 25962 12484 25986 12486
rect 26042 12484 26048 12486
rect 25740 12475 26048 12484
rect 26400 11996 26708 12005
rect 26400 11994 26406 11996
rect 26462 11994 26486 11996
rect 26542 11994 26566 11996
rect 26622 11994 26646 11996
rect 26702 11994 26708 11996
rect 26462 11942 26464 11994
rect 26644 11942 26646 11994
rect 26400 11940 26406 11942
rect 26462 11940 26486 11942
rect 26542 11940 26566 11942
rect 26622 11940 26646 11942
rect 26702 11940 26708 11942
rect 26400 11931 26708 11940
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 25516 10690 25544 11834
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 25740 11452 26048 11461
rect 25740 11450 25746 11452
rect 25802 11450 25826 11452
rect 25882 11450 25906 11452
rect 25962 11450 25986 11452
rect 26042 11450 26048 11452
rect 25802 11398 25804 11450
rect 25984 11398 25986 11450
rect 25740 11396 25746 11398
rect 25802 11396 25826 11398
rect 25882 11396 25906 11398
rect 25962 11396 25986 11398
rect 26042 11396 26048 11398
rect 25740 11387 26048 11396
rect 25780 10736 25832 10742
rect 25516 10684 25780 10690
rect 25516 10678 25832 10684
rect 25516 10662 25820 10678
rect 26160 10674 26188 11494
rect 26712 11354 26740 11698
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 27068 11076 27120 11082
rect 27068 11018 27120 11024
rect 26792 11008 26844 11014
rect 26792 10950 26844 10956
rect 26400 10908 26708 10917
rect 26400 10906 26406 10908
rect 26462 10906 26486 10908
rect 26542 10906 26566 10908
rect 26622 10906 26646 10908
rect 26702 10906 26708 10908
rect 26462 10854 26464 10906
rect 26644 10854 26646 10906
rect 26400 10852 26406 10854
rect 26462 10852 26486 10854
rect 26542 10852 26566 10854
rect 26622 10852 26646 10854
rect 26702 10852 26708 10854
rect 26400 10843 26708 10852
rect 26148 10668 26200 10674
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24688 7886 24716 8230
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24688 7562 24716 7822
rect 24596 7534 24716 7562
rect 24596 7478 24624 7534
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24964 7410 24992 9114
rect 25516 8956 25544 10662
rect 26148 10610 26200 10616
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26608 10668 26660 10674
rect 26804 10656 26832 10950
rect 26660 10628 26832 10656
rect 26608 10610 26660 10616
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25608 10266 25636 10542
rect 25740 10364 26048 10373
rect 25740 10362 25746 10364
rect 25802 10362 25826 10364
rect 25882 10362 25906 10364
rect 25962 10362 25986 10364
rect 26042 10362 26048 10364
rect 25802 10310 25804 10362
rect 25984 10310 25986 10362
rect 25740 10308 25746 10310
rect 25802 10308 25826 10310
rect 25882 10308 25906 10310
rect 25962 10308 25986 10310
rect 26042 10308 26048 10310
rect 25740 10299 26048 10308
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 26160 9926 26188 10610
rect 26436 10062 26464 10610
rect 26528 10130 26556 10610
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26148 9920 26200 9926
rect 26148 9862 26200 9868
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 26148 9444 26200 9450
rect 26148 9386 26200 9392
rect 25596 9376 25648 9382
rect 25596 9318 25648 9324
rect 25608 9110 25636 9318
rect 25740 9276 26048 9285
rect 25740 9274 25746 9276
rect 25802 9274 25826 9276
rect 25882 9274 25906 9276
rect 25962 9274 25986 9276
rect 26042 9274 26048 9276
rect 25802 9222 25804 9274
rect 25984 9222 25986 9274
rect 25740 9220 25746 9222
rect 25802 9220 25826 9222
rect 25882 9220 25906 9222
rect 25962 9220 25986 9222
rect 26042 9220 26048 9222
rect 25740 9211 26048 9220
rect 25596 9104 25648 9110
rect 25596 9046 25648 9052
rect 25688 9104 25740 9110
rect 25688 9046 25740 9052
rect 25700 8956 25728 9046
rect 26160 8974 26188 9386
rect 25516 8928 25728 8956
rect 26148 8968 26200 8974
rect 25516 7954 25544 8928
rect 26148 8910 26200 8916
rect 25780 8900 25832 8906
rect 25780 8842 25832 8848
rect 25872 8900 25924 8906
rect 25872 8842 25924 8848
rect 25792 8566 25820 8842
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25884 8294 25912 8842
rect 26252 8566 26280 9862
rect 26400 9820 26708 9829
rect 26400 9818 26406 9820
rect 26462 9818 26486 9820
rect 26542 9818 26566 9820
rect 26622 9818 26646 9820
rect 26702 9818 26708 9820
rect 26462 9766 26464 9818
rect 26644 9766 26646 9818
rect 26400 9764 26406 9766
rect 26462 9764 26486 9766
rect 26542 9764 26566 9766
rect 26622 9764 26646 9766
rect 26702 9764 26708 9766
rect 26400 9755 26708 9764
rect 26896 9654 26924 10066
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 26240 8560 26292 8566
rect 26240 8502 26292 8508
rect 26344 8514 26372 9522
rect 26896 9518 26924 9590
rect 26884 9512 26936 9518
rect 26884 9454 26936 9460
rect 26792 8900 26844 8906
rect 26792 8842 26844 8848
rect 26400 8732 26708 8741
rect 26400 8730 26406 8732
rect 26462 8730 26486 8732
rect 26542 8730 26566 8732
rect 26622 8730 26646 8732
rect 26702 8730 26708 8732
rect 26462 8678 26464 8730
rect 26644 8678 26646 8730
rect 26400 8676 26406 8678
rect 26462 8676 26486 8678
rect 26542 8676 26566 8678
rect 26622 8676 26646 8678
rect 26702 8676 26708 8678
rect 26400 8667 26708 8676
rect 26344 8498 26464 8514
rect 26344 8492 26476 8498
rect 26344 8486 26424 8492
rect 26424 8434 26476 8440
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 25884 8266 26280 8294
rect 25740 8188 26048 8197
rect 25740 8186 25746 8188
rect 25802 8186 25826 8188
rect 25882 8186 25906 8188
rect 25962 8186 25986 8188
rect 26042 8186 26048 8188
rect 25802 8134 25804 8186
rect 25984 8134 25986 8186
rect 25740 8132 25746 8134
rect 25802 8132 25826 8134
rect 25882 8132 25906 8134
rect 25962 8132 25986 8134
rect 26042 8132 26048 8134
rect 25740 8123 26048 8132
rect 26148 8016 26200 8022
rect 26252 8004 26280 8266
rect 26344 8022 26372 8366
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 26608 8356 26660 8362
rect 26804 8344 26832 8842
rect 26896 8498 26924 9454
rect 27080 8906 27108 11018
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 26884 8492 26936 8498
rect 26884 8434 26936 8440
rect 26884 8356 26936 8362
rect 26804 8316 26884 8344
rect 26608 8298 26660 8304
rect 26884 8298 26936 8304
rect 26200 7976 26280 8004
rect 26148 7958 26200 7964
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 26252 7818 26280 7976
rect 26332 8016 26384 8022
rect 26332 7958 26384 7964
rect 26528 7886 26556 8298
rect 26620 8090 26648 8298
rect 26608 8084 26660 8090
rect 26608 8026 26660 8032
rect 26620 7886 26648 8026
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 25872 7812 25924 7818
rect 25872 7754 25924 7760
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 26792 7812 26844 7818
rect 26792 7754 26844 7760
rect 25596 7744 25648 7750
rect 25596 7686 25648 7692
rect 25608 7546 25636 7686
rect 25884 7546 25912 7754
rect 26400 7644 26708 7653
rect 26400 7642 26406 7644
rect 26462 7642 26486 7644
rect 26542 7642 26566 7644
rect 26622 7642 26646 7644
rect 26702 7642 26708 7644
rect 26462 7590 26464 7642
rect 26644 7590 26646 7642
rect 26400 7588 26406 7590
rect 26462 7588 26486 7590
rect 26542 7588 26566 7590
rect 26622 7588 26646 7590
rect 26702 7588 26708 7590
rect 26400 7579 26708 7588
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 25332 6730 25360 7278
rect 26804 7274 26832 7754
rect 26896 7410 26924 8298
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 26988 7410 27016 7822
rect 27080 7410 27108 8842
rect 26884 7404 26936 7410
rect 26884 7346 26936 7352
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 27068 7404 27120 7410
rect 27068 7346 27120 7352
rect 26792 7268 26844 7274
rect 26792 7210 26844 7216
rect 25740 7100 26048 7109
rect 25740 7098 25746 7100
rect 25802 7098 25826 7100
rect 25882 7098 25906 7100
rect 25962 7098 25986 7100
rect 26042 7098 26048 7100
rect 25802 7046 25804 7098
rect 25984 7046 25986 7098
rect 25740 7044 25746 7046
rect 25802 7044 25826 7046
rect 25882 7044 25906 7046
rect 25962 7044 25986 7046
rect 26042 7044 26048 7046
rect 25740 7035 26048 7044
rect 25320 6724 25372 6730
rect 25320 6666 25372 6672
rect 26400 6556 26708 6565
rect 26400 6554 26406 6556
rect 26462 6554 26486 6556
rect 26542 6554 26566 6556
rect 26622 6554 26646 6556
rect 26702 6554 26708 6556
rect 26462 6502 26464 6554
rect 26644 6502 26646 6554
rect 26400 6500 26406 6502
rect 26462 6500 26486 6502
rect 26542 6500 26566 6502
rect 26622 6500 26646 6502
rect 26702 6500 26708 6502
rect 26400 6491 26708 6500
rect 25740 6012 26048 6021
rect 25740 6010 25746 6012
rect 25802 6010 25826 6012
rect 25882 6010 25906 6012
rect 25962 6010 25986 6012
rect 26042 6010 26048 6012
rect 25802 5958 25804 6010
rect 25984 5958 25986 6010
rect 25740 5956 25746 5958
rect 25802 5956 25826 5958
rect 25882 5956 25906 5958
rect 25962 5956 25986 5958
rect 26042 5956 26048 5958
rect 25740 5947 26048 5956
rect 26400 5468 26708 5477
rect 26400 5466 26406 5468
rect 26462 5466 26486 5468
rect 26542 5466 26566 5468
rect 26622 5466 26646 5468
rect 26702 5466 26708 5468
rect 26462 5414 26464 5466
rect 26644 5414 26646 5466
rect 26400 5412 26406 5414
rect 26462 5412 26486 5414
rect 26542 5412 26566 5414
rect 26622 5412 26646 5414
rect 26702 5412 26708 5414
rect 26400 5403 26708 5412
rect 25740 4924 26048 4933
rect 25740 4922 25746 4924
rect 25802 4922 25826 4924
rect 25882 4922 25906 4924
rect 25962 4922 25986 4924
rect 26042 4922 26048 4924
rect 25802 4870 25804 4922
rect 25984 4870 25986 4922
rect 25740 4868 25746 4870
rect 25802 4868 25826 4870
rect 25882 4868 25906 4870
rect 25962 4868 25986 4870
rect 26042 4868 26048 4870
rect 25740 4859 26048 4868
rect 26400 4380 26708 4389
rect 26400 4378 26406 4380
rect 26462 4378 26486 4380
rect 26542 4378 26566 4380
rect 26622 4378 26646 4380
rect 26702 4378 26708 4380
rect 26462 4326 26464 4378
rect 26644 4326 26646 4378
rect 26400 4324 26406 4326
rect 26462 4324 26486 4326
rect 26542 4324 26566 4326
rect 26622 4324 26646 4326
rect 26702 4324 26708 4326
rect 26400 4315 26708 4324
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 23938 4040 23994 4049
rect 23938 3975 23994 3984
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 20180 3602 20208 3878
rect 24412 3738 24440 3878
rect 24964 3738 24992 3878
rect 25740 3836 26048 3845
rect 25740 3834 25746 3836
rect 25802 3834 25826 3836
rect 25882 3834 25906 3836
rect 25962 3834 25986 3836
rect 26042 3834 26048 3836
rect 25802 3782 25804 3834
rect 25984 3782 25986 3834
rect 25740 3780 25746 3782
rect 25802 3780 25826 3782
rect 25882 3780 25906 3782
rect 25962 3780 25986 3782
rect 26042 3780 26048 3782
rect 25740 3771 26048 3780
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 21928 2366 22048 2394
rect 22112 2378 22140 3402
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 25240 2446 25268 3334
rect 26400 3292 26708 3301
rect 26400 3290 26406 3292
rect 26462 3290 26486 3292
rect 26542 3290 26566 3292
rect 26622 3290 26646 3292
rect 26702 3290 26708 3292
rect 26462 3238 26464 3290
rect 26644 3238 26646 3290
rect 26400 3236 26406 3238
rect 26462 3236 26486 3238
rect 26542 3236 26566 3238
rect 26622 3236 26646 3238
rect 26702 3236 26708 3238
rect 26400 3227 26708 3236
rect 27172 2774 27200 15014
rect 27264 14958 27292 15302
rect 27252 14952 27304 14958
rect 27252 14894 27304 14900
rect 27356 14822 27384 15438
rect 27540 14958 27568 15982
rect 27620 15700 27672 15706
rect 27620 15642 27672 15648
rect 27632 15162 27660 15642
rect 27712 15564 27764 15570
rect 27712 15506 27764 15512
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27724 14890 27752 15506
rect 27894 15464 27950 15473
rect 27894 15399 27896 15408
rect 27948 15399 27950 15408
rect 27896 15370 27948 15376
rect 27712 14884 27764 14890
rect 27712 14826 27764 14832
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27528 14340 27580 14346
rect 27528 14282 27580 14288
rect 27540 13870 27568 14282
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27632 13326 27660 14010
rect 28000 13938 28028 17167
rect 28092 16590 28120 17478
rect 28080 16584 28132 16590
rect 28080 16526 28132 16532
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 28080 9648 28132 9654
rect 28080 9590 28132 9596
rect 27804 9580 27856 9586
rect 27804 9522 27856 9528
rect 27816 9178 27844 9522
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 28092 8498 28120 9590
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 28184 8498 28212 9522
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 27632 8378 27660 8434
rect 27540 8362 27660 8378
rect 27528 8356 27660 8362
rect 27580 8350 27660 8356
rect 27528 8298 27580 8304
rect 27540 8090 27568 8298
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 27356 7410 27384 8026
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27540 7274 27568 7890
rect 27528 7268 27580 7274
rect 27528 7210 27580 7216
rect 28276 5370 28304 26930
rect 29000 26784 29052 26790
rect 29000 26726 29052 26732
rect 29012 26625 29040 26726
rect 28998 26616 29054 26625
rect 28998 26551 29054 26560
rect 28816 22636 28868 22642
rect 28816 22578 28868 22584
rect 28828 22030 28856 22578
rect 28998 22536 29054 22545
rect 28998 22471 29000 22480
rect 29052 22471 29054 22480
rect 29000 22442 29052 22448
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28908 21004 28960 21010
rect 28908 20946 28960 20952
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 28552 20534 28580 20742
rect 28540 20528 28592 20534
rect 28540 20470 28592 20476
rect 28920 20466 28948 20946
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28356 20256 28408 20262
rect 28356 20198 28408 20204
rect 28368 18442 28396 20198
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28368 18414 28580 18442
rect 28448 18216 28500 18222
rect 28448 18158 28500 18164
rect 28460 17610 28488 18158
rect 28448 17604 28500 17610
rect 28448 17546 28500 17552
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28368 17134 28396 17478
rect 28460 17202 28488 17546
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28356 17128 28408 17134
rect 28356 17070 28408 17076
rect 28368 16590 28396 17070
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28368 15162 28396 16526
rect 28356 15156 28408 15162
rect 28356 15098 28408 15104
rect 28448 9376 28500 9382
rect 28448 9318 28500 9324
rect 28460 8906 28488 9318
rect 28448 8900 28500 8906
rect 28448 8842 28500 8848
rect 28460 8566 28488 8842
rect 28448 8560 28500 8566
rect 28448 8502 28500 8508
rect 28264 5364 28316 5370
rect 28264 5306 28316 5312
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 28092 4826 28120 5170
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 25740 2748 26048 2757
rect 25740 2746 25746 2748
rect 25802 2746 25826 2748
rect 25882 2746 25906 2748
rect 25962 2746 25986 2748
rect 26042 2746 26048 2748
rect 25802 2694 25804 2746
rect 25984 2694 25986 2746
rect 25740 2692 25746 2694
rect 25802 2692 25826 2694
rect 25882 2692 25906 2694
rect 25962 2692 25986 2694
rect 26042 2692 26048 2694
rect 25740 2683 26048 2692
rect 27080 2746 27200 2774
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 27080 2378 27108 2746
rect 28552 2446 28580 18414
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28644 16590 28672 16934
rect 28632 16584 28684 16590
rect 28632 16526 28684 16532
rect 28736 11150 28764 19654
rect 29000 18624 29052 18630
rect 29000 18566 29052 18572
rect 29012 18465 29040 18566
rect 28998 18456 29054 18465
rect 28998 18391 29054 18400
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 28828 14482 28856 14962
rect 28816 14476 28868 14482
rect 28816 14418 28868 14424
rect 28906 14376 28962 14385
rect 28906 14311 28962 14320
rect 28920 13530 28948 14311
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 28908 11212 28960 11218
rect 28908 11154 28960 11160
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 28920 10985 28948 11154
rect 28906 10976 28962 10985
rect 28906 10911 28962 10920
rect 28724 7404 28776 7410
rect 28724 7346 28776 7352
rect 28736 6458 28764 7346
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 28920 6905 28948 7142
rect 28906 6896 28962 6905
rect 28906 6831 28962 6840
rect 28724 6452 28776 6458
rect 28724 6394 28776 6400
rect 29000 2848 29052 2854
rect 28998 2816 29000 2825
rect 29052 2816 29054 2825
rect 28998 2751 29054 2760
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 20 2304 72 2310
rect 3424 2304 3476 2310
rect 20 2246 72 2252
rect 3252 2264 3424 2292
rect 32 800 60 2246
rect 3252 800 3280 2264
rect 3424 2246 3476 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 5151 2204 5459 2213
rect 5151 2202 5157 2204
rect 5213 2202 5237 2204
rect 5293 2202 5317 2204
rect 5373 2202 5397 2204
rect 5453 2202 5459 2204
rect 5213 2150 5215 2202
rect 5395 2150 5397 2202
rect 5151 2148 5157 2150
rect 5213 2148 5237 2150
rect 5293 2148 5317 2150
rect 5373 2148 5397 2150
rect 5453 2148 5459 2150
rect 5151 2139 5459 2148
rect 7116 800 7144 2246
rect 11164 1442 11192 2246
rect 12234 2204 12542 2213
rect 12234 2202 12240 2204
rect 12296 2202 12320 2204
rect 12376 2202 12400 2204
rect 12456 2202 12480 2204
rect 12536 2202 12542 2204
rect 12296 2150 12298 2202
rect 12478 2150 12480 2202
rect 12234 2148 12240 2150
rect 12296 2148 12320 2150
rect 12376 2148 12400 2150
rect 12456 2148 12480 2150
rect 12536 2148 12542 2150
rect 12234 2139 12542 2148
rect 10980 1414 11192 1442
rect 10980 800 11008 1414
rect 14936 1170 14964 2246
rect 18892 1170 18920 2246
rect 19317 2204 19625 2213
rect 19317 2202 19323 2204
rect 19379 2202 19403 2204
rect 19459 2202 19483 2204
rect 19539 2202 19563 2204
rect 19619 2202 19625 2204
rect 19379 2150 19381 2202
rect 19561 2150 19563 2202
rect 19317 2148 19323 2150
rect 19379 2148 19403 2150
rect 19459 2148 19483 2150
rect 19539 2148 19563 2150
rect 19619 2148 19625 2150
rect 19317 2139 19625 2148
rect 14844 1142 14964 1170
rect 18708 1142 18920 1170
rect 14844 800 14872 1142
rect 18708 800 18736 1142
rect 21928 800 21956 2366
rect 22020 2310 22048 2366
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 29644 2372 29696 2378
rect 29644 2314 29696 2320
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 25792 870 25912 898
rect 25792 800 25820 870
rect 18 0 74 800
rect 3238 0 3294 800
rect 7102 0 7158 800
rect 10966 0 11022 800
rect 14830 0 14886 800
rect 18694 0 18750 800
rect 21914 0 21970 800
rect 25778 0 25834 800
rect 25884 762 25912 870
rect 26160 762 26188 2246
rect 26400 2204 26708 2213
rect 26400 2202 26406 2204
rect 26462 2202 26486 2204
rect 26542 2202 26566 2204
rect 26622 2202 26646 2204
rect 26702 2202 26708 2204
rect 26462 2150 26464 2202
rect 26644 2150 26646 2202
rect 26400 2148 26406 2150
rect 26462 2148 26486 2150
rect 26542 2148 26566 2150
rect 26622 2148 26646 2150
rect 26702 2148 26708 2150
rect 26400 2139 26708 2148
rect 29656 800 29684 2314
rect 25884 734 26188 762
rect 29642 0 29698 800
<< via2 >>
rect 1582 30912 1638 30968
rect 5157 30490 5213 30492
rect 5237 30490 5293 30492
rect 5317 30490 5373 30492
rect 5397 30490 5453 30492
rect 5157 30438 5203 30490
rect 5203 30438 5213 30490
rect 5237 30438 5267 30490
rect 5267 30438 5279 30490
rect 5279 30438 5293 30490
rect 5317 30438 5331 30490
rect 5331 30438 5343 30490
rect 5343 30438 5373 30490
rect 5397 30438 5407 30490
rect 5407 30438 5453 30490
rect 5157 30436 5213 30438
rect 5237 30436 5293 30438
rect 5317 30436 5373 30438
rect 5397 30436 5453 30438
rect 12240 30490 12296 30492
rect 12320 30490 12376 30492
rect 12400 30490 12456 30492
rect 12480 30490 12536 30492
rect 12240 30438 12286 30490
rect 12286 30438 12296 30490
rect 12320 30438 12350 30490
rect 12350 30438 12362 30490
rect 12362 30438 12376 30490
rect 12400 30438 12414 30490
rect 12414 30438 12426 30490
rect 12426 30438 12456 30490
rect 12480 30438 12490 30490
rect 12490 30438 12536 30490
rect 12240 30436 12296 30438
rect 12320 30436 12376 30438
rect 12400 30436 12456 30438
rect 12480 30436 12536 30438
rect 938 27276 940 27296
rect 940 27276 992 27296
rect 992 27276 994 27296
rect 938 27240 994 27276
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 1490 23024 1546 23080
rect 1582 19508 1638 19544
rect 1582 19488 1584 19508
rect 1584 19488 1636 19508
rect 1636 19488 1638 19508
rect 938 15680 994 15736
rect 938 11600 994 11656
rect 4497 29946 4553 29948
rect 4577 29946 4633 29948
rect 4657 29946 4713 29948
rect 4737 29946 4793 29948
rect 4497 29894 4543 29946
rect 4543 29894 4553 29946
rect 4577 29894 4607 29946
rect 4607 29894 4619 29946
rect 4619 29894 4633 29946
rect 4657 29894 4671 29946
rect 4671 29894 4683 29946
rect 4683 29894 4713 29946
rect 4737 29894 4747 29946
rect 4747 29894 4793 29946
rect 4497 29892 4553 29894
rect 4577 29892 4633 29894
rect 4657 29892 4713 29894
rect 4737 29892 4793 29894
rect 4497 28858 4553 28860
rect 4577 28858 4633 28860
rect 4657 28858 4713 28860
rect 4737 28858 4793 28860
rect 4497 28806 4543 28858
rect 4543 28806 4553 28858
rect 4577 28806 4607 28858
rect 4607 28806 4619 28858
rect 4619 28806 4633 28858
rect 4657 28806 4671 28858
rect 4671 28806 4683 28858
rect 4683 28806 4713 28858
rect 4737 28806 4747 28858
rect 4747 28806 4793 28858
rect 4497 28804 4553 28806
rect 4577 28804 4633 28806
rect 4657 28804 4713 28806
rect 4737 28804 4793 28806
rect 5157 29402 5213 29404
rect 5237 29402 5293 29404
rect 5317 29402 5373 29404
rect 5397 29402 5453 29404
rect 5157 29350 5203 29402
rect 5203 29350 5213 29402
rect 5237 29350 5267 29402
rect 5267 29350 5279 29402
rect 5279 29350 5293 29402
rect 5317 29350 5331 29402
rect 5331 29350 5343 29402
rect 5343 29350 5373 29402
rect 5397 29350 5407 29402
rect 5407 29350 5453 29402
rect 5157 29348 5213 29350
rect 5237 29348 5293 29350
rect 5317 29348 5373 29350
rect 5397 29348 5453 29350
rect 4497 27770 4553 27772
rect 4577 27770 4633 27772
rect 4657 27770 4713 27772
rect 4737 27770 4793 27772
rect 4497 27718 4543 27770
rect 4543 27718 4553 27770
rect 4577 27718 4607 27770
rect 4607 27718 4619 27770
rect 4619 27718 4633 27770
rect 4657 27718 4671 27770
rect 4671 27718 4683 27770
rect 4683 27718 4713 27770
rect 4737 27718 4747 27770
rect 4747 27718 4793 27770
rect 4497 27716 4553 27718
rect 4577 27716 4633 27718
rect 4657 27716 4713 27718
rect 4737 27716 4793 27718
rect 5157 28314 5213 28316
rect 5237 28314 5293 28316
rect 5317 28314 5373 28316
rect 5397 28314 5453 28316
rect 5157 28262 5203 28314
rect 5203 28262 5213 28314
rect 5237 28262 5267 28314
rect 5267 28262 5279 28314
rect 5279 28262 5293 28314
rect 5317 28262 5331 28314
rect 5331 28262 5343 28314
rect 5343 28262 5373 28314
rect 5397 28262 5407 28314
rect 5407 28262 5453 28314
rect 5157 28260 5213 28262
rect 5237 28260 5293 28262
rect 5317 28260 5373 28262
rect 5397 28260 5453 28262
rect 4497 26682 4553 26684
rect 4577 26682 4633 26684
rect 4657 26682 4713 26684
rect 4737 26682 4793 26684
rect 4497 26630 4543 26682
rect 4543 26630 4553 26682
rect 4577 26630 4607 26682
rect 4607 26630 4619 26682
rect 4619 26630 4633 26682
rect 4657 26630 4671 26682
rect 4671 26630 4683 26682
rect 4683 26630 4713 26682
rect 4737 26630 4747 26682
rect 4747 26630 4793 26682
rect 4497 26628 4553 26630
rect 4577 26628 4633 26630
rect 4657 26628 4713 26630
rect 4737 26628 4793 26630
rect 5157 27226 5213 27228
rect 5237 27226 5293 27228
rect 5317 27226 5373 27228
rect 5397 27226 5453 27228
rect 5157 27174 5203 27226
rect 5203 27174 5213 27226
rect 5237 27174 5267 27226
rect 5267 27174 5279 27226
rect 5279 27174 5293 27226
rect 5317 27174 5331 27226
rect 5331 27174 5343 27226
rect 5343 27174 5373 27226
rect 5397 27174 5407 27226
rect 5407 27174 5453 27226
rect 5157 27172 5213 27174
rect 5237 27172 5293 27174
rect 5317 27172 5373 27174
rect 5397 27172 5453 27174
rect 5157 26138 5213 26140
rect 5237 26138 5293 26140
rect 5317 26138 5373 26140
rect 5397 26138 5453 26140
rect 5157 26086 5203 26138
rect 5203 26086 5213 26138
rect 5237 26086 5267 26138
rect 5267 26086 5279 26138
rect 5279 26086 5293 26138
rect 5317 26086 5331 26138
rect 5331 26086 5343 26138
rect 5343 26086 5373 26138
rect 5397 26086 5407 26138
rect 5407 26086 5453 26138
rect 5157 26084 5213 26086
rect 5237 26084 5293 26086
rect 5317 26084 5373 26086
rect 5397 26084 5453 26086
rect 4497 25594 4553 25596
rect 4577 25594 4633 25596
rect 4657 25594 4713 25596
rect 4737 25594 4793 25596
rect 4497 25542 4543 25594
rect 4543 25542 4553 25594
rect 4577 25542 4607 25594
rect 4607 25542 4619 25594
rect 4619 25542 4633 25594
rect 4657 25542 4671 25594
rect 4671 25542 4683 25594
rect 4683 25542 4713 25594
rect 4737 25542 4747 25594
rect 4747 25542 4793 25594
rect 4497 25540 4553 25542
rect 4577 25540 4633 25542
rect 4657 25540 4713 25542
rect 4737 25540 4793 25542
rect 4497 24506 4553 24508
rect 4577 24506 4633 24508
rect 4657 24506 4713 24508
rect 4737 24506 4793 24508
rect 4497 24454 4543 24506
rect 4543 24454 4553 24506
rect 4577 24454 4607 24506
rect 4607 24454 4619 24506
rect 4619 24454 4633 24506
rect 4657 24454 4671 24506
rect 4671 24454 4683 24506
rect 4683 24454 4713 24506
rect 4737 24454 4747 24506
rect 4747 24454 4793 24506
rect 4497 24452 4553 24454
rect 4577 24452 4633 24454
rect 4657 24452 4713 24454
rect 4737 24452 4793 24454
rect 5157 25050 5213 25052
rect 5237 25050 5293 25052
rect 5317 25050 5373 25052
rect 5397 25050 5453 25052
rect 5157 24998 5203 25050
rect 5203 24998 5213 25050
rect 5237 24998 5267 25050
rect 5267 24998 5279 25050
rect 5279 24998 5293 25050
rect 5317 24998 5331 25050
rect 5331 24998 5343 25050
rect 5343 24998 5373 25050
rect 5397 24998 5407 25050
rect 5407 24998 5453 25050
rect 5157 24996 5213 24998
rect 5237 24996 5293 24998
rect 5317 24996 5373 24998
rect 5397 24996 5453 24998
rect 4497 23418 4553 23420
rect 4577 23418 4633 23420
rect 4657 23418 4713 23420
rect 4737 23418 4793 23420
rect 4497 23366 4543 23418
rect 4543 23366 4553 23418
rect 4577 23366 4607 23418
rect 4607 23366 4619 23418
rect 4619 23366 4633 23418
rect 4657 23366 4671 23418
rect 4671 23366 4683 23418
rect 4683 23366 4713 23418
rect 4737 23366 4747 23418
rect 4747 23366 4793 23418
rect 4497 23364 4553 23366
rect 4577 23364 4633 23366
rect 4657 23364 4713 23366
rect 4737 23364 4793 23366
rect 2226 11756 2282 11792
rect 2226 11736 2228 11756
rect 2228 11736 2280 11756
rect 2280 11736 2282 11756
rect 2134 10648 2190 10704
rect 3054 12280 3110 12336
rect 3146 11092 3148 11112
rect 3148 11092 3200 11112
rect 3200 11092 3202 11112
rect 3146 11056 3202 11092
rect 1490 6296 1546 6352
rect 2410 3984 2466 4040
rect 4497 22330 4553 22332
rect 4577 22330 4633 22332
rect 4657 22330 4713 22332
rect 4737 22330 4793 22332
rect 4497 22278 4543 22330
rect 4543 22278 4553 22330
rect 4577 22278 4607 22330
rect 4607 22278 4619 22330
rect 4619 22278 4633 22330
rect 4657 22278 4671 22330
rect 4671 22278 4683 22330
rect 4683 22278 4713 22330
rect 4737 22278 4747 22330
rect 4747 22278 4793 22330
rect 4497 22276 4553 22278
rect 4577 22276 4633 22278
rect 4657 22276 4713 22278
rect 4737 22276 4793 22278
rect 5157 23962 5213 23964
rect 5237 23962 5293 23964
rect 5317 23962 5373 23964
rect 5397 23962 5453 23964
rect 5157 23910 5203 23962
rect 5203 23910 5213 23962
rect 5237 23910 5267 23962
rect 5267 23910 5279 23962
rect 5279 23910 5293 23962
rect 5317 23910 5331 23962
rect 5331 23910 5343 23962
rect 5343 23910 5373 23962
rect 5397 23910 5407 23962
rect 5407 23910 5453 23962
rect 5157 23908 5213 23910
rect 5237 23908 5293 23910
rect 5317 23908 5373 23910
rect 5397 23908 5453 23910
rect 4710 21528 4766 21584
rect 4497 21242 4553 21244
rect 4577 21242 4633 21244
rect 4657 21242 4713 21244
rect 4737 21242 4793 21244
rect 4497 21190 4543 21242
rect 4543 21190 4553 21242
rect 4577 21190 4607 21242
rect 4607 21190 4619 21242
rect 4619 21190 4633 21242
rect 4657 21190 4671 21242
rect 4671 21190 4683 21242
rect 4683 21190 4713 21242
rect 4737 21190 4747 21242
rect 4747 21190 4793 21242
rect 4497 21188 4553 21190
rect 4577 21188 4633 21190
rect 4657 21188 4713 21190
rect 4737 21188 4793 21190
rect 4894 20340 4896 20360
rect 4896 20340 4948 20360
rect 4948 20340 4950 20360
rect 4894 20304 4950 20340
rect 4497 20154 4553 20156
rect 4577 20154 4633 20156
rect 4657 20154 4713 20156
rect 4737 20154 4793 20156
rect 4497 20102 4543 20154
rect 4543 20102 4553 20154
rect 4577 20102 4607 20154
rect 4607 20102 4619 20154
rect 4619 20102 4633 20154
rect 4657 20102 4671 20154
rect 4671 20102 4683 20154
rect 4683 20102 4713 20154
rect 4737 20102 4747 20154
rect 4747 20102 4793 20154
rect 4497 20100 4553 20102
rect 4577 20100 4633 20102
rect 4657 20100 4713 20102
rect 4737 20100 4793 20102
rect 4497 19066 4553 19068
rect 4577 19066 4633 19068
rect 4657 19066 4713 19068
rect 4737 19066 4793 19068
rect 4497 19014 4543 19066
rect 4543 19014 4553 19066
rect 4577 19014 4607 19066
rect 4607 19014 4619 19066
rect 4619 19014 4633 19066
rect 4657 19014 4671 19066
rect 4671 19014 4683 19066
rect 4683 19014 4713 19066
rect 4737 19014 4747 19066
rect 4747 19014 4793 19066
rect 4497 19012 4553 19014
rect 4577 19012 4633 19014
rect 4657 19012 4713 19014
rect 4737 19012 4793 19014
rect 4497 17978 4553 17980
rect 4577 17978 4633 17980
rect 4657 17978 4713 17980
rect 4737 17978 4793 17980
rect 4497 17926 4543 17978
rect 4543 17926 4553 17978
rect 4577 17926 4607 17978
rect 4607 17926 4619 17978
rect 4619 17926 4633 17978
rect 4657 17926 4671 17978
rect 4671 17926 4683 17978
rect 4683 17926 4713 17978
rect 4737 17926 4747 17978
rect 4747 17926 4793 17978
rect 4497 17924 4553 17926
rect 4577 17924 4633 17926
rect 4657 17924 4713 17926
rect 4737 17924 4793 17926
rect 4250 17720 4306 17776
rect 3698 11328 3754 11384
rect 3882 11212 3938 11248
rect 3882 11192 3884 11212
rect 3884 11192 3936 11212
rect 3936 11192 3938 11212
rect 4497 16890 4553 16892
rect 4577 16890 4633 16892
rect 4657 16890 4713 16892
rect 4737 16890 4793 16892
rect 4497 16838 4543 16890
rect 4543 16838 4553 16890
rect 4577 16838 4607 16890
rect 4607 16838 4619 16890
rect 4619 16838 4633 16890
rect 4657 16838 4671 16890
rect 4671 16838 4683 16890
rect 4683 16838 4713 16890
rect 4737 16838 4747 16890
rect 4747 16838 4793 16890
rect 4497 16836 4553 16838
rect 4577 16836 4633 16838
rect 4657 16836 4713 16838
rect 4737 16836 4793 16838
rect 5157 22874 5213 22876
rect 5237 22874 5293 22876
rect 5317 22874 5373 22876
rect 5397 22874 5453 22876
rect 5157 22822 5203 22874
rect 5203 22822 5213 22874
rect 5237 22822 5267 22874
rect 5267 22822 5279 22874
rect 5279 22822 5293 22874
rect 5317 22822 5331 22874
rect 5331 22822 5343 22874
rect 5343 22822 5373 22874
rect 5397 22822 5407 22874
rect 5407 22822 5453 22874
rect 5157 22820 5213 22822
rect 5237 22820 5293 22822
rect 5317 22820 5373 22822
rect 5397 22820 5453 22822
rect 5446 21936 5502 21992
rect 5157 21786 5213 21788
rect 5237 21786 5293 21788
rect 5317 21786 5373 21788
rect 5397 21786 5453 21788
rect 5157 21734 5203 21786
rect 5203 21734 5213 21786
rect 5237 21734 5267 21786
rect 5267 21734 5279 21786
rect 5279 21734 5293 21786
rect 5317 21734 5331 21786
rect 5331 21734 5343 21786
rect 5343 21734 5373 21786
rect 5397 21734 5407 21786
rect 5407 21734 5453 21786
rect 5157 21732 5213 21734
rect 5237 21732 5293 21734
rect 5317 21732 5373 21734
rect 5397 21732 5453 21734
rect 5630 21684 5686 21720
rect 5630 21664 5632 21684
rect 5632 21664 5684 21684
rect 5684 21664 5686 21684
rect 5157 20698 5213 20700
rect 5237 20698 5293 20700
rect 5317 20698 5373 20700
rect 5397 20698 5453 20700
rect 5157 20646 5203 20698
rect 5203 20646 5213 20698
rect 5237 20646 5267 20698
rect 5267 20646 5279 20698
rect 5279 20646 5293 20698
rect 5317 20646 5331 20698
rect 5331 20646 5343 20698
rect 5343 20646 5373 20698
rect 5397 20646 5407 20698
rect 5407 20646 5453 20698
rect 5157 20644 5213 20646
rect 5237 20644 5293 20646
rect 5317 20644 5373 20646
rect 5397 20644 5453 20646
rect 5157 19610 5213 19612
rect 5237 19610 5293 19612
rect 5317 19610 5373 19612
rect 5397 19610 5453 19612
rect 5157 19558 5203 19610
rect 5203 19558 5213 19610
rect 5237 19558 5267 19610
rect 5267 19558 5279 19610
rect 5279 19558 5293 19610
rect 5317 19558 5331 19610
rect 5331 19558 5343 19610
rect 5343 19558 5373 19610
rect 5397 19558 5407 19610
rect 5407 19558 5453 19610
rect 5157 19556 5213 19558
rect 5237 19556 5293 19558
rect 5317 19556 5373 19558
rect 5397 19556 5453 19558
rect 5157 18522 5213 18524
rect 5237 18522 5293 18524
rect 5317 18522 5373 18524
rect 5397 18522 5453 18524
rect 5157 18470 5203 18522
rect 5203 18470 5213 18522
rect 5237 18470 5267 18522
rect 5267 18470 5279 18522
rect 5279 18470 5293 18522
rect 5317 18470 5331 18522
rect 5331 18470 5343 18522
rect 5343 18470 5373 18522
rect 5397 18470 5407 18522
rect 5407 18470 5453 18522
rect 5157 18468 5213 18470
rect 5237 18468 5293 18470
rect 5317 18468 5373 18470
rect 5397 18468 5453 18470
rect 5157 17434 5213 17436
rect 5237 17434 5293 17436
rect 5317 17434 5373 17436
rect 5397 17434 5453 17436
rect 5157 17382 5203 17434
rect 5203 17382 5213 17434
rect 5237 17382 5267 17434
rect 5267 17382 5279 17434
rect 5279 17382 5293 17434
rect 5317 17382 5331 17434
rect 5331 17382 5343 17434
rect 5343 17382 5373 17434
rect 5397 17382 5407 17434
rect 5407 17382 5453 17434
rect 5157 17380 5213 17382
rect 5237 17380 5293 17382
rect 5317 17380 5373 17382
rect 5397 17380 5453 17382
rect 4497 15802 4553 15804
rect 4577 15802 4633 15804
rect 4657 15802 4713 15804
rect 4737 15802 4793 15804
rect 4497 15750 4543 15802
rect 4543 15750 4553 15802
rect 4577 15750 4607 15802
rect 4607 15750 4619 15802
rect 4619 15750 4633 15802
rect 4657 15750 4671 15802
rect 4671 15750 4683 15802
rect 4683 15750 4713 15802
rect 4737 15750 4747 15802
rect 4747 15750 4793 15802
rect 4497 15748 4553 15750
rect 4577 15748 4633 15750
rect 4657 15748 4713 15750
rect 4737 15748 4793 15750
rect 4497 14714 4553 14716
rect 4577 14714 4633 14716
rect 4657 14714 4713 14716
rect 4737 14714 4793 14716
rect 4497 14662 4543 14714
rect 4543 14662 4553 14714
rect 4577 14662 4607 14714
rect 4607 14662 4619 14714
rect 4619 14662 4633 14714
rect 4657 14662 4671 14714
rect 4671 14662 4683 14714
rect 4683 14662 4713 14714
rect 4737 14662 4747 14714
rect 4747 14662 4793 14714
rect 4497 14660 4553 14662
rect 4577 14660 4633 14662
rect 4657 14660 4713 14662
rect 4737 14660 4793 14662
rect 4497 13626 4553 13628
rect 4577 13626 4633 13628
rect 4657 13626 4713 13628
rect 4737 13626 4793 13628
rect 4497 13574 4543 13626
rect 4543 13574 4553 13626
rect 4577 13574 4607 13626
rect 4607 13574 4619 13626
rect 4619 13574 4633 13626
rect 4657 13574 4671 13626
rect 4671 13574 4683 13626
rect 4683 13574 4713 13626
rect 4737 13574 4747 13626
rect 4747 13574 4793 13626
rect 4497 13572 4553 13574
rect 4577 13572 4633 13574
rect 4657 13572 4713 13574
rect 4737 13572 4793 13574
rect 4066 10804 4122 10840
rect 5157 16346 5213 16348
rect 5237 16346 5293 16348
rect 5317 16346 5373 16348
rect 5397 16346 5453 16348
rect 5157 16294 5203 16346
rect 5203 16294 5213 16346
rect 5237 16294 5267 16346
rect 5267 16294 5279 16346
rect 5279 16294 5293 16346
rect 5317 16294 5331 16346
rect 5331 16294 5343 16346
rect 5343 16294 5373 16346
rect 5397 16294 5407 16346
rect 5407 16294 5453 16346
rect 5157 16292 5213 16294
rect 5237 16292 5293 16294
rect 5317 16292 5373 16294
rect 5397 16292 5453 16294
rect 5157 15258 5213 15260
rect 5237 15258 5293 15260
rect 5317 15258 5373 15260
rect 5397 15258 5453 15260
rect 5157 15206 5203 15258
rect 5203 15206 5213 15258
rect 5237 15206 5267 15258
rect 5267 15206 5279 15258
rect 5279 15206 5293 15258
rect 5317 15206 5331 15258
rect 5331 15206 5343 15258
rect 5343 15206 5373 15258
rect 5397 15206 5407 15258
rect 5407 15206 5453 15258
rect 5157 15204 5213 15206
rect 5237 15204 5293 15206
rect 5317 15204 5373 15206
rect 5397 15204 5453 15206
rect 7102 28464 7158 28520
rect 8758 28484 8814 28520
rect 8758 28464 8760 28484
rect 8760 28464 8812 28484
rect 8812 28464 8814 28484
rect 6918 22072 6974 22128
rect 6918 21936 6974 21992
rect 7194 21528 7250 21584
rect 5157 14170 5213 14172
rect 5237 14170 5293 14172
rect 5317 14170 5373 14172
rect 5397 14170 5453 14172
rect 5157 14118 5203 14170
rect 5203 14118 5213 14170
rect 5237 14118 5267 14170
rect 5267 14118 5279 14170
rect 5279 14118 5293 14170
rect 5317 14118 5331 14170
rect 5331 14118 5343 14170
rect 5343 14118 5373 14170
rect 5397 14118 5407 14170
rect 5407 14118 5453 14170
rect 5157 14116 5213 14118
rect 5237 14116 5293 14118
rect 5317 14116 5373 14118
rect 5397 14116 5453 14118
rect 5157 13082 5213 13084
rect 5237 13082 5293 13084
rect 5317 13082 5373 13084
rect 5397 13082 5453 13084
rect 5157 13030 5203 13082
rect 5203 13030 5213 13082
rect 5237 13030 5267 13082
rect 5267 13030 5279 13082
rect 5279 13030 5293 13082
rect 5317 13030 5331 13082
rect 5331 13030 5343 13082
rect 5343 13030 5373 13082
rect 5397 13030 5407 13082
rect 5407 13030 5453 13082
rect 5157 13028 5213 13030
rect 5237 13028 5293 13030
rect 5317 13028 5373 13030
rect 5397 13028 5453 13030
rect 4497 12538 4553 12540
rect 4577 12538 4633 12540
rect 4657 12538 4713 12540
rect 4737 12538 4793 12540
rect 4497 12486 4543 12538
rect 4543 12486 4553 12538
rect 4577 12486 4607 12538
rect 4607 12486 4619 12538
rect 4619 12486 4633 12538
rect 4657 12486 4671 12538
rect 4671 12486 4683 12538
rect 4683 12486 4713 12538
rect 4737 12486 4747 12538
rect 4747 12486 4793 12538
rect 4497 12484 4553 12486
rect 4577 12484 4633 12486
rect 4657 12484 4713 12486
rect 4737 12484 4793 12486
rect 4250 11328 4306 11384
rect 4497 11450 4553 11452
rect 4577 11450 4633 11452
rect 4657 11450 4713 11452
rect 4737 11450 4793 11452
rect 4497 11398 4543 11450
rect 4543 11398 4553 11450
rect 4577 11398 4607 11450
rect 4607 11398 4619 11450
rect 4619 11398 4633 11450
rect 4657 11398 4671 11450
rect 4671 11398 4683 11450
rect 4683 11398 4713 11450
rect 4737 11398 4747 11450
rect 4747 11398 4793 11450
rect 4497 11396 4553 11398
rect 4577 11396 4633 11398
rect 4657 11396 4713 11398
rect 4737 11396 4793 11398
rect 4894 11192 4950 11248
rect 4066 10784 4068 10804
rect 4068 10784 4120 10804
rect 4120 10784 4122 10804
rect 4250 10512 4306 10568
rect 8390 21664 8446 21720
rect 7378 17720 7434 17776
rect 7102 17604 7158 17640
rect 7102 17584 7104 17604
rect 7104 17584 7156 17604
rect 7156 17584 7158 17604
rect 5157 11994 5213 11996
rect 5237 11994 5293 11996
rect 5317 11994 5373 11996
rect 5397 11994 5453 11996
rect 5157 11942 5203 11994
rect 5203 11942 5213 11994
rect 5237 11942 5267 11994
rect 5267 11942 5279 11994
rect 5279 11942 5293 11994
rect 5317 11942 5331 11994
rect 5331 11942 5343 11994
rect 5343 11942 5373 11994
rect 5397 11942 5407 11994
rect 5407 11942 5453 11994
rect 5157 11940 5213 11942
rect 5237 11940 5293 11942
rect 5317 11940 5373 11942
rect 5397 11940 5453 11942
rect 5157 10906 5213 10908
rect 5237 10906 5293 10908
rect 5317 10906 5373 10908
rect 5397 10906 5453 10908
rect 5157 10854 5203 10906
rect 5203 10854 5213 10906
rect 5237 10854 5267 10906
rect 5267 10854 5279 10906
rect 5279 10854 5293 10906
rect 5317 10854 5331 10906
rect 5331 10854 5343 10906
rect 5343 10854 5373 10906
rect 5397 10854 5407 10906
rect 5407 10854 5453 10906
rect 5157 10852 5213 10854
rect 5237 10852 5293 10854
rect 5317 10852 5373 10854
rect 5397 10852 5453 10854
rect 4986 10784 5042 10840
rect 4618 10512 4674 10568
rect 5262 10684 5264 10704
rect 5264 10684 5316 10704
rect 5316 10684 5318 10704
rect 5262 10648 5318 10684
rect 4497 10362 4553 10364
rect 4577 10362 4633 10364
rect 4657 10362 4713 10364
rect 4737 10362 4793 10364
rect 4497 10310 4543 10362
rect 4543 10310 4553 10362
rect 4577 10310 4607 10362
rect 4607 10310 4619 10362
rect 4619 10310 4633 10362
rect 4657 10310 4671 10362
rect 4671 10310 4683 10362
rect 4683 10310 4713 10362
rect 4737 10310 4747 10362
rect 4747 10310 4793 10362
rect 4497 10308 4553 10310
rect 4577 10308 4633 10310
rect 4657 10308 4713 10310
rect 4737 10308 4793 10310
rect 4497 9274 4553 9276
rect 4577 9274 4633 9276
rect 4657 9274 4713 9276
rect 4737 9274 4793 9276
rect 4497 9222 4543 9274
rect 4543 9222 4553 9274
rect 4577 9222 4607 9274
rect 4607 9222 4619 9274
rect 4619 9222 4633 9274
rect 4657 9222 4671 9274
rect 4671 9222 4683 9274
rect 4683 9222 4713 9274
rect 4737 9222 4747 9274
rect 4747 9222 4793 9274
rect 4497 9220 4553 9222
rect 4577 9220 4633 9222
rect 4657 9220 4713 9222
rect 4737 9220 4793 9222
rect 5157 9818 5213 9820
rect 5237 9818 5293 9820
rect 5317 9818 5373 9820
rect 5397 9818 5453 9820
rect 5157 9766 5203 9818
rect 5203 9766 5213 9818
rect 5237 9766 5267 9818
rect 5267 9766 5279 9818
rect 5279 9766 5293 9818
rect 5317 9766 5331 9818
rect 5331 9766 5343 9818
rect 5343 9766 5373 9818
rect 5397 9766 5407 9818
rect 5407 9766 5453 9818
rect 5157 9764 5213 9766
rect 5237 9764 5293 9766
rect 5317 9764 5373 9766
rect 5397 9764 5453 9766
rect 5446 9580 5502 9616
rect 5446 9560 5448 9580
rect 5448 9560 5500 9580
rect 5500 9560 5502 9580
rect 4497 8186 4553 8188
rect 4577 8186 4633 8188
rect 4657 8186 4713 8188
rect 4737 8186 4793 8188
rect 4497 8134 4543 8186
rect 4543 8134 4553 8186
rect 4577 8134 4607 8186
rect 4607 8134 4619 8186
rect 4619 8134 4633 8186
rect 4657 8134 4671 8186
rect 4671 8134 4683 8186
rect 4683 8134 4713 8186
rect 4737 8134 4747 8186
rect 4747 8134 4793 8186
rect 4497 8132 4553 8134
rect 4577 8132 4633 8134
rect 4657 8132 4713 8134
rect 4737 8132 4793 8134
rect 5157 8730 5213 8732
rect 5237 8730 5293 8732
rect 5317 8730 5373 8732
rect 5397 8730 5453 8732
rect 5157 8678 5203 8730
rect 5203 8678 5213 8730
rect 5237 8678 5267 8730
rect 5267 8678 5279 8730
rect 5279 8678 5293 8730
rect 5317 8678 5331 8730
rect 5331 8678 5343 8730
rect 5343 8678 5373 8730
rect 5397 8678 5407 8730
rect 5407 8678 5453 8730
rect 5157 8676 5213 8678
rect 5237 8676 5293 8678
rect 5317 8676 5373 8678
rect 5397 8676 5453 8678
rect 5446 8492 5502 8528
rect 5446 8472 5448 8492
rect 5448 8472 5500 8492
rect 5500 8472 5502 8492
rect 4066 7520 4122 7576
rect 4497 7098 4553 7100
rect 4577 7098 4633 7100
rect 4657 7098 4713 7100
rect 4737 7098 4793 7100
rect 4497 7046 4543 7098
rect 4543 7046 4553 7098
rect 4577 7046 4607 7098
rect 4607 7046 4619 7098
rect 4619 7046 4633 7098
rect 4657 7046 4671 7098
rect 4671 7046 4683 7098
rect 4683 7046 4713 7098
rect 4737 7046 4747 7098
rect 4747 7046 4793 7098
rect 4497 7044 4553 7046
rect 4577 7044 4633 7046
rect 4657 7044 4713 7046
rect 4737 7044 4793 7046
rect 5157 7642 5213 7644
rect 5237 7642 5293 7644
rect 5317 7642 5373 7644
rect 5397 7642 5453 7644
rect 5157 7590 5203 7642
rect 5203 7590 5213 7642
rect 5237 7590 5267 7642
rect 5267 7590 5279 7642
rect 5279 7590 5293 7642
rect 5317 7590 5331 7642
rect 5331 7590 5343 7642
rect 5343 7590 5373 7642
rect 5397 7590 5407 7642
rect 5407 7590 5453 7642
rect 5157 7588 5213 7590
rect 5237 7588 5293 7590
rect 5317 7588 5373 7590
rect 5397 7588 5453 7590
rect 5157 6554 5213 6556
rect 5237 6554 5293 6556
rect 5317 6554 5373 6556
rect 5397 6554 5453 6556
rect 5157 6502 5203 6554
rect 5203 6502 5213 6554
rect 5237 6502 5267 6554
rect 5267 6502 5279 6554
rect 5279 6502 5293 6554
rect 5317 6502 5331 6554
rect 5331 6502 5343 6554
rect 5343 6502 5373 6554
rect 5397 6502 5407 6554
rect 5407 6502 5453 6554
rect 5157 6500 5213 6502
rect 5237 6500 5293 6502
rect 5317 6500 5373 6502
rect 5397 6500 5453 6502
rect 6182 11076 6238 11112
rect 6182 11056 6184 11076
rect 6184 11056 6236 11076
rect 6236 11056 6238 11076
rect 4497 6010 4553 6012
rect 4577 6010 4633 6012
rect 4657 6010 4713 6012
rect 4737 6010 4793 6012
rect 4497 5958 4543 6010
rect 4543 5958 4553 6010
rect 4577 5958 4607 6010
rect 4607 5958 4619 6010
rect 4619 5958 4633 6010
rect 4657 5958 4671 6010
rect 4671 5958 4683 6010
rect 4683 5958 4713 6010
rect 4737 5958 4747 6010
rect 4747 5958 4793 6010
rect 4497 5956 4553 5958
rect 4577 5956 4633 5958
rect 4657 5956 4713 5958
rect 4737 5956 4793 5958
rect 5157 5466 5213 5468
rect 5237 5466 5293 5468
rect 5317 5466 5373 5468
rect 5397 5466 5453 5468
rect 5157 5414 5203 5466
rect 5203 5414 5213 5466
rect 5237 5414 5267 5466
rect 5267 5414 5279 5466
rect 5279 5414 5293 5466
rect 5317 5414 5331 5466
rect 5331 5414 5343 5466
rect 5343 5414 5373 5466
rect 5397 5414 5407 5466
rect 5407 5414 5453 5466
rect 5157 5412 5213 5414
rect 5237 5412 5293 5414
rect 5317 5412 5373 5414
rect 5397 5412 5453 5414
rect 4497 4922 4553 4924
rect 4577 4922 4633 4924
rect 4657 4922 4713 4924
rect 4737 4922 4793 4924
rect 4497 4870 4543 4922
rect 4543 4870 4553 4922
rect 4577 4870 4607 4922
rect 4607 4870 4619 4922
rect 4619 4870 4633 4922
rect 4657 4870 4671 4922
rect 4671 4870 4683 4922
rect 4683 4870 4713 4922
rect 4737 4870 4747 4922
rect 4747 4870 4793 4922
rect 4497 4868 4553 4870
rect 4577 4868 4633 4870
rect 4657 4868 4713 4870
rect 4737 4868 4793 4870
rect 11580 29946 11636 29948
rect 11660 29946 11716 29948
rect 11740 29946 11796 29948
rect 11820 29946 11876 29948
rect 11580 29894 11626 29946
rect 11626 29894 11636 29946
rect 11660 29894 11690 29946
rect 11690 29894 11702 29946
rect 11702 29894 11716 29946
rect 11740 29894 11754 29946
rect 11754 29894 11766 29946
rect 11766 29894 11796 29946
rect 11820 29894 11830 29946
rect 11830 29894 11876 29946
rect 11580 29892 11636 29894
rect 11660 29892 11716 29894
rect 11740 29892 11796 29894
rect 11820 29892 11876 29894
rect 11058 28056 11114 28112
rect 12240 29402 12296 29404
rect 12320 29402 12376 29404
rect 12400 29402 12456 29404
rect 12480 29402 12536 29404
rect 12240 29350 12286 29402
rect 12286 29350 12296 29402
rect 12320 29350 12350 29402
rect 12350 29350 12362 29402
rect 12362 29350 12376 29402
rect 12400 29350 12414 29402
rect 12414 29350 12426 29402
rect 12426 29350 12456 29402
rect 12480 29350 12490 29402
rect 12490 29350 12536 29402
rect 12240 29348 12296 29350
rect 12320 29348 12376 29350
rect 12400 29348 12456 29350
rect 12480 29348 12536 29350
rect 11580 28858 11636 28860
rect 11660 28858 11716 28860
rect 11740 28858 11796 28860
rect 11820 28858 11876 28860
rect 11580 28806 11626 28858
rect 11626 28806 11636 28858
rect 11660 28806 11690 28858
rect 11690 28806 11702 28858
rect 11702 28806 11716 28858
rect 11740 28806 11754 28858
rect 11754 28806 11766 28858
rect 11766 28806 11796 28858
rect 11820 28806 11830 28858
rect 11830 28806 11876 28858
rect 11580 28804 11636 28806
rect 11660 28804 11716 28806
rect 11740 28804 11796 28806
rect 11820 28804 11876 28806
rect 12070 28056 12126 28112
rect 11580 27770 11636 27772
rect 11660 27770 11716 27772
rect 11740 27770 11796 27772
rect 11820 27770 11876 27772
rect 11580 27718 11626 27770
rect 11626 27718 11636 27770
rect 11660 27718 11690 27770
rect 11690 27718 11702 27770
rect 11702 27718 11716 27770
rect 11740 27718 11754 27770
rect 11754 27718 11766 27770
rect 11766 27718 11796 27770
rect 11820 27718 11830 27770
rect 11830 27718 11876 27770
rect 11580 27716 11636 27718
rect 11660 27716 11716 27718
rect 11740 27716 11796 27718
rect 11820 27716 11876 27718
rect 12070 27920 12126 27976
rect 12240 28314 12296 28316
rect 12320 28314 12376 28316
rect 12400 28314 12456 28316
rect 12480 28314 12536 28316
rect 12240 28262 12286 28314
rect 12286 28262 12296 28314
rect 12320 28262 12350 28314
rect 12350 28262 12362 28314
rect 12362 28262 12376 28314
rect 12400 28262 12414 28314
rect 12414 28262 12426 28314
rect 12426 28262 12456 28314
rect 12480 28262 12490 28314
rect 12490 28262 12536 28314
rect 12240 28260 12296 28262
rect 12320 28260 12376 28262
rect 12400 28260 12456 28262
rect 12480 28260 12536 28262
rect 13634 28620 13690 28656
rect 13634 28600 13636 28620
rect 13636 28600 13688 28620
rect 13688 28600 13690 28620
rect 11580 26682 11636 26684
rect 11660 26682 11716 26684
rect 11740 26682 11796 26684
rect 11820 26682 11876 26684
rect 11580 26630 11626 26682
rect 11626 26630 11636 26682
rect 11660 26630 11690 26682
rect 11690 26630 11702 26682
rect 11702 26630 11716 26682
rect 11740 26630 11754 26682
rect 11754 26630 11766 26682
rect 11766 26630 11796 26682
rect 11820 26630 11830 26682
rect 11830 26630 11876 26682
rect 11580 26628 11636 26630
rect 11660 26628 11716 26630
rect 11740 26628 11796 26630
rect 11820 26628 11876 26630
rect 12240 27226 12296 27228
rect 12320 27226 12376 27228
rect 12400 27226 12456 27228
rect 12480 27226 12536 27228
rect 12240 27174 12286 27226
rect 12286 27174 12296 27226
rect 12320 27174 12350 27226
rect 12350 27174 12362 27226
rect 12362 27174 12376 27226
rect 12400 27174 12414 27226
rect 12414 27174 12426 27226
rect 12426 27174 12456 27226
rect 12480 27174 12490 27226
rect 12490 27174 12536 27226
rect 12240 27172 12296 27174
rect 12320 27172 12376 27174
rect 12400 27172 12456 27174
rect 12480 27172 12536 27174
rect 12240 26138 12296 26140
rect 12320 26138 12376 26140
rect 12400 26138 12456 26140
rect 12480 26138 12536 26140
rect 12240 26086 12286 26138
rect 12286 26086 12296 26138
rect 12320 26086 12350 26138
rect 12350 26086 12362 26138
rect 12362 26086 12376 26138
rect 12400 26086 12414 26138
rect 12414 26086 12426 26138
rect 12426 26086 12456 26138
rect 12480 26086 12490 26138
rect 12490 26086 12536 26138
rect 12240 26084 12296 26086
rect 12320 26084 12376 26086
rect 12400 26084 12456 26086
rect 12480 26084 12536 26086
rect 11580 25594 11636 25596
rect 11660 25594 11716 25596
rect 11740 25594 11796 25596
rect 11820 25594 11876 25596
rect 11580 25542 11626 25594
rect 11626 25542 11636 25594
rect 11660 25542 11690 25594
rect 11690 25542 11702 25594
rect 11702 25542 11716 25594
rect 11740 25542 11754 25594
rect 11754 25542 11766 25594
rect 11766 25542 11796 25594
rect 11820 25542 11830 25594
rect 11830 25542 11876 25594
rect 11580 25540 11636 25542
rect 11660 25540 11716 25542
rect 11740 25540 11796 25542
rect 11820 25540 11876 25542
rect 13634 28192 13690 28248
rect 13542 27920 13598 27976
rect 12240 25050 12296 25052
rect 12320 25050 12376 25052
rect 12400 25050 12456 25052
rect 12480 25050 12536 25052
rect 12240 24998 12286 25050
rect 12286 24998 12296 25050
rect 12320 24998 12350 25050
rect 12350 24998 12362 25050
rect 12362 24998 12376 25050
rect 12400 24998 12414 25050
rect 12414 24998 12426 25050
rect 12426 24998 12456 25050
rect 12480 24998 12490 25050
rect 12490 24998 12536 25050
rect 12240 24996 12296 24998
rect 12320 24996 12376 24998
rect 12400 24996 12456 24998
rect 12480 24996 12536 24998
rect 9862 21936 9918 21992
rect 9862 20304 9918 20360
rect 7562 11192 7618 11248
rect 10322 20304 10378 20360
rect 10690 22072 10746 22128
rect 11580 24506 11636 24508
rect 11660 24506 11716 24508
rect 11740 24506 11796 24508
rect 11820 24506 11876 24508
rect 11580 24454 11626 24506
rect 11626 24454 11636 24506
rect 11660 24454 11690 24506
rect 11690 24454 11702 24506
rect 11702 24454 11716 24506
rect 11740 24454 11754 24506
rect 11754 24454 11766 24506
rect 11766 24454 11796 24506
rect 11820 24454 11830 24506
rect 11830 24454 11876 24506
rect 11580 24452 11636 24454
rect 11660 24452 11716 24454
rect 11740 24452 11796 24454
rect 11820 24452 11876 24454
rect 12240 23962 12296 23964
rect 12320 23962 12376 23964
rect 12400 23962 12456 23964
rect 12480 23962 12536 23964
rect 12240 23910 12286 23962
rect 12286 23910 12296 23962
rect 12320 23910 12350 23962
rect 12350 23910 12362 23962
rect 12362 23910 12376 23962
rect 12400 23910 12414 23962
rect 12414 23910 12426 23962
rect 12426 23910 12456 23962
rect 12480 23910 12490 23962
rect 12490 23910 12536 23962
rect 12240 23908 12296 23910
rect 12320 23908 12376 23910
rect 12400 23908 12456 23910
rect 12480 23908 12536 23910
rect 11580 23418 11636 23420
rect 11660 23418 11716 23420
rect 11740 23418 11796 23420
rect 11820 23418 11876 23420
rect 11580 23366 11626 23418
rect 11626 23366 11636 23418
rect 11660 23366 11690 23418
rect 11690 23366 11702 23418
rect 11702 23366 11716 23418
rect 11740 23366 11754 23418
rect 11754 23366 11766 23418
rect 11766 23366 11796 23418
rect 11820 23366 11830 23418
rect 11830 23366 11876 23418
rect 11580 23364 11636 23366
rect 11660 23364 11716 23366
rect 11740 23364 11796 23366
rect 11820 23364 11876 23366
rect 12240 22874 12296 22876
rect 12320 22874 12376 22876
rect 12400 22874 12456 22876
rect 12480 22874 12536 22876
rect 12240 22822 12286 22874
rect 12286 22822 12296 22874
rect 12320 22822 12350 22874
rect 12350 22822 12362 22874
rect 12362 22822 12376 22874
rect 12400 22822 12414 22874
rect 12414 22822 12426 22874
rect 12426 22822 12456 22874
rect 12480 22822 12490 22874
rect 12490 22822 12536 22874
rect 12240 22820 12296 22822
rect 12320 22820 12376 22822
rect 12400 22820 12456 22822
rect 12480 22820 12536 22822
rect 11580 22330 11636 22332
rect 11660 22330 11716 22332
rect 11740 22330 11796 22332
rect 11820 22330 11876 22332
rect 11580 22278 11626 22330
rect 11626 22278 11636 22330
rect 11660 22278 11690 22330
rect 11690 22278 11702 22330
rect 11702 22278 11716 22330
rect 11740 22278 11754 22330
rect 11754 22278 11766 22330
rect 11766 22278 11796 22330
rect 11820 22278 11830 22330
rect 11830 22278 11876 22330
rect 11580 22276 11636 22278
rect 11660 22276 11716 22278
rect 11740 22276 11796 22278
rect 11820 22276 11876 22278
rect 11580 21242 11636 21244
rect 11660 21242 11716 21244
rect 11740 21242 11796 21244
rect 11820 21242 11876 21244
rect 11580 21190 11626 21242
rect 11626 21190 11636 21242
rect 11660 21190 11690 21242
rect 11690 21190 11702 21242
rect 11702 21190 11716 21242
rect 11740 21190 11754 21242
rect 11754 21190 11766 21242
rect 11766 21190 11796 21242
rect 11820 21190 11830 21242
rect 11830 21190 11876 21242
rect 11580 21188 11636 21190
rect 11660 21188 11716 21190
rect 11740 21188 11796 21190
rect 11820 21188 11876 21190
rect 10506 19916 10562 19952
rect 10506 19896 10508 19916
rect 10508 19896 10560 19916
rect 10560 19896 10562 19916
rect 10966 19760 11022 19816
rect 10506 15564 10562 15600
rect 10506 15544 10508 15564
rect 10508 15544 10560 15564
rect 10560 15544 10562 15564
rect 10506 14492 10508 14512
rect 10508 14492 10560 14512
rect 10560 14492 10562 14512
rect 10506 14456 10562 14492
rect 10230 13368 10286 13424
rect 10506 13776 10562 13832
rect 12240 21786 12296 21788
rect 12320 21786 12376 21788
rect 12400 21786 12456 21788
rect 12480 21786 12536 21788
rect 12240 21734 12286 21786
rect 12286 21734 12296 21786
rect 12320 21734 12350 21786
rect 12350 21734 12362 21786
rect 12362 21734 12376 21786
rect 12400 21734 12414 21786
rect 12414 21734 12426 21786
rect 12426 21734 12456 21786
rect 12480 21734 12490 21786
rect 12490 21734 12536 21786
rect 12240 21732 12296 21734
rect 12320 21732 12376 21734
rect 12400 21732 12456 21734
rect 12480 21732 12536 21734
rect 11580 20154 11636 20156
rect 11660 20154 11716 20156
rect 11740 20154 11796 20156
rect 11820 20154 11876 20156
rect 11580 20102 11626 20154
rect 11626 20102 11636 20154
rect 11660 20102 11690 20154
rect 11690 20102 11702 20154
rect 11702 20102 11716 20154
rect 11740 20102 11754 20154
rect 11754 20102 11766 20154
rect 11766 20102 11796 20154
rect 11820 20102 11830 20154
rect 11830 20102 11876 20154
rect 11580 20100 11636 20102
rect 11660 20100 11716 20102
rect 11740 20100 11796 20102
rect 11820 20100 11876 20102
rect 11580 19066 11636 19068
rect 11660 19066 11716 19068
rect 11740 19066 11796 19068
rect 11820 19066 11876 19068
rect 11580 19014 11626 19066
rect 11626 19014 11636 19066
rect 11660 19014 11690 19066
rect 11690 19014 11702 19066
rect 11702 19014 11716 19066
rect 11740 19014 11754 19066
rect 11754 19014 11766 19066
rect 11766 19014 11796 19066
rect 11820 19014 11830 19066
rect 11830 19014 11876 19066
rect 11580 19012 11636 19014
rect 11660 19012 11716 19014
rect 11740 19012 11796 19014
rect 11820 19012 11876 19014
rect 11580 17978 11636 17980
rect 11660 17978 11716 17980
rect 11740 17978 11796 17980
rect 11820 17978 11876 17980
rect 11580 17926 11626 17978
rect 11626 17926 11636 17978
rect 11660 17926 11690 17978
rect 11690 17926 11702 17978
rect 11702 17926 11716 17978
rect 11740 17926 11754 17978
rect 11754 17926 11766 17978
rect 11766 17926 11796 17978
rect 11820 17926 11830 17978
rect 11830 17926 11876 17978
rect 11580 17924 11636 17926
rect 11660 17924 11716 17926
rect 11740 17924 11796 17926
rect 11820 17924 11876 17926
rect 12240 20698 12296 20700
rect 12320 20698 12376 20700
rect 12400 20698 12456 20700
rect 12480 20698 12536 20700
rect 12240 20646 12286 20698
rect 12286 20646 12296 20698
rect 12320 20646 12350 20698
rect 12350 20646 12362 20698
rect 12362 20646 12376 20698
rect 12400 20646 12414 20698
rect 12414 20646 12426 20698
rect 12426 20646 12456 20698
rect 12480 20646 12490 20698
rect 12490 20646 12536 20698
rect 12240 20644 12296 20646
rect 12320 20644 12376 20646
rect 12400 20644 12456 20646
rect 12480 20644 12536 20646
rect 19323 30490 19379 30492
rect 19403 30490 19459 30492
rect 19483 30490 19539 30492
rect 19563 30490 19619 30492
rect 19323 30438 19369 30490
rect 19369 30438 19379 30490
rect 19403 30438 19433 30490
rect 19433 30438 19445 30490
rect 19445 30438 19459 30490
rect 19483 30438 19497 30490
rect 19497 30438 19509 30490
rect 19509 30438 19539 30490
rect 19563 30438 19573 30490
rect 19573 30438 19619 30490
rect 19323 30436 19379 30438
rect 19403 30436 19459 30438
rect 19483 30436 19539 30438
rect 19563 30436 19619 30438
rect 28906 30640 28962 30696
rect 26406 30490 26462 30492
rect 26486 30490 26542 30492
rect 26566 30490 26622 30492
rect 26646 30490 26702 30492
rect 26406 30438 26452 30490
rect 26452 30438 26462 30490
rect 26486 30438 26516 30490
rect 26516 30438 26528 30490
rect 26528 30438 26542 30490
rect 26566 30438 26580 30490
rect 26580 30438 26592 30490
rect 26592 30438 26622 30490
rect 26646 30438 26656 30490
rect 26656 30438 26702 30490
rect 26406 30436 26462 30438
rect 26486 30436 26542 30438
rect 26566 30436 26622 30438
rect 26646 30436 26702 30438
rect 12714 20440 12770 20496
rect 12240 19610 12296 19612
rect 12320 19610 12376 19612
rect 12400 19610 12456 19612
rect 12480 19610 12536 19612
rect 12240 19558 12286 19610
rect 12286 19558 12296 19610
rect 12320 19558 12350 19610
rect 12350 19558 12362 19610
rect 12362 19558 12376 19610
rect 12400 19558 12414 19610
rect 12414 19558 12426 19610
rect 12426 19558 12456 19610
rect 12480 19558 12490 19610
rect 12490 19558 12536 19610
rect 12240 19556 12296 19558
rect 12320 19556 12376 19558
rect 12400 19556 12456 19558
rect 12480 19556 12536 19558
rect 13174 19796 13176 19816
rect 13176 19796 13228 19816
rect 13228 19796 13230 19816
rect 13174 19760 13230 19796
rect 12240 18522 12296 18524
rect 12320 18522 12376 18524
rect 12400 18522 12456 18524
rect 12480 18522 12536 18524
rect 12240 18470 12286 18522
rect 12286 18470 12296 18522
rect 12320 18470 12350 18522
rect 12350 18470 12362 18522
rect 12362 18470 12376 18522
rect 12400 18470 12414 18522
rect 12414 18470 12426 18522
rect 12426 18470 12456 18522
rect 12480 18470 12490 18522
rect 12490 18470 12536 18522
rect 12240 18468 12296 18470
rect 12320 18468 12376 18470
rect 12400 18468 12456 18470
rect 12480 18468 12536 18470
rect 7010 6704 7066 6760
rect 8850 9460 8852 9480
rect 8852 9460 8904 9480
rect 8904 9460 8906 9480
rect 8850 9424 8906 9460
rect 8298 6740 8300 6760
rect 8300 6740 8352 6760
rect 8352 6740 8354 6760
rect 8298 6704 8354 6740
rect 9034 8508 9036 8528
rect 9036 8508 9088 8528
rect 9088 8508 9090 8528
rect 9034 8472 9090 8508
rect 9954 9832 10010 9888
rect 11580 16890 11636 16892
rect 11660 16890 11716 16892
rect 11740 16890 11796 16892
rect 11820 16890 11876 16892
rect 11580 16838 11626 16890
rect 11626 16838 11636 16890
rect 11660 16838 11690 16890
rect 11690 16838 11702 16890
rect 11702 16838 11716 16890
rect 11740 16838 11754 16890
rect 11754 16838 11766 16890
rect 11766 16838 11796 16890
rect 11820 16838 11830 16890
rect 11830 16838 11876 16890
rect 11580 16836 11636 16838
rect 11660 16836 11716 16838
rect 11740 16836 11796 16838
rect 11820 16836 11876 16838
rect 11580 15802 11636 15804
rect 11660 15802 11716 15804
rect 11740 15802 11796 15804
rect 11820 15802 11876 15804
rect 11580 15750 11626 15802
rect 11626 15750 11636 15802
rect 11660 15750 11690 15802
rect 11690 15750 11702 15802
rect 11702 15750 11716 15802
rect 11740 15750 11754 15802
rect 11754 15750 11766 15802
rect 11766 15750 11796 15802
rect 11820 15750 11830 15802
rect 11830 15750 11876 15802
rect 11580 15748 11636 15750
rect 11660 15748 11716 15750
rect 11740 15748 11796 15750
rect 11820 15748 11876 15750
rect 11978 15408 12034 15464
rect 12240 17434 12296 17436
rect 12320 17434 12376 17436
rect 12400 17434 12456 17436
rect 12480 17434 12536 17436
rect 12240 17382 12286 17434
rect 12286 17382 12296 17434
rect 12320 17382 12350 17434
rect 12350 17382 12362 17434
rect 12362 17382 12376 17434
rect 12400 17382 12414 17434
rect 12414 17382 12426 17434
rect 12426 17382 12456 17434
rect 12480 17382 12490 17434
rect 12490 17382 12536 17434
rect 12240 17380 12296 17382
rect 12320 17380 12376 17382
rect 12400 17380 12456 17382
rect 12480 17380 12536 17382
rect 12240 16346 12296 16348
rect 12320 16346 12376 16348
rect 12400 16346 12456 16348
rect 12480 16346 12536 16348
rect 12240 16294 12286 16346
rect 12286 16294 12296 16346
rect 12320 16294 12350 16346
rect 12350 16294 12362 16346
rect 12362 16294 12376 16346
rect 12400 16294 12414 16346
rect 12414 16294 12426 16346
rect 12426 16294 12456 16346
rect 12480 16294 12490 16346
rect 12490 16294 12536 16346
rect 12240 16292 12296 16294
rect 12320 16292 12376 16294
rect 12400 16292 12456 16294
rect 12480 16292 12536 16294
rect 13818 19236 13874 19272
rect 13818 19216 13820 19236
rect 13820 19216 13872 19236
rect 13872 19216 13874 19236
rect 12240 15258 12296 15260
rect 12320 15258 12376 15260
rect 12400 15258 12456 15260
rect 12480 15258 12536 15260
rect 12240 15206 12286 15258
rect 12286 15206 12296 15258
rect 12320 15206 12350 15258
rect 12350 15206 12362 15258
rect 12362 15206 12376 15258
rect 12400 15206 12414 15258
rect 12414 15206 12426 15258
rect 12426 15206 12456 15258
rect 12480 15206 12490 15258
rect 12490 15206 12536 15258
rect 12240 15204 12296 15206
rect 12320 15204 12376 15206
rect 12400 15204 12456 15206
rect 12480 15204 12536 15206
rect 11580 14714 11636 14716
rect 11660 14714 11716 14716
rect 11740 14714 11796 14716
rect 11820 14714 11876 14716
rect 11580 14662 11626 14714
rect 11626 14662 11636 14714
rect 11660 14662 11690 14714
rect 11690 14662 11702 14714
rect 11702 14662 11716 14714
rect 11740 14662 11754 14714
rect 11754 14662 11766 14714
rect 11766 14662 11796 14714
rect 11820 14662 11830 14714
rect 11830 14662 11876 14714
rect 11580 14660 11636 14662
rect 11660 14660 11716 14662
rect 11740 14660 11796 14662
rect 11820 14660 11876 14662
rect 12162 14456 12218 14512
rect 11580 13626 11636 13628
rect 11660 13626 11716 13628
rect 11740 13626 11796 13628
rect 11820 13626 11876 13628
rect 11580 13574 11626 13626
rect 11626 13574 11636 13626
rect 11660 13574 11690 13626
rect 11690 13574 11702 13626
rect 11702 13574 11716 13626
rect 11740 13574 11754 13626
rect 11754 13574 11766 13626
rect 11766 13574 11796 13626
rect 11820 13574 11830 13626
rect 11830 13574 11876 13626
rect 11580 13572 11636 13574
rect 11660 13572 11716 13574
rect 11740 13572 11796 13574
rect 11820 13572 11876 13574
rect 12240 14170 12296 14172
rect 12320 14170 12376 14172
rect 12400 14170 12456 14172
rect 12480 14170 12536 14172
rect 12240 14118 12286 14170
rect 12286 14118 12296 14170
rect 12320 14118 12350 14170
rect 12350 14118 12362 14170
rect 12362 14118 12376 14170
rect 12400 14118 12414 14170
rect 12414 14118 12426 14170
rect 12426 14118 12456 14170
rect 12480 14118 12490 14170
rect 12490 14118 12536 14170
rect 12240 14116 12296 14118
rect 12320 14116 12376 14118
rect 12400 14116 12456 14118
rect 12480 14116 12536 14118
rect 11518 13232 11574 13288
rect 12240 13082 12296 13084
rect 12320 13082 12376 13084
rect 12400 13082 12456 13084
rect 12480 13082 12536 13084
rect 12240 13030 12286 13082
rect 12286 13030 12296 13082
rect 12320 13030 12350 13082
rect 12350 13030 12362 13082
rect 12362 13030 12376 13082
rect 12400 13030 12414 13082
rect 12414 13030 12426 13082
rect 12426 13030 12456 13082
rect 12480 13030 12490 13082
rect 12490 13030 12536 13082
rect 12240 13028 12296 13030
rect 12320 13028 12376 13030
rect 12400 13028 12456 13030
rect 12480 13028 12536 13030
rect 13542 15408 13598 15464
rect 11580 12538 11636 12540
rect 11660 12538 11716 12540
rect 11740 12538 11796 12540
rect 11820 12538 11876 12540
rect 11580 12486 11626 12538
rect 11626 12486 11636 12538
rect 11660 12486 11690 12538
rect 11690 12486 11702 12538
rect 11702 12486 11716 12538
rect 11740 12486 11754 12538
rect 11754 12486 11766 12538
rect 11766 12486 11796 12538
rect 11820 12486 11830 12538
rect 11830 12486 11876 12538
rect 11580 12484 11636 12486
rect 11660 12484 11716 12486
rect 11740 12484 11796 12486
rect 11820 12484 11876 12486
rect 12240 11994 12296 11996
rect 12320 11994 12376 11996
rect 12400 11994 12456 11996
rect 12480 11994 12536 11996
rect 12240 11942 12286 11994
rect 12286 11942 12296 11994
rect 12320 11942 12350 11994
rect 12350 11942 12362 11994
rect 12362 11942 12376 11994
rect 12400 11942 12414 11994
rect 12414 11942 12426 11994
rect 12426 11942 12456 11994
rect 12480 11942 12490 11994
rect 12490 11942 12536 11994
rect 12240 11940 12296 11942
rect 12320 11940 12376 11942
rect 12400 11940 12456 11942
rect 12480 11940 12536 11942
rect 18663 29946 18719 29948
rect 18743 29946 18799 29948
rect 18823 29946 18879 29948
rect 18903 29946 18959 29948
rect 18663 29894 18709 29946
rect 18709 29894 18719 29946
rect 18743 29894 18773 29946
rect 18773 29894 18785 29946
rect 18785 29894 18799 29946
rect 18823 29894 18837 29946
rect 18837 29894 18849 29946
rect 18849 29894 18879 29946
rect 18903 29894 18913 29946
rect 18913 29894 18959 29946
rect 18663 29892 18719 29894
rect 18743 29892 18799 29894
rect 18823 29892 18879 29894
rect 18903 29892 18959 29894
rect 19323 29402 19379 29404
rect 19403 29402 19459 29404
rect 19483 29402 19539 29404
rect 19563 29402 19619 29404
rect 19323 29350 19369 29402
rect 19369 29350 19379 29402
rect 19403 29350 19433 29402
rect 19433 29350 19445 29402
rect 19445 29350 19459 29402
rect 19483 29350 19497 29402
rect 19497 29350 19509 29402
rect 19509 29350 19539 29402
rect 19563 29350 19573 29402
rect 19573 29350 19619 29402
rect 19323 29348 19379 29350
rect 19403 29348 19459 29350
rect 19483 29348 19539 29350
rect 19563 29348 19619 29350
rect 17958 28192 18014 28248
rect 15106 24248 15162 24304
rect 15014 20304 15070 20360
rect 16302 24248 16358 24304
rect 14094 15544 14150 15600
rect 11580 11450 11636 11452
rect 11660 11450 11716 11452
rect 11740 11450 11796 11452
rect 11820 11450 11876 11452
rect 11580 11398 11626 11450
rect 11626 11398 11636 11450
rect 11660 11398 11690 11450
rect 11690 11398 11702 11450
rect 11702 11398 11716 11450
rect 11740 11398 11754 11450
rect 11754 11398 11766 11450
rect 11766 11398 11796 11450
rect 11820 11398 11830 11450
rect 11830 11398 11876 11450
rect 11580 11396 11636 11398
rect 11660 11396 11716 11398
rect 11740 11396 11796 11398
rect 11820 11396 11876 11398
rect 11334 10512 11390 10568
rect 11580 10362 11636 10364
rect 11660 10362 11716 10364
rect 11740 10362 11796 10364
rect 11820 10362 11876 10364
rect 11580 10310 11626 10362
rect 11626 10310 11636 10362
rect 11660 10310 11690 10362
rect 11690 10310 11702 10362
rect 11702 10310 11716 10362
rect 11740 10310 11754 10362
rect 11754 10310 11766 10362
rect 11766 10310 11796 10362
rect 11820 10310 11830 10362
rect 11830 10310 11876 10362
rect 11580 10308 11636 10310
rect 11660 10308 11716 10310
rect 11740 10308 11796 10310
rect 11820 10308 11876 10310
rect 11334 9832 11390 9888
rect 9954 9016 10010 9072
rect 11242 9036 11298 9072
rect 11242 9016 11244 9036
rect 11244 9016 11296 9036
rect 11296 9016 11298 9036
rect 10782 8200 10838 8256
rect 10598 8064 10654 8120
rect 11580 9274 11636 9276
rect 11660 9274 11716 9276
rect 11740 9274 11796 9276
rect 11820 9274 11876 9276
rect 11580 9222 11626 9274
rect 11626 9222 11636 9274
rect 11660 9222 11690 9274
rect 11690 9222 11702 9274
rect 11702 9222 11716 9274
rect 11740 9222 11754 9274
rect 11754 9222 11766 9274
rect 11766 9222 11796 9274
rect 11820 9222 11830 9274
rect 11830 9222 11876 9274
rect 11580 9220 11636 9222
rect 11660 9220 11716 9222
rect 11740 9220 11796 9222
rect 11820 9220 11876 9222
rect 11580 8186 11636 8188
rect 11660 8186 11716 8188
rect 11740 8186 11796 8188
rect 11820 8186 11876 8188
rect 11580 8134 11626 8186
rect 11626 8134 11636 8186
rect 11660 8134 11690 8186
rect 11690 8134 11702 8186
rect 11702 8134 11716 8186
rect 11740 8134 11754 8186
rect 11754 8134 11766 8186
rect 11766 8134 11796 8186
rect 11820 8134 11830 8186
rect 11830 8134 11876 8186
rect 11580 8132 11636 8134
rect 11660 8132 11716 8134
rect 11740 8132 11796 8134
rect 11820 8132 11876 8134
rect 12240 10906 12296 10908
rect 12320 10906 12376 10908
rect 12400 10906 12456 10908
rect 12480 10906 12536 10908
rect 12240 10854 12286 10906
rect 12286 10854 12296 10906
rect 12320 10854 12350 10906
rect 12350 10854 12362 10906
rect 12362 10854 12376 10906
rect 12400 10854 12414 10906
rect 12414 10854 12426 10906
rect 12426 10854 12456 10906
rect 12480 10854 12490 10906
rect 12490 10854 12536 10906
rect 12240 10852 12296 10854
rect 12320 10852 12376 10854
rect 12400 10852 12456 10854
rect 12480 10852 12536 10854
rect 12622 10784 12678 10840
rect 13266 10648 13322 10704
rect 13358 9988 13414 10024
rect 13358 9968 13360 9988
rect 13360 9968 13412 9988
rect 13412 9968 13414 9988
rect 12240 9818 12296 9820
rect 12320 9818 12376 9820
rect 12400 9818 12456 9820
rect 12480 9818 12536 9820
rect 12240 9766 12286 9818
rect 12286 9766 12296 9818
rect 12320 9766 12350 9818
rect 12350 9766 12362 9818
rect 12362 9766 12376 9818
rect 12400 9766 12414 9818
rect 12414 9766 12426 9818
rect 12426 9766 12456 9818
rect 12480 9766 12490 9818
rect 12490 9766 12536 9818
rect 12240 9764 12296 9766
rect 12320 9764 12376 9766
rect 12400 9764 12456 9766
rect 12480 9764 12536 9766
rect 12162 9560 12218 9616
rect 11580 7098 11636 7100
rect 11660 7098 11716 7100
rect 11740 7098 11796 7100
rect 11820 7098 11876 7100
rect 11580 7046 11626 7098
rect 11626 7046 11636 7098
rect 11660 7046 11690 7098
rect 11690 7046 11702 7098
rect 11702 7046 11716 7098
rect 11740 7046 11754 7098
rect 11754 7046 11766 7098
rect 11766 7046 11796 7098
rect 11820 7046 11830 7098
rect 11830 7046 11876 7098
rect 11580 7044 11636 7046
rect 11660 7044 11716 7046
rect 11740 7044 11796 7046
rect 11820 7044 11876 7046
rect 10966 6704 11022 6760
rect 13174 9596 13176 9616
rect 13176 9596 13228 9616
rect 13228 9596 13230 9616
rect 13174 9560 13230 9596
rect 12240 8730 12296 8732
rect 12320 8730 12376 8732
rect 12400 8730 12456 8732
rect 12480 8730 12536 8732
rect 12240 8678 12286 8730
rect 12286 8678 12296 8730
rect 12320 8678 12350 8730
rect 12350 8678 12362 8730
rect 12362 8678 12376 8730
rect 12400 8678 12414 8730
rect 12414 8678 12426 8730
rect 12426 8678 12456 8730
rect 12480 8678 12490 8730
rect 12490 8678 12536 8730
rect 12240 8676 12296 8678
rect 12320 8676 12376 8678
rect 12400 8676 12456 8678
rect 12480 8676 12536 8678
rect 14094 12144 14150 12200
rect 12240 7642 12296 7644
rect 12320 7642 12376 7644
rect 12400 7642 12456 7644
rect 12480 7642 12536 7644
rect 12240 7590 12286 7642
rect 12286 7590 12296 7642
rect 12320 7590 12350 7642
rect 12350 7590 12362 7642
rect 12362 7590 12376 7642
rect 12400 7590 12414 7642
rect 12414 7590 12426 7642
rect 12426 7590 12456 7642
rect 12480 7590 12490 7642
rect 12490 7590 12536 7642
rect 12240 7588 12296 7590
rect 12320 7588 12376 7590
rect 12400 7588 12456 7590
rect 12480 7588 12536 7590
rect 12240 6554 12296 6556
rect 12320 6554 12376 6556
rect 12400 6554 12456 6556
rect 12480 6554 12536 6556
rect 12240 6502 12286 6554
rect 12286 6502 12296 6554
rect 12320 6502 12350 6554
rect 12350 6502 12362 6554
rect 12362 6502 12376 6554
rect 12400 6502 12414 6554
rect 12414 6502 12426 6554
rect 12426 6502 12456 6554
rect 12480 6502 12490 6554
rect 12490 6502 12536 6554
rect 12240 6500 12296 6502
rect 12320 6500 12376 6502
rect 12400 6500 12456 6502
rect 12480 6500 12536 6502
rect 11580 6010 11636 6012
rect 11660 6010 11716 6012
rect 11740 6010 11796 6012
rect 11820 6010 11876 6012
rect 11580 5958 11626 6010
rect 11626 5958 11636 6010
rect 11660 5958 11690 6010
rect 11690 5958 11702 6010
rect 11702 5958 11716 6010
rect 11740 5958 11754 6010
rect 11754 5958 11766 6010
rect 11766 5958 11796 6010
rect 11820 5958 11830 6010
rect 11830 5958 11876 6010
rect 11580 5956 11636 5958
rect 11660 5956 11716 5958
rect 11740 5956 11796 5958
rect 11820 5956 11876 5958
rect 12240 5466 12296 5468
rect 12320 5466 12376 5468
rect 12400 5466 12456 5468
rect 12480 5466 12536 5468
rect 12240 5414 12286 5466
rect 12286 5414 12296 5466
rect 12320 5414 12350 5466
rect 12350 5414 12362 5466
rect 12362 5414 12376 5466
rect 12400 5414 12414 5466
rect 12414 5414 12426 5466
rect 12426 5414 12456 5466
rect 12480 5414 12490 5466
rect 12490 5414 12536 5466
rect 12240 5412 12296 5414
rect 12320 5412 12376 5414
rect 12400 5412 12456 5414
rect 12480 5412 12536 5414
rect 15106 19896 15162 19952
rect 14278 12280 14334 12336
rect 13910 6740 13912 6760
rect 13912 6740 13964 6760
rect 13964 6740 13966 6760
rect 13910 6704 13966 6740
rect 11580 4922 11636 4924
rect 11660 4922 11716 4924
rect 11740 4922 11796 4924
rect 11820 4922 11876 4924
rect 11580 4870 11626 4922
rect 11626 4870 11636 4922
rect 11660 4870 11690 4922
rect 11690 4870 11702 4922
rect 11702 4870 11716 4922
rect 11740 4870 11754 4922
rect 11754 4870 11766 4922
rect 11766 4870 11796 4922
rect 11820 4870 11830 4922
rect 11830 4870 11876 4922
rect 11580 4868 11636 4870
rect 11660 4868 11716 4870
rect 11740 4868 11796 4870
rect 11820 4868 11876 4870
rect 5157 4378 5213 4380
rect 5237 4378 5293 4380
rect 5317 4378 5373 4380
rect 5397 4378 5453 4380
rect 5157 4326 5203 4378
rect 5203 4326 5213 4378
rect 5237 4326 5267 4378
rect 5267 4326 5279 4378
rect 5279 4326 5293 4378
rect 5317 4326 5331 4378
rect 5331 4326 5343 4378
rect 5343 4326 5373 4378
rect 5397 4326 5407 4378
rect 5407 4326 5453 4378
rect 5157 4324 5213 4326
rect 5237 4324 5293 4326
rect 5317 4324 5373 4326
rect 5397 4324 5453 4326
rect 12240 4378 12296 4380
rect 12320 4378 12376 4380
rect 12400 4378 12456 4380
rect 12480 4378 12536 4380
rect 12240 4326 12286 4378
rect 12286 4326 12296 4378
rect 12320 4326 12350 4378
rect 12350 4326 12362 4378
rect 12362 4326 12376 4378
rect 12400 4326 12414 4378
rect 12414 4326 12426 4378
rect 12426 4326 12456 4378
rect 12480 4326 12490 4378
rect 12490 4326 12536 4378
rect 12240 4324 12296 4326
rect 12320 4324 12376 4326
rect 12400 4324 12456 4326
rect 12480 4324 12536 4326
rect 4497 3834 4553 3836
rect 4577 3834 4633 3836
rect 4657 3834 4713 3836
rect 4737 3834 4793 3836
rect 4497 3782 4543 3834
rect 4543 3782 4553 3834
rect 4577 3782 4607 3834
rect 4607 3782 4619 3834
rect 4619 3782 4633 3834
rect 4657 3782 4671 3834
rect 4671 3782 4683 3834
rect 4683 3782 4713 3834
rect 4737 3782 4747 3834
rect 4747 3782 4793 3834
rect 4497 3780 4553 3782
rect 4577 3780 4633 3782
rect 4657 3780 4713 3782
rect 4737 3780 4793 3782
rect 11580 3834 11636 3836
rect 11660 3834 11716 3836
rect 11740 3834 11796 3836
rect 11820 3834 11876 3836
rect 11580 3782 11626 3834
rect 11626 3782 11636 3834
rect 11660 3782 11690 3834
rect 11690 3782 11702 3834
rect 11702 3782 11716 3834
rect 11740 3782 11754 3834
rect 11754 3782 11766 3834
rect 11766 3782 11796 3834
rect 11820 3782 11830 3834
rect 11830 3782 11876 3834
rect 11580 3780 11636 3782
rect 11660 3780 11716 3782
rect 11740 3780 11796 3782
rect 11820 3780 11876 3782
rect 12898 3596 12954 3632
rect 12898 3576 12900 3596
rect 12900 3576 12952 3596
rect 12952 3576 12954 3596
rect 938 3440 994 3496
rect 5157 3290 5213 3292
rect 5237 3290 5293 3292
rect 5317 3290 5373 3292
rect 5397 3290 5453 3292
rect 5157 3238 5203 3290
rect 5203 3238 5213 3290
rect 5237 3238 5267 3290
rect 5267 3238 5279 3290
rect 5279 3238 5293 3290
rect 5317 3238 5331 3290
rect 5331 3238 5343 3290
rect 5343 3238 5373 3290
rect 5397 3238 5407 3290
rect 5407 3238 5453 3290
rect 5157 3236 5213 3238
rect 5237 3236 5293 3238
rect 5317 3236 5373 3238
rect 5397 3236 5453 3238
rect 12240 3290 12296 3292
rect 12320 3290 12376 3292
rect 12400 3290 12456 3292
rect 12480 3290 12536 3292
rect 12240 3238 12286 3290
rect 12286 3238 12296 3290
rect 12320 3238 12350 3290
rect 12350 3238 12362 3290
rect 12362 3238 12376 3290
rect 12400 3238 12414 3290
rect 12414 3238 12426 3290
rect 12426 3238 12456 3290
rect 12480 3238 12490 3290
rect 12490 3238 12536 3290
rect 12240 3236 12296 3238
rect 12320 3236 12376 3238
rect 12400 3236 12456 3238
rect 12480 3236 12536 3238
rect 4497 2746 4553 2748
rect 4577 2746 4633 2748
rect 4657 2746 4713 2748
rect 4737 2746 4793 2748
rect 4497 2694 4543 2746
rect 4543 2694 4553 2746
rect 4577 2694 4607 2746
rect 4607 2694 4619 2746
rect 4619 2694 4633 2746
rect 4657 2694 4671 2746
rect 4671 2694 4683 2746
rect 4683 2694 4713 2746
rect 4737 2694 4747 2746
rect 4747 2694 4793 2746
rect 4497 2692 4553 2694
rect 4577 2692 4633 2694
rect 4657 2692 4713 2694
rect 4737 2692 4793 2694
rect 11580 2746 11636 2748
rect 11660 2746 11716 2748
rect 11740 2746 11796 2748
rect 11820 2746 11876 2748
rect 11580 2694 11626 2746
rect 11626 2694 11636 2746
rect 11660 2694 11690 2746
rect 11690 2694 11702 2746
rect 11702 2694 11716 2746
rect 11740 2694 11754 2746
rect 11754 2694 11766 2746
rect 11766 2694 11796 2746
rect 11820 2694 11830 2746
rect 11830 2694 11876 2746
rect 11580 2692 11636 2694
rect 11660 2692 11716 2694
rect 11740 2692 11796 2694
rect 11820 2692 11876 2694
rect 14646 4140 14702 4176
rect 14646 4120 14648 4140
rect 14648 4120 14700 4140
rect 14700 4120 14702 4140
rect 16118 12688 16174 12744
rect 18663 28858 18719 28860
rect 18743 28858 18799 28860
rect 18823 28858 18879 28860
rect 18903 28858 18959 28860
rect 18663 28806 18709 28858
rect 18709 28806 18719 28858
rect 18743 28806 18773 28858
rect 18773 28806 18785 28858
rect 18785 28806 18799 28858
rect 18823 28806 18837 28858
rect 18837 28806 18849 28858
rect 18849 28806 18879 28858
rect 18903 28806 18913 28858
rect 18913 28806 18959 28858
rect 18663 28804 18719 28806
rect 18743 28804 18799 28806
rect 18823 28804 18879 28806
rect 18903 28804 18959 28806
rect 19323 28314 19379 28316
rect 19403 28314 19459 28316
rect 19483 28314 19539 28316
rect 19563 28314 19619 28316
rect 19323 28262 19369 28314
rect 19369 28262 19379 28314
rect 19403 28262 19433 28314
rect 19433 28262 19445 28314
rect 19445 28262 19459 28314
rect 19483 28262 19497 28314
rect 19497 28262 19509 28314
rect 19509 28262 19539 28314
rect 19563 28262 19573 28314
rect 19573 28262 19619 28314
rect 19323 28260 19379 28262
rect 19403 28260 19459 28262
rect 19483 28260 19539 28262
rect 19563 28260 19619 28262
rect 18663 27770 18719 27772
rect 18743 27770 18799 27772
rect 18823 27770 18879 27772
rect 18903 27770 18959 27772
rect 18663 27718 18709 27770
rect 18709 27718 18719 27770
rect 18743 27718 18773 27770
rect 18773 27718 18785 27770
rect 18785 27718 18799 27770
rect 18823 27718 18837 27770
rect 18837 27718 18849 27770
rect 18849 27718 18879 27770
rect 18903 27718 18913 27770
rect 18913 27718 18959 27770
rect 18663 27716 18719 27718
rect 18743 27716 18799 27718
rect 18823 27716 18879 27718
rect 18903 27716 18959 27718
rect 19798 28056 19854 28112
rect 19323 27226 19379 27228
rect 19403 27226 19459 27228
rect 19483 27226 19539 27228
rect 19563 27226 19619 27228
rect 19323 27174 19369 27226
rect 19369 27174 19379 27226
rect 19403 27174 19433 27226
rect 19433 27174 19445 27226
rect 19445 27174 19459 27226
rect 19483 27174 19497 27226
rect 19497 27174 19509 27226
rect 19509 27174 19539 27226
rect 19563 27174 19573 27226
rect 19573 27174 19619 27226
rect 19323 27172 19379 27174
rect 19403 27172 19459 27174
rect 19483 27172 19539 27174
rect 19563 27172 19619 27174
rect 18663 26682 18719 26684
rect 18743 26682 18799 26684
rect 18823 26682 18879 26684
rect 18903 26682 18959 26684
rect 18663 26630 18709 26682
rect 18709 26630 18719 26682
rect 18743 26630 18773 26682
rect 18773 26630 18785 26682
rect 18785 26630 18799 26682
rect 18823 26630 18837 26682
rect 18837 26630 18849 26682
rect 18849 26630 18879 26682
rect 18903 26630 18913 26682
rect 18913 26630 18959 26682
rect 18663 26628 18719 26630
rect 18743 26628 18799 26630
rect 18823 26628 18879 26630
rect 18903 26628 18959 26630
rect 19323 26138 19379 26140
rect 19403 26138 19459 26140
rect 19483 26138 19539 26140
rect 19563 26138 19619 26140
rect 19323 26086 19369 26138
rect 19369 26086 19379 26138
rect 19403 26086 19433 26138
rect 19433 26086 19445 26138
rect 19445 26086 19459 26138
rect 19483 26086 19497 26138
rect 19497 26086 19509 26138
rect 19509 26086 19539 26138
rect 19563 26086 19573 26138
rect 19573 26086 19619 26138
rect 19323 26084 19379 26086
rect 19403 26084 19459 26086
rect 19483 26084 19539 26086
rect 19563 26084 19619 26086
rect 17682 21936 17738 21992
rect 18663 25594 18719 25596
rect 18743 25594 18799 25596
rect 18823 25594 18879 25596
rect 18903 25594 18959 25596
rect 18663 25542 18709 25594
rect 18709 25542 18719 25594
rect 18743 25542 18773 25594
rect 18773 25542 18785 25594
rect 18785 25542 18799 25594
rect 18823 25542 18837 25594
rect 18837 25542 18849 25594
rect 18849 25542 18879 25594
rect 18903 25542 18913 25594
rect 18913 25542 18959 25594
rect 18663 25540 18719 25542
rect 18743 25540 18799 25542
rect 18823 25540 18879 25542
rect 18903 25540 18959 25542
rect 18663 24506 18719 24508
rect 18743 24506 18799 24508
rect 18823 24506 18879 24508
rect 18903 24506 18959 24508
rect 18663 24454 18709 24506
rect 18709 24454 18719 24506
rect 18743 24454 18773 24506
rect 18773 24454 18785 24506
rect 18785 24454 18799 24506
rect 18823 24454 18837 24506
rect 18837 24454 18849 24506
rect 18849 24454 18879 24506
rect 18903 24454 18913 24506
rect 18913 24454 18959 24506
rect 18663 24452 18719 24454
rect 18743 24452 18799 24454
rect 18823 24452 18879 24454
rect 18903 24452 18959 24454
rect 19323 25050 19379 25052
rect 19403 25050 19459 25052
rect 19483 25050 19539 25052
rect 19563 25050 19619 25052
rect 19323 24998 19369 25050
rect 19369 24998 19379 25050
rect 19403 24998 19433 25050
rect 19433 24998 19445 25050
rect 19445 24998 19459 25050
rect 19483 24998 19497 25050
rect 19497 24998 19509 25050
rect 19509 24998 19539 25050
rect 19563 24998 19573 25050
rect 19573 24998 19619 25050
rect 19323 24996 19379 24998
rect 19403 24996 19459 24998
rect 19483 24996 19539 24998
rect 19563 24996 19619 24998
rect 22006 28600 22062 28656
rect 21914 27956 21916 27976
rect 21916 27956 21968 27976
rect 21968 27956 21970 27976
rect 19323 23962 19379 23964
rect 19403 23962 19459 23964
rect 19483 23962 19539 23964
rect 19563 23962 19619 23964
rect 19323 23910 19369 23962
rect 19369 23910 19379 23962
rect 19403 23910 19433 23962
rect 19433 23910 19445 23962
rect 19445 23910 19459 23962
rect 19483 23910 19497 23962
rect 19497 23910 19509 23962
rect 19509 23910 19539 23962
rect 19563 23910 19573 23962
rect 19573 23910 19619 23962
rect 19323 23908 19379 23910
rect 19403 23908 19459 23910
rect 19483 23908 19539 23910
rect 19563 23908 19619 23910
rect 18663 23418 18719 23420
rect 18743 23418 18799 23420
rect 18823 23418 18879 23420
rect 18903 23418 18959 23420
rect 18663 23366 18709 23418
rect 18709 23366 18719 23418
rect 18743 23366 18773 23418
rect 18773 23366 18785 23418
rect 18785 23366 18799 23418
rect 18823 23366 18837 23418
rect 18837 23366 18849 23418
rect 18849 23366 18879 23418
rect 18903 23366 18913 23418
rect 18913 23366 18959 23418
rect 18663 23364 18719 23366
rect 18743 23364 18799 23366
rect 18823 23364 18879 23366
rect 18903 23364 18959 23366
rect 19323 22874 19379 22876
rect 19403 22874 19459 22876
rect 19483 22874 19539 22876
rect 19563 22874 19619 22876
rect 19323 22822 19369 22874
rect 19369 22822 19379 22874
rect 19403 22822 19433 22874
rect 19433 22822 19445 22874
rect 19445 22822 19459 22874
rect 19483 22822 19497 22874
rect 19497 22822 19509 22874
rect 19509 22822 19539 22874
rect 19563 22822 19573 22874
rect 19573 22822 19619 22874
rect 19323 22820 19379 22822
rect 19403 22820 19459 22822
rect 19483 22820 19539 22822
rect 19563 22820 19619 22822
rect 18663 22330 18719 22332
rect 18743 22330 18799 22332
rect 18823 22330 18879 22332
rect 18903 22330 18959 22332
rect 18663 22278 18709 22330
rect 18709 22278 18719 22330
rect 18743 22278 18773 22330
rect 18773 22278 18785 22330
rect 18785 22278 18799 22330
rect 18823 22278 18837 22330
rect 18837 22278 18849 22330
rect 18849 22278 18879 22330
rect 18903 22278 18913 22330
rect 18913 22278 18959 22330
rect 18663 22276 18719 22278
rect 18743 22276 18799 22278
rect 18823 22276 18879 22278
rect 18903 22276 18959 22278
rect 19323 21786 19379 21788
rect 19403 21786 19459 21788
rect 19483 21786 19539 21788
rect 19563 21786 19619 21788
rect 19323 21734 19369 21786
rect 19369 21734 19379 21786
rect 19403 21734 19433 21786
rect 19433 21734 19445 21786
rect 19445 21734 19459 21786
rect 19483 21734 19497 21786
rect 19497 21734 19509 21786
rect 19509 21734 19539 21786
rect 19563 21734 19573 21786
rect 19573 21734 19619 21786
rect 19323 21732 19379 21734
rect 19403 21732 19459 21734
rect 19483 21732 19539 21734
rect 19563 21732 19619 21734
rect 21914 27920 21970 27956
rect 18663 21242 18719 21244
rect 18743 21242 18799 21244
rect 18823 21242 18879 21244
rect 18903 21242 18959 21244
rect 18663 21190 18709 21242
rect 18709 21190 18719 21242
rect 18743 21190 18773 21242
rect 18773 21190 18785 21242
rect 18785 21190 18799 21242
rect 18823 21190 18837 21242
rect 18837 21190 18849 21242
rect 18849 21190 18879 21242
rect 18903 21190 18913 21242
rect 18913 21190 18959 21242
rect 18663 21188 18719 21190
rect 18743 21188 18799 21190
rect 18823 21188 18879 21190
rect 18903 21188 18959 21190
rect 18234 20576 18290 20632
rect 17958 19216 18014 19272
rect 19338 20848 19394 20904
rect 18234 19352 18290 19408
rect 19062 20460 19118 20496
rect 19062 20440 19064 20460
rect 19064 20440 19116 20460
rect 19116 20440 19118 20460
rect 19323 20698 19379 20700
rect 19403 20698 19459 20700
rect 19483 20698 19539 20700
rect 19563 20698 19619 20700
rect 19323 20646 19369 20698
rect 19369 20646 19379 20698
rect 19403 20646 19433 20698
rect 19433 20646 19445 20698
rect 19445 20646 19459 20698
rect 19483 20646 19497 20698
rect 19497 20646 19509 20698
rect 19509 20646 19539 20698
rect 19563 20646 19573 20698
rect 19573 20646 19619 20698
rect 19323 20644 19379 20646
rect 19403 20644 19459 20646
rect 19483 20644 19539 20646
rect 19563 20644 19619 20646
rect 18663 20154 18719 20156
rect 18743 20154 18799 20156
rect 18823 20154 18879 20156
rect 18903 20154 18959 20156
rect 18663 20102 18709 20154
rect 18709 20102 18719 20154
rect 18743 20102 18773 20154
rect 18773 20102 18785 20154
rect 18785 20102 18799 20154
rect 18823 20102 18837 20154
rect 18837 20102 18849 20154
rect 18849 20102 18879 20154
rect 18903 20102 18913 20154
rect 18913 20102 18959 20154
rect 18663 20100 18719 20102
rect 18743 20100 18799 20102
rect 18823 20100 18879 20102
rect 18903 20100 18959 20102
rect 18878 19216 18934 19272
rect 18663 19066 18719 19068
rect 18743 19066 18799 19068
rect 18823 19066 18879 19068
rect 18903 19066 18959 19068
rect 18663 19014 18709 19066
rect 18709 19014 18719 19066
rect 18743 19014 18773 19066
rect 18773 19014 18785 19066
rect 18785 19014 18799 19066
rect 18823 19014 18837 19066
rect 18837 19014 18849 19066
rect 18849 19014 18879 19066
rect 18903 19014 18913 19066
rect 18913 19014 18959 19066
rect 18663 19012 18719 19014
rect 18743 19012 18799 19014
rect 18823 19012 18879 19014
rect 18903 19012 18959 19014
rect 19154 19352 19210 19408
rect 19323 19610 19379 19612
rect 19403 19610 19459 19612
rect 19483 19610 19539 19612
rect 19563 19610 19619 19612
rect 19323 19558 19369 19610
rect 19369 19558 19379 19610
rect 19403 19558 19433 19610
rect 19433 19558 19445 19610
rect 19445 19558 19459 19610
rect 19483 19558 19497 19610
rect 19497 19558 19509 19610
rect 19509 19558 19539 19610
rect 19563 19558 19573 19610
rect 19573 19558 19619 19610
rect 19323 19556 19379 19558
rect 19403 19556 19459 19558
rect 19483 19556 19539 19558
rect 19563 19556 19619 19558
rect 18663 17978 18719 17980
rect 18743 17978 18799 17980
rect 18823 17978 18879 17980
rect 18903 17978 18959 17980
rect 18663 17926 18709 17978
rect 18709 17926 18719 17978
rect 18743 17926 18773 17978
rect 18773 17926 18785 17978
rect 18785 17926 18799 17978
rect 18823 17926 18837 17978
rect 18837 17926 18849 17978
rect 18849 17926 18879 17978
rect 18903 17926 18913 17978
rect 18913 17926 18959 17978
rect 18663 17924 18719 17926
rect 18743 17924 18799 17926
rect 18823 17924 18879 17926
rect 18903 17924 18959 17926
rect 19323 18522 19379 18524
rect 19403 18522 19459 18524
rect 19483 18522 19539 18524
rect 19563 18522 19619 18524
rect 19323 18470 19369 18522
rect 19369 18470 19379 18522
rect 19403 18470 19433 18522
rect 19433 18470 19445 18522
rect 19445 18470 19459 18522
rect 19483 18470 19497 18522
rect 19497 18470 19509 18522
rect 19509 18470 19539 18522
rect 19563 18470 19573 18522
rect 19573 18470 19619 18522
rect 19323 18468 19379 18470
rect 19403 18468 19459 18470
rect 19483 18468 19539 18470
rect 19563 18468 19619 18470
rect 19522 17720 19578 17776
rect 21178 23044 21234 23080
rect 21178 23024 21180 23044
rect 21180 23024 21232 23044
rect 21232 23024 21234 23044
rect 20350 21836 20352 21856
rect 20352 21836 20404 21856
rect 20404 21836 20406 21856
rect 20350 21800 20406 21836
rect 19982 19352 20038 19408
rect 20258 19216 20314 19272
rect 19430 17584 19486 17640
rect 22190 22208 22246 22264
rect 21822 21528 21878 21584
rect 22190 20984 22246 21040
rect 19323 17434 19379 17436
rect 19403 17434 19459 17436
rect 19483 17434 19539 17436
rect 19563 17434 19619 17436
rect 19323 17382 19369 17434
rect 19369 17382 19379 17434
rect 19403 17382 19433 17434
rect 19433 17382 19445 17434
rect 19445 17382 19459 17434
rect 19483 17382 19497 17434
rect 19497 17382 19509 17434
rect 19509 17382 19539 17434
rect 19563 17382 19573 17434
rect 19573 17382 19619 17434
rect 19323 17380 19379 17382
rect 19403 17380 19459 17382
rect 19483 17380 19539 17382
rect 19563 17380 19619 17382
rect 18663 16890 18719 16892
rect 18743 16890 18799 16892
rect 18823 16890 18879 16892
rect 18903 16890 18959 16892
rect 18663 16838 18709 16890
rect 18709 16838 18719 16890
rect 18743 16838 18773 16890
rect 18773 16838 18785 16890
rect 18785 16838 18799 16890
rect 18823 16838 18837 16890
rect 18837 16838 18849 16890
rect 18849 16838 18879 16890
rect 18903 16838 18913 16890
rect 18913 16838 18959 16890
rect 18663 16836 18719 16838
rect 18743 16836 18799 16838
rect 18823 16836 18879 16838
rect 18903 16836 18959 16838
rect 19323 16346 19379 16348
rect 19403 16346 19459 16348
rect 19483 16346 19539 16348
rect 19563 16346 19619 16348
rect 19323 16294 19369 16346
rect 19369 16294 19379 16346
rect 19403 16294 19433 16346
rect 19433 16294 19445 16346
rect 19445 16294 19459 16346
rect 19483 16294 19497 16346
rect 19497 16294 19509 16346
rect 19509 16294 19539 16346
rect 19563 16294 19573 16346
rect 19573 16294 19619 16346
rect 19323 16292 19379 16294
rect 19403 16292 19459 16294
rect 19483 16292 19539 16294
rect 19563 16292 19619 16294
rect 18663 15802 18719 15804
rect 18743 15802 18799 15804
rect 18823 15802 18879 15804
rect 18903 15802 18959 15804
rect 18663 15750 18709 15802
rect 18709 15750 18719 15802
rect 18743 15750 18773 15802
rect 18773 15750 18785 15802
rect 18785 15750 18799 15802
rect 18823 15750 18837 15802
rect 18837 15750 18849 15802
rect 18849 15750 18879 15802
rect 18903 15750 18913 15802
rect 18913 15750 18959 15802
rect 18663 15748 18719 15750
rect 18743 15748 18799 15750
rect 18823 15748 18879 15750
rect 18903 15748 18959 15750
rect 16670 12280 16726 12336
rect 16026 9560 16082 9616
rect 18663 14714 18719 14716
rect 18743 14714 18799 14716
rect 18823 14714 18879 14716
rect 18903 14714 18959 14716
rect 18663 14662 18709 14714
rect 18709 14662 18719 14714
rect 18743 14662 18773 14714
rect 18773 14662 18785 14714
rect 18785 14662 18799 14714
rect 18823 14662 18837 14714
rect 18837 14662 18849 14714
rect 18849 14662 18879 14714
rect 18903 14662 18913 14714
rect 18913 14662 18959 14714
rect 18663 14660 18719 14662
rect 18743 14660 18799 14662
rect 18823 14660 18879 14662
rect 18903 14660 18959 14662
rect 17038 9288 17094 9344
rect 16486 5364 16542 5400
rect 16486 5344 16488 5364
rect 16488 5344 16540 5364
rect 16540 5344 16542 5364
rect 16210 5072 16266 5128
rect 16394 4664 16450 4720
rect 17222 7384 17278 7440
rect 17406 7928 17462 7984
rect 17406 7656 17462 7712
rect 19323 15258 19379 15260
rect 19403 15258 19459 15260
rect 19483 15258 19539 15260
rect 19563 15258 19619 15260
rect 19323 15206 19369 15258
rect 19369 15206 19379 15258
rect 19403 15206 19433 15258
rect 19433 15206 19445 15258
rect 19445 15206 19459 15258
rect 19483 15206 19497 15258
rect 19497 15206 19509 15258
rect 19509 15206 19539 15258
rect 19563 15206 19573 15258
rect 19573 15206 19619 15258
rect 19323 15204 19379 15206
rect 19403 15204 19459 15206
rect 19483 15204 19539 15206
rect 19563 15204 19619 15206
rect 19062 14320 19118 14376
rect 18663 13626 18719 13628
rect 18743 13626 18799 13628
rect 18823 13626 18879 13628
rect 18903 13626 18959 13628
rect 18663 13574 18709 13626
rect 18709 13574 18719 13626
rect 18743 13574 18773 13626
rect 18773 13574 18785 13626
rect 18785 13574 18799 13626
rect 18823 13574 18837 13626
rect 18837 13574 18849 13626
rect 18849 13574 18879 13626
rect 18903 13574 18913 13626
rect 18913 13574 18959 13626
rect 18663 13572 18719 13574
rect 18743 13572 18799 13574
rect 18823 13572 18879 13574
rect 18903 13572 18959 13574
rect 19323 14170 19379 14172
rect 19403 14170 19459 14172
rect 19483 14170 19539 14172
rect 19563 14170 19619 14172
rect 19323 14118 19369 14170
rect 19369 14118 19379 14170
rect 19403 14118 19433 14170
rect 19433 14118 19445 14170
rect 19445 14118 19459 14170
rect 19483 14118 19497 14170
rect 19497 14118 19509 14170
rect 19509 14118 19539 14170
rect 19563 14118 19573 14170
rect 19573 14118 19619 14170
rect 19323 14116 19379 14118
rect 19403 14116 19459 14118
rect 19483 14116 19539 14118
rect 19563 14116 19619 14118
rect 19706 14048 19762 14104
rect 20166 14048 20222 14104
rect 19323 13082 19379 13084
rect 19403 13082 19459 13084
rect 19483 13082 19539 13084
rect 19563 13082 19619 13084
rect 19323 13030 19369 13082
rect 19369 13030 19379 13082
rect 19403 13030 19433 13082
rect 19433 13030 19445 13082
rect 19445 13030 19459 13082
rect 19483 13030 19497 13082
rect 19497 13030 19509 13082
rect 19509 13030 19539 13082
rect 19563 13030 19573 13082
rect 19573 13030 19619 13082
rect 19323 13028 19379 13030
rect 19403 13028 19459 13030
rect 19483 13028 19539 13030
rect 19563 13028 19619 13030
rect 19062 12688 19118 12744
rect 18663 12538 18719 12540
rect 18743 12538 18799 12540
rect 18823 12538 18879 12540
rect 18903 12538 18959 12540
rect 18663 12486 18709 12538
rect 18709 12486 18719 12538
rect 18743 12486 18773 12538
rect 18773 12486 18785 12538
rect 18785 12486 18799 12538
rect 18823 12486 18837 12538
rect 18837 12486 18849 12538
rect 18849 12486 18879 12538
rect 18903 12486 18913 12538
rect 18913 12486 18959 12538
rect 18663 12484 18719 12486
rect 18743 12484 18799 12486
rect 18823 12484 18879 12486
rect 18903 12484 18959 12486
rect 18234 12144 18290 12200
rect 17774 9560 17830 9616
rect 18663 11450 18719 11452
rect 18743 11450 18799 11452
rect 18823 11450 18879 11452
rect 18903 11450 18959 11452
rect 18663 11398 18709 11450
rect 18709 11398 18719 11450
rect 18743 11398 18773 11450
rect 18773 11398 18785 11450
rect 18785 11398 18799 11450
rect 18823 11398 18837 11450
rect 18837 11398 18849 11450
rect 18849 11398 18879 11450
rect 18903 11398 18913 11450
rect 18913 11398 18959 11450
rect 18663 11396 18719 11398
rect 18743 11396 18799 11398
rect 18823 11396 18879 11398
rect 18903 11396 18959 11398
rect 18694 10648 18750 10704
rect 18970 10784 19026 10840
rect 18878 10512 18934 10568
rect 18663 10362 18719 10364
rect 18743 10362 18799 10364
rect 18823 10362 18879 10364
rect 18903 10362 18959 10364
rect 18663 10310 18709 10362
rect 18709 10310 18719 10362
rect 18743 10310 18773 10362
rect 18773 10310 18785 10362
rect 18785 10310 18799 10362
rect 18823 10310 18837 10362
rect 18837 10310 18849 10362
rect 18849 10310 18879 10362
rect 18903 10310 18913 10362
rect 18913 10310 18959 10362
rect 18663 10308 18719 10310
rect 18743 10308 18799 10310
rect 18823 10308 18879 10310
rect 18903 10308 18959 10310
rect 19323 11994 19379 11996
rect 19403 11994 19459 11996
rect 19483 11994 19539 11996
rect 19563 11994 19619 11996
rect 19323 11942 19369 11994
rect 19369 11942 19379 11994
rect 19403 11942 19433 11994
rect 19433 11942 19445 11994
rect 19445 11942 19459 11994
rect 19483 11942 19497 11994
rect 19497 11942 19509 11994
rect 19509 11942 19539 11994
rect 19563 11942 19573 11994
rect 19573 11942 19619 11994
rect 19323 11940 19379 11942
rect 19403 11940 19459 11942
rect 19483 11940 19539 11942
rect 19563 11940 19619 11942
rect 18970 9560 19026 9616
rect 18418 9424 18474 9480
rect 18326 9288 18382 9344
rect 18663 9274 18719 9276
rect 18743 9274 18799 9276
rect 18823 9274 18879 9276
rect 18903 9274 18959 9276
rect 18663 9222 18709 9274
rect 18709 9222 18719 9274
rect 18743 9222 18773 9274
rect 18773 9222 18785 9274
rect 18785 9222 18799 9274
rect 18823 9222 18837 9274
rect 18837 9222 18849 9274
rect 18849 9222 18879 9274
rect 18903 9222 18913 9274
rect 18913 9222 18959 9274
rect 18663 9220 18719 9222
rect 18743 9220 18799 9222
rect 18823 9220 18879 9222
rect 18903 9220 18959 9222
rect 20902 14320 20958 14376
rect 23110 22208 23166 22264
rect 22926 20984 22982 21040
rect 23938 22344 23994 22400
rect 23754 21564 23756 21584
rect 23756 21564 23808 21584
rect 23808 21564 23810 21584
rect 23754 21528 23810 21564
rect 19323 10906 19379 10908
rect 19403 10906 19459 10908
rect 19483 10906 19539 10908
rect 19563 10906 19619 10908
rect 19323 10854 19369 10906
rect 19369 10854 19379 10906
rect 19403 10854 19433 10906
rect 19433 10854 19445 10906
rect 19445 10854 19459 10906
rect 19483 10854 19497 10906
rect 19497 10854 19509 10906
rect 19509 10854 19539 10906
rect 19563 10854 19573 10906
rect 19573 10854 19619 10906
rect 19323 10852 19379 10854
rect 19403 10852 19459 10854
rect 19483 10852 19539 10854
rect 19563 10852 19619 10854
rect 19798 10240 19854 10296
rect 19323 9818 19379 9820
rect 19403 9818 19459 9820
rect 19483 9818 19539 9820
rect 19563 9818 19619 9820
rect 19323 9766 19369 9818
rect 19369 9766 19379 9818
rect 19403 9766 19433 9818
rect 19433 9766 19445 9818
rect 19445 9766 19459 9818
rect 19483 9766 19497 9818
rect 19497 9766 19509 9818
rect 19509 9766 19539 9818
rect 19563 9766 19573 9818
rect 19573 9766 19619 9818
rect 19323 9764 19379 9766
rect 19403 9764 19459 9766
rect 19483 9764 19539 9766
rect 19563 9764 19619 9766
rect 19323 8730 19379 8732
rect 19403 8730 19459 8732
rect 19483 8730 19539 8732
rect 19563 8730 19619 8732
rect 19323 8678 19369 8730
rect 19369 8678 19379 8730
rect 19403 8678 19433 8730
rect 19433 8678 19445 8730
rect 19445 8678 19459 8730
rect 19483 8678 19497 8730
rect 19497 8678 19509 8730
rect 19509 8678 19539 8730
rect 19563 8678 19573 8730
rect 19573 8678 19619 8730
rect 19323 8676 19379 8678
rect 19403 8676 19459 8678
rect 19483 8676 19539 8678
rect 19563 8676 19619 8678
rect 18663 8186 18719 8188
rect 18743 8186 18799 8188
rect 18823 8186 18879 8188
rect 18903 8186 18959 8188
rect 18663 8134 18709 8186
rect 18709 8134 18719 8186
rect 18743 8134 18773 8186
rect 18773 8134 18785 8186
rect 18785 8134 18799 8186
rect 18823 8134 18837 8186
rect 18837 8134 18849 8186
rect 18849 8134 18879 8186
rect 18903 8134 18913 8186
rect 18913 8134 18959 8186
rect 18663 8132 18719 8134
rect 18743 8132 18799 8134
rect 18823 8132 18879 8134
rect 18903 8132 18959 8134
rect 17958 7656 18014 7712
rect 17866 7404 17922 7440
rect 19323 7642 19379 7644
rect 19403 7642 19459 7644
rect 19483 7642 19539 7644
rect 19563 7642 19619 7644
rect 19323 7590 19369 7642
rect 19369 7590 19379 7642
rect 19403 7590 19433 7642
rect 19433 7590 19445 7642
rect 19445 7590 19459 7642
rect 19483 7590 19497 7642
rect 19497 7590 19509 7642
rect 19509 7590 19539 7642
rect 19563 7590 19573 7642
rect 19573 7590 19619 7642
rect 19323 7588 19379 7590
rect 19403 7588 19459 7590
rect 19483 7588 19539 7590
rect 19563 7588 19619 7590
rect 17866 7384 17868 7404
rect 17868 7384 17920 7404
rect 17920 7384 17922 7404
rect 18663 7098 18719 7100
rect 18743 7098 18799 7100
rect 18823 7098 18879 7100
rect 18903 7098 18959 7100
rect 18663 7046 18709 7098
rect 18709 7046 18719 7098
rect 18743 7046 18773 7098
rect 18773 7046 18785 7098
rect 18785 7046 18799 7098
rect 18823 7046 18837 7098
rect 18837 7046 18849 7098
rect 18849 7046 18879 7098
rect 18903 7046 18913 7098
rect 18913 7046 18959 7098
rect 18663 7044 18719 7046
rect 18743 7044 18799 7046
rect 18823 7044 18879 7046
rect 18903 7044 18959 7046
rect 22650 7928 22706 7984
rect 22926 10260 22982 10296
rect 22926 10240 22928 10260
rect 22928 10240 22980 10260
rect 22980 10240 22982 10260
rect 24398 22344 24454 22400
rect 25746 29946 25802 29948
rect 25826 29946 25882 29948
rect 25906 29946 25962 29948
rect 25986 29946 26042 29948
rect 25746 29894 25792 29946
rect 25792 29894 25802 29946
rect 25826 29894 25856 29946
rect 25856 29894 25868 29946
rect 25868 29894 25882 29946
rect 25906 29894 25920 29946
rect 25920 29894 25932 29946
rect 25932 29894 25962 29946
rect 25986 29894 25996 29946
rect 25996 29894 26042 29946
rect 25746 29892 25802 29894
rect 25826 29892 25882 29894
rect 25906 29892 25962 29894
rect 25986 29892 26042 29894
rect 26406 29402 26462 29404
rect 26486 29402 26542 29404
rect 26566 29402 26622 29404
rect 26646 29402 26702 29404
rect 26406 29350 26452 29402
rect 26452 29350 26462 29402
rect 26486 29350 26516 29402
rect 26516 29350 26528 29402
rect 26528 29350 26542 29402
rect 26566 29350 26580 29402
rect 26580 29350 26592 29402
rect 26592 29350 26622 29402
rect 26646 29350 26656 29402
rect 26656 29350 26702 29402
rect 26406 29348 26462 29350
rect 26486 29348 26542 29350
rect 26566 29348 26622 29350
rect 26646 29348 26702 29350
rect 28722 29008 28778 29064
rect 25746 28858 25802 28860
rect 25826 28858 25882 28860
rect 25906 28858 25962 28860
rect 25986 28858 26042 28860
rect 25746 28806 25792 28858
rect 25792 28806 25802 28858
rect 25826 28806 25856 28858
rect 25856 28806 25868 28858
rect 25868 28806 25882 28858
rect 25906 28806 25920 28858
rect 25920 28806 25932 28858
rect 25932 28806 25962 28858
rect 25986 28806 25996 28858
rect 25996 28806 26042 28858
rect 25746 28804 25802 28806
rect 25826 28804 25882 28806
rect 25906 28804 25962 28806
rect 25986 28804 26042 28806
rect 26406 28314 26462 28316
rect 26486 28314 26542 28316
rect 26566 28314 26622 28316
rect 26646 28314 26702 28316
rect 26406 28262 26452 28314
rect 26452 28262 26462 28314
rect 26486 28262 26516 28314
rect 26516 28262 26528 28314
rect 26528 28262 26542 28314
rect 26566 28262 26580 28314
rect 26580 28262 26592 28314
rect 26592 28262 26622 28314
rect 26646 28262 26656 28314
rect 26656 28262 26702 28314
rect 26406 28260 26462 28262
rect 26486 28260 26542 28262
rect 26566 28260 26622 28262
rect 26646 28260 26702 28262
rect 25746 27770 25802 27772
rect 25826 27770 25882 27772
rect 25906 27770 25962 27772
rect 25986 27770 26042 27772
rect 25746 27718 25792 27770
rect 25792 27718 25802 27770
rect 25826 27718 25856 27770
rect 25856 27718 25868 27770
rect 25868 27718 25882 27770
rect 25906 27718 25920 27770
rect 25920 27718 25932 27770
rect 25932 27718 25962 27770
rect 25986 27718 25996 27770
rect 25996 27718 26042 27770
rect 25746 27716 25802 27718
rect 25826 27716 25882 27718
rect 25906 27716 25962 27718
rect 25986 27716 26042 27718
rect 26406 27226 26462 27228
rect 26486 27226 26542 27228
rect 26566 27226 26622 27228
rect 26646 27226 26702 27228
rect 26406 27174 26452 27226
rect 26452 27174 26462 27226
rect 26486 27174 26516 27226
rect 26516 27174 26528 27226
rect 26528 27174 26542 27226
rect 26566 27174 26580 27226
rect 26580 27174 26592 27226
rect 26592 27174 26622 27226
rect 26646 27174 26656 27226
rect 26656 27174 26702 27226
rect 26406 27172 26462 27174
rect 26486 27172 26542 27174
rect 26566 27172 26622 27174
rect 26646 27172 26702 27174
rect 25746 26682 25802 26684
rect 25826 26682 25882 26684
rect 25906 26682 25962 26684
rect 25986 26682 26042 26684
rect 25746 26630 25792 26682
rect 25792 26630 25802 26682
rect 25826 26630 25856 26682
rect 25856 26630 25868 26682
rect 25868 26630 25882 26682
rect 25906 26630 25920 26682
rect 25920 26630 25932 26682
rect 25932 26630 25962 26682
rect 25986 26630 25996 26682
rect 25996 26630 26042 26682
rect 25746 26628 25802 26630
rect 25826 26628 25882 26630
rect 25906 26628 25962 26630
rect 25986 26628 26042 26630
rect 26406 26138 26462 26140
rect 26486 26138 26542 26140
rect 26566 26138 26622 26140
rect 26646 26138 26702 26140
rect 26406 26086 26452 26138
rect 26452 26086 26462 26138
rect 26486 26086 26516 26138
rect 26516 26086 26528 26138
rect 26528 26086 26542 26138
rect 26566 26086 26580 26138
rect 26580 26086 26592 26138
rect 26592 26086 26622 26138
rect 26646 26086 26656 26138
rect 26656 26086 26702 26138
rect 26406 26084 26462 26086
rect 26486 26084 26542 26086
rect 26566 26084 26622 26086
rect 26646 26084 26702 26086
rect 25746 25594 25802 25596
rect 25826 25594 25882 25596
rect 25906 25594 25962 25596
rect 25986 25594 26042 25596
rect 25746 25542 25792 25594
rect 25792 25542 25802 25594
rect 25826 25542 25856 25594
rect 25856 25542 25868 25594
rect 25868 25542 25882 25594
rect 25906 25542 25920 25594
rect 25920 25542 25932 25594
rect 25932 25542 25962 25594
rect 25986 25542 25996 25594
rect 25996 25542 26042 25594
rect 25746 25540 25802 25542
rect 25826 25540 25882 25542
rect 25906 25540 25962 25542
rect 25986 25540 26042 25542
rect 26406 25050 26462 25052
rect 26486 25050 26542 25052
rect 26566 25050 26622 25052
rect 26646 25050 26702 25052
rect 26406 24998 26452 25050
rect 26452 24998 26462 25050
rect 26486 24998 26516 25050
rect 26516 24998 26528 25050
rect 26528 24998 26542 25050
rect 26566 24998 26580 25050
rect 26580 24998 26592 25050
rect 26592 24998 26622 25050
rect 26646 24998 26656 25050
rect 26656 24998 26702 25050
rect 26406 24996 26462 24998
rect 26486 24996 26542 24998
rect 26566 24996 26622 24998
rect 26646 24996 26702 24998
rect 25746 24506 25802 24508
rect 25826 24506 25882 24508
rect 25906 24506 25962 24508
rect 25986 24506 26042 24508
rect 25746 24454 25792 24506
rect 25792 24454 25802 24506
rect 25826 24454 25856 24506
rect 25856 24454 25868 24506
rect 25868 24454 25882 24506
rect 25906 24454 25920 24506
rect 25920 24454 25932 24506
rect 25932 24454 25962 24506
rect 25986 24454 25996 24506
rect 25996 24454 26042 24506
rect 25746 24452 25802 24454
rect 25826 24452 25882 24454
rect 25906 24452 25962 24454
rect 25986 24452 26042 24454
rect 26406 23962 26462 23964
rect 26486 23962 26542 23964
rect 26566 23962 26622 23964
rect 26646 23962 26702 23964
rect 26406 23910 26452 23962
rect 26452 23910 26462 23962
rect 26486 23910 26516 23962
rect 26516 23910 26528 23962
rect 26528 23910 26542 23962
rect 26566 23910 26580 23962
rect 26580 23910 26592 23962
rect 26592 23910 26622 23962
rect 26646 23910 26656 23962
rect 26656 23910 26702 23962
rect 26406 23908 26462 23910
rect 26486 23908 26542 23910
rect 26566 23908 26622 23910
rect 26646 23908 26702 23910
rect 25746 23418 25802 23420
rect 25826 23418 25882 23420
rect 25906 23418 25962 23420
rect 25986 23418 26042 23420
rect 25746 23366 25792 23418
rect 25792 23366 25802 23418
rect 25826 23366 25856 23418
rect 25856 23366 25868 23418
rect 25868 23366 25882 23418
rect 25906 23366 25920 23418
rect 25920 23366 25932 23418
rect 25932 23366 25962 23418
rect 25986 23366 25996 23418
rect 25996 23366 26042 23418
rect 25746 23364 25802 23366
rect 25826 23364 25882 23366
rect 25906 23364 25962 23366
rect 25986 23364 26042 23366
rect 24766 22636 24822 22672
rect 24766 22616 24768 22636
rect 24768 22616 24820 22636
rect 24820 22616 24822 22636
rect 24858 22208 24914 22264
rect 26406 22874 26462 22876
rect 26486 22874 26542 22876
rect 26566 22874 26622 22876
rect 26646 22874 26702 22876
rect 26406 22822 26452 22874
rect 26452 22822 26462 22874
rect 26486 22822 26516 22874
rect 26516 22822 26528 22874
rect 26528 22822 26542 22874
rect 26566 22822 26580 22874
rect 26580 22822 26592 22874
rect 26592 22822 26622 22874
rect 26646 22822 26656 22874
rect 26656 22822 26702 22874
rect 26406 22820 26462 22822
rect 26486 22820 26542 22822
rect 26566 22820 26622 22822
rect 26646 22820 26702 22822
rect 25746 22330 25802 22332
rect 25826 22330 25882 22332
rect 25906 22330 25962 22332
rect 25986 22330 26042 22332
rect 25746 22278 25792 22330
rect 25792 22278 25802 22330
rect 25826 22278 25856 22330
rect 25856 22278 25868 22330
rect 25868 22278 25882 22330
rect 25906 22278 25920 22330
rect 25920 22278 25932 22330
rect 25932 22278 25962 22330
rect 25986 22278 25996 22330
rect 25996 22278 26042 22330
rect 25746 22276 25802 22278
rect 25826 22276 25882 22278
rect 25906 22276 25962 22278
rect 25986 22276 26042 22278
rect 25042 21800 25098 21856
rect 26146 21936 26202 21992
rect 25746 21242 25802 21244
rect 25826 21242 25882 21244
rect 25906 21242 25962 21244
rect 25986 21242 26042 21244
rect 25746 21190 25792 21242
rect 25792 21190 25802 21242
rect 25826 21190 25856 21242
rect 25856 21190 25868 21242
rect 25868 21190 25882 21242
rect 25906 21190 25920 21242
rect 25920 21190 25932 21242
rect 25932 21190 25962 21242
rect 25986 21190 25996 21242
rect 25996 21190 26042 21242
rect 25746 21188 25802 21190
rect 25826 21188 25882 21190
rect 25906 21188 25962 21190
rect 25986 21188 26042 21190
rect 26406 21786 26462 21788
rect 26486 21786 26542 21788
rect 26566 21786 26622 21788
rect 26646 21786 26702 21788
rect 26406 21734 26452 21786
rect 26452 21734 26462 21786
rect 26486 21734 26516 21786
rect 26516 21734 26528 21786
rect 26528 21734 26542 21786
rect 26566 21734 26580 21786
rect 26580 21734 26592 21786
rect 26592 21734 26622 21786
rect 26646 21734 26656 21786
rect 26656 21734 26702 21786
rect 26406 21732 26462 21734
rect 26486 21732 26542 21734
rect 26566 21732 26622 21734
rect 26646 21732 26702 21734
rect 27066 21412 27122 21448
rect 27066 21392 27068 21412
rect 27068 21392 27120 21412
rect 27120 21392 27122 21412
rect 26406 20698 26462 20700
rect 26486 20698 26542 20700
rect 26566 20698 26622 20700
rect 26646 20698 26702 20700
rect 26406 20646 26452 20698
rect 26452 20646 26462 20698
rect 26486 20646 26516 20698
rect 26516 20646 26528 20698
rect 26528 20646 26542 20698
rect 26566 20646 26580 20698
rect 26580 20646 26592 20698
rect 26592 20646 26622 20698
rect 26646 20646 26656 20698
rect 26656 20646 26702 20698
rect 26406 20644 26462 20646
rect 26486 20644 26542 20646
rect 26566 20644 26622 20646
rect 26646 20644 26702 20646
rect 25746 20154 25802 20156
rect 25826 20154 25882 20156
rect 25906 20154 25962 20156
rect 25986 20154 26042 20156
rect 25746 20102 25792 20154
rect 25792 20102 25802 20154
rect 25826 20102 25856 20154
rect 25856 20102 25868 20154
rect 25868 20102 25882 20154
rect 25906 20102 25920 20154
rect 25920 20102 25932 20154
rect 25932 20102 25962 20154
rect 25986 20102 25996 20154
rect 25996 20102 26042 20154
rect 25746 20100 25802 20102
rect 25826 20100 25882 20102
rect 25906 20100 25962 20102
rect 25986 20100 26042 20102
rect 25746 19066 25802 19068
rect 25826 19066 25882 19068
rect 25906 19066 25962 19068
rect 25986 19066 26042 19068
rect 25746 19014 25792 19066
rect 25792 19014 25802 19066
rect 25826 19014 25856 19066
rect 25856 19014 25868 19066
rect 25868 19014 25882 19066
rect 25906 19014 25920 19066
rect 25920 19014 25932 19066
rect 25932 19014 25962 19066
rect 25986 19014 25996 19066
rect 25996 19014 26042 19066
rect 25746 19012 25802 19014
rect 25826 19012 25882 19014
rect 25906 19012 25962 19014
rect 25986 19012 26042 19014
rect 24950 17176 25006 17232
rect 25746 17978 25802 17980
rect 25826 17978 25882 17980
rect 25906 17978 25962 17980
rect 25986 17978 26042 17980
rect 25746 17926 25792 17978
rect 25792 17926 25802 17978
rect 25826 17926 25856 17978
rect 25856 17926 25868 17978
rect 25868 17926 25882 17978
rect 25906 17926 25920 17978
rect 25920 17926 25932 17978
rect 25932 17926 25962 17978
rect 25986 17926 25996 17978
rect 25996 17926 26042 17978
rect 25746 17924 25802 17926
rect 25826 17924 25882 17926
rect 25906 17924 25962 17926
rect 25986 17924 26042 17926
rect 25594 17720 25650 17776
rect 25746 16890 25802 16892
rect 25826 16890 25882 16892
rect 25906 16890 25962 16892
rect 25986 16890 26042 16892
rect 25746 16838 25792 16890
rect 25792 16838 25802 16890
rect 25826 16838 25856 16890
rect 25856 16838 25868 16890
rect 25868 16838 25882 16890
rect 25906 16838 25920 16890
rect 25920 16838 25932 16890
rect 25932 16838 25962 16890
rect 25986 16838 25996 16890
rect 25996 16838 26042 16890
rect 25746 16836 25802 16838
rect 25826 16836 25882 16838
rect 25906 16836 25962 16838
rect 25986 16836 26042 16838
rect 26406 19610 26462 19612
rect 26486 19610 26542 19612
rect 26566 19610 26622 19612
rect 26646 19610 26702 19612
rect 26406 19558 26452 19610
rect 26452 19558 26462 19610
rect 26486 19558 26516 19610
rect 26516 19558 26528 19610
rect 26528 19558 26542 19610
rect 26566 19558 26580 19610
rect 26580 19558 26592 19610
rect 26592 19558 26622 19610
rect 26646 19558 26656 19610
rect 26656 19558 26702 19610
rect 26406 19556 26462 19558
rect 26486 19556 26542 19558
rect 26566 19556 26622 19558
rect 26646 19556 26702 19558
rect 26406 18522 26462 18524
rect 26486 18522 26542 18524
rect 26566 18522 26622 18524
rect 26646 18522 26702 18524
rect 26406 18470 26452 18522
rect 26452 18470 26462 18522
rect 26486 18470 26516 18522
rect 26516 18470 26528 18522
rect 26528 18470 26542 18522
rect 26566 18470 26580 18522
rect 26580 18470 26592 18522
rect 26592 18470 26622 18522
rect 26646 18470 26656 18522
rect 26656 18470 26702 18522
rect 26406 18468 26462 18470
rect 26486 18468 26542 18470
rect 26566 18468 26622 18470
rect 26646 18468 26702 18470
rect 26406 17434 26462 17436
rect 26486 17434 26542 17436
rect 26566 17434 26622 17436
rect 26646 17434 26702 17436
rect 26406 17382 26452 17434
rect 26452 17382 26462 17434
rect 26486 17382 26516 17434
rect 26516 17382 26528 17434
rect 26528 17382 26542 17434
rect 26566 17382 26580 17434
rect 26580 17382 26592 17434
rect 26592 17382 26622 17434
rect 26646 17382 26656 17434
rect 26656 17382 26702 17434
rect 26406 17380 26462 17382
rect 26486 17380 26542 17382
rect 26566 17380 26622 17382
rect 26646 17380 26702 17382
rect 26330 17040 26386 17096
rect 26406 16346 26462 16348
rect 26486 16346 26542 16348
rect 26566 16346 26622 16348
rect 26646 16346 26702 16348
rect 26406 16294 26452 16346
rect 26452 16294 26462 16346
rect 26486 16294 26516 16346
rect 26516 16294 26528 16346
rect 26528 16294 26542 16346
rect 26566 16294 26580 16346
rect 26580 16294 26592 16346
rect 26592 16294 26622 16346
rect 26646 16294 26656 16346
rect 26656 16294 26702 16346
rect 26406 16292 26462 16294
rect 26486 16292 26542 16294
rect 26566 16292 26622 16294
rect 26646 16292 26702 16294
rect 25746 15802 25802 15804
rect 25826 15802 25882 15804
rect 25906 15802 25962 15804
rect 25986 15802 26042 15804
rect 25746 15750 25792 15802
rect 25792 15750 25802 15802
rect 25826 15750 25856 15802
rect 25856 15750 25868 15802
rect 25868 15750 25882 15802
rect 25906 15750 25920 15802
rect 25920 15750 25932 15802
rect 25932 15750 25962 15802
rect 25986 15750 25996 15802
rect 25996 15750 26042 15802
rect 25746 15748 25802 15750
rect 25826 15748 25882 15750
rect 25906 15748 25962 15750
rect 25986 15748 26042 15750
rect 26606 15408 26662 15464
rect 26406 15258 26462 15260
rect 26486 15258 26542 15260
rect 26566 15258 26622 15260
rect 26646 15258 26702 15260
rect 26406 15206 26452 15258
rect 26452 15206 26462 15258
rect 26486 15206 26516 15258
rect 26516 15206 26528 15258
rect 26528 15206 26542 15258
rect 26566 15206 26580 15258
rect 26580 15206 26592 15258
rect 26592 15206 26622 15258
rect 26646 15206 26656 15258
rect 26656 15206 26702 15258
rect 26406 15204 26462 15206
rect 26486 15204 26542 15206
rect 26566 15204 26622 15206
rect 26646 15204 26702 15206
rect 25746 14714 25802 14716
rect 25826 14714 25882 14716
rect 25906 14714 25962 14716
rect 25986 14714 26042 14716
rect 25746 14662 25792 14714
rect 25792 14662 25802 14714
rect 25826 14662 25856 14714
rect 25856 14662 25868 14714
rect 25868 14662 25882 14714
rect 25906 14662 25920 14714
rect 25920 14662 25932 14714
rect 25932 14662 25962 14714
rect 25986 14662 25996 14714
rect 25996 14662 26042 14714
rect 25746 14660 25802 14662
rect 25826 14660 25882 14662
rect 25906 14660 25962 14662
rect 25986 14660 26042 14662
rect 27802 17992 27858 18048
rect 27986 17176 28042 17232
rect 27894 17040 27950 17096
rect 26406 14170 26462 14172
rect 26486 14170 26542 14172
rect 26566 14170 26622 14172
rect 26646 14170 26702 14172
rect 26406 14118 26452 14170
rect 26452 14118 26462 14170
rect 26486 14118 26516 14170
rect 26516 14118 26528 14170
rect 26528 14118 26542 14170
rect 26566 14118 26580 14170
rect 26580 14118 26592 14170
rect 26592 14118 26622 14170
rect 26646 14118 26656 14170
rect 26656 14118 26702 14170
rect 26406 14116 26462 14118
rect 26486 14116 26542 14118
rect 26566 14116 26622 14118
rect 26646 14116 26702 14118
rect 23110 9968 23166 10024
rect 20074 6704 20130 6760
rect 19323 6554 19379 6556
rect 19403 6554 19459 6556
rect 19483 6554 19539 6556
rect 19563 6554 19619 6556
rect 19323 6502 19369 6554
rect 19369 6502 19379 6554
rect 19403 6502 19433 6554
rect 19433 6502 19445 6554
rect 19445 6502 19459 6554
rect 19483 6502 19497 6554
rect 19497 6502 19509 6554
rect 19509 6502 19539 6554
rect 19563 6502 19573 6554
rect 19573 6502 19619 6554
rect 19323 6500 19379 6502
rect 19403 6500 19459 6502
rect 19483 6500 19539 6502
rect 19563 6500 19619 6502
rect 20258 6316 20314 6352
rect 20258 6296 20260 6316
rect 20260 6296 20312 6316
rect 20312 6296 20314 6316
rect 18663 6010 18719 6012
rect 18743 6010 18799 6012
rect 18823 6010 18879 6012
rect 18903 6010 18959 6012
rect 18663 5958 18709 6010
rect 18709 5958 18719 6010
rect 18743 5958 18773 6010
rect 18773 5958 18785 6010
rect 18785 5958 18799 6010
rect 18823 5958 18837 6010
rect 18837 5958 18849 6010
rect 18849 5958 18879 6010
rect 18903 5958 18913 6010
rect 18913 5958 18959 6010
rect 18663 5956 18719 5958
rect 18743 5956 18799 5958
rect 18823 5956 18879 5958
rect 18903 5956 18959 5958
rect 18326 5344 18382 5400
rect 18234 5092 18290 5128
rect 18234 5072 18236 5092
rect 18236 5072 18288 5092
rect 18288 5072 18290 5092
rect 17774 4936 17830 4992
rect 17774 4820 17830 4856
rect 17774 4800 17776 4820
rect 17776 4800 17828 4820
rect 17828 4800 17830 4820
rect 17498 4120 17554 4176
rect 17866 4684 17922 4720
rect 17866 4664 17868 4684
rect 17868 4664 17920 4684
rect 17920 4664 17922 4684
rect 19323 5466 19379 5468
rect 19403 5466 19459 5468
rect 19483 5466 19539 5468
rect 19563 5466 19619 5468
rect 19323 5414 19369 5466
rect 19369 5414 19379 5466
rect 19403 5414 19433 5466
rect 19433 5414 19445 5466
rect 19445 5414 19459 5466
rect 19483 5414 19497 5466
rect 19497 5414 19509 5466
rect 19509 5414 19539 5466
rect 19563 5414 19573 5466
rect 19573 5414 19619 5466
rect 19323 5412 19379 5414
rect 19403 5412 19459 5414
rect 19483 5412 19539 5414
rect 19563 5412 19619 5414
rect 18418 4936 18474 4992
rect 18663 4922 18719 4924
rect 18743 4922 18799 4924
rect 18823 4922 18879 4924
rect 18903 4922 18959 4924
rect 18663 4870 18709 4922
rect 18709 4870 18719 4922
rect 18743 4870 18773 4922
rect 18773 4870 18785 4922
rect 18785 4870 18799 4922
rect 18823 4870 18837 4922
rect 18837 4870 18849 4922
rect 18849 4870 18879 4922
rect 18903 4870 18913 4922
rect 18913 4870 18959 4922
rect 18663 4868 18719 4870
rect 18743 4868 18799 4870
rect 18823 4868 18879 4870
rect 18903 4868 18959 4870
rect 18602 4664 18658 4720
rect 18663 3834 18719 3836
rect 18743 3834 18799 3836
rect 18823 3834 18879 3836
rect 18903 3834 18959 3836
rect 18663 3782 18709 3834
rect 18709 3782 18719 3834
rect 18743 3782 18773 3834
rect 18773 3782 18785 3834
rect 18785 3782 18799 3834
rect 18823 3782 18837 3834
rect 18837 3782 18849 3834
rect 18849 3782 18879 3834
rect 18903 3782 18913 3834
rect 18913 3782 18959 3834
rect 18663 3780 18719 3782
rect 18743 3780 18799 3782
rect 18823 3780 18879 3782
rect 18903 3780 18959 3782
rect 18878 3612 18880 3632
rect 18880 3612 18932 3632
rect 18932 3612 18934 3632
rect 18878 3576 18934 3612
rect 19323 4378 19379 4380
rect 19403 4378 19459 4380
rect 19483 4378 19539 4380
rect 19563 4378 19619 4380
rect 19323 4326 19369 4378
rect 19369 4326 19379 4378
rect 19403 4326 19433 4378
rect 19433 4326 19445 4378
rect 19445 4326 19459 4378
rect 19483 4326 19497 4378
rect 19497 4326 19509 4378
rect 19509 4326 19539 4378
rect 19563 4326 19573 4378
rect 19573 4326 19619 4378
rect 19323 4324 19379 4326
rect 19403 4324 19459 4326
rect 19483 4324 19539 4326
rect 19563 4324 19619 4326
rect 19323 3290 19379 3292
rect 19403 3290 19459 3292
rect 19483 3290 19539 3292
rect 19563 3290 19619 3292
rect 19323 3238 19369 3290
rect 19369 3238 19379 3290
rect 19403 3238 19433 3290
rect 19433 3238 19445 3290
rect 19445 3238 19459 3290
rect 19483 3238 19497 3290
rect 19497 3238 19509 3290
rect 19509 3238 19539 3290
rect 19563 3238 19573 3290
rect 19573 3238 19619 3290
rect 19323 3236 19379 3238
rect 19403 3236 19459 3238
rect 19483 3236 19539 3238
rect 19563 3236 19619 3238
rect 18663 2746 18719 2748
rect 18743 2746 18799 2748
rect 18823 2746 18879 2748
rect 18903 2746 18959 2748
rect 18663 2694 18709 2746
rect 18709 2694 18719 2746
rect 18743 2694 18773 2746
rect 18773 2694 18785 2746
rect 18785 2694 18799 2746
rect 18823 2694 18837 2746
rect 18837 2694 18849 2746
rect 18849 2694 18879 2746
rect 18903 2694 18913 2746
rect 18913 2694 18959 2746
rect 18663 2692 18719 2694
rect 18743 2692 18799 2694
rect 18823 2692 18879 2694
rect 18903 2692 18959 2694
rect 24306 5480 24362 5536
rect 25746 13626 25802 13628
rect 25826 13626 25882 13628
rect 25906 13626 25962 13628
rect 25986 13626 26042 13628
rect 25746 13574 25792 13626
rect 25792 13574 25802 13626
rect 25826 13574 25856 13626
rect 25856 13574 25868 13626
rect 25868 13574 25882 13626
rect 25906 13574 25920 13626
rect 25920 13574 25932 13626
rect 25932 13574 25962 13626
rect 25986 13574 25996 13626
rect 25996 13574 26042 13626
rect 25746 13572 25802 13574
rect 25826 13572 25882 13574
rect 25906 13572 25962 13574
rect 25986 13572 26042 13574
rect 26406 13082 26462 13084
rect 26486 13082 26542 13084
rect 26566 13082 26622 13084
rect 26646 13082 26702 13084
rect 26406 13030 26452 13082
rect 26452 13030 26462 13082
rect 26486 13030 26516 13082
rect 26516 13030 26528 13082
rect 26528 13030 26542 13082
rect 26566 13030 26580 13082
rect 26580 13030 26592 13082
rect 26592 13030 26622 13082
rect 26646 13030 26656 13082
rect 26656 13030 26702 13082
rect 26406 13028 26462 13030
rect 26486 13028 26542 13030
rect 26566 13028 26622 13030
rect 26646 13028 26702 13030
rect 25746 12538 25802 12540
rect 25826 12538 25882 12540
rect 25906 12538 25962 12540
rect 25986 12538 26042 12540
rect 25746 12486 25792 12538
rect 25792 12486 25802 12538
rect 25826 12486 25856 12538
rect 25856 12486 25868 12538
rect 25868 12486 25882 12538
rect 25906 12486 25920 12538
rect 25920 12486 25932 12538
rect 25932 12486 25962 12538
rect 25986 12486 25996 12538
rect 25996 12486 26042 12538
rect 25746 12484 25802 12486
rect 25826 12484 25882 12486
rect 25906 12484 25962 12486
rect 25986 12484 26042 12486
rect 26406 11994 26462 11996
rect 26486 11994 26542 11996
rect 26566 11994 26622 11996
rect 26646 11994 26702 11996
rect 26406 11942 26452 11994
rect 26452 11942 26462 11994
rect 26486 11942 26516 11994
rect 26516 11942 26528 11994
rect 26528 11942 26542 11994
rect 26566 11942 26580 11994
rect 26580 11942 26592 11994
rect 26592 11942 26622 11994
rect 26646 11942 26656 11994
rect 26656 11942 26702 11994
rect 26406 11940 26462 11942
rect 26486 11940 26542 11942
rect 26566 11940 26622 11942
rect 26646 11940 26702 11942
rect 25746 11450 25802 11452
rect 25826 11450 25882 11452
rect 25906 11450 25962 11452
rect 25986 11450 26042 11452
rect 25746 11398 25792 11450
rect 25792 11398 25802 11450
rect 25826 11398 25856 11450
rect 25856 11398 25868 11450
rect 25868 11398 25882 11450
rect 25906 11398 25920 11450
rect 25920 11398 25932 11450
rect 25932 11398 25962 11450
rect 25986 11398 25996 11450
rect 25996 11398 26042 11450
rect 25746 11396 25802 11398
rect 25826 11396 25882 11398
rect 25906 11396 25962 11398
rect 25986 11396 26042 11398
rect 26406 10906 26462 10908
rect 26486 10906 26542 10908
rect 26566 10906 26622 10908
rect 26646 10906 26702 10908
rect 26406 10854 26452 10906
rect 26452 10854 26462 10906
rect 26486 10854 26516 10906
rect 26516 10854 26528 10906
rect 26528 10854 26542 10906
rect 26566 10854 26580 10906
rect 26580 10854 26592 10906
rect 26592 10854 26622 10906
rect 26646 10854 26656 10906
rect 26656 10854 26702 10906
rect 26406 10852 26462 10854
rect 26486 10852 26542 10854
rect 26566 10852 26622 10854
rect 26646 10852 26702 10854
rect 25746 10362 25802 10364
rect 25826 10362 25882 10364
rect 25906 10362 25962 10364
rect 25986 10362 26042 10364
rect 25746 10310 25792 10362
rect 25792 10310 25802 10362
rect 25826 10310 25856 10362
rect 25856 10310 25868 10362
rect 25868 10310 25882 10362
rect 25906 10310 25920 10362
rect 25920 10310 25932 10362
rect 25932 10310 25962 10362
rect 25986 10310 25996 10362
rect 25996 10310 26042 10362
rect 25746 10308 25802 10310
rect 25826 10308 25882 10310
rect 25906 10308 25962 10310
rect 25986 10308 26042 10310
rect 25746 9274 25802 9276
rect 25826 9274 25882 9276
rect 25906 9274 25962 9276
rect 25986 9274 26042 9276
rect 25746 9222 25792 9274
rect 25792 9222 25802 9274
rect 25826 9222 25856 9274
rect 25856 9222 25868 9274
rect 25868 9222 25882 9274
rect 25906 9222 25920 9274
rect 25920 9222 25932 9274
rect 25932 9222 25962 9274
rect 25986 9222 25996 9274
rect 25996 9222 26042 9274
rect 25746 9220 25802 9222
rect 25826 9220 25882 9222
rect 25906 9220 25962 9222
rect 25986 9220 26042 9222
rect 26406 9818 26462 9820
rect 26486 9818 26542 9820
rect 26566 9818 26622 9820
rect 26646 9818 26702 9820
rect 26406 9766 26452 9818
rect 26452 9766 26462 9818
rect 26486 9766 26516 9818
rect 26516 9766 26528 9818
rect 26528 9766 26542 9818
rect 26566 9766 26580 9818
rect 26580 9766 26592 9818
rect 26592 9766 26622 9818
rect 26646 9766 26656 9818
rect 26656 9766 26702 9818
rect 26406 9764 26462 9766
rect 26486 9764 26542 9766
rect 26566 9764 26622 9766
rect 26646 9764 26702 9766
rect 26406 8730 26462 8732
rect 26486 8730 26542 8732
rect 26566 8730 26622 8732
rect 26646 8730 26702 8732
rect 26406 8678 26452 8730
rect 26452 8678 26462 8730
rect 26486 8678 26516 8730
rect 26516 8678 26528 8730
rect 26528 8678 26542 8730
rect 26566 8678 26580 8730
rect 26580 8678 26592 8730
rect 26592 8678 26622 8730
rect 26646 8678 26656 8730
rect 26656 8678 26702 8730
rect 26406 8676 26462 8678
rect 26486 8676 26542 8678
rect 26566 8676 26622 8678
rect 26646 8676 26702 8678
rect 25746 8186 25802 8188
rect 25826 8186 25882 8188
rect 25906 8186 25962 8188
rect 25986 8186 26042 8188
rect 25746 8134 25792 8186
rect 25792 8134 25802 8186
rect 25826 8134 25856 8186
rect 25856 8134 25868 8186
rect 25868 8134 25882 8186
rect 25906 8134 25920 8186
rect 25920 8134 25932 8186
rect 25932 8134 25962 8186
rect 25986 8134 25996 8186
rect 25996 8134 26042 8186
rect 25746 8132 25802 8134
rect 25826 8132 25882 8134
rect 25906 8132 25962 8134
rect 25986 8132 26042 8134
rect 26406 7642 26462 7644
rect 26486 7642 26542 7644
rect 26566 7642 26622 7644
rect 26646 7642 26702 7644
rect 26406 7590 26452 7642
rect 26452 7590 26462 7642
rect 26486 7590 26516 7642
rect 26516 7590 26528 7642
rect 26528 7590 26542 7642
rect 26566 7590 26580 7642
rect 26580 7590 26592 7642
rect 26592 7590 26622 7642
rect 26646 7590 26656 7642
rect 26656 7590 26702 7642
rect 26406 7588 26462 7590
rect 26486 7588 26542 7590
rect 26566 7588 26622 7590
rect 26646 7588 26702 7590
rect 25746 7098 25802 7100
rect 25826 7098 25882 7100
rect 25906 7098 25962 7100
rect 25986 7098 26042 7100
rect 25746 7046 25792 7098
rect 25792 7046 25802 7098
rect 25826 7046 25856 7098
rect 25856 7046 25868 7098
rect 25868 7046 25882 7098
rect 25906 7046 25920 7098
rect 25920 7046 25932 7098
rect 25932 7046 25962 7098
rect 25986 7046 25996 7098
rect 25996 7046 26042 7098
rect 25746 7044 25802 7046
rect 25826 7044 25882 7046
rect 25906 7044 25962 7046
rect 25986 7044 26042 7046
rect 26406 6554 26462 6556
rect 26486 6554 26542 6556
rect 26566 6554 26622 6556
rect 26646 6554 26702 6556
rect 26406 6502 26452 6554
rect 26452 6502 26462 6554
rect 26486 6502 26516 6554
rect 26516 6502 26528 6554
rect 26528 6502 26542 6554
rect 26566 6502 26580 6554
rect 26580 6502 26592 6554
rect 26592 6502 26622 6554
rect 26646 6502 26656 6554
rect 26656 6502 26702 6554
rect 26406 6500 26462 6502
rect 26486 6500 26542 6502
rect 26566 6500 26622 6502
rect 26646 6500 26702 6502
rect 25746 6010 25802 6012
rect 25826 6010 25882 6012
rect 25906 6010 25962 6012
rect 25986 6010 26042 6012
rect 25746 5958 25792 6010
rect 25792 5958 25802 6010
rect 25826 5958 25856 6010
rect 25856 5958 25868 6010
rect 25868 5958 25882 6010
rect 25906 5958 25920 6010
rect 25920 5958 25932 6010
rect 25932 5958 25962 6010
rect 25986 5958 25996 6010
rect 25996 5958 26042 6010
rect 25746 5956 25802 5958
rect 25826 5956 25882 5958
rect 25906 5956 25962 5958
rect 25986 5956 26042 5958
rect 26406 5466 26462 5468
rect 26486 5466 26542 5468
rect 26566 5466 26622 5468
rect 26646 5466 26702 5468
rect 26406 5414 26452 5466
rect 26452 5414 26462 5466
rect 26486 5414 26516 5466
rect 26516 5414 26528 5466
rect 26528 5414 26542 5466
rect 26566 5414 26580 5466
rect 26580 5414 26592 5466
rect 26592 5414 26622 5466
rect 26646 5414 26656 5466
rect 26656 5414 26702 5466
rect 26406 5412 26462 5414
rect 26486 5412 26542 5414
rect 26566 5412 26622 5414
rect 26646 5412 26702 5414
rect 25746 4922 25802 4924
rect 25826 4922 25882 4924
rect 25906 4922 25962 4924
rect 25986 4922 26042 4924
rect 25746 4870 25792 4922
rect 25792 4870 25802 4922
rect 25826 4870 25856 4922
rect 25856 4870 25868 4922
rect 25868 4870 25882 4922
rect 25906 4870 25920 4922
rect 25920 4870 25932 4922
rect 25932 4870 25962 4922
rect 25986 4870 25996 4922
rect 25996 4870 26042 4922
rect 25746 4868 25802 4870
rect 25826 4868 25882 4870
rect 25906 4868 25962 4870
rect 25986 4868 26042 4870
rect 26406 4378 26462 4380
rect 26486 4378 26542 4380
rect 26566 4378 26622 4380
rect 26646 4378 26702 4380
rect 26406 4326 26452 4378
rect 26452 4326 26462 4378
rect 26486 4326 26516 4378
rect 26516 4326 26528 4378
rect 26528 4326 26542 4378
rect 26566 4326 26580 4378
rect 26580 4326 26592 4378
rect 26592 4326 26622 4378
rect 26646 4326 26656 4378
rect 26656 4326 26702 4378
rect 26406 4324 26462 4326
rect 26486 4324 26542 4326
rect 26566 4324 26622 4326
rect 26646 4324 26702 4326
rect 23938 3984 23994 4040
rect 25746 3834 25802 3836
rect 25826 3834 25882 3836
rect 25906 3834 25962 3836
rect 25986 3834 26042 3836
rect 25746 3782 25792 3834
rect 25792 3782 25802 3834
rect 25826 3782 25856 3834
rect 25856 3782 25868 3834
rect 25868 3782 25882 3834
rect 25906 3782 25920 3834
rect 25920 3782 25932 3834
rect 25932 3782 25962 3834
rect 25986 3782 25996 3834
rect 25996 3782 26042 3834
rect 25746 3780 25802 3782
rect 25826 3780 25882 3782
rect 25906 3780 25962 3782
rect 25986 3780 26042 3782
rect 26406 3290 26462 3292
rect 26486 3290 26542 3292
rect 26566 3290 26622 3292
rect 26646 3290 26702 3292
rect 26406 3238 26452 3290
rect 26452 3238 26462 3290
rect 26486 3238 26516 3290
rect 26516 3238 26528 3290
rect 26528 3238 26542 3290
rect 26566 3238 26580 3290
rect 26580 3238 26592 3290
rect 26592 3238 26622 3290
rect 26646 3238 26656 3290
rect 26656 3238 26702 3290
rect 26406 3236 26462 3238
rect 26486 3236 26542 3238
rect 26566 3236 26622 3238
rect 26646 3236 26702 3238
rect 27894 15428 27950 15464
rect 27894 15408 27896 15428
rect 27896 15408 27948 15428
rect 27948 15408 27950 15428
rect 28998 26560 29054 26616
rect 28998 22500 29054 22536
rect 28998 22480 29000 22500
rect 29000 22480 29052 22500
rect 29052 22480 29054 22500
rect 25746 2746 25802 2748
rect 25826 2746 25882 2748
rect 25906 2746 25962 2748
rect 25986 2746 26042 2748
rect 25746 2694 25792 2746
rect 25792 2694 25802 2746
rect 25826 2694 25856 2746
rect 25856 2694 25868 2746
rect 25868 2694 25882 2746
rect 25906 2694 25920 2746
rect 25920 2694 25932 2746
rect 25932 2694 25962 2746
rect 25986 2694 25996 2746
rect 25996 2694 26042 2746
rect 25746 2692 25802 2694
rect 25826 2692 25882 2694
rect 25906 2692 25962 2694
rect 25986 2692 26042 2694
rect 28998 18400 29054 18456
rect 28906 14320 28962 14376
rect 28906 10920 28962 10976
rect 28906 6840 28962 6896
rect 28998 2796 29000 2816
rect 29000 2796 29052 2816
rect 29052 2796 29054 2816
rect 28998 2760 29054 2796
rect 5157 2202 5213 2204
rect 5237 2202 5293 2204
rect 5317 2202 5373 2204
rect 5397 2202 5453 2204
rect 5157 2150 5203 2202
rect 5203 2150 5213 2202
rect 5237 2150 5267 2202
rect 5267 2150 5279 2202
rect 5279 2150 5293 2202
rect 5317 2150 5331 2202
rect 5331 2150 5343 2202
rect 5343 2150 5373 2202
rect 5397 2150 5407 2202
rect 5407 2150 5453 2202
rect 5157 2148 5213 2150
rect 5237 2148 5293 2150
rect 5317 2148 5373 2150
rect 5397 2148 5453 2150
rect 12240 2202 12296 2204
rect 12320 2202 12376 2204
rect 12400 2202 12456 2204
rect 12480 2202 12536 2204
rect 12240 2150 12286 2202
rect 12286 2150 12296 2202
rect 12320 2150 12350 2202
rect 12350 2150 12362 2202
rect 12362 2150 12376 2202
rect 12400 2150 12414 2202
rect 12414 2150 12426 2202
rect 12426 2150 12456 2202
rect 12480 2150 12490 2202
rect 12490 2150 12536 2202
rect 12240 2148 12296 2150
rect 12320 2148 12376 2150
rect 12400 2148 12456 2150
rect 12480 2148 12536 2150
rect 19323 2202 19379 2204
rect 19403 2202 19459 2204
rect 19483 2202 19539 2204
rect 19563 2202 19619 2204
rect 19323 2150 19369 2202
rect 19369 2150 19379 2202
rect 19403 2150 19433 2202
rect 19433 2150 19445 2202
rect 19445 2150 19459 2202
rect 19483 2150 19497 2202
rect 19497 2150 19509 2202
rect 19509 2150 19539 2202
rect 19563 2150 19573 2202
rect 19573 2150 19619 2202
rect 19323 2148 19379 2150
rect 19403 2148 19459 2150
rect 19483 2148 19539 2150
rect 19563 2148 19619 2150
rect 26406 2202 26462 2204
rect 26486 2202 26542 2204
rect 26566 2202 26622 2204
rect 26646 2202 26702 2204
rect 26406 2150 26452 2202
rect 26452 2150 26462 2202
rect 26486 2150 26516 2202
rect 26516 2150 26528 2202
rect 26528 2150 26542 2202
rect 26566 2150 26580 2202
rect 26580 2150 26592 2202
rect 26592 2150 26622 2202
rect 26646 2150 26656 2202
rect 26656 2150 26702 2202
rect 26406 2148 26462 2150
rect 26486 2148 26542 2150
rect 26566 2148 26622 2150
rect 26646 2148 26702 2150
<< metal3 >>
rect 0 31378 800 31408
rect 0 31288 858 31378
rect 798 30970 858 31288
rect 1577 30970 1643 30973
rect 798 30968 1643 30970
rect 798 30912 1582 30968
rect 1638 30912 1643 30968
rect 798 30910 1643 30912
rect 1577 30907 1643 30910
rect 28901 30698 28967 30701
rect 29781 30698 30581 30728
rect 28901 30696 30581 30698
rect 28901 30640 28906 30696
rect 28962 30640 30581 30696
rect 28901 30638 30581 30640
rect 28901 30635 28967 30638
rect 29781 30608 30581 30638
rect 5147 30496 5463 30497
rect 5147 30432 5153 30496
rect 5217 30432 5233 30496
rect 5297 30432 5313 30496
rect 5377 30432 5393 30496
rect 5457 30432 5463 30496
rect 5147 30431 5463 30432
rect 12230 30496 12546 30497
rect 12230 30432 12236 30496
rect 12300 30432 12316 30496
rect 12380 30432 12396 30496
rect 12460 30432 12476 30496
rect 12540 30432 12546 30496
rect 12230 30431 12546 30432
rect 19313 30496 19629 30497
rect 19313 30432 19319 30496
rect 19383 30432 19399 30496
rect 19463 30432 19479 30496
rect 19543 30432 19559 30496
rect 19623 30432 19629 30496
rect 19313 30431 19629 30432
rect 26396 30496 26712 30497
rect 26396 30432 26402 30496
rect 26466 30432 26482 30496
rect 26546 30432 26562 30496
rect 26626 30432 26642 30496
rect 26706 30432 26712 30496
rect 26396 30431 26712 30432
rect 4487 29952 4803 29953
rect 4487 29888 4493 29952
rect 4557 29888 4573 29952
rect 4637 29888 4653 29952
rect 4717 29888 4733 29952
rect 4797 29888 4803 29952
rect 4487 29887 4803 29888
rect 11570 29952 11886 29953
rect 11570 29888 11576 29952
rect 11640 29888 11656 29952
rect 11720 29888 11736 29952
rect 11800 29888 11816 29952
rect 11880 29888 11886 29952
rect 11570 29887 11886 29888
rect 18653 29952 18969 29953
rect 18653 29888 18659 29952
rect 18723 29888 18739 29952
rect 18803 29888 18819 29952
rect 18883 29888 18899 29952
rect 18963 29888 18969 29952
rect 18653 29887 18969 29888
rect 25736 29952 26052 29953
rect 25736 29888 25742 29952
rect 25806 29888 25822 29952
rect 25886 29888 25902 29952
rect 25966 29888 25982 29952
rect 26046 29888 26052 29952
rect 25736 29887 26052 29888
rect 5147 29408 5463 29409
rect 5147 29344 5153 29408
rect 5217 29344 5233 29408
rect 5297 29344 5313 29408
rect 5377 29344 5393 29408
rect 5457 29344 5463 29408
rect 5147 29343 5463 29344
rect 12230 29408 12546 29409
rect 12230 29344 12236 29408
rect 12300 29344 12316 29408
rect 12380 29344 12396 29408
rect 12460 29344 12476 29408
rect 12540 29344 12546 29408
rect 12230 29343 12546 29344
rect 19313 29408 19629 29409
rect 19313 29344 19319 29408
rect 19383 29344 19399 29408
rect 19463 29344 19479 29408
rect 19543 29344 19559 29408
rect 19623 29344 19629 29408
rect 19313 29343 19629 29344
rect 26396 29408 26712 29409
rect 26396 29344 26402 29408
rect 26466 29344 26482 29408
rect 26546 29344 26562 29408
rect 26626 29344 26642 29408
rect 26706 29344 26712 29408
rect 26396 29343 26712 29344
rect 28717 29068 28783 29069
rect 28717 29064 28764 29068
rect 28828 29066 28834 29068
rect 28717 29008 28722 29064
rect 28717 29004 28764 29008
rect 28828 29006 28874 29066
rect 28828 29004 28834 29006
rect 28717 29003 28783 29004
rect 4487 28864 4803 28865
rect 4487 28800 4493 28864
rect 4557 28800 4573 28864
rect 4637 28800 4653 28864
rect 4717 28800 4733 28864
rect 4797 28800 4803 28864
rect 4487 28799 4803 28800
rect 11570 28864 11886 28865
rect 11570 28800 11576 28864
rect 11640 28800 11656 28864
rect 11720 28800 11736 28864
rect 11800 28800 11816 28864
rect 11880 28800 11886 28864
rect 11570 28799 11886 28800
rect 18653 28864 18969 28865
rect 18653 28800 18659 28864
rect 18723 28800 18739 28864
rect 18803 28800 18819 28864
rect 18883 28800 18899 28864
rect 18963 28800 18969 28864
rect 18653 28799 18969 28800
rect 25736 28864 26052 28865
rect 25736 28800 25742 28864
rect 25806 28800 25822 28864
rect 25886 28800 25902 28864
rect 25966 28800 25982 28864
rect 26046 28800 26052 28864
rect 25736 28799 26052 28800
rect 13629 28658 13695 28661
rect 22001 28658 22067 28661
rect 13629 28656 22067 28658
rect 13629 28600 13634 28656
rect 13690 28600 22006 28656
rect 22062 28600 22067 28656
rect 13629 28598 22067 28600
rect 13629 28595 13695 28598
rect 22001 28595 22067 28598
rect 7097 28522 7163 28525
rect 8753 28522 8819 28525
rect 7097 28520 8819 28522
rect 7097 28464 7102 28520
rect 7158 28464 8758 28520
rect 8814 28464 8819 28520
rect 7097 28462 8819 28464
rect 7097 28459 7163 28462
rect 8753 28459 8819 28462
rect 5147 28320 5463 28321
rect 5147 28256 5153 28320
rect 5217 28256 5233 28320
rect 5297 28256 5313 28320
rect 5377 28256 5393 28320
rect 5457 28256 5463 28320
rect 5147 28255 5463 28256
rect 12230 28320 12546 28321
rect 12230 28256 12236 28320
rect 12300 28256 12316 28320
rect 12380 28256 12396 28320
rect 12460 28256 12476 28320
rect 12540 28256 12546 28320
rect 12230 28255 12546 28256
rect 19313 28320 19629 28321
rect 19313 28256 19319 28320
rect 19383 28256 19399 28320
rect 19463 28256 19479 28320
rect 19543 28256 19559 28320
rect 19623 28256 19629 28320
rect 19313 28255 19629 28256
rect 26396 28320 26712 28321
rect 26396 28256 26402 28320
rect 26466 28256 26482 28320
rect 26546 28256 26562 28320
rect 26626 28256 26642 28320
rect 26706 28256 26712 28320
rect 26396 28255 26712 28256
rect 13629 28250 13695 28253
rect 17953 28250 18019 28253
rect 13629 28248 18019 28250
rect 13629 28192 13634 28248
rect 13690 28192 17958 28248
rect 18014 28192 18019 28248
rect 13629 28190 18019 28192
rect 13629 28187 13695 28190
rect 17953 28187 18019 28190
rect 11053 28114 11119 28117
rect 12065 28114 12131 28117
rect 19793 28114 19859 28117
rect 11053 28112 19859 28114
rect 11053 28056 11058 28112
rect 11114 28056 12070 28112
rect 12126 28056 19798 28112
rect 19854 28056 19859 28112
rect 11053 28054 19859 28056
rect 11053 28051 11119 28054
rect 12065 28051 12131 28054
rect 19793 28051 19859 28054
rect 12065 27978 12131 27981
rect 13537 27978 13603 27981
rect 21909 27978 21975 27981
rect 12065 27976 21975 27978
rect 12065 27920 12070 27976
rect 12126 27920 13542 27976
rect 13598 27920 21914 27976
rect 21970 27920 21975 27976
rect 12065 27918 21975 27920
rect 12065 27915 12131 27918
rect 13537 27915 13603 27918
rect 21909 27915 21975 27918
rect 4487 27776 4803 27777
rect 4487 27712 4493 27776
rect 4557 27712 4573 27776
rect 4637 27712 4653 27776
rect 4717 27712 4733 27776
rect 4797 27712 4803 27776
rect 4487 27711 4803 27712
rect 11570 27776 11886 27777
rect 11570 27712 11576 27776
rect 11640 27712 11656 27776
rect 11720 27712 11736 27776
rect 11800 27712 11816 27776
rect 11880 27712 11886 27776
rect 11570 27711 11886 27712
rect 18653 27776 18969 27777
rect 18653 27712 18659 27776
rect 18723 27712 18739 27776
rect 18803 27712 18819 27776
rect 18883 27712 18899 27776
rect 18963 27712 18969 27776
rect 18653 27711 18969 27712
rect 25736 27776 26052 27777
rect 25736 27712 25742 27776
rect 25806 27712 25822 27776
rect 25886 27712 25902 27776
rect 25966 27712 25982 27776
rect 26046 27712 26052 27776
rect 25736 27711 26052 27712
rect 0 27298 800 27328
rect 933 27298 999 27301
rect 0 27296 999 27298
rect 0 27240 938 27296
rect 994 27240 999 27296
rect 0 27238 999 27240
rect 0 27208 800 27238
rect 933 27235 999 27238
rect 5147 27232 5463 27233
rect 5147 27168 5153 27232
rect 5217 27168 5233 27232
rect 5297 27168 5313 27232
rect 5377 27168 5393 27232
rect 5457 27168 5463 27232
rect 5147 27167 5463 27168
rect 12230 27232 12546 27233
rect 12230 27168 12236 27232
rect 12300 27168 12316 27232
rect 12380 27168 12396 27232
rect 12460 27168 12476 27232
rect 12540 27168 12546 27232
rect 12230 27167 12546 27168
rect 19313 27232 19629 27233
rect 19313 27168 19319 27232
rect 19383 27168 19399 27232
rect 19463 27168 19479 27232
rect 19543 27168 19559 27232
rect 19623 27168 19629 27232
rect 19313 27167 19629 27168
rect 26396 27232 26712 27233
rect 26396 27168 26402 27232
rect 26466 27168 26482 27232
rect 26546 27168 26562 27232
rect 26626 27168 26642 27232
rect 26706 27168 26712 27232
rect 26396 27167 26712 27168
rect 4487 26688 4803 26689
rect 4487 26624 4493 26688
rect 4557 26624 4573 26688
rect 4637 26624 4653 26688
rect 4717 26624 4733 26688
rect 4797 26624 4803 26688
rect 4487 26623 4803 26624
rect 11570 26688 11886 26689
rect 11570 26624 11576 26688
rect 11640 26624 11656 26688
rect 11720 26624 11736 26688
rect 11800 26624 11816 26688
rect 11880 26624 11886 26688
rect 11570 26623 11886 26624
rect 18653 26688 18969 26689
rect 18653 26624 18659 26688
rect 18723 26624 18739 26688
rect 18803 26624 18819 26688
rect 18883 26624 18899 26688
rect 18963 26624 18969 26688
rect 18653 26623 18969 26624
rect 25736 26688 26052 26689
rect 25736 26624 25742 26688
rect 25806 26624 25822 26688
rect 25886 26624 25902 26688
rect 25966 26624 25982 26688
rect 26046 26624 26052 26688
rect 25736 26623 26052 26624
rect 28993 26618 29059 26621
rect 29781 26618 30581 26648
rect 28993 26616 30581 26618
rect 28993 26560 28998 26616
rect 29054 26560 30581 26616
rect 28993 26558 30581 26560
rect 28993 26555 29059 26558
rect 29781 26528 30581 26558
rect 5147 26144 5463 26145
rect 5147 26080 5153 26144
rect 5217 26080 5233 26144
rect 5297 26080 5313 26144
rect 5377 26080 5393 26144
rect 5457 26080 5463 26144
rect 5147 26079 5463 26080
rect 12230 26144 12546 26145
rect 12230 26080 12236 26144
rect 12300 26080 12316 26144
rect 12380 26080 12396 26144
rect 12460 26080 12476 26144
rect 12540 26080 12546 26144
rect 12230 26079 12546 26080
rect 19313 26144 19629 26145
rect 19313 26080 19319 26144
rect 19383 26080 19399 26144
rect 19463 26080 19479 26144
rect 19543 26080 19559 26144
rect 19623 26080 19629 26144
rect 19313 26079 19629 26080
rect 26396 26144 26712 26145
rect 26396 26080 26402 26144
rect 26466 26080 26482 26144
rect 26546 26080 26562 26144
rect 26626 26080 26642 26144
rect 26706 26080 26712 26144
rect 26396 26079 26712 26080
rect 4487 25600 4803 25601
rect 4487 25536 4493 25600
rect 4557 25536 4573 25600
rect 4637 25536 4653 25600
rect 4717 25536 4733 25600
rect 4797 25536 4803 25600
rect 4487 25535 4803 25536
rect 11570 25600 11886 25601
rect 11570 25536 11576 25600
rect 11640 25536 11656 25600
rect 11720 25536 11736 25600
rect 11800 25536 11816 25600
rect 11880 25536 11886 25600
rect 11570 25535 11886 25536
rect 18653 25600 18969 25601
rect 18653 25536 18659 25600
rect 18723 25536 18739 25600
rect 18803 25536 18819 25600
rect 18883 25536 18899 25600
rect 18963 25536 18969 25600
rect 18653 25535 18969 25536
rect 25736 25600 26052 25601
rect 25736 25536 25742 25600
rect 25806 25536 25822 25600
rect 25886 25536 25902 25600
rect 25966 25536 25982 25600
rect 26046 25536 26052 25600
rect 25736 25535 26052 25536
rect 5147 25056 5463 25057
rect 5147 24992 5153 25056
rect 5217 24992 5233 25056
rect 5297 24992 5313 25056
rect 5377 24992 5393 25056
rect 5457 24992 5463 25056
rect 5147 24991 5463 24992
rect 12230 25056 12546 25057
rect 12230 24992 12236 25056
rect 12300 24992 12316 25056
rect 12380 24992 12396 25056
rect 12460 24992 12476 25056
rect 12540 24992 12546 25056
rect 12230 24991 12546 24992
rect 19313 25056 19629 25057
rect 19313 24992 19319 25056
rect 19383 24992 19399 25056
rect 19463 24992 19479 25056
rect 19543 24992 19559 25056
rect 19623 24992 19629 25056
rect 19313 24991 19629 24992
rect 26396 25056 26712 25057
rect 26396 24992 26402 25056
rect 26466 24992 26482 25056
rect 26546 24992 26562 25056
rect 26626 24992 26642 25056
rect 26706 24992 26712 25056
rect 26396 24991 26712 24992
rect 4487 24512 4803 24513
rect 4487 24448 4493 24512
rect 4557 24448 4573 24512
rect 4637 24448 4653 24512
rect 4717 24448 4733 24512
rect 4797 24448 4803 24512
rect 4487 24447 4803 24448
rect 11570 24512 11886 24513
rect 11570 24448 11576 24512
rect 11640 24448 11656 24512
rect 11720 24448 11736 24512
rect 11800 24448 11816 24512
rect 11880 24448 11886 24512
rect 11570 24447 11886 24448
rect 18653 24512 18969 24513
rect 18653 24448 18659 24512
rect 18723 24448 18739 24512
rect 18803 24448 18819 24512
rect 18883 24448 18899 24512
rect 18963 24448 18969 24512
rect 18653 24447 18969 24448
rect 25736 24512 26052 24513
rect 25736 24448 25742 24512
rect 25806 24448 25822 24512
rect 25886 24448 25902 24512
rect 25966 24448 25982 24512
rect 26046 24448 26052 24512
rect 25736 24447 26052 24448
rect 15101 24306 15167 24309
rect 16297 24306 16363 24309
rect 15101 24304 16363 24306
rect 15101 24248 15106 24304
rect 15162 24248 16302 24304
rect 16358 24248 16363 24304
rect 15101 24246 16363 24248
rect 15101 24243 15167 24246
rect 16297 24243 16363 24246
rect 5147 23968 5463 23969
rect 5147 23904 5153 23968
rect 5217 23904 5233 23968
rect 5297 23904 5313 23968
rect 5377 23904 5393 23968
rect 5457 23904 5463 23968
rect 5147 23903 5463 23904
rect 12230 23968 12546 23969
rect 12230 23904 12236 23968
rect 12300 23904 12316 23968
rect 12380 23904 12396 23968
rect 12460 23904 12476 23968
rect 12540 23904 12546 23968
rect 12230 23903 12546 23904
rect 19313 23968 19629 23969
rect 19313 23904 19319 23968
rect 19383 23904 19399 23968
rect 19463 23904 19479 23968
rect 19543 23904 19559 23968
rect 19623 23904 19629 23968
rect 19313 23903 19629 23904
rect 26396 23968 26712 23969
rect 26396 23904 26402 23968
rect 26466 23904 26482 23968
rect 26546 23904 26562 23968
rect 26626 23904 26642 23968
rect 26706 23904 26712 23968
rect 26396 23903 26712 23904
rect 1577 23490 1643 23493
rect 798 23488 1643 23490
rect 798 23432 1582 23488
rect 1638 23432 1643 23488
rect 798 23430 1643 23432
rect 798 23248 858 23430
rect 1577 23427 1643 23430
rect 4487 23424 4803 23425
rect 4487 23360 4493 23424
rect 4557 23360 4573 23424
rect 4637 23360 4653 23424
rect 4717 23360 4733 23424
rect 4797 23360 4803 23424
rect 4487 23359 4803 23360
rect 11570 23424 11886 23425
rect 11570 23360 11576 23424
rect 11640 23360 11656 23424
rect 11720 23360 11736 23424
rect 11800 23360 11816 23424
rect 11880 23360 11886 23424
rect 11570 23359 11886 23360
rect 18653 23424 18969 23425
rect 18653 23360 18659 23424
rect 18723 23360 18739 23424
rect 18803 23360 18819 23424
rect 18883 23360 18899 23424
rect 18963 23360 18969 23424
rect 18653 23359 18969 23360
rect 25736 23424 26052 23425
rect 25736 23360 25742 23424
rect 25806 23360 25822 23424
rect 25886 23360 25902 23424
rect 25966 23360 25982 23424
rect 26046 23360 26052 23424
rect 25736 23359 26052 23360
rect 0 23158 858 23248
rect 0 23128 800 23158
rect 1485 23082 1551 23085
rect 21173 23082 21239 23085
rect 1485 23080 21239 23082
rect 1485 23024 1490 23080
rect 1546 23024 21178 23080
rect 21234 23024 21239 23080
rect 1485 23022 21239 23024
rect 1485 23019 1551 23022
rect 21173 23019 21239 23022
rect 5147 22880 5463 22881
rect 5147 22816 5153 22880
rect 5217 22816 5233 22880
rect 5297 22816 5313 22880
rect 5377 22816 5393 22880
rect 5457 22816 5463 22880
rect 5147 22815 5463 22816
rect 12230 22880 12546 22881
rect 12230 22816 12236 22880
rect 12300 22816 12316 22880
rect 12380 22816 12396 22880
rect 12460 22816 12476 22880
rect 12540 22816 12546 22880
rect 12230 22815 12546 22816
rect 19313 22880 19629 22881
rect 19313 22816 19319 22880
rect 19383 22816 19399 22880
rect 19463 22816 19479 22880
rect 19543 22816 19559 22880
rect 19623 22816 19629 22880
rect 19313 22815 19629 22816
rect 26396 22880 26712 22881
rect 26396 22816 26402 22880
rect 26466 22816 26482 22880
rect 26546 22816 26562 22880
rect 26626 22816 26642 22880
rect 26706 22816 26712 22880
rect 26396 22815 26712 22816
rect 24761 22674 24827 22677
rect 24350 22672 24827 22674
rect 24350 22616 24766 22672
rect 24822 22616 24827 22672
rect 24350 22614 24827 22616
rect 24350 22540 24410 22614
rect 24761 22611 24827 22614
rect 24342 22476 24348 22540
rect 24412 22476 24418 22540
rect 28993 22538 29059 22541
rect 29781 22538 30581 22568
rect 28993 22536 30581 22538
rect 28993 22480 28998 22536
rect 29054 22480 30581 22536
rect 28993 22478 30581 22480
rect 28993 22475 29059 22478
rect 29781 22448 30581 22478
rect 23933 22402 23999 22405
rect 24393 22402 24459 22405
rect 23933 22400 24459 22402
rect 23933 22344 23938 22400
rect 23994 22344 24398 22400
rect 24454 22344 24459 22400
rect 23933 22342 24459 22344
rect 23933 22339 23999 22342
rect 24393 22339 24459 22342
rect 4487 22336 4803 22337
rect 4487 22272 4493 22336
rect 4557 22272 4573 22336
rect 4637 22272 4653 22336
rect 4717 22272 4733 22336
rect 4797 22272 4803 22336
rect 4487 22271 4803 22272
rect 11570 22336 11886 22337
rect 11570 22272 11576 22336
rect 11640 22272 11656 22336
rect 11720 22272 11736 22336
rect 11800 22272 11816 22336
rect 11880 22272 11886 22336
rect 11570 22271 11886 22272
rect 18653 22336 18969 22337
rect 18653 22272 18659 22336
rect 18723 22272 18739 22336
rect 18803 22272 18819 22336
rect 18883 22272 18899 22336
rect 18963 22272 18969 22336
rect 18653 22271 18969 22272
rect 25736 22336 26052 22337
rect 25736 22272 25742 22336
rect 25806 22272 25822 22336
rect 25886 22272 25902 22336
rect 25966 22272 25982 22336
rect 26046 22272 26052 22336
rect 25736 22271 26052 22272
rect 22185 22266 22251 22269
rect 23105 22266 23171 22269
rect 24853 22266 24919 22269
rect 22185 22264 24919 22266
rect 22185 22208 22190 22264
rect 22246 22208 23110 22264
rect 23166 22208 24858 22264
rect 24914 22208 24919 22264
rect 22185 22206 24919 22208
rect 22185 22203 22251 22206
rect 23105 22203 23171 22206
rect 24853 22203 24919 22206
rect 6913 22130 6979 22133
rect 10685 22130 10751 22133
rect 6913 22128 10751 22130
rect 6913 22072 6918 22128
rect 6974 22072 10690 22128
rect 10746 22072 10751 22128
rect 6913 22070 10751 22072
rect 6913 22067 6979 22070
rect 10685 22067 10751 22070
rect 5441 21994 5507 21997
rect 6913 21994 6979 21997
rect 5441 21992 6979 21994
rect 5441 21936 5446 21992
rect 5502 21936 6918 21992
rect 6974 21936 6979 21992
rect 5441 21934 6979 21936
rect 5441 21931 5507 21934
rect 6913 21931 6979 21934
rect 9857 21994 9923 21997
rect 17677 21994 17743 21997
rect 26141 21994 26207 21997
rect 9857 21992 10058 21994
rect 9857 21936 9862 21992
rect 9918 21936 10058 21992
rect 9857 21934 10058 21936
rect 9857 21931 9923 21934
rect 5147 21792 5463 21793
rect 5147 21728 5153 21792
rect 5217 21728 5233 21792
rect 5297 21728 5313 21792
rect 5377 21728 5393 21792
rect 5457 21728 5463 21792
rect 5147 21727 5463 21728
rect 5625 21722 5691 21725
rect 8385 21722 8451 21725
rect 5625 21720 8451 21722
rect 5625 21664 5630 21720
rect 5686 21664 8390 21720
rect 8446 21664 8451 21720
rect 5625 21662 8451 21664
rect 5625 21659 5691 21662
rect 8385 21659 8451 21662
rect 4705 21586 4771 21589
rect 7189 21586 7255 21589
rect 4705 21584 7255 21586
rect 4705 21528 4710 21584
rect 4766 21528 7194 21584
rect 7250 21528 7255 21584
rect 4705 21526 7255 21528
rect 9998 21586 10058 21934
rect 17677 21992 26207 21994
rect 17677 21936 17682 21992
rect 17738 21936 26146 21992
rect 26202 21936 26207 21992
rect 17677 21934 26207 21936
rect 17677 21931 17743 21934
rect 26141 21931 26207 21934
rect 20345 21858 20411 21861
rect 25037 21858 25103 21861
rect 20345 21856 25103 21858
rect 20345 21800 20350 21856
rect 20406 21800 25042 21856
rect 25098 21800 25103 21856
rect 20345 21798 25103 21800
rect 20345 21795 20411 21798
rect 25037 21795 25103 21798
rect 12230 21792 12546 21793
rect 12230 21728 12236 21792
rect 12300 21728 12316 21792
rect 12380 21728 12396 21792
rect 12460 21728 12476 21792
rect 12540 21728 12546 21792
rect 12230 21727 12546 21728
rect 19313 21792 19629 21793
rect 19313 21728 19319 21792
rect 19383 21728 19399 21792
rect 19463 21728 19479 21792
rect 19543 21728 19559 21792
rect 19623 21728 19629 21792
rect 19313 21727 19629 21728
rect 26396 21792 26712 21793
rect 26396 21728 26402 21792
rect 26466 21728 26482 21792
rect 26546 21728 26562 21792
rect 26626 21728 26642 21792
rect 26706 21728 26712 21792
rect 26396 21727 26712 21728
rect 21817 21586 21883 21589
rect 23749 21586 23815 21589
rect 9998 21526 12450 21586
rect 4705 21523 4771 21526
rect 7189 21523 7255 21526
rect 12390 21450 12450 21526
rect 21817 21584 23815 21586
rect 21817 21528 21822 21584
rect 21878 21528 23754 21584
rect 23810 21528 23815 21584
rect 21817 21526 23815 21528
rect 21817 21523 21883 21526
rect 23749 21523 23815 21526
rect 27061 21450 27127 21453
rect 12390 21448 27127 21450
rect 12390 21392 27066 21448
rect 27122 21392 27127 21448
rect 12390 21390 27127 21392
rect 27061 21387 27127 21390
rect 4487 21248 4803 21249
rect 4487 21184 4493 21248
rect 4557 21184 4573 21248
rect 4637 21184 4653 21248
rect 4717 21184 4733 21248
rect 4797 21184 4803 21248
rect 4487 21183 4803 21184
rect 11570 21248 11886 21249
rect 11570 21184 11576 21248
rect 11640 21184 11656 21248
rect 11720 21184 11736 21248
rect 11800 21184 11816 21248
rect 11880 21184 11886 21248
rect 11570 21183 11886 21184
rect 18653 21248 18969 21249
rect 18653 21184 18659 21248
rect 18723 21184 18739 21248
rect 18803 21184 18819 21248
rect 18883 21184 18899 21248
rect 18963 21184 18969 21248
rect 18653 21183 18969 21184
rect 25736 21248 26052 21249
rect 25736 21184 25742 21248
rect 25806 21184 25822 21248
rect 25886 21184 25902 21248
rect 25966 21184 25982 21248
rect 26046 21184 26052 21248
rect 25736 21183 26052 21184
rect 22185 21042 22251 21045
rect 22921 21042 22987 21045
rect 22185 21040 22987 21042
rect 22185 20984 22190 21040
rect 22246 20984 22926 21040
rect 22982 20984 22987 21040
rect 22185 20982 22987 20984
rect 22185 20979 22251 20982
rect 22921 20979 22987 20982
rect 19333 20906 19399 20909
rect 19014 20904 19399 20906
rect 19014 20848 19338 20904
rect 19394 20848 19399 20904
rect 19014 20846 19399 20848
rect 5147 20704 5463 20705
rect 5147 20640 5153 20704
rect 5217 20640 5233 20704
rect 5297 20640 5313 20704
rect 5377 20640 5393 20704
rect 5457 20640 5463 20704
rect 5147 20639 5463 20640
rect 12230 20704 12546 20705
rect 12230 20640 12236 20704
rect 12300 20640 12316 20704
rect 12380 20640 12396 20704
rect 12460 20640 12476 20704
rect 12540 20640 12546 20704
rect 12230 20639 12546 20640
rect 18229 20634 18295 20637
rect 19014 20634 19074 20846
rect 19333 20843 19399 20846
rect 19313 20704 19629 20705
rect 19313 20640 19319 20704
rect 19383 20640 19399 20704
rect 19463 20640 19479 20704
rect 19543 20640 19559 20704
rect 19623 20640 19629 20704
rect 19313 20639 19629 20640
rect 26396 20704 26712 20705
rect 26396 20640 26402 20704
rect 26466 20640 26482 20704
rect 26546 20640 26562 20704
rect 26626 20640 26642 20704
rect 26706 20640 26712 20704
rect 26396 20639 26712 20640
rect 18229 20632 19074 20634
rect 18229 20576 18234 20632
rect 18290 20576 19074 20632
rect 18229 20574 19074 20576
rect 18229 20571 18295 20574
rect 12709 20498 12775 20501
rect 19057 20498 19123 20501
rect 12709 20496 19123 20498
rect 12709 20440 12714 20496
rect 12770 20440 19062 20496
rect 19118 20440 19123 20496
rect 12709 20438 19123 20440
rect 12709 20435 12775 20438
rect 19057 20435 19123 20438
rect 4889 20362 4955 20365
rect 9857 20362 9923 20365
rect 4889 20360 9923 20362
rect 4889 20304 4894 20360
rect 4950 20304 9862 20360
rect 9918 20304 9923 20360
rect 4889 20302 9923 20304
rect 4889 20299 4955 20302
rect 9857 20299 9923 20302
rect 10317 20362 10383 20365
rect 15009 20362 15075 20365
rect 10317 20360 15075 20362
rect 10317 20304 10322 20360
rect 10378 20304 15014 20360
rect 15070 20304 15075 20360
rect 10317 20302 15075 20304
rect 10317 20299 10383 20302
rect 15009 20299 15075 20302
rect 4487 20160 4803 20161
rect 4487 20096 4493 20160
rect 4557 20096 4573 20160
rect 4637 20096 4653 20160
rect 4717 20096 4733 20160
rect 4797 20096 4803 20160
rect 4487 20095 4803 20096
rect 11570 20160 11886 20161
rect 11570 20096 11576 20160
rect 11640 20096 11656 20160
rect 11720 20096 11736 20160
rect 11800 20096 11816 20160
rect 11880 20096 11886 20160
rect 11570 20095 11886 20096
rect 18653 20160 18969 20161
rect 18653 20096 18659 20160
rect 18723 20096 18739 20160
rect 18803 20096 18819 20160
rect 18883 20096 18899 20160
rect 18963 20096 18969 20160
rect 18653 20095 18969 20096
rect 25736 20160 26052 20161
rect 25736 20096 25742 20160
rect 25806 20096 25822 20160
rect 25886 20096 25902 20160
rect 25966 20096 25982 20160
rect 26046 20096 26052 20160
rect 25736 20095 26052 20096
rect 10501 19954 10567 19957
rect 15101 19954 15167 19957
rect 10501 19952 15167 19954
rect 10501 19896 10506 19952
rect 10562 19896 15106 19952
rect 15162 19896 15167 19952
rect 10501 19894 15167 19896
rect 10501 19891 10567 19894
rect 15101 19891 15167 19894
rect 0 19818 800 19848
rect 10961 19818 11027 19821
rect 13169 19818 13235 19821
rect 0 19728 858 19818
rect 10961 19816 13235 19818
rect 10961 19760 10966 19816
rect 11022 19760 13174 19816
rect 13230 19760 13235 19816
rect 10961 19758 13235 19760
rect 10961 19755 11027 19758
rect 13169 19755 13235 19758
rect 798 19546 858 19728
rect 5147 19616 5463 19617
rect 5147 19552 5153 19616
rect 5217 19552 5233 19616
rect 5297 19552 5313 19616
rect 5377 19552 5393 19616
rect 5457 19552 5463 19616
rect 5147 19551 5463 19552
rect 12230 19616 12546 19617
rect 12230 19552 12236 19616
rect 12300 19552 12316 19616
rect 12380 19552 12396 19616
rect 12460 19552 12476 19616
rect 12540 19552 12546 19616
rect 12230 19551 12546 19552
rect 19313 19616 19629 19617
rect 19313 19552 19319 19616
rect 19383 19552 19399 19616
rect 19463 19552 19479 19616
rect 19543 19552 19559 19616
rect 19623 19552 19629 19616
rect 19313 19551 19629 19552
rect 26396 19616 26712 19617
rect 26396 19552 26402 19616
rect 26466 19552 26482 19616
rect 26546 19552 26562 19616
rect 26626 19552 26642 19616
rect 26706 19552 26712 19616
rect 26396 19551 26712 19552
rect 1577 19546 1643 19549
rect 798 19544 1643 19546
rect 798 19488 1582 19544
rect 1638 19488 1643 19544
rect 798 19486 1643 19488
rect 1577 19483 1643 19486
rect 18229 19410 18295 19413
rect 19149 19410 19215 19413
rect 19977 19410 20043 19413
rect 18229 19408 20043 19410
rect 18229 19352 18234 19408
rect 18290 19352 19154 19408
rect 19210 19352 19982 19408
rect 20038 19352 20043 19408
rect 18229 19350 20043 19352
rect 18229 19347 18295 19350
rect 19149 19347 19215 19350
rect 19977 19347 20043 19350
rect 13813 19274 13879 19277
rect 17953 19274 18019 19277
rect 13813 19272 18019 19274
rect 13813 19216 13818 19272
rect 13874 19216 17958 19272
rect 18014 19216 18019 19272
rect 13813 19214 18019 19216
rect 13813 19211 13879 19214
rect 17953 19211 18019 19214
rect 18873 19274 18939 19277
rect 20253 19274 20319 19277
rect 18873 19272 20319 19274
rect 18873 19216 18878 19272
rect 18934 19216 20258 19272
rect 20314 19216 20319 19272
rect 18873 19214 20319 19216
rect 18873 19211 18939 19214
rect 20253 19211 20319 19214
rect 4487 19072 4803 19073
rect 4487 19008 4493 19072
rect 4557 19008 4573 19072
rect 4637 19008 4653 19072
rect 4717 19008 4733 19072
rect 4797 19008 4803 19072
rect 4487 19007 4803 19008
rect 11570 19072 11886 19073
rect 11570 19008 11576 19072
rect 11640 19008 11656 19072
rect 11720 19008 11736 19072
rect 11800 19008 11816 19072
rect 11880 19008 11886 19072
rect 11570 19007 11886 19008
rect 18653 19072 18969 19073
rect 18653 19008 18659 19072
rect 18723 19008 18739 19072
rect 18803 19008 18819 19072
rect 18883 19008 18899 19072
rect 18963 19008 18969 19072
rect 18653 19007 18969 19008
rect 25736 19072 26052 19073
rect 25736 19008 25742 19072
rect 25806 19008 25822 19072
rect 25886 19008 25902 19072
rect 25966 19008 25982 19072
rect 26046 19008 26052 19072
rect 25736 19007 26052 19008
rect 5147 18528 5463 18529
rect 5147 18464 5153 18528
rect 5217 18464 5233 18528
rect 5297 18464 5313 18528
rect 5377 18464 5393 18528
rect 5457 18464 5463 18528
rect 5147 18463 5463 18464
rect 12230 18528 12546 18529
rect 12230 18464 12236 18528
rect 12300 18464 12316 18528
rect 12380 18464 12396 18528
rect 12460 18464 12476 18528
rect 12540 18464 12546 18528
rect 12230 18463 12546 18464
rect 19313 18528 19629 18529
rect 19313 18464 19319 18528
rect 19383 18464 19399 18528
rect 19463 18464 19479 18528
rect 19543 18464 19559 18528
rect 19623 18464 19629 18528
rect 19313 18463 19629 18464
rect 26396 18528 26712 18529
rect 26396 18464 26402 18528
rect 26466 18464 26482 18528
rect 26546 18464 26562 18528
rect 26626 18464 26642 18528
rect 26706 18464 26712 18528
rect 26396 18463 26712 18464
rect 28993 18458 29059 18461
rect 29781 18458 30581 18488
rect 28993 18456 30581 18458
rect 28993 18400 28998 18456
rect 29054 18400 30581 18456
rect 28993 18398 30581 18400
rect 28993 18395 29059 18398
rect 29781 18368 30581 18398
rect 27654 17988 27660 18052
rect 27724 18050 27730 18052
rect 27797 18050 27863 18053
rect 27724 18048 27863 18050
rect 27724 17992 27802 18048
rect 27858 17992 27863 18048
rect 27724 17990 27863 17992
rect 27724 17988 27730 17990
rect 27797 17987 27863 17990
rect 4487 17984 4803 17985
rect 4487 17920 4493 17984
rect 4557 17920 4573 17984
rect 4637 17920 4653 17984
rect 4717 17920 4733 17984
rect 4797 17920 4803 17984
rect 4487 17919 4803 17920
rect 11570 17984 11886 17985
rect 11570 17920 11576 17984
rect 11640 17920 11656 17984
rect 11720 17920 11736 17984
rect 11800 17920 11816 17984
rect 11880 17920 11886 17984
rect 11570 17919 11886 17920
rect 18653 17984 18969 17985
rect 18653 17920 18659 17984
rect 18723 17920 18739 17984
rect 18803 17920 18819 17984
rect 18883 17920 18899 17984
rect 18963 17920 18969 17984
rect 18653 17919 18969 17920
rect 25736 17984 26052 17985
rect 25736 17920 25742 17984
rect 25806 17920 25822 17984
rect 25886 17920 25902 17984
rect 25966 17920 25982 17984
rect 26046 17920 26052 17984
rect 25736 17919 26052 17920
rect 4245 17778 4311 17781
rect 7373 17778 7439 17781
rect 4245 17776 7439 17778
rect 4245 17720 4250 17776
rect 4306 17720 7378 17776
rect 7434 17720 7439 17776
rect 4245 17718 7439 17720
rect 4245 17715 4311 17718
rect 7373 17715 7439 17718
rect 19517 17778 19583 17781
rect 25589 17778 25655 17781
rect 19517 17776 25655 17778
rect 19517 17720 19522 17776
rect 19578 17720 25594 17776
rect 25650 17720 25655 17776
rect 19517 17718 25655 17720
rect 19517 17715 19583 17718
rect 25589 17715 25655 17718
rect 7097 17642 7163 17645
rect 19425 17642 19491 17645
rect 7097 17640 19491 17642
rect 7097 17584 7102 17640
rect 7158 17584 19430 17640
rect 19486 17584 19491 17640
rect 7097 17582 19491 17584
rect 7097 17579 7163 17582
rect 19425 17579 19491 17582
rect 5147 17440 5463 17441
rect 5147 17376 5153 17440
rect 5217 17376 5233 17440
rect 5297 17376 5313 17440
rect 5377 17376 5393 17440
rect 5457 17376 5463 17440
rect 5147 17375 5463 17376
rect 12230 17440 12546 17441
rect 12230 17376 12236 17440
rect 12300 17376 12316 17440
rect 12380 17376 12396 17440
rect 12460 17376 12476 17440
rect 12540 17376 12546 17440
rect 12230 17375 12546 17376
rect 19313 17440 19629 17441
rect 19313 17376 19319 17440
rect 19383 17376 19399 17440
rect 19463 17376 19479 17440
rect 19543 17376 19559 17440
rect 19623 17376 19629 17440
rect 19313 17375 19629 17376
rect 26396 17440 26712 17441
rect 26396 17376 26402 17440
rect 26466 17376 26482 17440
rect 26546 17376 26562 17440
rect 26626 17376 26642 17440
rect 26706 17376 26712 17440
rect 26396 17375 26712 17376
rect 24945 17234 25011 17237
rect 27981 17234 28047 17237
rect 24945 17232 28047 17234
rect 24945 17176 24950 17232
rect 25006 17176 27986 17232
rect 28042 17176 28047 17232
rect 24945 17174 28047 17176
rect 24945 17171 25011 17174
rect 27981 17171 28047 17174
rect 26325 17098 26391 17101
rect 27889 17098 27955 17101
rect 26325 17096 27955 17098
rect 26325 17040 26330 17096
rect 26386 17040 27894 17096
rect 27950 17040 27955 17096
rect 26325 17038 27955 17040
rect 26325 17035 26391 17038
rect 27889 17035 27955 17038
rect 4487 16896 4803 16897
rect 4487 16832 4493 16896
rect 4557 16832 4573 16896
rect 4637 16832 4653 16896
rect 4717 16832 4733 16896
rect 4797 16832 4803 16896
rect 4487 16831 4803 16832
rect 11570 16896 11886 16897
rect 11570 16832 11576 16896
rect 11640 16832 11656 16896
rect 11720 16832 11736 16896
rect 11800 16832 11816 16896
rect 11880 16832 11886 16896
rect 11570 16831 11886 16832
rect 18653 16896 18969 16897
rect 18653 16832 18659 16896
rect 18723 16832 18739 16896
rect 18803 16832 18819 16896
rect 18883 16832 18899 16896
rect 18963 16832 18969 16896
rect 18653 16831 18969 16832
rect 25736 16896 26052 16897
rect 25736 16832 25742 16896
rect 25806 16832 25822 16896
rect 25886 16832 25902 16896
rect 25966 16832 25982 16896
rect 26046 16832 26052 16896
rect 25736 16831 26052 16832
rect 5147 16352 5463 16353
rect 5147 16288 5153 16352
rect 5217 16288 5233 16352
rect 5297 16288 5313 16352
rect 5377 16288 5393 16352
rect 5457 16288 5463 16352
rect 5147 16287 5463 16288
rect 12230 16352 12546 16353
rect 12230 16288 12236 16352
rect 12300 16288 12316 16352
rect 12380 16288 12396 16352
rect 12460 16288 12476 16352
rect 12540 16288 12546 16352
rect 12230 16287 12546 16288
rect 19313 16352 19629 16353
rect 19313 16288 19319 16352
rect 19383 16288 19399 16352
rect 19463 16288 19479 16352
rect 19543 16288 19559 16352
rect 19623 16288 19629 16352
rect 19313 16287 19629 16288
rect 26396 16352 26712 16353
rect 26396 16288 26402 16352
rect 26466 16288 26482 16352
rect 26546 16288 26562 16352
rect 26626 16288 26642 16352
rect 26706 16288 26712 16352
rect 26396 16287 26712 16288
rect 4487 15808 4803 15809
rect 0 15738 800 15768
rect 4487 15744 4493 15808
rect 4557 15744 4573 15808
rect 4637 15744 4653 15808
rect 4717 15744 4733 15808
rect 4797 15744 4803 15808
rect 4487 15743 4803 15744
rect 11570 15808 11886 15809
rect 11570 15744 11576 15808
rect 11640 15744 11656 15808
rect 11720 15744 11736 15808
rect 11800 15744 11816 15808
rect 11880 15744 11886 15808
rect 11570 15743 11886 15744
rect 18653 15808 18969 15809
rect 18653 15744 18659 15808
rect 18723 15744 18739 15808
rect 18803 15744 18819 15808
rect 18883 15744 18899 15808
rect 18963 15744 18969 15808
rect 18653 15743 18969 15744
rect 25736 15808 26052 15809
rect 25736 15744 25742 15808
rect 25806 15744 25822 15808
rect 25886 15744 25902 15808
rect 25966 15744 25982 15808
rect 26046 15744 26052 15808
rect 25736 15743 26052 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 10501 15602 10567 15605
rect 14089 15602 14155 15605
rect 10501 15600 14155 15602
rect 10501 15544 10506 15600
rect 10562 15544 14094 15600
rect 14150 15544 14155 15600
rect 10501 15542 14155 15544
rect 10501 15539 10567 15542
rect 14089 15539 14155 15542
rect 11973 15466 12039 15469
rect 13537 15466 13603 15469
rect 11973 15464 13603 15466
rect 11973 15408 11978 15464
rect 12034 15408 13542 15464
rect 13598 15408 13603 15464
rect 11973 15406 13603 15408
rect 11973 15403 12039 15406
rect 13537 15403 13603 15406
rect 26601 15466 26667 15469
rect 27889 15466 27955 15469
rect 26601 15464 27955 15466
rect 26601 15408 26606 15464
rect 26662 15408 27894 15464
rect 27950 15408 27955 15464
rect 26601 15406 27955 15408
rect 26601 15403 26667 15406
rect 27889 15403 27955 15406
rect 5147 15264 5463 15265
rect 5147 15200 5153 15264
rect 5217 15200 5233 15264
rect 5297 15200 5313 15264
rect 5377 15200 5393 15264
rect 5457 15200 5463 15264
rect 5147 15199 5463 15200
rect 12230 15264 12546 15265
rect 12230 15200 12236 15264
rect 12300 15200 12316 15264
rect 12380 15200 12396 15264
rect 12460 15200 12476 15264
rect 12540 15200 12546 15264
rect 12230 15199 12546 15200
rect 19313 15264 19629 15265
rect 19313 15200 19319 15264
rect 19383 15200 19399 15264
rect 19463 15200 19479 15264
rect 19543 15200 19559 15264
rect 19623 15200 19629 15264
rect 19313 15199 19629 15200
rect 26396 15264 26712 15265
rect 26396 15200 26402 15264
rect 26466 15200 26482 15264
rect 26546 15200 26562 15264
rect 26626 15200 26642 15264
rect 26706 15200 26712 15264
rect 26396 15199 26712 15200
rect 4487 14720 4803 14721
rect 4487 14656 4493 14720
rect 4557 14656 4573 14720
rect 4637 14656 4653 14720
rect 4717 14656 4733 14720
rect 4797 14656 4803 14720
rect 4487 14655 4803 14656
rect 11570 14720 11886 14721
rect 11570 14656 11576 14720
rect 11640 14656 11656 14720
rect 11720 14656 11736 14720
rect 11800 14656 11816 14720
rect 11880 14656 11886 14720
rect 11570 14655 11886 14656
rect 18653 14720 18969 14721
rect 18653 14656 18659 14720
rect 18723 14656 18739 14720
rect 18803 14656 18819 14720
rect 18883 14656 18899 14720
rect 18963 14656 18969 14720
rect 18653 14655 18969 14656
rect 25736 14720 26052 14721
rect 25736 14656 25742 14720
rect 25806 14656 25822 14720
rect 25886 14656 25902 14720
rect 25966 14656 25982 14720
rect 26046 14656 26052 14720
rect 25736 14655 26052 14656
rect 10501 14514 10567 14517
rect 12157 14514 12223 14517
rect 10501 14512 12223 14514
rect 10501 14456 10506 14512
rect 10562 14456 12162 14512
rect 12218 14456 12223 14512
rect 10501 14454 12223 14456
rect 10501 14451 10567 14454
rect 12157 14451 12223 14454
rect 19057 14378 19123 14381
rect 20897 14378 20963 14381
rect 19057 14376 20963 14378
rect 19057 14320 19062 14376
rect 19118 14320 20902 14376
rect 20958 14320 20963 14376
rect 19057 14318 20963 14320
rect 19057 14315 19123 14318
rect 20897 14315 20963 14318
rect 28901 14378 28967 14381
rect 29781 14378 30581 14408
rect 28901 14376 30581 14378
rect 28901 14320 28906 14376
rect 28962 14320 30581 14376
rect 28901 14318 30581 14320
rect 28901 14315 28967 14318
rect 29781 14288 30581 14318
rect 5147 14176 5463 14177
rect 5147 14112 5153 14176
rect 5217 14112 5233 14176
rect 5297 14112 5313 14176
rect 5377 14112 5393 14176
rect 5457 14112 5463 14176
rect 5147 14111 5463 14112
rect 12230 14176 12546 14177
rect 12230 14112 12236 14176
rect 12300 14112 12316 14176
rect 12380 14112 12396 14176
rect 12460 14112 12476 14176
rect 12540 14112 12546 14176
rect 12230 14111 12546 14112
rect 19313 14176 19629 14177
rect 19313 14112 19319 14176
rect 19383 14112 19399 14176
rect 19463 14112 19479 14176
rect 19543 14112 19559 14176
rect 19623 14112 19629 14176
rect 19313 14111 19629 14112
rect 26396 14176 26712 14177
rect 26396 14112 26402 14176
rect 26466 14112 26482 14176
rect 26546 14112 26562 14176
rect 26626 14112 26642 14176
rect 26706 14112 26712 14176
rect 26396 14111 26712 14112
rect 19701 14106 19767 14109
rect 20161 14106 20227 14109
rect 19701 14104 20227 14106
rect 19701 14048 19706 14104
rect 19762 14048 20166 14104
rect 20222 14048 20227 14104
rect 19701 14046 20227 14048
rect 19701 14043 19767 14046
rect 20161 14043 20227 14046
rect 10501 13836 10567 13837
rect 10501 13834 10548 13836
rect 10456 13832 10548 13834
rect 10456 13776 10506 13832
rect 10456 13774 10548 13776
rect 10501 13772 10548 13774
rect 10612 13772 10618 13836
rect 10501 13771 10567 13772
rect 4487 13632 4803 13633
rect 4487 13568 4493 13632
rect 4557 13568 4573 13632
rect 4637 13568 4653 13632
rect 4717 13568 4733 13632
rect 4797 13568 4803 13632
rect 4487 13567 4803 13568
rect 11570 13632 11886 13633
rect 11570 13568 11576 13632
rect 11640 13568 11656 13632
rect 11720 13568 11736 13632
rect 11800 13568 11816 13632
rect 11880 13568 11886 13632
rect 11570 13567 11886 13568
rect 18653 13632 18969 13633
rect 18653 13568 18659 13632
rect 18723 13568 18739 13632
rect 18803 13568 18819 13632
rect 18883 13568 18899 13632
rect 18963 13568 18969 13632
rect 18653 13567 18969 13568
rect 25736 13632 26052 13633
rect 25736 13568 25742 13632
rect 25806 13568 25822 13632
rect 25886 13568 25902 13632
rect 25966 13568 25982 13632
rect 26046 13568 26052 13632
rect 25736 13567 26052 13568
rect 10225 13426 10291 13429
rect 10225 13424 10794 13426
rect 10225 13368 10230 13424
rect 10286 13368 10794 13424
rect 10225 13366 10794 13368
rect 10225 13363 10291 13366
rect 10734 13292 10794 13366
rect 10726 13228 10732 13292
rect 10796 13290 10802 13292
rect 11513 13290 11579 13293
rect 10796 13288 11579 13290
rect 10796 13232 11518 13288
rect 11574 13232 11579 13288
rect 10796 13230 11579 13232
rect 10796 13228 10802 13230
rect 11513 13227 11579 13230
rect 5147 13088 5463 13089
rect 5147 13024 5153 13088
rect 5217 13024 5233 13088
rect 5297 13024 5313 13088
rect 5377 13024 5393 13088
rect 5457 13024 5463 13088
rect 5147 13023 5463 13024
rect 12230 13088 12546 13089
rect 12230 13024 12236 13088
rect 12300 13024 12316 13088
rect 12380 13024 12396 13088
rect 12460 13024 12476 13088
rect 12540 13024 12546 13088
rect 12230 13023 12546 13024
rect 19313 13088 19629 13089
rect 19313 13024 19319 13088
rect 19383 13024 19399 13088
rect 19463 13024 19479 13088
rect 19543 13024 19559 13088
rect 19623 13024 19629 13088
rect 19313 13023 19629 13024
rect 26396 13088 26712 13089
rect 26396 13024 26402 13088
rect 26466 13024 26482 13088
rect 26546 13024 26562 13088
rect 26626 13024 26642 13088
rect 26706 13024 26712 13088
rect 26396 13023 26712 13024
rect 16113 12746 16179 12749
rect 19057 12746 19123 12749
rect 16113 12744 19123 12746
rect 16113 12688 16118 12744
rect 16174 12688 19062 12744
rect 19118 12688 19123 12744
rect 16113 12686 19123 12688
rect 16113 12683 16179 12686
rect 19057 12683 19123 12686
rect 4487 12544 4803 12545
rect 4487 12480 4493 12544
rect 4557 12480 4573 12544
rect 4637 12480 4653 12544
rect 4717 12480 4733 12544
rect 4797 12480 4803 12544
rect 4487 12479 4803 12480
rect 11570 12544 11886 12545
rect 11570 12480 11576 12544
rect 11640 12480 11656 12544
rect 11720 12480 11736 12544
rect 11800 12480 11816 12544
rect 11880 12480 11886 12544
rect 11570 12479 11886 12480
rect 18653 12544 18969 12545
rect 18653 12480 18659 12544
rect 18723 12480 18739 12544
rect 18803 12480 18819 12544
rect 18883 12480 18899 12544
rect 18963 12480 18969 12544
rect 18653 12479 18969 12480
rect 25736 12544 26052 12545
rect 25736 12480 25742 12544
rect 25806 12480 25822 12544
rect 25886 12480 25902 12544
rect 25966 12480 25982 12544
rect 26046 12480 26052 12544
rect 25736 12479 26052 12480
rect 3049 12338 3115 12341
rect 14273 12338 14339 12341
rect 16665 12338 16731 12341
rect 3049 12336 16731 12338
rect 3049 12280 3054 12336
rect 3110 12280 14278 12336
rect 14334 12280 16670 12336
rect 16726 12280 16731 12336
rect 3049 12278 16731 12280
rect 3049 12275 3115 12278
rect 14273 12275 14339 12278
rect 16665 12275 16731 12278
rect 14089 12202 14155 12205
rect 18229 12202 18295 12205
rect 14089 12200 18295 12202
rect 14089 12144 14094 12200
rect 14150 12144 18234 12200
rect 18290 12144 18295 12200
rect 14089 12142 18295 12144
rect 14089 12139 14155 12142
rect 18229 12139 18295 12142
rect 5147 12000 5463 12001
rect 5147 11936 5153 12000
rect 5217 11936 5233 12000
rect 5297 11936 5313 12000
rect 5377 11936 5393 12000
rect 5457 11936 5463 12000
rect 5147 11935 5463 11936
rect 12230 12000 12546 12001
rect 12230 11936 12236 12000
rect 12300 11936 12316 12000
rect 12380 11936 12396 12000
rect 12460 11936 12476 12000
rect 12540 11936 12546 12000
rect 12230 11935 12546 11936
rect 19313 12000 19629 12001
rect 19313 11936 19319 12000
rect 19383 11936 19399 12000
rect 19463 11936 19479 12000
rect 19543 11936 19559 12000
rect 19623 11936 19629 12000
rect 19313 11935 19629 11936
rect 26396 12000 26712 12001
rect 26396 11936 26402 12000
rect 26466 11936 26482 12000
rect 26546 11936 26562 12000
rect 26626 11936 26642 12000
rect 26706 11936 26712 12000
rect 26396 11935 26712 11936
rect 2221 11794 2287 11797
rect 27654 11794 27660 11796
rect 2221 11792 27660 11794
rect 2221 11736 2226 11792
rect 2282 11736 27660 11792
rect 2221 11734 27660 11736
rect 2221 11731 2287 11734
rect 27654 11732 27660 11734
rect 27724 11732 27730 11796
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 4487 11456 4803 11457
rect 4487 11392 4493 11456
rect 4557 11392 4573 11456
rect 4637 11392 4653 11456
rect 4717 11392 4733 11456
rect 4797 11392 4803 11456
rect 4487 11391 4803 11392
rect 11570 11456 11886 11457
rect 11570 11392 11576 11456
rect 11640 11392 11656 11456
rect 11720 11392 11736 11456
rect 11800 11392 11816 11456
rect 11880 11392 11886 11456
rect 11570 11391 11886 11392
rect 18653 11456 18969 11457
rect 18653 11392 18659 11456
rect 18723 11392 18739 11456
rect 18803 11392 18819 11456
rect 18883 11392 18899 11456
rect 18963 11392 18969 11456
rect 18653 11391 18969 11392
rect 25736 11456 26052 11457
rect 25736 11392 25742 11456
rect 25806 11392 25822 11456
rect 25886 11392 25902 11456
rect 25966 11392 25982 11456
rect 26046 11392 26052 11456
rect 25736 11391 26052 11392
rect 3693 11386 3759 11389
rect 4245 11386 4311 11389
rect 3693 11384 4311 11386
rect 3693 11328 3698 11384
rect 3754 11328 4250 11384
rect 4306 11328 4311 11384
rect 3693 11326 4311 11328
rect 3693 11323 3759 11326
rect 4245 11323 4311 11326
rect 3877 11250 3943 11253
rect 4889 11250 4955 11253
rect 7557 11250 7623 11253
rect 3877 11248 7623 11250
rect 3877 11192 3882 11248
rect 3938 11192 4894 11248
rect 4950 11192 7562 11248
rect 7618 11192 7623 11248
rect 3877 11190 7623 11192
rect 3877 11187 3943 11190
rect 4889 11187 4955 11190
rect 7557 11187 7623 11190
rect 3141 11114 3207 11117
rect 6177 11114 6243 11117
rect 3141 11112 6243 11114
rect 3141 11056 3146 11112
rect 3202 11056 6182 11112
rect 6238 11056 6243 11112
rect 3141 11054 6243 11056
rect 3141 11051 3207 11054
rect 6177 11051 6243 11054
rect 28901 10978 28967 10981
rect 29781 10978 30581 11008
rect 28901 10976 30581 10978
rect 28901 10920 28906 10976
rect 28962 10920 30581 10976
rect 28901 10918 30581 10920
rect 28901 10915 28967 10918
rect 5147 10912 5463 10913
rect 5147 10848 5153 10912
rect 5217 10848 5233 10912
rect 5297 10848 5313 10912
rect 5377 10848 5393 10912
rect 5457 10848 5463 10912
rect 5147 10847 5463 10848
rect 12230 10912 12546 10913
rect 12230 10848 12236 10912
rect 12300 10848 12316 10912
rect 12380 10848 12396 10912
rect 12460 10848 12476 10912
rect 12540 10848 12546 10912
rect 12230 10847 12546 10848
rect 19313 10912 19629 10913
rect 19313 10848 19319 10912
rect 19383 10848 19399 10912
rect 19463 10848 19479 10912
rect 19543 10848 19559 10912
rect 19623 10848 19629 10912
rect 19313 10847 19629 10848
rect 26396 10912 26712 10913
rect 26396 10848 26402 10912
rect 26466 10848 26482 10912
rect 26546 10848 26562 10912
rect 26626 10848 26642 10912
rect 26706 10848 26712 10912
rect 29781 10888 30581 10918
rect 26396 10847 26712 10848
rect 4061 10842 4127 10845
rect 4981 10842 5047 10845
rect 4061 10840 5047 10842
rect 4061 10784 4066 10840
rect 4122 10784 4986 10840
rect 5042 10784 5047 10840
rect 4061 10782 5047 10784
rect 4061 10779 4127 10782
rect 4981 10779 5047 10782
rect 12617 10842 12683 10845
rect 18965 10842 19031 10845
rect 12617 10840 19031 10842
rect 12617 10784 12622 10840
rect 12678 10784 18970 10840
rect 19026 10784 19031 10840
rect 12617 10782 19031 10784
rect 12617 10779 12683 10782
rect 18965 10779 19031 10782
rect 2129 10706 2195 10709
rect 5257 10706 5323 10709
rect 2129 10704 5323 10706
rect 2129 10648 2134 10704
rect 2190 10648 5262 10704
rect 5318 10648 5323 10704
rect 2129 10646 5323 10648
rect 2129 10643 2195 10646
rect 5257 10643 5323 10646
rect 13261 10706 13327 10709
rect 18689 10706 18755 10709
rect 13261 10704 18755 10706
rect 13261 10648 13266 10704
rect 13322 10648 18694 10704
rect 18750 10648 18755 10704
rect 13261 10646 18755 10648
rect 13261 10643 13327 10646
rect 18689 10643 18755 10646
rect 4245 10570 4311 10573
rect 4613 10570 4679 10573
rect 4245 10568 4679 10570
rect 4245 10512 4250 10568
rect 4306 10512 4618 10568
rect 4674 10512 4679 10568
rect 4245 10510 4679 10512
rect 4245 10507 4311 10510
rect 4613 10507 4679 10510
rect 11329 10570 11395 10573
rect 18873 10570 18939 10573
rect 11329 10568 18939 10570
rect 11329 10512 11334 10568
rect 11390 10512 18878 10568
rect 18934 10512 18939 10568
rect 11329 10510 18939 10512
rect 11329 10507 11395 10510
rect 18873 10507 18939 10510
rect 4487 10368 4803 10369
rect 4487 10304 4493 10368
rect 4557 10304 4573 10368
rect 4637 10304 4653 10368
rect 4717 10304 4733 10368
rect 4797 10304 4803 10368
rect 4487 10303 4803 10304
rect 11570 10368 11886 10369
rect 11570 10304 11576 10368
rect 11640 10304 11656 10368
rect 11720 10304 11736 10368
rect 11800 10304 11816 10368
rect 11880 10304 11886 10368
rect 11570 10303 11886 10304
rect 18653 10368 18969 10369
rect 18653 10304 18659 10368
rect 18723 10304 18739 10368
rect 18803 10304 18819 10368
rect 18883 10304 18899 10368
rect 18963 10304 18969 10368
rect 18653 10303 18969 10304
rect 25736 10368 26052 10369
rect 25736 10304 25742 10368
rect 25806 10304 25822 10368
rect 25886 10304 25902 10368
rect 25966 10304 25982 10368
rect 26046 10304 26052 10368
rect 25736 10303 26052 10304
rect 19793 10298 19859 10301
rect 22921 10298 22987 10301
rect 19793 10296 22987 10298
rect 19793 10240 19798 10296
rect 19854 10240 22926 10296
rect 22982 10240 22987 10296
rect 19793 10238 22987 10240
rect 19793 10235 19859 10238
rect 22921 10235 22987 10238
rect 13353 10026 13419 10029
rect 23105 10026 23171 10029
rect 13353 10024 23171 10026
rect 13353 9968 13358 10024
rect 13414 9968 23110 10024
rect 23166 9968 23171 10024
rect 13353 9966 23171 9968
rect 13353 9963 13419 9966
rect 23105 9963 23171 9966
rect 9949 9890 10015 9893
rect 11329 9890 11395 9893
rect 9949 9888 11395 9890
rect 9949 9832 9954 9888
rect 10010 9832 11334 9888
rect 11390 9832 11395 9888
rect 9949 9830 11395 9832
rect 9949 9827 10015 9830
rect 11329 9827 11395 9830
rect 5147 9824 5463 9825
rect 5147 9760 5153 9824
rect 5217 9760 5233 9824
rect 5297 9760 5313 9824
rect 5377 9760 5393 9824
rect 5457 9760 5463 9824
rect 5147 9759 5463 9760
rect 12230 9824 12546 9825
rect 12230 9760 12236 9824
rect 12300 9760 12316 9824
rect 12380 9760 12396 9824
rect 12460 9760 12476 9824
rect 12540 9760 12546 9824
rect 12230 9759 12546 9760
rect 19313 9824 19629 9825
rect 19313 9760 19319 9824
rect 19383 9760 19399 9824
rect 19463 9760 19479 9824
rect 19543 9760 19559 9824
rect 19623 9760 19629 9824
rect 19313 9759 19629 9760
rect 26396 9824 26712 9825
rect 26396 9760 26402 9824
rect 26466 9760 26482 9824
rect 26546 9760 26562 9824
rect 26626 9760 26642 9824
rect 26706 9760 26712 9824
rect 26396 9759 26712 9760
rect 5441 9618 5507 9621
rect 12157 9618 12223 9621
rect 5441 9616 12223 9618
rect 5441 9560 5446 9616
rect 5502 9560 12162 9616
rect 12218 9560 12223 9616
rect 5441 9558 12223 9560
rect 5441 9555 5507 9558
rect 12157 9555 12223 9558
rect 13169 9618 13235 9621
rect 16021 9618 16087 9621
rect 13169 9616 16087 9618
rect 13169 9560 13174 9616
rect 13230 9560 16026 9616
rect 16082 9560 16087 9616
rect 13169 9558 16087 9560
rect 13169 9555 13235 9558
rect 16021 9555 16087 9558
rect 17769 9618 17835 9621
rect 18965 9618 19031 9621
rect 17769 9616 19031 9618
rect 17769 9560 17774 9616
rect 17830 9560 18970 9616
rect 19026 9560 19031 9616
rect 17769 9558 19031 9560
rect 17769 9555 17835 9558
rect 18965 9555 19031 9558
rect 8845 9482 8911 9485
rect 18413 9482 18479 9485
rect 8845 9480 18479 9482
rect 8845 9424 8850 9480
rect 8906 9424 18418 9480
rect 18474 9424 18479 9480
rect 8845 9422 18479 9424
rect 8845 9419 8911 9422
rect 18413 9419 18479 9422
rect 17033 9346 17099 9349
rect 18321 9346 18387 9349
rect 17033 9344 18387 9346
rect 17033 9288 17038 9344
rect 17094 9288 18326 9344
rect 18382 9288 18387 9344
rect 17033 9286 18387 9288
rect 17033 9283 17099 9286
rect 18321 9283 18387 9286
rect 4487 9280 4803 9281
rect 4487 9216 4493 9280
rect 4557 9216 4573 9280
rect 4637 9216 4653 9280
rect 4717 9216 4733 9280
rect 4797 9216 4803 9280
rect 4487 9215 4803 9216
rect 11570 9280 11886 9281
rect 11570 9216 11576 9280
rect 11640 9216 11656 9280
rect 11720 9216 11736 9280
rect 11800 9216 11816 9280
rect 11880 9216 11886 9280
rect 11570 9215 11886 9216
rect 18653 9280 18969 9281
rect 18653 9216 18659 9280
rect 18723 9216 18739 9280
rect 18803 9216 18819 9280
rect 18883 9216 18899 9280
rect 18963 9216 18969 9280
rect 18653 9215 18969 9216
rect 25736 9280 26052 9281
rect 25736 9216 25742 9280
rect 25806 9216 25822 9280
rect 25886 9216 25902 9280
rect 25966 9216 25982 9280
rect 26046 9216 26052 9280
rect 25736 9215 26052 9216
rect 9949 9074 10015 9077
rect 11237 9074 11303 9077
rect 9949 9072 11303 9074
rect 9949 9016 9954 9072
rect 10010 9016 11242 9072
rect 11298 9016 11303 9072
rect 9949 9014 11303 9016
rect 9949 9011 10015 9014
rect 11237 9011 11303 9014
rect 5147 8736 5463 8737
rect 5147 8672 5153 8736
rect 5217 8672 5233 8736
rect 5297 8672 5313 8736
rect 5377 8672 5393 8736
rect 5457 8672 5463 8736
rect 5147 8671 5463 8672
rect 12230 8736 12546 8737
rect 12230 8672 12236 8736
rect 12300 8672 12316 8736
rect 12380 8672 12396 8736
rect 12460 8672 12476 8736
rect 12540 8672 12546 8736
rect 12230 8671 12546 8672
rect 19313 8736 19629 8737
rect 19313 8672 19319 8736
rect 19383 8672 19399 8736
rect 19463 8672 19479 8736
rect 19543 8672 19559 8736
rect 19623 8672 19629 8736
rect 19313 8671 19629 8672
rect 26396 8736 26712 8737
rect 26396 8672 26402 8736
rect 26466 8672 26482 8736
rect 26546 8672 26562 8736
rect 26626 8672 26642 8736
rect 26706 8672 26712 8736
rect 26396 8671 26712 8672
rect 5441 8530 5507 8533
rect 9029 8530 9095 8533
rect 5441 8528 9095 8530
rect 5441 8472 5446 8528
rect 5502 8472 9034 8528
rect 9090 8472 9095 8528
rect 5441 8470 9095 8472
rect 5441 8467 5507 8470
rect 9029 8467 9095 8470
rect 10542 8196 10548 8260
rect 10612 8258 10618 8260
rect 10777 8258 10843 8261
rect 10612 8256 10843 8258
rect 10612 8200 10782 8256
rect 10838 8200 10843 8256
rect 10612 8198 10843 8200
rect 10612 8196 10618 8198
rect 10777 8195 10843 8198
rect 4487 8192 4803 8193
rect 4487 8128 4493 8192
rect 4557 8128 4573 8192
rect 4637 8128 4653 8192
rect 4717 8128 4733 8192
rect 4797 8128 4803 8192
rect 4487 8127 4803 8128
rect 11570 8192 11886 8193
rect 11570 8128 11576 8192
rect 11640 8128 11656 8192
rect 11720 8128 11736 8192
rect 11800 8128 11816 8192
rect 11880 8128 11886 8192
rect 11570 8127 11886 8128
rect 18653 8192 18969 8193
rect 18653 8128 18659 8192
rect 18723 8128 18739 8192
rect 18803 8128 18819 8192
rect 18883 8128 18899 8192
rect 18963 8128 18969 8192
rect 18653 8127 18969 8128
rect 25736 8192 26052 8193
rect 25736 8128 25742 8192
rect 25806 8128 25822 8192
rect 25886 8128 25902 8192
rect 25966 8128 25982 8192
rect 26046 8128 26052 8192
rect 25736 8127 26052 8128
rect 10593 8122 10659 8125
rect 10726 8122 10732 8124
rect 10593 8120 10732 8122
rect 10593 8064 10598 8120
rect 10654 8064 10732 8120
rect 10593 8062 10732 8064
rect 10593 8059 10659 8062
rect 10726 8060 10732 8062
rect 10796 8060 10802 8124
rect 17401 7986 17467 7989
rect 22645 7986 22711 7989
rect 17401 7984 22711 7986
rect 17401 7928 17406 7984
rect 17462 7928 22650 7984
rect 22706 7928 22711 7984
rect 17401 7926 22711 7928
rect 17401 7923 17467 7926
rect 22645 7923 22711 7926
rect 17401 7714 17467 7717
rect 17953 7714 18019 7717
rect 17401 7712 18019 7714
rect 17401 7656 17406 7712
rect 17462 7656 17958 7712
rect 18014 7656 18019 7712
rect 17401 7654 18019 7656
rect 17401 7651 17467 7654
rect 17953 7651 18019 7654
rect 5147 7648 5463 7649
rect 0 7578 800 7608
rect 5147 7584 5153 7648
rect 5217 7584 5233 7648
rect 5297 7584 5313 7648
rect 5377 7584 5393 7648
rect 5457 7584 5463 7648
rect 5147 7583 5463 7584
rect 12230 7648 12546 7649
rect 12230 7584 12236 7648
rect 12300 7584 12316 7648
rect 12380 7584 12396 7648
rect 12460 7584 12476 7648
rect 12540 7584 12546 7648
rect 12230 7583 12546 7584
rect 19313 7648 19629 7649
rect 19313 7584 19319 7648
rect 19383 7584 19399 7648
rect 19463 7584 19479 7648
rect 19543 7584 19559 7648
rect 19623 7584 19629 7648
rect 19313 7583 19629 7584
rect 26396 7648 26712 7649
rect 26396 7584 26402 7648
rect 26466 7584 26482 7648
rect 26546 7584 26562 7648
rect 26626 7584 26642 7648
rect 26706 7584 26712 7648
rect 26396 7583 26712 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 800 7518
rect 4061 7515 4127 7518
rect 17217 7442 17283 7445
rect 17861 7442 17927 7445
rect 17217 7440 17927 7442
rect 17217 7384 17222 7440
rect 17278 7384 17866 7440
rect 17922 7384 17927 7440
rect 17217 7382 17927 7384
rect 17217 7379 17283 7382
rect 17861 7379 17927 7382
rect 4487 7104 4803 7105
rect 4487 7040 4493 7104
rect 4557 7040 4573 7104
rect 4637 7040 4653 7104
rect 4717 7040 4733 7104
rect 4797 7040 4803 7104
rect 4487 7039 4803 7040
rect 11570 7104 11886 7105
rect 11570 7040 11576 7104
rect 11640 7040 11656 7104
rect 11720 7040 11736 7104
rect 11800 7040 11816 7104
rect 11880 7040 11886 7104
rect 11570 7039 11886 7040
rect 18653 7104 18969 7105
rect 18653 7040 18659 7104
rect 18723 7040 18739 7104
rect 18803 7040 18819 7104
rect 18883 7040 18899 7104
rect 18963 7040 18969 7104
rect 18653 7039 18969 7040
rect 25736 7104 26052 7105
rect 25736 7040 25742 7104
rect 25806 7040 25822 7104
rect 25886 7040 25902 7104
rect 25966 7040 25982 7104
rect 26046 7040 26052 7104
rect 25736 7039 26052 7040
rect 28901 6898 28967 6901
rect 29781 6898 30581 6928
rect 28901 6896 30581 6898
rect 28901 6840 28906 6896
rect 28962 6840 30581 6896
rect 28901 6838 30581 6840
rect 28901 6835 28967 6838
rect 29781 6808 30581 6838
rect 7005 6762 7071 6765
rect 8293 6762 8359 6765
rect 7005 6760 8359 6762
rect 7005 6704 7010 6760
rect 7066 6704 8298 6760
rect 8354 6704 8359 6760
rect 7005 6702 8359 6704
rect 7005 6699 7071 6702
rect 8293 6699 8359 6702
rect 10961 6762 11027 6765
rect 13905 6762 13971 6765
rect 10961 6760 13971 6762
rect 10961 6704 10966 6760
rect 11022 6704 13910 6760
rect 13966 6704 13971 6760
rect 10961 6702 13971 6704
rect 10961 6699 11027 6702
rect 13905 6699 13971 6702
rect 20069 6762 20135 6765
rect 28758 6762 28764 6764
rect 20069 6760 28764 6762
rect 20069 6704 20074 6760
rect 20130 6704 28764 6760
rect 20069 6702 28764 6704
rect 20069 6699 20135 6702
rect 28758 6700 28764 6702
rect 28828 6700 28834 6764
rect 5147 6560 5463 6561
rect 5147 6496 5153 6560
rect 5217 6496 5233 6560
rect 5297 6496 5313 6560
rect 5377 6496 5393 6560
rect 5457 6496 5463 6560
rect 5147 6495 5463 6496
rect 12230 6560 12546 6561
rect 12230 6496 12236 6560
rect 12300 6496 12316 6560
rect 12380 6496 12396 6560
rect 12460 6496 12476 6560
rect 12540 6496 12546 6560
rect 12230 6495 12546 6496
rect 19313 6560 19629 6561
rect 19313 6496 19319 6560
rect 19383 6496 19399 6560
rect 19463 6496 19479 6560
rect 19543 6496 19559 6560
rect 19623 6496 19629 6560
rect 19313 6495 19629 6496
rect 26396 6560 26712 6561
rect 26396 6496 26402 6560
rect 26466 6496 26482 6560
rect 26546 6496 26562 6560
rect 26626 6496 26642 6560
rect 26706 6496 26712 6560
rect 26396 6495 26712 6496
rect 1485 6354 1551 6357
rect 20253 6354 20319 6357
rect 1485 6352 20319 6354
rect 1485 6296 1490 6352
rect 1546 6296 20258 6352
rect 20314 6296 20319 6352
rect 1485 6294 20319 6296
rect 1485 6291 1551 6294
rect 20253 6291 20319 6294
rect 4487 6016 4803 6017
rect 4487 5952 4493 6016
rect 4557 5952 4573 6016
rect 4637 5952 4653 6016
rect 4717 5952 4733 6016
rect 4797 5952 4803 6016
rect 4487 5951 4803 5952
rect 11570 6016 11886 6017
rect 11570 5952 11576 6016
rect 11640 5952 11656 6016
rect 11720 5952 11736 6016
rect 11800 5952 11816 6016
rect 11880 5952 11886 6016
rect 11570 5951 11886 5952
rect 18653 6016 18969 6017
rect 18653 5952 18659 6016
rect 18723 5952 18739 6016
rect 18803 5952 18819 6016
rect 18883 5952 18899 6016
rect 18963 5952 18969 6016
rect 18653 5951 18969 5952
rect 25736 6016 26052 6017
rect 25736 5952 25742 6016
rect 25806 5952 25822 6016
rect 25886 5952 25902 6016
rect 25966 5952 25982 6016
rect 26046 5952 26052 6016
rect 25736 5951 26052 5952
rect 24301 5540 24367 5541
rect 24301 5538 24348 5540
rect 24256 5536 24348 5538
rect 24256 5480 24306 5536
rect 24256 5478 24348 5480
rect 24301 5476 24348 5478
rect 24412 5476 24418 5540
rect 24301 5475 24367 5476
rect 5147 5472 5463 5473
rect 5147 5408 5153 5472
rect 5217 5408 5233 5472
rect 5297 5408 5313 5472
rect 5377 5408 5393 5472
rect 5457 5408 5463 5472
rect 5147 5407 5463 5408
rect 12230 5472 12546 5473
rect 12230 5408 12236 5472
rect 12300 5408 12316 5472
rect 12380 5408 12396 5472
rect 12460 5408 12476 5472
rect 12540 5408 12546 5472
rect 12230 5407 12546 5408
rect 19313 5472 19629 5473
rect 19313 5408 19319 5472
rect 19383 5408 19399 5472
rect 19463 5408 19479 5472
rect 19543 5408 19559 5472
rect 19623 5408 19629 5472
rect 19313 5407 19629 5408
rect 26396 5472 26712 5473
rect 26396 5408 26402 5472
rect 26466 5408 26482 5472
rect 26546 5408 26562 5472
rect 26626 5408 26642 5472
rect 26706 5408 26712 5472
rect 26396 5407 26712 5408
rect 16481 5402 16547 5405
rect 18321 5402 18387 5405
rect 16481 5400 18387 5402
rect 16481 5344 16486 5400
rect 16542 5344 18326 5400
rect 18382 5344 18387 5400
rect 16481 5342 18387 5344
rect 16481 5339 16547 5342
rect 18321 5339 18387 5342
rect 16205 5130 16271 5133
rect 18229 5130 18295 5133
rect 16205 5128 18295 5130
rect 16205 5072 16210 5128
rect 16266 5072 18234 5128
rect 18290 5072 18295 5128
rect 16205 5070 18295 5072
rect 16205 5067 16271 5070
rect 18229 5067 18295 5070
rect 17769 4994 17835 4997
rect 18413 4994 18479 4997
rect 17769 4992 18479 4994
rect 17769 4936 17774 4992
rect 17830 4936 18418 4992
rect 18474 4936 18479 4992
rect 17769 4934 18479 4936
rect 17769 4931 17835 4934
rect 18413 4931 18479 4934
rect 4487 4928 4803 4929
rect 4487 4864 4493 4928
rect 4557 4864 4573 4928
rect 4637 4864 4653 4928
rect 4717 4864 4733 4928
rect 4797 4864 4803 4928
rect 4487 4863 4803 4864
rect 11570 4928 11886 4929
rect 11570 4864 11576 4928
rect 11640 4864 11656 4928
rect 11720 4864 11736 4928
rect 11800 4864 11816 4928
rect 11880 4864 11886 4928
rect 11570 4863 11886 4864
rect 18653 4928 18969 4929
rect 18653 4864 18659 4928
rect 18723 4864 18739 4928
rect 18803 4864 18819 4928
rect 18883 4864 18899 4928
rect 18963 4864 18969 4928
rect 18653 4863 18969 4864
rect 25736 4928 26052 4929
rect 25736 4864 25742 4928
rect 25806 4864 25822 4928
rect 25886 4864 25902 4928
rect 25966 4864 25982 4928
rect 26046 4864 26052 4928
rect 25736 4863 26052 4864
rect 17769 4858 17835 4861
rect 17769 4856 18522 4858
rect 17769 4800 17774 4856
rect 17830 4800 18522 4856
rect 17769 4798 18522 4800
rect 17769 4795 17835 4798
rect 16389 4722 16455 4725
rect 17861 4722 17927 4725
rect 16389 4720 17927 4722
rect 16389 4664 16394 4720
rect 16450 4664 17866 4720
rect 17922 4664 17927 4720
rect 16389 4662 17927 4664
rect 18462 4722 18522 4798
rect 18597 4722 18663 4725
rect 18462 4720 18663 4722
rect 18462 4664 18602 4720
rect 18658 4664 18663 4720
rect 18462 4662 18663 4664
rect 16389 4659 16455 4662
rect 17861 4659 17927 4662
rect 18597 4659 18663 4662
rect 5147 4384 5463 4385
rect 5147 4320 5153 4384
rect 5217 4320 5233 4384
rect 5297 4320 5313 4384
rect 5377 4320 5393 4384
rect 5457 4320 5463 4384
rect 5147 4319 5463 4320
rect 12230 4384 12546 4385
rect 12230 4320 12236 4384
rect 12300 4320 12316 4384
rect 12380 4320 12396 4384
rect 12460 4320 12476 4384
rect 12540 4320 12546 4384
rect 12230 4319 12546 4320
rect 19313 4384 19629 4385
rect 19313 4320 19319 4384
rect 19383 4320 19399 4384
rect 19463 4320 19479 4384
rect 19543 4320 19559 4384
rect 19623 4320 19629 4384
rect 19313 4319 19629 4320
rect 26396 4384 26712 4385
rect 26396 4320 26402 4384
rect 26466 4320 26482 4384
rect 26546 4320 26562 4384
rect 26626 4320 26642 4384
rect 26706 4320 26712 4384
rect 26396 4319 26712 4320
rect 14641 4178 14707 4181
rect 17493 4178 17559 4181
rect 14641 4176 17559 4178
rect 14641 4120 14646 4176
rect 14702 4120 17498 4176
rect 17554 4120 17559 4176
rect 14641 4118 17559 4120
rect 14641 4115 14707 4118
rect 17493 4115 17559 4118
rect 2405 4042 2471 4045
rect 23933 4042 23999 4045
rect 2405 4040 23999 4042
rect 2405 3984 2410 4040
rect 2466 3984 23938 4040
rect 23994 3984 23999 4040
rect 2405 3982 23999 3984
rect 2405 3979 2471 3982
rect 23933 3979 23999 3982
rect 4487 3840 4803 3841
rect 4487 3776 4493 3840
rect 4557 3776 4573 3840
rect 4637 3776 4653 3840
rect 4717 3776 4733 3840
rect 4797 3776 4803 3840
rect 4487 3775 4803 3776
rect 11570 3840 11886 3841
rect 11570 3776 11576 3840
rect 11640 3776 11656 3840
rect 11720 3776 11736 3840
rect 11800 3776 11816 3840
rect 11880 3776 11886 3840
rect 11570 3775 11886 3776
rect 18653 3840 18969 3841
rect 18653 3776 18659 3840
rect 18723 3776 18739 3840
rect 18803 3776 18819 3840
rect 18883 3776 18899 3840
rect 18963 3776 18969 3840
rect 18653 3775 18969 3776
rect 25736 3840 26052 3841
rect 25736 3776 25742 3840
rect 25806 3776 25822 3840
rect 25886 3776 25902 3840
rect 25966 3776 25982 3840
rect 26046 3776 26052 3840
rect 25736 3775 26052 3776
rect 12893 3634 12959 3637
rect 18873 3634 18939 3637
rect 12893 3632 18939 3634
rect 12893 3576 12898 3632
rect 12954 3576 18878 3632
rect 18934 3576 18939 3632
rect 12893 3574 18939 3576
rect 12893 3571 12959 3574
rect 18873 3571 18939 3574
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 5147 3296 5463 3297
rect 5147 3232 5153 3296
rect 5217 3232 5233 3296
rect 5297 3232 5313 3296
rect 5377 3232 5393 3296
rect 5457 3232 5463 3296
rect 5147 3231 5463 3232
rect 12230 3296 12546 3297
rect 12230 3232 12236 3296
rect 12300 3232 12316 3296
rect 12380 3232 12396 3296
rect 12460 3232 12476 3296
rect 12540 3232 12546 3296
rect 12230 3231 12546 3232
rect 19313 3296 19629 3297
rect 19313 3232 19319 3296
rect 19383 3232 19399 3296
rect 19463 3232 19479 3296
rect 19543 3232 19559 3296
rect 19623 3232 19629 3296
rect 19313 3231 19629 3232
rect 26396 3296 26712 3297
rect 26396 3232 26402 3296
rect 26466 3232 26482 3296
rect 26546 3232 26562 3296
rect 26626 3232 26642 3296
rect 26706 3232 26712 3296
rect 26396 3231 26712 3232
rect 28993 2818 29059 2821
rect 29781 2818 30581 2848
rect 28993 2816 30581 2818
rect 28993 2760 28998 2816
rect 29054 2760 30581 2816
rect 28993 2758 30581 2760
rect 28993 2755 29059 2758
rect 4487 2752 4803 2753
rect 4487 2688 4493 2752
rect 4557 2688 4573 2752
rect 4637 2688 4653 2752
rect 4717 2688 4733 2752
rect 4797 2688 4803 2752
rect 4487 2687 4803 2688
rect 11570 2752 11886 2753
rect 11570 2688 11576 2752
rect 11640 2688 11656 2752
rect 11720 2688 11736 2752
rect 11800 2688 11816 2752
rect 11880 2688 11886 2752
rect 11570 2687 11886 2688
rect 18653 2752 18969 2753
rect 18653 2688 18659 2752
rect 18723 2688 18739 2752
rect 18803 2688 18819 2752
rect 18883 2688 18899 2752
rect 18963 2688 18969 2752
rect 18653 2687 18969 2688
rect 25736 2752 26052 2753
rect 25736 2688 25742 2752
rect 25806 2688 25822 2752
rect 25886 2688 25902 2752
rect 25966 2688 25982 2752
rect 26046 2688 26052 2752
rect 29781 2728 30581 2758
rect 25736 2687 26052 2688
rect 5147 2208 5463 2209
rect 5147 2144 5153 2208
rect 5217 2144 5233 2208
rect 5297 2144 5313 2208
rect 5377 2144 5393 2208
rect 5457 2144 5463 2208
rect 5147 2143 5463 2144
rect 12230 2208 12546 2209
rect 12230 2144 12236 2208
rect 12300 2144 12316 2208
rect 12380 2144 12396 2208
rect 12460 2144 12476 2208
rect 12540 2144 12546 2208
rect 12230 2143 12546 2144
rect 19313 2208 19629 2209
rect 19313 2144 19319 2208
rect 19383 2144 19399 2208
rect 19463 2144 19479 2208
rect 19543 2144 19559 2208
rect 19623 2144 19629 2208
rect 19313 2143 19629 2144
rect 26396 2208 26712 2209
rect 26396 2144 26402 2208
rect 26466 2144 26482 2208
rect 26546 2144 26562 2208
rect 26626 2144 26642 2208
rect 26706 2144 26712 2208
rect 26396 2143 26712 2144
<< via3 >>
rect 5153 30492 5217 30496
rect 5153 30436 5157 30492
rect 5157 30436 5213 30492
rect 5213 30436 5217 30492
rect 5153 30432 5217 30436
rect 5233 30492 5297 30496
rect 5233 30436 5237 30492
rect 5237 30436 5293 30492
rect 5293 30436 5297 30492
rect 5233 30432 5297 30436
rect 5313 30492 5377 30496
rect 5313 30436 5317 30492
rect 5317 30436 5373 30492
rect 5373 30436 5377 30492
rect 5313 30432 5377 30436
rect 5393 30492 5457 30496
rect 5393 30436 5397 30492
rect 5397 30436 5453 30492
rect 5453 30436 5457 30492
rect 5393 30432 5457 30436
rect 12236 30492 12300 30496
rect 12236 30436 12240 30492
rect 12240 30436 12296 30492
rect 12296 30436 12300 30492
rect 12236 30432 12300 30436
rect 12316 30492 12380 30496
rect 12316 30436 12320 30492
rect 12320 30436 12376 30492
rect 12376 30436 12380 30492
rect 12316 30432 12380 30436
rect 12396 30492 12460 30496
rect 12396 30436 12400 30492
rect 12400 30436 12456 30492
rect 12456 30436 12460 30492
rect 12396 30432 12460 30436
rect 12476 30492 12540 30496
rect 12476 30436 12480 30492
rect 12480 30436 12536 30492
rect 12536 30436 12540 30492
rect 12476 30432 12540 30436
rect 19319 30492 19383 30496
rect 19319 30436 19323 30492
rect 19323 30436 19379 30492
rect 19379 30436 19383 30492
rect 19319 30432 19383 30436
rect 19399 30492 19463 30496
rect 19399 30436 19403 30492
rect 19403 30436 19459 30492
rect 19459 30436 19463 30492
rect 19399 30432 19463 30436
rect 19479 30492 19543 30496
rect 19479 30436 19483 30492
rect 19483 30436 19539 30492
rect 19539 30436 19543 30492
rect 19479 30432 19543 30436
rect 19559 30492 19623 30496
rect 19559 30436 19563 30492
rect 19563 30436 19619 30492
rect 19619 30436 19623 30492
rect 19559 30432 19623 30436
rect 26402 30492 26466 30496
rect 26402 30436 26406 30492
rect 26406 30436 26462 30492
rect 26462 30436 26466 30492
rect 26402 30432 26466 30436
rect 26482 30492 26546 30496
rect 26482 30436 26486 30492
rect 26486 30436 26542 30492
rect 26542 30436 26546 30492
rect 26482 30432 26546 30436
rect 26562 30492 26626 30496
rect 26562 30436 26566 30492
rect 26566 30436 26622 30492
rect 26622 30436 26626 30492
rect 26562 30432 26626 30436
rect 26642 30492 26706 30496
rect 26642 30436 26646 30492
rect 26646 30436 26702 30492
rect 26702 30436 26706 30492
rect 26642 30432 26706 30436
rect 4493 29948 4557 29952
rect 4493 29892 4497 29948
rect 4497 29892 4553 29948
rect 4553 29892 4557 29948
rect 4493 29888 4557 29892
rect 4573 29948 4637 29952
rect 4573 29892 4577 29948
rect 4577 29892 4633 29948
rect 4633 29892 4637 29948
rect 4573 29888 4637 29892
rect 4653 29948 4717 29952
rect 4653 29892 4657 29948
rect 4657 29892 4713 29948
rect 4713 29892 4717 29948
rect 4653 29888 4717 29892
rect 4733 29948 4797 29952
rect 4733 29892 4737 29948
rect 4737 29892 4793 29948
rect 4793 29892 4797 29948
rect 4733 29888 4797 29892
rect 11576 29948 11640 29952
rect 11576 29892 11580 29948
rect 11580 29892 11636 29948
rect 11636 29892 11640 29948
rect 11576 29888 11640 29892
rect 11656 29948 11720 29952
rect 11656 29892 11660 29948
rect 11660 29892 11716 29948
rect 11716 29892 11720 29948
rect 11656 29888 11720 29892
rect 11736 29948 11800 29952
rect 11736 29892 11740 29948
rect 11740 29892 11796 29948
rect 11796 29892 11800 29948
rect 11736 29888 11800 29892
rect 11816 29948 11880 29952
rect 11816 29892 11820 29948
rect 11820 29892 11876 29948
rect 11876 29892 11880 29948
rect 11816 29888 11880 29892
rect 18659 29948 18723 29952
rect 18659 29892 18663 29948
rect 18663 29892 18719 29948
rect 18719 29892 18723 29948
rect 18659 29888 18723 29892
rect 18739 29948 18803 29952
rect 18739 29892 18743 29948
rect 18743 29892 18799 29948
rect 18799 29892 18803 29948
rect 18739 29888 18803 29892
rect 18819 29948 18883 29952
rect 18819 29892 18823 29948
rect 18823 29892 18879 29948
rect 18879 29892 18883 29948
rect 18819 29888 18883 29892
rect 18899 29948 18963 29952
rect 18899 29892 18903 29948
rect 18903 29892 18959 29948
rect 18959 29892 18963 29948
rect 18899 29888 18963 29892
rect 25742 29948 25806 29952
rect 25742 29892 25746 29948
rect 25746 29892 25802 29948
rect 25802 29892 25806 29948
rect 25742 29888 25806 29892
rect 25822 29948 25886 29952
rect 25822 29892 25826 29948
rect 25826 29892 25882 29948
rect 25882 29892 25886 29948
rect 25822 29888 25886 29892
rect 25902 29948 25966 29952
rect 25902 29892 25906 29948
rect 25906 29892 25962 29948
rect 25962 29892 25966 29948
rect 25902 29888 25966 29892
rect 25982 29948 26046 29952
rect 25982 29892 25986 29948
rect 25986 29892 26042 29948
rect 26042 29892 26046 29948
rect 25982 29888 26046 29892
rect 5153 29404 5217 29408
rect 5153 29348 5157 29404
rect 5157 29348 5213 29404
rect 5213 29348 5217 29404
rect 5153 29344 5217 29348
rect 5233 29404 5297 29408
rect 5233 29348 5237 29404
rect 5237 29348 5293 29404
rect 5293 29348 5297 29404
rect 5233 29344 5297 29348
rect 5313 29404 5377 29408
rect 5313 29348 5317 29404
rect 5317 29348 5373 29404
rect 5373 29348 5377 29404
rect 5313 29344 5377 29348
rect 5393 29404 5457 29408
rect 5393 29348 5397 29404
rect 5397 29348 5453 29404
rect 5453 29348 5457 29404
rect 5393 29344 5457 29348
rect 12236 29404 12300 29408
rect 12236 29348 12240 29404
rect 12240 29348 12296 29404
rect 12296 29348 12300 29404
rect 12236 29344 12300 29348
rect 12316 29404 12380 29408
rect 12316 29348 12320 29404
rect 12320 29348 12376 29404
rect 12376 29348 12380 29404
rect 12316 29344 12380 29348
rect 12396 29404 12460 29408
rect 12396 29348 12400 29404
rect 12400 29348 12456 29404
rect 12456 29348 12460 29404
rect 12396 29344 12460 29348
rect 12476 29404 12540 29408
rect 12476 29348 12480 29404
rect 12480 29348 12536 29404
rect 12536 29348 12540 29404
rect 12476 29344 12540 29348
rect 19319 29404 19383 29408
rect 19319 29348 19323 29404
rect 19323 29348 19379 29404
rect 19379 29348 19383 29404
rect 19319 29344 19383 29348
rect 19399 29404 19463 29408
rect 19399 29348 19403 29404
rect 19403 29348 19459 29404
rect 19459 29348 19463 29404
rect 19399 29344 19463 29348
rect 19479 29404 19543 29408
rect 19479 29348 19483 29404
rect 19483 29348 19539 29404
rect 19539 29348 19543 29404
rect 19479 29344 19543 29348
rect 19559 29404 19623 29408
rect 19559 29348 19563 29404
rect 19563 29348 19619 29404
rect 19619 29348 19623 29404
rect 19559 29344 19623 29348
rect 26402 29404 26466 29408
rect 26402 29348 26406 29404
rect 26406 29348 26462 29404
rect 26462 29348 26466 29404
rect 26402 29344 26466 29348
rect 26482 29404 26546 29408
rect 26482 29348 26486 29404
rect 26486 29348 26542 29404
rect 26542 29348 26546 29404
rect 26482 29344 26546 29348
rect 26562 29404 26626 29408
rect 26562 29348 26566 29404
rect 26566 29348 26622 29404
rect 26622 29348 26626 29404
rect 26562 29344 26626 29348
rect 26642 29404 26706 29408
rect 26642 29348 26646 29404
rect 26646 29348 26702 29404
rect 26702 29348 26706 29404
rect 26642 29344 26706 29348
rect 28764 29064 28828 29068
rect 28764 29008 28778 29064
rect 28778 29008 28828 29064
rect 28764 29004 28828 29008
rect 4493 28860 4557 28864
rect 4493 28804 4497 28860
rect 4497 28804 4553 28860
rect 4553 28804 4557 28860
rect 4493 28800 4557 28804
rect 4573 28860 4637 28864
rect 4573 28804 4577 28860
rect 4577 28804 4633 28860
rect 4633 28804 4637 28860
rect 4573 28800 4637 28804
rect 4653 28860 4717 28864
rect 4653 28804 4657 28860
rect 4657 28804 4713 28860
rect 4713 28804 4717 28860
rect 4653 28800 4717 28804
rect 4733 28860 4797 28864
rect 4733 28804 4737 28860
rect 4737 28804 4793 28860
rect 4793 28804 4797 28860
rect 4733 28800 4797 28804
rect 11576 28860 11640 28864
rect 11576 28804 11580 28860
rect 11580 28804 11636 28860
rect 11636 28804 11640 28860
rect 11576 28800 11640 28804
rect 11656 28860 11720 28864
rect 11656 28804 11660 28860
rect 11660 28804 11716 28860
rect 11716 28804 11720 28860
rect 11656 28800 11720 28804
rect 11736 28860 11800 28864
rect 11736 28804 11740 28860
rect 11740 28804 11796 28860
rect 11796 28804 11800 28860
rect 11736 28800 11800 28804
rect 11816 28860 11880 28864
rect 11816 28804 11820 28860
rect 11820 28804 11876 28860
rect 11876 28804 11880 28860
rect 11816 28800 11880 28804
rect 18659 28860 18723 28864
rect 18659 28804 18663 28860
rect 18663 28804 18719 28860
rect 18719 28804 18723 28860
rect 18659 28800 18723 28804
rect 18739 28860 18803 28864
rect 18739 28804 18743 28860
rect 18743 28804 18799 28860
rect 18799 28804 18803 28860
rect 18739 28800 18803 28804
rect 18819 28860 18883 28864
rect 18819 28804 18823 28860
rect 18823 28804 18879 28860
rect 18879 28804 18883 28860
rect 18819 28800 18883 28804
rect 18899 28860 18963 28864
rect 18899 28804 18903 28860
rect 18903 28804 18959 28860
rect 18959 28804 18963 28860
rect 18899 28800 18963 28804
rect 25742 28860 25806 28864
rect 25742 28804 25746 28860
rect 25746 28804 25802 28860
rect 25802 28804 25806 28860
rect 25742 28800 25806 28804
rect 25822 28860 25886 28864
rect 25822 28804 25826 28860
rect 25826 28804 25882 28860
rect 25882 28804 25886 28860
rect 25822 28800 25886 28804
rect 25902 28860 25966 28864
rect 25902 28804 25906 28860
rect 25906 28804 25962 28860
rect 25962 28804 25966 28860
rect 25902 28800 25966 28804
rect 25982 28860 26046 28864
rect 25982 28804 25986 28860
rect 25986 28804 26042 28860
rect 26042 28804 26046 28860
rect 25982 28800 26046 28804
rect 5153 28316 5217 28320
rect 5153 28260 5157 28316
rect 5157 28260 5213 28316
rect 5213 28260 5217 28316
rect 5153 28256 5217 28260
rect 5233 28316 5297 28320
rect 5233 28260 5237 28316
rect 5237 28260 5293 28316
rect 5293 28260 5297 28316
rect 5233 28256 5297 28260
rect 5313 28316 5377 28320
rect 5313 28260 5317 28316
rect 5317 28260 5373 28316
rect 5373 28260 5377 28316
rect 5313 28256 5377 28260
rect 5393 28316 5457 28320
rect 5393 28260 5397 28316
rect 5397 28260 5453 28316
rect 5453 28260 5457 28316
rect 5393 28256 5457 28260
rect 12236 28316 12300 28320
rect 12236 28260 12240 28316
rect 12240 28260 12296 28316
rect 12296 28260 12300 28316
rect 12236 28256 12300 28260
rect 12316 28316 12380 28320
rect 12316 28260 12320 28316
rect 12320 28260 12376 28316
rect 12376 28260 12380 28316
rect 12316 28256 12380 28260
rect 12396 28316 12460 28320
rect 12396 28260 12400 28316
rect 12400 28260 12456 28316
rect 12456 28260 12460 28316
rect 12396 28256 12460 28260
rect 12476 28316 12540 28320
rect 12476 28260 12480 28316
rect 12480 28260 12536 28316
rect 12536 28260 12540 28316
rect 12476 28256 12540 28260
rect 19319 28316 19383 28320
rect 19319 28260 19323 28316
rect 19323 28260 19379 28316
rect 19379 28260 19383 28316
rect 19319 28256 19383 28260
rect 19399 28316 19463 28320
rect 19399 28260 19403 28316
rect 19403 28260 19459 28316
rect 19459 28260 19463 28316
rect 19399 28256 19463 28260
rect 19479 28316 19543 28320
rect 19479 28260 19483 28316
rect 19483 28260 19539 28316
rect 19539 28260 19543 28316
rect 19479 28256 19543 28260
rect 19559 28316 19623 28320
rect 19559 28260 19563 28316
rect 19563 28260 19619 28316
rect 19619 28260 19623 28316
rect 19559 28256 19623 28260
rect 26402 28316 26466 28320
rect 26402 28260 26406 28316
rect 26406 28260 26462 28316
rect 26462 28260 26466 28316
rect 26402 28256 26466 28260
rect 26482 28316 26546 28320
rect 26482 28260 26486 28316
rect 26486 28260 26542 28316
rect 26542 28260 26546 28316
rect 26482 28256 26546 28260
rect 26562 28316 26626 28320
rect 26562 28260 26566 28316
rect 26566 28260 26622 28316
rect 26622 28260 26626 28316
rect 26562 28256 26626 28260
rect 26642 28316 26706 28320
rect 26642 28260 26646 28316
rect 26646 28260 26702 28316
rect 26702 28260 26706 28316
rect 26642 28256 26706 28260
rect 4493 27772 4557 27776
rect 4493 27716 4497 27772
rect 4497 27716 4553 27772
rect 4553 27716 4557 27772
rect 4493 27712 4557 27716
rect 4573 27772 4637 27776
rect 4573 27716 4577 27772
rect 4577 27716 4633 27772
rect 4633 27716 4637 27772
rect 4573 27712 4637 27716
rect 4653 27772 4717 27776
rect 4653 27716 4657 27772
rect 4657 27716 4713 27772
rect 4713 27716 4717 27772
rect 4653 27712 4717 27716
rect 4733 27772 4797 27776
rect 4733 27716 4737 27772
rect 4737 27716 4793 27772
rect 4793 27716 4797 27772
rect 4733 27712 4797 27716
rect 11576 27772 11640 27776
rect 11576 27716 11580 27772
rect 11580 27716 11636 27772
rect 11636 27716 11640 27772
rect 11576 27712 11640 27716
rect 11656 27772 11720 27776
rect 11656 27716 11660 27772
rect 11660 27716 11716 27772
rect 11716 27716 11720 27772
rect 11656 27712 11720 27716
rect 11736 27772 11800 27776
rect 11736 27716 11740 27772
rect 11740 27716 11796 27772
rect 11796 27716 11800 27772
rect 11736 27712 11800 27716
rect 11816 27772 11880 27776
rect 11816 27716 11820 27772
rect 11820 27716 11876 27772
rect 11876 27716 11880 27772
rect 11816 27712 11880 27716
rect 18659 27772 18723 27776
rect 18659 27716 18663 27772
rect 18663 27716 18719 27772
rect 18719 27716 18723 27772
rect 18659 27712 18723 27716
rect 18739 27772 18803 27776
rect 18739 27716 18743 27772
rect 18743 27716 18799 27772
rect 18799 27716 18803 27772
rect 18739 27712 18803 27716
rect 18819 27772 18883 27776
rect 18819 27716 18823 27772
rect 18823 27716 18879 27772
rect 18879 27716 18883 27772
rect 18819 27712 18883 27716
rect 18899 27772 18963 27776
rect 18899 27716 18903 27772
rect 18903 27716 18959 27772
rect 18959 27716 18963 27772
rect 18899 27712 18963 27716
rect 25742 27772 25806 27776
rect 25742 27716 25746 27772
rect 25746 27716 25802 27772
rect 25802 27716 25806 27772
rect 25742 27712 25806 27716
rect 25822 27772 25886 27776
rect 25822 27716 25826 27772
rect 25826 27716 25882 27772
rect 25882 27716 25886 27772
rect 25822 27712 25886 27716
rect 25902 27772 25966 27776
rect 25902 27716 25906 27772
rect 25906 27716 25962 27772
rect 25962 27716 25966 27772
rect 25902 27712 25966 27716
rect 25982 27772 26046 27776
rect 25982 27716 25986 27772
rect 25986 27716 26042 27772
rect 26042 27716 26046 27772
rect 25982 27712 26046 27716
rect 5153 27228 5217 27232
rect 5153 27172 5157 27228
rect 5157 27172 5213 27228
rect 5213 27172 5217 27228
rect 5153 27168 5217 27172
rect 5233 27228 5297 27232
rect 5233 27172 5237 27228
rect 5237 27172 5293 27228
rect 5293 27172 5297 27228
rect 5233 27168 5297 27172
rect 5313 27228 5377 27232
rect 5313 27172 5317 27228
rect 5317 27172 5373 27228
rect 5373 27172 5377 27228
rect 5313 27168 5377 27172
rect 5393 27228 5457 27232
rect 5393 27172 5397 27228
rect 5397 27172 5453 27228
rect 5453 27172 5457 27228
rect 5393 27168 5457 27172
rect 12236 27228 12300 27232
rect 12236 27172 12240 27228
rect 12240 27172 12296 27228
rect 12296 27172 12300 27228
rect 12236 27168 12300 27172
rect 12316 27228 12380 27232
rect 12316 27172 12320 27228
rect 12320 27172 12376 27228
rect 12376 27172 12380 27228
rect 12316 27168 12380 27172
rect 12396 27228 12460 27232
rect 12396 27172 12400 27228
rect 12400 27172 12456 27228
rect 12456 27172 12460 27228
rect 12396 27168 12460 27172
rect 12476 27228 12540 27232
rect 12476 27172 12480 27228
rect 12480 27172 12536 27228
rect 12536 27172 12540 27228
rect 12476 27168 12540 27172
rect 19319 27228 19383 27232
rect 19319 27172 19323 27228
rect 19323 27172 19379 27228
rect 19379 27172 19383 27228
rect 19319 27168 19383 27172
rect 19399 27228 19463 27232
rect 19399 27172 19403 27228
rect 19403 27172 19459 27228
rect 19459 27172 19463 27228
rect 19399 27168 19463 27172
rect 19479 27228 19543 27232
rect 19479 27172 19483 27228
rect 19483 27172 19539 27228
rect 19539 27172 19543 27228
rect 19479 27168 19543 27172
rect 19559 27228 19623 27232
rect 19559 27172 19563 27228
rect 19563 27172 19619 27228
rect 19619 27172 19623 27228
rect 19559 27168 19623 27172
rect 26402 27228 26466 27232
rect 26402 27172 26406 27228
rect 26406 27172 26462 27228
rect 26462 27172 26466 27228
rect 26402 27168 26466 27172
rect 26482 27228 26546 27232
rect 26482 27172 26486 27228
rect 26486 27172 26542 27228
rect 26542 27172 26546 27228
rect 26482 27168 26546 27172
rect 26562 27228 26626 27232
rect 26562 27172 26566 27228
rect 26566 27172 26622 27228
rect 26622 27172 26626 27228
rect 26562 27168 26626 27172
rect 26642 27228 26706 27232
rect 26642 27172 26646 27228
rect 26646 27172 26702 27228
rect 26702 27172 26706 27228
rect 26642 27168 26706 27172
rect 4493 26684 4557 26688
rect 4493 26628 4497 26684
rect 4497 26628 4553 26684
rect 4553 26628 4557 26684
rect 4493 26624 4557 26628
rect 4573 26684 4637 26688
rect 4573 26628 4577 26684
rect 4577 26628 4633 26684
rect 4633 26628 4637 26684
rect 4573 26624 4637 26628
rect 4653 26684 4717 26688
rect 4653 26628 4657 26684
rect 4657 26628 4713 26684
rect 4713 26628 4717 26684
rect 4653 26624 4717 26628
rect 4733 26684 4797 26688
rect 4733 26628 4737 26684
rect 4737 26628 4793 26684
rect 4793 26628 4797 26684
rect 4733 26624 4797 26628
rect 11576 26684 11640 26688
rect 11576 26628 11580 26684
rect 11580 26628 11636 26684
rect 11636 26628 11640 26684
rect 11576 26624 11640 26628
rect 11656 26684 11720 26688
rect 11656 26628 11660 26684
rect 11660 26628 11716 26684
rect 11716 26628 11720 26684
rect 11656 26624 11720 26628
rect 11736 26684 11800 26688
rect 11736 26628 11740 26684
rect 11740 26628 11796 26684
rect 11796 26628 11800 26684
rect 11736 26624 11800 26628
rect 11816 26684 11880 26688
rect 11816 26628 11820 26684
rect 11820 26628 11876 26684
rect 11876 26628 11880 26684
rect 11816 26624 11880 26628
rect 18659 26684 18723 26688
rect 18659 26628 18663 26684
rect 18663 26628 18719 26684
rect 18719 26628 18723 26684
rect 18659 26624 18723 26628
rect 18739 26684 18803 26688
rect 18739 26628 18743 26684
rect 18743 26628 18799 26684
rect 18799 26628 18803 26684
rect 18739 26624 18803 26628
rect 18819 26684 18883 26688
rect 18819 26628 18823 26684
rect 18823 26628 18879 26684
rect 18879 26628 18883 26684
rect 18819 26624 18883 26628
rect 18899 26684 18963 26688
rect 18899 26628 18903 26684
rect 18903 26628 18959 26684
rect 18959 26628 18963 26684
rect 18899 26624 18963 26628
rect 25742 26684 25806 26688
rect 25742 26628 25746 26684
rect 25746 26628 25802 26684
rect 25802 26628 25806 26684
rect 25742 26624 25806 26628
rect 25822 26684 25886 26688
rect 25822 26628 25826 26684
rect 25826 26628 25882 26684
rect 25882 26628 25886 26684
rect 25822 26624 25886 26628
rect 25902 26684 25966 26688
rect 25902 26628 25906 26684
rect 25906 26628 25962 26684
rect 25962 26628 25966 26684
rect 25902 26624 25966 26628
rect 25982 26684 26046 26688
rect 25982 26628 25986 26684
rect 25986 26628 26042 26684
rect 26042 26628 26046 26684
rect 25982 26624 26046 26628
rect 5153 26140 5217 26144
rect 5153 26084 5157 26140
rect 5157 26084 5213 26140
rect 5213 26084 5217 26140
rect 5153 26080 5217 26084
rect 5233 26140 5297 26144
rect 5233 26084 5237 26140
rect 5237 26084 5293 26140
rect 5293 26084 5297 26140
rect 5233 26080 5297 26084
rect 5313 26140 5377 26144
rect 5313 26084 5317 26140
rect 5317 26084 5373 26140
rect 5373 26084 5377 26140
rect 5313 26080 5377 26084
rect 5393 26140 5457 26144
rect 5393 26084 5397 26140
rect 5397 26084 5453 26140
rect 5453 26084 5457 26140
rect 5393 26080 5457 26084
rect 12236 26140 12300 26144
rect 12236 26084 12240 26140
rect 12240 26084 12296 26140
rect 12296 26084 12300 26140
rect 12236 26080 12300 26084
rect 12316 26140 12380 26144
rect 12316 26084 12320 26140
rect 12320 26084 12376 26140
rect 12376 26084 12380 26140
rect 12316 26080 12380 26084
rect 12396 26140 12460 26144
rect 12396 26084 12400 26140
rect 12400 26084 12456 26140
rect 12456 26084 12460 26140
rect 12396 26080 12460 26084
rect 12476 26140 12540 26144
rect 12476 26084 12480 26140
rect 12480 26084 12536 26140
rect 12536 26084 12540 26140
rect 12476 26080 12540 26084
rect 19319 26140 19383 26144
rect 19319 26084 19323 26140
rect 19323 26084 19379 26140
rect 19379 26084 19383 26140
rect 19319 26080 19383 26084
rect 19399 26140 19463 26144
rect 19399 26084 19403 26140
rect 19403 26084 19459 26140
rect 19459 26084 19463 26140
rect 19399 26080 19463 26084
rect 19479 26140 19543 26144
rect 19479 26084 19483 26140
rect 19483 26084 19539 26140
rect 19539 26084 19543 26140
rect 19479 26080 19543 26084
rect 19559 26140 19623 26144
rect 19559 26084 19563 26140
rect 19563 26084 19619 26140
rect 19619 26084 19623 26140
rect 19559 26080 19623 26084
rect 26402 26140 26466 26144
rect 26402 26084 26406 26140
rect 26406 26084 26462 26140
rect 26462 26084 26466 26140
rect 26402 26080 26466 26084
rect 26482 26140 26546 26144
rect 26482 26084 26486 26140
rect 26486 26084 26542 26140
rect 26542 26084 26546 26140
rect 26482 26080 26546 26084
rect 26562 26140 26626 26144
rect 26562 26084 26566 26140
rect 26566 26084 26622 26140
rect 26622 26084 26626 26140
rect 26562 26080 26626 26084
rect 26642 26140 26706 26144
rect 26642 26084 26646 26140
rect 26646 26084 26702 26140
rect 26702 26084 26706 26140
rect 26642 26080 26706 26084
rect 4493 25596 4557 25600
rect 4493 25540 4497 25596
rect 4497 25540 4553 25596
rect 4553 25540 4557 25596
rect 4493 25536 4557 25540
rect 4573 25596 4637 25600
rect 4573 25540 4577 25596
rect 4577 25540 4633 25596
rect 4633 25540 4637 25596
rect 4573 25536 4637 25540
rect 4653 25596 4717 25600
rect 4653 25540 4657 25596
rect 4657 25540 4713 25596
rect 4713 25540 4717 25596
rect 4653 25536 4717 25540
rect 4733 25596 4797 25600
rect 4733 25540 4737 25596
rect 4737 25540 4793 25596
rect 4793 25540 4797 25596
rect 4733 25536 4797 25540
rect 11576 25596 11640 25600
rect 11576 25540 11580 25596
rect 11580 25540 11636 25596
rect 11636 25540 11640 25596
rect 11576 25536 11640 25540
rect 11656 25596 11720 25600
rect 11656 25540 11660 25596
rect 11660 25540 11716 25596
rect 11716 25540 11720 25596
rect 11656 25536 11720 25540
rect 11736 25596 11800 25600
rect 11736 25540 11740 25596
rect 11740 25540 11796 25596
rect 11796 25540 11800 25596
rect 11736 25536 11800 25540
rect 11816 25596 11880 25600
rect 11816 25540 11820 25596
rect 11820 25540 11876 25596
rect 11876 25540 11880 25596
rect 11816 25536 11880 25540
rect 18659 25596 18723 25600
rect 18659 25540 18663 25596
rect 18663 25540 18719 25596
rect 18719 25540 18723 25596
rect 18659 25536 18723 25540
rect 18739 25596 18803 25600
rect 18739 25540 18743 25596
rect 18743 25540 18799 25596
rect 18799 25540 18803 25596
rect 18739 25536 18803 25540
rect 18819 25596 18883 25600
rect 18819 25540 18823 25596
rect 18823 25540 18879 25596
rect 18879 25540 18883 25596
rect 18819 25536 18883 25540
rect 18899 25596 18963 25600
rect 18899 25540 18903 25596
rect 18903 25540 18959 25596
rect 18959 25540 18963 25596
rect 18899 25536 18963 25540
rect 25742 25596 25806 25600
rect 25742 25540 25746 25596
rect 25746 25540 25802 25596
rect 25802 25540 25806 25596
rect 25742 25536 25806 25540
rect 25822 25596 25886 25600
rect 25822 25540 25826 25596
rect 25826 25540 25882 25596
rect 25882 25540 25886 25596
rect 25822 25536 25886 25540
rect 25902 25596 25966 25600
rect 25902 25540 25906 25596
rect 25906 25540 25962 25596
rect 25962 25540 25966 25596
rect 25902 25536 25966 25540
rect 25982 25596 26046 25600
rect 25982 25540 25986 25596
rect 25986 25540 26042 25596
rect 26042 25540 26046 25596
rect 25982 25536 26046 25540
rect 5153 25052 5217 25056
rect 5153 24996 5157 25052
rect 5157 24996 5213 25052
rect 5213 24996 5217 25052
rect 5153 24992 5217 24996
rect 5233 25052 5297 25056
rect 5233 24996 5237 25052
rect 5237 24996 5293 25052
rect 5293 24996 5297 25052
rect 5233 24992 5297 24996
rect 5313 25052 5377 25056
rect 5313 24996 5317 25052
rect 5317 24996 5373 25052
rect 5373 24996 5377 25052
rect 5313 24992 5377 24996
rect 5393 25052 5457 25056
rect 5393 24996 5397 25052
rect 5397 24996 5453 25052
rect 5453 24996 5457 25052
rect 5393 24992 5457 24996
rect 12236 25052 12300 25056
rect 12236 24996 12240 25052
rect 12240 24996 12296 25052
rect 12296 24996 12300 25052
rect 12236 24992 12300 24996
rect 12316 25052 12380 25056
rect 12316 24996 12320 25052
rect 12320 24996 12376 25052
rect 12376 24996 12380 25052
rect 12316 24992 12380 24996
rect 12396 25052 12460 25056
rect 12396 24996 12400 25052
rect 12400 24996 12456 25052
rect 12456 24996 12460 25052
rect 12396 24992 12460 24996
rect 12476 25052 12540 25056
rect 12476 24996 12480 25052
rect 12480 24996 12536 25052
rect 12536 24996 12540 25052
rect 12476 24992 12540 24996
rect 19319 25052 19383 25056
rect 19319 24996 19323 25052
rect 19323 24996 19379 25052
rect 19379 24996 19383 25052
rect 19319 24992 19383 24996
rect 19399 25052 19463 25056
rect 19399 24996 19403 25052
rect 19403 24996 19459 25052
rect 19459 24996 19463 25052
rect 19399 24992 19463 24996
rect 19479 25052 19543 25056
rect 19479 24996 19483 25052
rect 19483 24996 19539 25052
rect 19539 24996 19543 25052
rect 19479 24992 19543 24996
rect 19559 25052 19623 25056
rect 19559 24996 19563 25052
rect 19563 24996 19619 25052
rect 19619 24996 19623 25052
rect 19559 24992 19623 24996
rect 26402 25052 26466 25056
rect 26402 24996 26406 25052
rect 26406 24996 26462 25052
rect 26462 24996 26466 25052
rect 26402 24992 26466 24996
rect 26482 25052 26546 25056
rect 26482 24996 26486 25052
rect 26486 24996 26542 25052
rect 26542 24996 26546 25052
rect 26482 24992 26546 24996
rect 26562 25052 26626 25056
rect 26562 24996 26566 25052
rect 26566 24996 26622 25052
rect 26622 24996 26626 25052
rect 26562 24992 26626 24996
rect 26642 25052 26706 25056
rect 26642 24996 26646 25052
rect 26646 24996 26702 25052
rect 26702 24996 26706 25052
rect 26642 24992 26706 24996
rect 4493 24508 4557 24512
rect 4493 24452 4497 24508
rect 4497 24452 4553 24508
rect 4553 24452 4557 24508
rect 4493 24448 4557 24452
rect 4573 24508 4637 24512
rect 4573 24452 4577 24508
rect 4577 24452 4633 24508
rect 4633 24452 4637 24508
rect 4573 24448 4637 24452
rect 4653 24508 4717 24512
rect 4653 24452 4657 24508
rect 4657 24452 4713 24508
rect 4713 24452 4717 24508
rect 4653 24448 4717 24452
rect 4733 24508 4797 24512
rect 4733 24452 4737 24508
rect 4737 24452 4793 24508
rect 4793 24452 4797 24508
rect 4733 24448 4797 24452
rect 11576 24508 11640 24512
rect 11576 24452 11580 24508
rect 11580 24452 11636 24508
rect 11636 24452 11640 24508
rect 11576 24448 11640 24452
rect 11656 24508 11720 24512
rect 11656 24452 11660 24508
rect 11660 24452 11716 24508
rect 11716 24452 11720 24508
rect 11656 24448 11720 24452
rect 11736 24508 11800 24512
rect 11736 24452 11740 24508
rect 11740 24452 11796 24508
rect 11796 24452 11800 24508
rect 11736 24448 11800 24452
rect 11816 24508 11880 24512
rect 11816 24452 11820 24508
rect 11820 24452 11876 24508
rect 11876 24452 11880 24508
rect 11816 24448 11880 24452
rect 18659 24508 18723 24512
rect 18659 24452 18663 24508
rect 18663 24452 18719 24508
rect 18719 24452 18723 24508
rect 18659 24448 18723 24452
rect 18739 24508 18803 24512
rect 18739 24452 18743 24508
rect 18743 24452 18799 24508
rect 18799 24452 18803 24508
rect 18739 24448 18803 24452
rect 18819 24508 18883 24512
rect 18819 24452 18823 24508
rect 18823 24452 18879 24508
rect 18879 24452 18883 24508
rect 18819 24448 18883 24452
rect 18899 24508 18963 24512
rect 18899 24452 18903 24508
rect 18903 24452 18959 24508
rect 18959 24452 18963 24508
rect 18899 24448 18963 24452
rect 25742 24508 25806 24512
rect 25742 24452 25746 24508
rect 25746 24452 25802 24508
rect 25802 24452 25806 24508
rect 25742 24448 25806 24452
rect 25822 24508 25886 24512
rect 25822 24452 25826 24508
rect 25826 24452 25882 24508
rect 25882 24452 25886 24508
rect 25822 24448 25886 24452
rect 25902 24508 25966 24512
rect 25902 24452 25906 24508
rect 25906 24452 25962 24508
rect 25962 24452 25966 24508
rect 25902 24448 25966 24452
rect 25982 24508 26046 24512
rect 25982 24452 25986 24508
rect 25986 24452 26042 24508
rect 26042 24452 26046 24508
rect 25982 24448 26046 24452
rect 5153 23964 5217 23968
rect 5153 23908 5157 23964
rect 5157 23908 5213 23964
rect 5213 23908 5217 23964
rect 5153 23904 5217 23908
rect 5233 23964 5297 23968
rect 5233 23908 5237 23964
rect 5237 23908 5293 23964
rect 5293 23908 5297 23964
rect 5233 23904 5297 23908
rect 5313 23964 5377 23968
rect 5313 23908 5317 23964
rect 5317 23908 5373 23964
rect 5373 23908 5377 23964
rect 5313 23904 5377 23908
rect 5393 23964 5457 23968
rect 5393 23908 5397 23964
rect 5397 23908 5453 23964
rect 5453 23908 5457 23964
rect 5393 23904 5457 23908
rect 12236 23964 12300 23968
rect 12236 23908 12240 23964
rect 12240 23908 12296 23964
rect 12296 23908 12300 23964
rect 12236 23904 12300 23908
rect 12316 23964 12380 23968
rect 12316 23908 12320 23964
rect 12320 23908 12376 23964
rect 12376 23908 12380 23964
rect 12316 23904 12380 23908
rect 12396 23964 12460 23968
rect 12396 23908 12400 23964
rect 12400 23908 12456 23964
rect 12456 23908 12460 23964
rect 12396 23904 12460 23908
rect 12476 23964 12540 23968
rect 12476 23908 12480 23964
rect 12480 23908 12536 23964
rect 12536 23908 12540 23964
rect 12476 23904 12540 23908
rect 19319 23964 19383 23968
rect 19319 23908 19323 23964
rect 19323 23908 19379 23964
rect 19379 23908 19383 23964
rect 19319 23904 19383 23908
rect 19399 23964 19463 23968
rect 19399 23908 19403 23964
rect 19403 23908 19459 23964
rect 19459 23908 19463 23964
rect 19399 23904 19463 23908
rect 19479 23964 19543 23968
rect 19479 23908 19483 23964
rect 19483 23908 19539 23964
rect 19539 23908 19543 23964
rect 19479 23904 19543 23908
rect 19559 23964 19623 23968
rect 19559 23908 19563 23964
rect 19563 23908 19619 23964
rect 19619 23908 19623 23964
rect 19559 23904 19623 23908
rect 26402 23964 26466 23968
rect 26402 23908 26406 23964
rect 26406 23908 26462 23964
rect 26462 23908 26466 23964
rect 26402 23904 26466 23908
rect 26482 23964 26546 23968
rect 26482 23908 26486 23964
rect 26486 23908 26542 23964
rect 26542 23908 26546 23964
rect 26482 23904 26546 23908
rect 26562 23964 26626 23968
rect 26562 23908 26566 23964
rect 26566 23908 26622 23964
rect 26622 23908 26626 23964
rect 26562 23904 26626 23908
rect 26642 23964 26706 23968
rect 26642 23908 26646 23964
rect 26646 23908 26702 23964
rect 26702 23908 26706 23964
rect 26642 23904 26706 23908
rect 4493 23420 4557 23424
rect 4493 23364 4497 23420
rect 4497 23364 4553 23420
rect 4553 23364 4557 23420
rect 4493 23360 4557 23364
rect 4573 23420 4637 23424
rect 4573 23364 4577 23420
rect 4577 23364 4633 23420
rect 4633 23364 4637 23420
rect 4573 23360 4637 23364
rect 4653 23420 4717 23424
rect 4653 23364 4657 23420
rect 4657 23364 4713 23420
rect 4713 23364 4717 23420
rect 4653 23360 4717 23364
rect 4733 23420 4797 23424
rect 4733 23364 4737 23420
rect 4737 23364 4793 23420
rect 4793 23364 4797 23420
rect 4733 23360 4797 23364
rect 11576 23420 11640 23424
rect 11576 23364 11580 23420
rect 11580 23364 11636 23420
rect 11636 23364 11640 23420
rect 11576 23360 11640 23364
rect 11656 23420 11720 23424
rect 11656 23364 11660 23420
rect 11660 23364 11716 23420
rect 11716 23364 11720 23420
rect 11656 23360 11720 23364
rect 11736 23420 11800 23424
rect 11736 23364 11740 23420
rect 11740 23364 11796 23420
rect 11796 23364 11800 23420
rect 11736 23360 11800 23364
rect 11816 23420 11880 23424
rect 11816 23364 11820 23420
rect 11820 23364 11876 23420
rect 11876 23364 11880 23420
rect 11816 23360 11880 23364
rect 18659 23420 18723 23424
rect 18659 23364 18663 23420
rect 18663 23364 18719 23420
rect 18719 23364 18723 23420
rect 18659 23360 18723 23364
rect 18739 23420 18803 23424
rect 18739 23364 18743 23420
rect 18743 23364 18799 23420
rect 18799 23364 18803 23420
rect 18739 23360 18803 23364
rect 18819 23420 18883 23424
rect 18819 23364 18823 23420
rect 18823 23364 18879 23420
rect 18879 23364 18883 23420
rect 18819 23360 18883 23364
rect 18899 23420 18963 23424
rect 18899 23364 18903 23420
rect 18903 23364 18959 23420
rect 18959 23364 18963 23420
rect 18899 23360 18963 23364
rect 25742 23420 25806 23424
rect 25742 23364 25746 23420
rect 25746 23364 25802 23420
rect 25802 23364 25806 23420
rect 25742 23360 25806 23364
rect 25822 23420 25886 23424
rect 25822 23364 25826 23420
rect 25826 23364 25882 23420
rect 25882 23364 25886 23420
rect 25822 23360 25886 23364
rect 25902 23420 25966 23424
rect 25902 23364 25906 23420
rect 25906 23364 25962 23420
rect 25962 23364 25966 23420
rect 25902 23360 25966 23364
rect 25982 23420 26046 23424
rect 25982 23364 25986 23420
rect 25986 23364 26042 23420
rect 26042 23364 26046 23420
rect 25982 23360 26046 23364
rect 5153 22876 5217 22880
rect 5153 22820 5157 22876
rect 5157 22820 5213 22876
rect 5213 22820 5217 22876
rect 5153 22816 5217 22820
rect 5233 22876 5297 22880
rect 5233 22820 5237 22876
rect 5237 22820 5293 22876
rect 5293 22820 5297 22876
rect 5233 22816 5297 22820
rect 5313 22876 5377 22880
rect 5313 22820 5317 22876
rect 5317 22820 5373 22876
rect 5373 22820 5377 22876
rect 5313 22816 5377 22820
rect 5393 22876 5457 22880
rect 5393 22820 5397 22876
rect 5397 22820 5453 22876
rect 5453 22820 5457 22876
rect 5393 22816 5457 22820
rect 12236 22876 12300 22880
rect 12236 22820 12240 22876
rect 12240 22820 12296 22876
rect 12296 22820 12300 22876
rect 12236 22816 12300 22820
rect 12316 22876 12380 22880
rect 12316 22820 12320 22876
rect 12320 22820 12376 22876
rect 12376 22820 12380 22876
rect 12316 22816 12380 22820
rect 12396 22876 12460 22880
rect 12396 22820 12400 22876
rect 12400 22820 12456 22876
rect 12456 22820 12460 22876
rect 12396 22816 12460 22820
rect 12476 22876 12540 22880
rect 12476 22820 12480 22876
rect 12480 22820 12536 22876
rect 12536 22820 12540 22876
rect 12476 22816 12540 22820
rect 19319 22876 19383 22880
rect 19319 22820 19323 22876
rect 19323 22820 19379 22876
rect 19379 22820 19383 22876
rect 19319 22816 19383 22820
rect 19399 22876 19463 22880
rect 19399 22820 19403 22876
rect 19403 22820 19459 22876
rect 19459 22820 19463 22876
rect 19399 22816 19463 22820
rect 19479 22876 19543 22880
rect 19479 22820 19483 22876
rect 19483 22820 19539 22876
rect 19539 22820 19543 22876
rect 19479 22816 19543 22820
rect 19559 22876 19623 22880
rect 19559 22820 19563 22876
rect 19563 22820 19619 22876
rect 19619 22820 19623 22876
rect 19559 22816 19623 22820
rect 26402 22876 26466 22880
rect 26402 22820 26406 22876
rect 26406 22820 26462 22876
rect 26462 22820 26466 22876
rect 26402 22816 26466 22820
rect 26482 22876 26546 22880
rect 26482 22820 26486 22876
rect 26486 22820 26542 22876
rect 26542 22820 26546 22876
rect 26482 22816 26546 22820
rect 26562 22876 26626 22880
rect 26562 22820 26566 22876
rect 26566 22820 26622 22876
rect 26622 22820 26626 22876
rect 26562 22816 26626 22820
rect 26642 22876 26706 22880
rect 26642 22820 26646 22876
rect 26646 22820 26702 22876
rect 26702 22820 26706 22876
rect 26642 22816 26706 22820
rect 24348 22476 24412 22540
rect 4493 22332 4557 22336
rect 4493 22276 4497 22332
rect 4497 22276 4553 22332
rect 4553 22276 4557 22332
rect 4493 22272 4557 22276
rect 4573 22332 4637 22336
rect 4573 22276 4577 22332
rect 4577 22276 4633 22332
rect 4633 22276 4637 22332
rect 4573 22272 4637 22276
rect 4653 22332 4717 22336
rect 4653 22276 4657 22332
rect 4657 22276 4713 22332
rect 4713 22276 4717 22332
rect 4653 22272 4717 22276
rect 4733 22332 4797 22336
rect 4733 22276 4737 22332
rect 4737 22276 4793 22332
rect 4793 22276 4797 22332
rect 4733 22272 4797 22276
rect 11576 22332 11640 22336
rect 11576 22276 11580 22332
rect 11580 22276 11636 22332
rect 11636 22276 11640 22332
rect 11576 22272 11640 22276
rect 11656 22332 11720 22336
rect 11656 22276 11660 22332
rect 11660 22276 11716 22332
rect 11716 22276 11720 22332
rect 11656 22272 11720 22276
rect 11736 22332 11800 22336
rect 11736 22276 11740 22332
rect 11740 22276 11796 22332
rect 11796 22276 11800 22332
rect 11736 22272 11800 22276
rect 11816 22332 11880 22336
rect 11816 22276 11820 22332
rect 11820 22276 11876 22332
rect 11876 22276 11880 22332
rect 11816 22272 11880 22276
rect 18659 22332 18723 22336
rect 18659 22276 18663 22332
rect 18663 22276 18719 22332
rect 18719 22276 18723 22332
rect 18659 22272 18723 22276
rect 18739 22332 18803 22336
rect 18739 22276 18743 22332
rect 18743 22276 18799 22332
rect 18799 22276 18803 22332
rect 18739 22272 18803 22276
rect 18819 22332 18883 22336
rect 18819 22276 18823 22332
rect 18823 22276 18879 22332
rect 18879 22276 18883 22332
rect 18819 22272 18883 22276
rect 18899 22332 18963 22336
rect 18899 22276 18903 22332
rect 18903 22276 18959 22332
rect 18959 22276 18963 22332
rect 18899 22272 18963 22276
rect 25742 22332 25806 22336
rect 25742 22276 25746 22332
rect 25746 22276 25802 22332
rect 25802 22276 25806 22332
rect 25742 22272 25806 22276
rect 25822 22332 25886 22336
rect 25822 22276 25826 22332
rect 25826 22276 25882 22332
rect 25882 22276 25886 22332
rect 25822 22272 25886 22276
rect 25902 22332 25966 22336
rect 25902 22276 25906 22332
rect 25906 22276 25962 22332
rect 25962 22276 25966 22332
rect 25902 22272 25966 22276
rect 25982 22332 26046 22336
rect 25982 22276 25986 22332
rect 25986 22276 26042 22332
rect 26042 22276 26046 22332
rect 25982 22272 26046 22276
rect 5153 21788 5217 21792
rect 5153 21732 5157 21788
rect 5157 21732 5213 21788
rect 5213 21732 5217 21788
rect 5153 21728 5217 21732
rect 5233 21788 5297 21792
rect 5233 21732 5237 21788
rect 5237 21732 5293 21788
rect 5293 21732 5297 21788
rect 5233 21728 5297 21732
rect 5313 21788 5377 21792
rect 5313 21732 5317 21788
rect 5317 21732 5373 21788
rect 5373 21732 5377 21788
rect 5313 21728 5377 21732
rect 5393 21788 5457 21792
rect 5393 21732 5397 21788
rect 5397 21732 5453 21788
rect 5453 21732 5457 21788
rect 5393 21728 5457 21732
rect 12236 21788 12300 21792
rect 12236 21732 12240 21788
rect 12240 21732 12296 21788
rect 12296 21732 12300 21788
rect 12236 21728 12300 21732
rect 12316 21788 12380 21792
rect 12316 21732 12320 21788
rect 12320 21732 12376 21788
rect 12376 21732 12380 21788
rect 12316 21728 12380 21732
rect 12396 21788 12460 21792
rect 12396 21732 12400 21788
rect 12400 21732 12456 21788
rect 12456 21732 12460 21788
rect 12396 21728 12460 21732
rect 12476 21788 12540 21792
rect 12476 21732 12480 21788
rect 12480 21732 12536 21788
rect 12536 21732 12540 21788
rect 12476 21728 12540 21732
rect 19319 21788 19383 21792
rect 19319 21732 19323 21788
rect 19323 21732 19379 21788
rect 19379 21732 19383 21788
rect 19319 21728 19383 21732
rect 19399 21788 19463 21792
rect 19399 21732 19403 21788
rect 19403 21732 19459 21788
rect 19459 21732 19463 21788
rect 19399 21728 19463 21732
rect 19479 21788 19543 21792
rect 19479 21732 19483 21788
rect 19483 21732 19539 21788
rect 19539 21732 19543 21788
rect 19479 21728 19543 21732
rect 19559 21788 19623 21792
rect 19559 21732 19563 21788
rect 19563 21732 19619 21788
rect 19619 21732 19623 21788
rect 19559 21728 19623 21732
rect 26402 21788 26466 21792
rect 26402 21732 26406 21788
rect 26406 21732 26462 21788
rect 26462 21732 26466 21788
rect 26402 21728 26466 21732
rect 26482 21788 26546 21792
rect 26482 21732 26486 21788
rect 26486 21732 26542 21788
rect 26542 21732 26546 21788
rect 26482 21728 26546 21732
rect 26562 21788 26626 21792
rect 26562 21732 26566 21788
rect 26566 21732 26622 21788
rect 26622 21732 26626 21788
rect 26562 21728 26626 21732
rect 26642 21788 26706 21792
rect 26642 21732 26646 21788
rect 26646 21732 26702 21788
rect 26702 21732 26706 21788
rect 26642 21728 26706 21732
rect 4493 21244 4557 21248
rect 4493 21188 4497 21244
rect 4497 21188 4553 21244
rect 4553 21188 4557 21244
rect 4493 21184 4557 21188
rect 4573 21244 4637 21248
rect 4573 21188 4577 21244
rect 4577 21188 4633 21244
rect 4633 21188 4637 21244
rect 4573 21184 4637 21188
rect 4653 21244 4717 21248
rect 4653 21188 4657 21244
rect 4657 21188 4713 21244
rect 4713 21188 4717 21244
rect 4653 21184 4717 21188
rect 4733 21244 4797 21248
rect 4733 21188 4737 21244
rect 4737 21188 4793 21244
rect 4793 21188 4797 21244
rect 4733 21184 4797 21188
rect 11576 21244 11640 21248
rect 11576 21188 11580 21244
rect 11580 21188 11636 21244
rect 11636 21188 11640 21244
rect 11576 21184 11640 21188
rect 11656 21244 11720 21248
rect 11656 21188 11660 21244
rect 11660 21188 11716 21244
rect 11716 21188 11720 21244
rect 11656 21184 11720 21188
rect 11736 21244 11800 21248
rect 11736 21188 11740 21244
rect 11740 21188 11796 21244
rect 11796 21188 11800 21244
rect 11736 21184 11800 21188
rect 11816 21244 11880 21248
rect 11816 21188 11820 21244
rect 11820 21188 11876 21244
rect 11876 21188 11880 21244
rect 11816 21184 11880 21188
rect 18659 21244 18723 21248
rect 18659 21188 18663 21244
rect 18663 21188 18719 21244
rect 18719 21188 18723 21244
rect 18659 21184 18723 21188
rect 18739 21244 18803 21248
rect 18739 21188 18743 21244
rect 18743 21188 18799 21244
rect 18799 21188 18803 21244
rect 18739 21184 18803 21188
rect 18819 21244 18883 21248
rect 18819 21188 18823 21244
rect 18823 21188 18879 21244
rect 18879 21188 18883 21244
rect 18819 21184 18883 21188
rect 18899 21244 18963 21248
rect 18899 21188 18903 21244
rect 18903 21188 18959 21244
rect 18959 21188 18963 21244
rect 18899 21184 18963 21188
rect 25742 21244 25806 21248
rect 25742 21188 25746 21244
rect 25746 21188 25802 21244
rect 25802 21188 25806 21244
rect 25742 21184 25806 21188
rect 25822 21244 25886 21248
rect 25822 21188 25826 21244
rect 25826 21188 25882 21244
rect 25882 21188 25886 21244
rect 25822 21184 25886 21188
rect 25902 21244 25966 21248
rect 25902 21188 25906 21244
rect 25906 21188 25962 21244
rect 25962 21188 25966 21244
rect 25902 21184 25966 21188
rect 25982 21244 26046 21248
rect 25982 21188 25986 21244
rect 25986 21188 26042 21244
rect 26042 21188 26046 21244
rect 25982 21184 26046 21188
rect 5153 20700 5217 20704
rect 5153 20644 5157 20700
rect 5157 20644 5213 20700
rect 5213 20644 5217 20700
rect 5153 20640 5217 20644
rect 5233 20700 5297 20704
rect 5233 20644 5237 20700
rect 5237 20644 5293 20700
rect 5293 20644 5297 20700
rect 5233 20640 5297 20644
rect 5313 20700 5377 20704
rect 5313 20644 5317 20700
rect 5317 20644 5373 20700
rect 5373 20644 5377 20700
rect 5313 20640 5377 20644
rect 5393 20700 5457 20704
rect 5393 20644 5397 20700
rect 5397 20644 5453 20700
rect 5453 20644 5457 20700
rect 5393 20640 5457 20644
rect 12236 20700 12300 20704
rect 12236 20644 12240 20700
rect 12240 20644 12296 20700
rect 12296 20644 12300 20700
rect 12236 20640 12300 20644
rect 12316 20700 12380 20704
rect 12316 20644 12320 20700
rect 12320 20644 12376 20700
rect 12376 20644 12380 20700
rect 12316 20640 12380 20644
rect 12396 20700 12460 20704
rect 12396 20644 12400 20700
rect 12400 20644 12456 20700
rect 12456 20644 12460 20700
rect 12396 20640 12460 20644
rect 12476 20700 12540 20704
rect 12476 20644 12480 20700
rect 12480 20644 12536 20700
rect 12536 20644 12540 20700
rect 12476 20640 12540 20644
rect 19319 20700 19383 20704
rect 19319 20644 19323 20700
rect 19323 20644 19379 20700
rect 19379 20644 19383 20700
rect 19319 20640 19383 20644
rect 19399 20700 19463 20704
rect 19399 20644 19403 20700
rect 19403 20644 19459 20700
rect 19459 20644 19463 20700
rect 19399 20640 19463 20644
rect 19479 20700 19543 20704
rect 19479 20644 19483 20700
rect 19483 20644 19539 20700
rect 19539 20644 19543 20700
rect 19479 20640 19543 20644
rect 19559 20700 19623 20704
rect 19559 20644 19563 20700
rect 19563 20644 19619 20700
rect 19619 20644 19623 20700
rect 19559 20640 19623 20644
rect 26402 20700 26466 20704
rect 26402 20644 26406 20700
rect 26406 20644 26462 20700
rect 26462 20644 26466 20700
rect 26402 20640 26466 20644
rect 26482 20700 26546 20704
rect 26482 20644 26486 20700
rect 26486 20644 26542 20700
rect 26542 20644 26546 20700
rect 26482 20640 26546 20644
rect 26562 20700 26626 20704
rect 26562 20644 26566 20700
rect 26566 20644 26622 20700
rect 26622 20644 26626 20700
rect 26562 20640 26626 20644
rect 26642 20700 26706 20704
rect 26642 20644 26646 20700
rect 26646 20644 26702 20700
rect 26702 20644 26706 20700
rect 26642 20640 26706 20644
rect 4493 20156 4557 20160
rect 4493 20100 4497 20156
rect 4497 20100 4553 20156
rect 4553 20100 4557 20156
rect 4493 20096 4557 20100
rect 4573 20156 4637 20160
rect 4573 20100 4577 20156
rect 4577 20100 4633 20156
rect 4633 20100 4637 20156
rect 4573 20096 4637 20100
rect 4653 20156 4717 20160
rect 4653 20100 4657 20156
rect 4657 20100 4713 20156
rect 4713 20100 4717 20156
rect 4653 20096 4717 20100
rect 4733 20156 4797 20160
rect 4733 20100 4737 20156
rect 4737 20100 4793 20156
rect 4793 20100 4797 20156
rect 4733 20096 4797 20100
rect 11576 20156 11640 20160
rect 11576 20100 11580 20156
rect 11580 20100 11636 20156
rect 11636 20100 11640 20156
rect 11576 20096 11640 20100
rect 11656 20156 11720 20160
rect 11656 20100 11660 20156
rect 11660 20100 11716 20156
rect 11716 20100 11720 20156
rect 11656 20096 11720 20100
rect 11736 20156 11800 20160
rect 11736 20100 11740 20156
rect 11740 20100 11796 20156
rect 11796 20100 11800 20156
rect 11736 20096 11800 20100
rect 11816 20156 11880 20160
rect 11816 20100 11820 20156
rect 11820 20100 11876 20156
rect 11876 20100 11880 20156
rect 11816 20096 11880 20100
rect 18659 20156 18723 20160
rect 18659 20100 18663 20156
rect 18663 20100 18719 20156
rect 18719 20100 18723 20156
rect 18659 20096 18723 20100
rect 18739 20156 18803 20160
rect 18739 20100 18743 20156
rect 18743 20100 18799 20156
rect 18799 20100 18803 20156
rect 18739 20096 18803 20100
rect 18819 20156 18883 20160
rect 18819 20100 18823 20156
rect 18823 20100 18879 20156
rect 18879 20100 18883 20156
rect 18819 20096 18883 20100
rect 18899 20156 18963 20160
rect 18899 20100 18903 20156
rect 18903 20100 18959 20156
rect 18959 20100 18963 20156
rect 18899 20096 18963 20100
rect 25742 20156 25806 20160
rect 25742 20100 25746 20156
rect 25746 20100 25802 20156
rect 25802 20100 25806 20156
rect 25742 20096 25806 20100
rect 25822 20156 25886 20160
rect 25822 20100 25826 20156
rect 25826 20100 25882 20156
rect 25882 20100 25886 20156
rect 25822 20096 25886 20100
rect 25902 20156 25966 20160
rect 25902 20100 25906 20156
rect 25906 20100 25962 20156
rect 25962 20100 25966 20156
rect 25902 20096 25966 20100
rect 25982 20156 26046 20160
rect 25982 20100 25986 20156
rect 25986 20100 26042 20156
rect 26042 20100 26046 20156
rect 25982 20096 26046 20100
rect 5153 19612 5217 19616
rect 5153 19556 5157 19612
rect 5157 19556 5213 19612
rect 5213 19556 5217 19612
rect 5153 19552 5217 19556
rect 5233 19612 5297 19616
rect 5233 19556 5237 19612
rect 5237 19556 5293 19612
rect 5293 19556 5297 19612
rect 5233 19552 5297 19556
rect 5313 19612 5377 19616
rect 5313 19556 5317 19612
rect 5317 19556 5373 19612
rect 5373 19556 5377 19612
rect 5313 19552 5377 19556
rect 5393 19612 5457 19616
rect 5393 19556 5397 19612
rect 5397 19556 5453 19612
rect 5453 19556 5457 19612
rect 5393 19552 5457 19556
rect 12236 19612 12300 19616
rect 12236 19556 12240 19612
rect 12240 19556 12296 19612
rect 12296 19556 12300 19612
rect 12236 19552 12300 19556
rect 12316 19612 12380 19616
rect 12316 19556 12320 19612
rect 12320 19556 12376 19612
rect 12376 19556 12380 19612
rect 12316 19552 12380 19556
rect 12396 19612 12460 19616
rect 12396 19556 12400 19612
rect 12400 19556 12456 19612
rect 12456 19556 12460 19612
rect 12396 19552 12460 19556
rect 12476 19612 12540 19616
rect 12476 19556 12480 19612
rect 12480 19556 12536 19612
rect 12536 19556 12540 19612
rect 12476 19552 12540 19556
rect 19319 19612 19383 19616
rect 19319 19556 19323 19612
rect 19323 19556 19379 19612
rect 19379 19556 19383 19612
rect 19319 19552 19383 19556
rect 19399 19612 19463 19616
rect 19399 19556 19403 19612
rect 19403 19556 19459 19612
rect 19459 19556 19463 19612
rect 19399 19552 19463 19556
rect 19479 19612 19543 19616
rect 19479 19556 19483 19612
rect 19483 19556 19539 19612
rect 19539 19556 19543 19612
rect 19479 19552 19543 19556
rect 19559 19612 19623 19616
rect 19559 19556 19563 19612
rect 19563 19556 19619 19612
rect 19619 19556 19623 19612
rect 19559 19552 19623 19556
rect 26402 19612 26466 19616
rect 26402 19556 26406 19612
rect 26406 19556 26462 19612
rect 26462 19556 26466 19612
rect 26402 19552 26466 19556
rect 26482 19612 26546 19616
rect 26482 19556 26486 19612
rect 26486 19556 26542 19612
rect 26542 19556 26546 19612
rect 26482 19552 26546 19556
rect 26562 19612 26626 19616
rect 26562 19556 26566 19612
rect 26566 19556 26622 19612
rect 26622 19556 26626 19612
rect 26562 19552 26626 19556
rect 26642 19612 26706 19616
rect 26642 19556 26646 19612
rect 26646 19556 26702 19612
rect 26702 19556 26706 19612
rect 26642 19552 26706 19556
rect 4493 19068 4557 19072
rect 4493 19012 4497 19068
rect 4497 19012 4553 19068
rect 4553 19012 4557 19068
rect 4493 19008 4557 19012
rect 4573 19068 4637 19072
rect 4573 19012 4577 19068
rect 4577 19012 4633 19068
rect 4633 19012 4637 19068
rect 4573 19008 4637 19012
rect 4653 19068 4717 19072
rect 4653 19012 4657 19068
rect 4657 19012 4713 19068
rect 4713 19012 4717 19068
rect 4653 19008 4717 19012
rect 4733 19068 4797 19072
rect 4733 19012 4737 19068
rect 4737 19012 4793 19068
rect 4793 19012 4797 19068
rect 4733 19008 4797 19012
rect 11576 19068 11640 19072
rect 11576 19012 11580 19068
rect 11580 19012 11636 19068
rect 11636 19012 11640 19068
rect 11576 19008 11640 19012
rect 11656 19068 11720 19072
rect 11656 19012 11660 19068
rect 11660 19012 11716 19068
rect 11716 19012 11720 19068
rect 11656 19008 11720 19012
rect 11736 19068 11800 19072
rect 11736 19012 11740 19068
rect 11740 19012 11796 19068
rect 11796 19012 11800 19068
rect 11736 19008 11800 19012
rect 11816 19068 11880 19072
rect 11816 19012 11820 19068
rect 11820 19012 11876 19068
rect 11876 19012 11880 19068
rect 11816 19008 11880 19012
rect 18659 19068 18723 19072
rect 18659 19012 18663 19068
rect 18663 19012 18719 19068
rect 18719 19012 18723 19068
rect 18659 19008 18723 19012
rect 18739 19068 18803 19072
rect 18739 19012 18743 19068
rect 18743 19012 18799 19068
rect 18799 19012 18803 19068
rect 18739 19008 18803 19012
rect 18819 19068 18883 19072
rect 18819 19012 18823 19068
rect 18823 19012 18879 19068
rect 18879 19012 18883 19068
rect 18819 19008 18883 19012
rect 18899 19068 18963 19072
rect 18899 19012 18903 19068
rect 18903 19012 18959 19068
rect 18959 19012 18963 19068
rect 18899 19008 18963 19012
rect 25742 19068 25806 19072
rect 25742 19012 25746 19068
rect 25746 19012 25802 19068
rect 25802 19012 25806 19068
rect 25742 19008 25806 19012
rect 25822 19068 25886 19072
rect 25822 19012 25826 19068
rect 25826 19012 25882 19068
rect 25882 19012 25886 19068
rect 25822 19008 25886 19012
rect 25902 19068 25966 19072
rect 25902 19012 25906 19068
rect 25906 19012 25962 19068
rect 25962 19012 25966 19068
rect 25902 19008 25966 19012
rect 25982 19068 26046 19072
rect 25982 19012 25986 19068
rect 25986 19012 26042 19068
rect 26042 19012 26046 19068
rect 25982 19008 26046 19012
rect 5153 18524 5217 18528
rect 5153 18468 5157 18524
rect 5157 18468 5213 18524
rect 5213 18468 5217 18524
rect 5153 18464 5217 18468
rect 5233 18524 5297 18528
rect 5233 18468 5237 18524
rect 5237 18468 5293 18524
rect 5293 18468 5297 18524
rect 5233 18464 5297 18468
rect 5313 18524 5377 18528
rect 5313 18468 5317 18524
rect 5317 18468 5373 18524
rect 5373 18468 5377 18524
rect 5313 18464 5377 18468
rect 5393 18524 5457 18528
rect 5393 18468 5397 18524
rect 5397 18468 5453 18524
rect 5453 18468 5457 18524
rect 5393 18464 5457 18468
rect 12236 18524 12300 18528
rect 12236 18468 12240 18524
rect 12240 18468 12296 18524
rect 12296 18468 12300 18524
rect 12236 18464 12300 18468
rect 12316 18524 12380 18528
rect 12316 18468 12320 18524
rect 12320 18468 12376 18524
rect 12376 18468 12380 18524
rect 12316 18464 12380 18468
rect 12396 18524 12460 18528
rect 12396 18468 12400 18524
rect 12400 18468 12456 18524
rect 12456 18468 12460 18524
rect 12396 18464 12460 18468
rect 12476 18524 12540 18528
rect 12476 18468 12480 18524
rect 12480 18468 12536 18524
rect 12536 18468 12540 18524
rect 12476 18464 12540 18468
rect 19319 18524 19383 18528
rect 19319 18468 19323 18524
rect 19323 18468 19379 18524
rect 19379 18468 19383 18524
rect 19319 18464 19383 18468
rect 19399 18524 19463 18528
rect 19399 18468 19403 18524
rect 19403 18468 19459 18524
rect 19459 18468 19463 18524
rect 19399 18464 19463 18468
rect 19479 18524 19543 18528
rect 19479 18468 19483 18524
rect 19483 18468 19539 18524
rect 19539 18468 19543 18524
rect 19479 18464 19543 18468
rect 19559 18524 19623 18528
rect 19559 18468 19563 18524
rect 19563 18468 19619 18524
rect 19619 18468 19623 18524
rect 19559 18464 19623 18468
rect 26402 18524 26466 18528
rect 26402 18468 26406 18524
rect 26406 18468 26462 18524
rect 26462 18468 26466 18524
rect 26402 18464 26466 18468
rect 26482 18524 26546 18528
rect 26482 18468 26486 18524
rect 26486 18468 26542 18524
rect 26542 18468 26546 18524
rect 26482 18464 26546 18468
rect 26562 18524 26626 18528
rect 26562 18468 26566 18524
rect 26566 18468 26622 18524
rect 26622 18468 26626 18524
rect 26562 18464 26626 18468
rect 26642 18524 26706 18528
rect 26642 18468 26646 18524
rect 26646 18468 26702 18524
rect 26702 18468 26706 18524
rect 26642 18464 26706 18468
rect 27660 17988 27724 18052
rect 4493 17980 4557 17984
rect 4493 17924 4497 17980
rect 4497 17924 4553 17980
rect 4553 17924 4557 17980
rect 4493 17920 4557 17924
rect 4573 17980 4637 17984
rect 4573 17924 4577 17980
rect 4577 17924 4633 17980
rect 4633 17924 4637 17980
rect 4573 17920 4637 17924
rect 4653 17980 4717 17984
rect 4653 17924 4657 17980
rect 4657 17924 4713 17980
rect 4713 17924 4717 17980
rect 4653 17920 4717 17924
rect 4733 17980 4797 17984
rect 4733 17924 4737 17980
rect 4737 17924 4793 17980
rect 4793 17924 4797 17980
rect 4733 17920 4797 17924
rect 11576 17980 11640 17984
rect 11576 17924 11580 17980
rect 11580 17924 11636 17980
rect 11636 17924 11640 17980
rect 11576 17920 11640 17924
rect 11656 17980 11720 17984
rect 11656 17924 11660 17980
rect 11660 17924 11716 17980
rect 11716 17924 11720 17980
rect 11656 17920 11720 17924
rect 11736 17980 11800 17984
rect 11736 17924 11740 17980
rect 11740 17924 11796 17980
rect 11796 17924 11800 17980
rect 11736 17920 11800 17924
rect 11816 17980 11880 17984
rect 11816 17924 11820 17980
rect 11820 17924 11876 17980
rect 11876 17924 11880 17980
rect 11816 17920 11880 17924
rect 18659 17980 18723 17984
rect 18659 17924 18663 17980
rect 18663 17924 18719 17980
rect 18719 17924 18723 17980
rect 18659 17920 18723 17924
rect 18739 17980 18803 17984
rect 18739 17924 18743 17980
rect 18743 17924 18799 17980
rect 18799 17924 18803 17980
rect 18739 17920 18803 17924
rect 18819 17980 18883 17984
rect 18819 17924 18823 17980
rect 18823 17924 18879 17980
rect 18879 17924 18883 17980
rect 18819 17920 18883 17924
rect 18899 17980 18963 17984
rect 18899 17924 18903 17980
rect 18903 17924 18959 17980
rect 18959 17924 18963 17980
rect 18899 17920 18963 17924
rect 25742 17980 25806 17984
rect 25742 17924 25746 17980
rect 25746 17924 25802 17980
rect 25802 17924 25806 17980
rect 25742 17920 25806 17924
rect 25822 17980 25886 17984
rect 25822 17924 25826 17980
rect 25826 17924 25882 17980
rect 25882 17924 25886 17980
rect 25822 17920 25886 17924
rect 25902 17980 25966 17984
rect 25902 17924 25906 17980
rect 25906 17924 25962 17980
rect 25962 17924 25966 17980
rect 25902 17920 25966 17924
rect 25982 17980 26046 17984
rect 25982 17924 25986 17980
rect 25986 17924 26042 17980
rect 26042 17924 26046 17980
rect 25982 17920 26046 17924
rect 5153 17436 5217 17440
rect 5153 17380 5157 17436
rect 5157 17380 5213 17436
rect 5213 17380 5217 17436
rect 5153 17376 5217 17380
rect 5233 17436 5297 17440
rect 5233 17380 5237 17436
rect 5237 17380 5293 17436
rect 5293 17380 5297 17436
rect 5233 17376 5297 17380
rect 5313 17436 5377 17440
rect 5313 17380 5317 17436
rect 5317 17380 5373 17436
rect 5373 17380 5377 17436
rect 5313 17376 5377 17380
rect 5393 17436 5457 17440
rect 5393 17380 5397 17436
rect 5397 17380 5453 17436
rect 5453 17380 5457 17436
rect 5393 17376 5457 17380
rect 12236 17436 12300 17440
rect 12236 17380 12240 17436
rect 12240 17380 12296 17436
rect 12296 17380 12300 17436
rect 12236 17376 12300 17380
rect 12316 17436 12380 17440
rect 12316 17380 12320 17436
rect 12320 17380 12376 17436
rect 12376 17380 12380 17436
rect 12316 17376 12380 17380
rect 12396 17436 12460 17440
rect 12396 17380 12400 17436
rect 12400 17380 12456 17436
rect 12456 17380 12460 17436
rect 12396 17376 12460 17380
rect 12476 17436 12540 17440
rect 12476 17380 12480 17436
rect 12480 17380 12536 17436
rect 12536 17380 12540 17436
rect 12476 17376 12540 17380
rect 19319 17436 19383 17440
rect 19319 17380 19323 17436
rect 19323 17380 19379 17436
rect 19379 17380 19383 17436
rect 19319 17376 19383 17380
rect 19399 17436 19463 17440
rect 19399 17380 19403 17436
rect 19403 17380 19459 17436
rect 19459 17380 19463 17436
rect 19399 17376 19463 17380
rect 19479 17436 19543 17440
rect 19479 17380 19483 17436
rect 19483 17380 19539 17436
rect 19539 17380 19543 17436
rect 19479 17376 19543 17380
rect 19559 17436 19623 17440
rect 19559 17380 19563 17436
rect 19563 17380 19619 17436
rect 19619 17380 19623 17436
rect 19559 17376 19623 17380
rect 26402 17436 26466 17440
rect 26402 17380 26406 17436
rect 26406 17380 26462 17436
rect 26462 17380 26466 17436
rect 26402 17376 26466 17380
rect 26482 17436 26546 17440
rect 26482 17380 26486 17436
rect 26486 17380 26542 17436
rect 26542 17380 26546 17436
rect 26482 17376 26546 17380
rect 26562 17436 26626 17440
rect 26562 17380 26566 17436
rect 26566 17380 26622 17436
rect 26622 17380 26626 17436
rect 26562 17376 26626 17380
rect 26642 17436 26706 17440
rect 26642 17380 26646 17436
rect 26646 17380 26702 17436
rect 26702 17380 26706 17436
rect 26642 17376 26706 17380
rect 4493 16892 4557 16896
rect 4493 16836 4497 16892
rect 4497 16836 4553 16892
rect 4553 16836 4557 16892
rect 4493 16832 4557 16836
rect 4573 16892 4637 16896
rect 4573 16836 4577 16892
rect 4577 16836 4633 16892
rect 4633 16836 4637 16892
rect 4573 16832 4637 16836
rect 4653 16892 4717 16896
rect 4653 16836 4657 16892
rect 4657 16836 4713 16892
rect 4713 16836 4717 16892
rect 4653 16832 4717 16836
rect 4733 16892 4797 16896
rect 4733 16836 4737 16892
rect 4737 16836 4793 16892
rect 4793 16836 4797 16892
rect 4733 16832 4797 16836
rect 11576 16892 11640 16896
rect 11576 16836 11580 16892
rect 11580 16836 11636 16892
rect 11636 16836 11640 16892
rect 11576 16832 11640 16836
rect 11656 16892 11720 16896
rect 11656 16836 11660 16892
rect 11660 16836 11716 16892
rect 11716 16836 11720 16892
rect 11656 16832 11720 16836
rect 11736 16892 11800 16896
rect 11736 16836 11740 16892
rect 11740 16836 11796 16892
rect 11796 16836 11800 16892
rect 11736 16832 11800 16836
rect 11816 16892 11880 16896
rect 11816 16836 11820 16892
rect 11820 16836 11876 16892
rect 11876 16836 11880 16892
rect 11816 16832 11880 16836
rect 18659 16892 18723 16896
rect 18659 16836 18663 16892
rect 18663 16836 18719 16892
rect 18719 16836 18723 16892
rect 18659 16832 18723 16836
rect 18739 16892 18803 16896
rect 18739 16836 18743 16892
rect 18743 16836 18799 16892
rect 18799 16836 18803 16892
rect 18739 16832 18803 16836
rect 18819 16892 18883 16896
rect 18819 16836 18823 16892
rect 18823 16836 18879 16892
rect 18879 16836 18883 16892
rect 18819 16832 18883 16836
rect 18899 16892 18963 16896
rect 18899 16836 18903 16892
rect 18903 16836 18959 16892
rect 18959 16836 18963 16892
rect 18899 16832 18963 16836
rect 25742 16892 25806 16896
rect 25742 16836 25746 16892
rect 25746 16836 25802 16892
rect 25802 16836 25806 16892
rect 25742 16832 25806 16836
rect 25822 16892 25886 16896
rect 25822 16836 25826 16892
rect 25826 16836 25882 16892
rect 25882 16836 25886 16892
rect 25822 16832 25886 16836
rect 25902 16892 25966 16896
rect 25902 16836 25906 16892
rect 25906 16836 25962 16892
rect 25962 16836 25966 16892
rect 25902 16832 25966 16836
rect 25982 16892 26046 16896
rect 25982 16836 25986 16892
rect 25986 16836 26042 16892
rect 26042 16836 26046 16892
rect 25982 16832 26046 16836
rect 5153 16348 5217 16352
rect 5153 16292 5157 16348
rect 5157 16292 5213 16348
rect 5213 16292 5217 16348
rect 5153 16288 5217 16292
rect 5233 16348 5297 16352
rect 5233 16292 5237 16348
rect 5237 16292 5293 16348
rect 5293 16292 5297 16348
rect 5233 16288 5297 16292
rect 5313 16348 5377 16352
rect 5313 16292 5317 16348
rect 5317 16292 5373 16348
rect 5373 16292 5377 16348
rect 5313 16288 5377 16292
rect 5393 16348 5457 16352
rect 5393 16292 5397 16348
rect 5397 16292 5453 16348
rect 5453 16292 5457 16348
rect 5393 16288 5457 16292
rect 12236 16348 12300 16352
rect 12236 16292 12240 16348
rect 12240 16292 12296 16348
rect 12296 16292 12300 16348
rect 12236 16288 12300 16292
rect 12316 16348 12380 16352
rect 12316 16292 12320 16348
rect 12320 16292 12376 16348
rect 12376 16292 12380 16348
rect 12316 16288 12380 16292
rect 12396 16348 12460 16352
rect 12396 16292 12400 16348
rect 12400 16292 12456 16348
rect 12456 16292 12460 16348
rect 12396 16288 12460 16292
rect 12476 16348 12540 16352
rect 12476 16292 12480 16348
rect 12480 16292 12536 16348
rect 12536 16292 12540 16348
rect 12476 16288 12540 16292
rect 19319 16348 19383 16352
rect 19319 16292 19323 16348
rect 19323 16292 19379 16348
rect 19379 16292 19383 16348
rect 19319 16288 19383 16292
rect 19399 16348 19463 16352
rect 19399 16292 19403 16348
rect 19403 16292 19459 16348
rect 19459 16292 19463 16348
rect 19399 16288 19463 16292
rect 19479 16348 19543 16352
rect 19479 16292 19483 16348
rect 19483 16292 19539 16348
rect 19539 16292 19543 16348
rect 19479 16288 19543 16292
rect 19559 16348 19623 16352
rect 19559 16292 19563 16348
rect 19563 16292 19619 16348
rect 19619 16292 19623 16348
rect 19559 16288 19623 16292
rect 26402 16348 26466 16352
rect 26402 16292 26406 16348
rect 26406 16292 26462 16348
rect 26462 16292 26466 16348
rect 26402 16288 26466 16292
rect 26482 16348 26546 16352
rect 26482 16292 26486 16348
rect 26486 16292 26542 16348
rect 26542 16292 26546 16348
rect 26482 16288 26546 16292
rect 26562 16348 26626 16352
rect 26562 16292 26566 16348
rect 26566 16292 26622 16348
rect 26622 16292 26626 16348
rect 26562 16288 26626 16292
rect 26642 16348 26706 16352
rect 26642 16292 26646 16348
rect 26646 16292 26702 16348
rect 26702 16292 26706 16348
rect 26642 16288 26706 16292
rect 4493 15804 4557 15808
rect 4493 15748 4497 15804
rect 4497 15748 4553 15804
rect 4553 15748 4557 15804
rect 4493 15744 4557 15748
rect 4573 15804 4637 15808
rect 4573 15748 4577 15804
rect 4577 15748 4633 15804
rect 4633 15748 4637 15804
rect 4573 15744 4637 15748
rect 4653 15804 4717 15808
rect 4653 15748 4657 15804
rect 4657 15748 4713 15804
rect 4713 15748 4717 15804
rect 4653 15744 4717 15748
rect 4733 15804 4797 15808
rect 4733 15748 4737 15804
rect 4737 15748 4793 15804
rect 4793 15748 4797 15804
rect 4733 15744 4797 15748
rect 11576 15804 11640 15808
rect 11576 15748 11580 15804
rect 11580 15748 11636 15804
rect 11636 15748 11640 15804
rect 11576 15744 11640 15748
rect 11656 15804 11720 15808
rect 11656 15748 11660 15804
rect 11660 15748 11716 15804
rect 11716 15748 11720 15804
rect 11656 15744 11720 15748
rect 11736 15804 11800 15808
rect 11736 15748 11740 15804
rect 11740 15748 11796 15804
rect 11796 15748 11800 15804
rect 11736 15744 11800 15748
rect 11816 15804 11880 15808
rect 11816 15748 11820 15804
rect 11820 15748 11876 15804
rect 11876 15748 11880 15804
rect 11816 15744 11880 15748
rect 18659 15804 18723 15808
rect 18659 15748 18663 15804
rect 18663 15748 18719 15804
rect 18719 15748 18723 15804
rect 18659 15744 18723 15748
rect 18739 15804 18803 15808
rect 18739 15748 18743 15804
rect 18743 15748 18799 15804
rect 18799 15748 18803 15804
rect 18739 15744 18803 15748
rect 18819 15804 18883 15808
rect 18819 15748 18823 15804
rect 18823 15748 18879 15804
rect 18879 15748 18883 15804
rect 18819 15744 18883 15748
rect 18899 15804 18963 15808
rect 18899 15748 18903 15804
rect 18903 15748 18959 15804
rect 18959 15748 18963 15804
rect 18899 15744 18963 15748
rect 25742 15804 25806 15808
rect 25742 15748 25746 15804
rect 25746 15748 25802 15804
rect 25802 15748 25806 15804
rect 25742 15744 25806 15748
rect 25822 15804 25886 15808
rect 25822 15748 25826 15804
rect 25826 15748 25882 15804
rect 25882 15748 25886 15804
rect 25822 15744 25886 15748
rect 25902 15804 25966 15808
rect 25902 15748 25906 15804
rect 25906 15748 25962 15804
rect 25962 15748 25966 15804
rect 25902 15744 25966 15748
rect 25982 15804 26046 15808
rect 25982 15748 25986 15804
rect 25986 15748 26042 15804
rect 26042 15748 26046 15804
rect 25982 15744 26046 15748
rect 5153 15260 5217 15264
rect 5153 15204 5157 15260
rect 5157 15204 5213 15260
rect 5213 15204 5217 15260
rect 5153 15200 5217 15204
rect 5233 15260 5297 15264
rect 5233 15204 5237 15260
rect 5237 15204 5293 15260
rect 5293 15204 5297 15260
rect 5233 15200 5297 15204
rect 5313 15260 5377 15264
rect 5313 15204 5317 15260
rect 5317 15204 5373 15260
rect 5373 15204 5377 15260
rect 5313 15200 5377 15204
rect 5393 15260 5457 15264
rect 5393 15204 5397 15260
rect 5397 15204 5453 15260
rect 5453 15204 5457 15260
rect 5393 15200 5457 15204
rect 12236 15260 12300 15264
rect 12236 15204 12240 15260
rect 12240 15204 12296 15260
rect 12296 15204 12300 15260
rect 12236 15200 12300 15204
rect 12316 15260 12380 15264
rect 12316 15204 12320 15260
rect 12320 15204 12376 15260
rect 12376 15204 12380 15260
rect 12316 15200 12380 15204
rect 12396 15260 12460 15264
rect 12396 15204 12400 15260
rect 12400 15204 12456 15260
rect 12456 15204 12460 15260
rect 12396 15200 12460 15204
rect 12476 15260 12540 15264
rect 12476 15204 12480 15260
rect 12480 15204 12536 15260
rect 12536 15204 12540 15260
rect 12476 15200 12540 15204
rect 19319 15260 19383 15264
rect 19319 15204 19323 15260
rect 19323 15204 19379 15260
rect 19379 15204 19383 15260
rect 19319 15200 19383 15204
rect 19399 15260 19463 15264
rect 19399 15204 19403 15260
rect 19403 15204 19459 15260
rect 19459 15204 19463 15260
rect 19399 15200 19463 15204
rect 19479 15260 19543 15264
rect 19479 15204 19483 15260
rect 19483 15204 19539 15260
rect 19539 15204 19543 15260
rect 19479 15200 19543 15204
rect 19559 15260 19623 15264
rect 19559 15204 19563 15260
rect 19563 15204 19619 15260
rect 19619 15204 19623 15260
rect 19559 15200 19623 15204
rect 26402 15260 26466 15264
rect 26402 15204 26406 15260
rect 26406 15204 26462 15260
rect 26462 15204 26466 15260
rect 26402 15200 26466 15204
rect 26482 15260 26546 15264
rect 26482 15204 26486 15260
rect 26486 15204 26542 15260
rect 26542 15204 26546 15260
rect 26482 15200 26546 15204
rect 26562 15260 26626 15264
rect 26562 15204 26566 15260
rect 26566 15204 26622 15260
rect 26622 15204 26626 15260
rect 26562 15200 26626 15204
rect 26642 15260 26706 15264
rect 26642 15204 26646 15260
rect 26646 15204 26702 15260
rect 26702 15204 26706 15260
rect 26642 15200 26706 15204
rect 4493 14716 4557 14720
rect 4493 14660 4497 14716
rect 4497 14660 4553 14716
rect 4553 14660 4557 14716
rect 4493 14656 4557 14660
rect 4573 14716 4637 14720
rect 4573 14660 4577 14716
rect 4577 14660 4633 14716
rect 4633 14660 4637 14716
rect 4573 14656 4637 14660
rect 4653 14716 4717 14720
rect 4653 14660 4657 14716
rect 4657 14660 4713 14716
rect 4713 14660 4717 14716
rect 4653 14656 4717 14660
rect 4733 14716 4797 14720
rect 4733 14660 4737 14716
rect 4737 14660 4793 14716
rect 4793 14660 4797 14716
rect 4733 14656 4797 14660
rect 11576 14716 11640 14720
rect 11576 14660 11580 14716
rect 11580 14660 11636 14716
rect 11636 14660 11640 14716
rect 11576 14656 11640 14660
rect 11656 14716 11720 14720
rect 11656 14660 11660 14716
rect 11660 14660 11716 14716
rect 11716 14660 11720 14716
rect 11656 14656 11720 14660
rect 11736 14716 11800 14720
rect 11736 14660 11740 14716
rect 11740 14660 11796 14716
rect 11796 14660 11800 14716
rect 11736 14656 11800 14660
rect 11816 14716 11880 14720
rect 11816 14660 11820 14716
rect 11820 14660 11876 14716
rect 11876 14660 11880 14716
rect 11816 14656 11880 14660
rect 18659 14716 18723 14720
rect 18659 14660 18663 14716
rect 18663 14660 18719 14716
rect 18719 14660 18723 14716
rect 18659 14656 18723 14660
rect 18739 14716 18803 14720
rect 18739 14660 18743 14716
rect 18743 14660 18799 14716
rect 18799 14660 18803 14716
rect 18739 14656 18803 14660
rect 18819 14716 18883 14720
rect 18819 14660 18823 14716
rect 18823 14660 18879 14716
rect 18879 14660 18883 14716
rect 18819 14656 18883 14660
rect 18899 14716 18963 14720
rect 18899 14660 18903 14716
rect 18903 14660 18959 14716
rect 18959 14660 18963 14716
rect 18899 14656 18963 14660
rect 25742 14716 25806 14720
rect 25742 14660 25746 14716
rect 25746 14660 25802 14716
rect 25802 14660 25806 14716
rect 25742 14656 25806 14660
rect 25822 14716 25886 14720
rect 25822 14660 25826 14716
rect 25826 14660 25882 14716
rect 25882 14660 25886 14716
rect 25822 14656 25886 14660
rect 25902 14716 25966 14720
rect 25902 14660 25906 14716
rect 25906 14660 25962 14716
rect 25962 14660 25966 14716
rect 25902 14656 25966 14660
rect 25982 14716 26046 14720
rect 25982 14660 25986 14716
rect 25986 14660 26042 14716
rect 26042 14660 26046 14716
rect 25982 14656 26046 14660
rect 5153 14172 5217 14176
rect 5153 14116 5157 14172
rect 5157 14116 5213 14172
rect 5213 14116 5217 14172
rect 5153 14112 5217 14116
rect 5233 14172 5297 14176
rect 5233 14116 5237 14172
rect 5237 14116 5293 14172
rect 5293 14116 5297 14172
rect 5233 14112 5297 14116
rect 5313 14172 5377 14176
rect 5313 14116 5317 14172
rect 5317 14116 5373 14172
rect 5373 14116 5377 14172
rect 5313 14112 5377 14116
rect 5393 14172 5457 14176
rect 5393 14116 5397 14172
rect 5397 14116 5453 14172
rect 5453 14116 5457 14172
rect 5393 14112 5457 14116
rect 12236 14172 12300 14176
rect 12236 14116 12240 14172
rect 12240 14116 12296 14172
rect 12296 14116 12300 14172
rect 12236 14112 12300 14116
rect 12316 14172 12380 14176
rect 12316 14116 12320 14172
rect 12320 14116 12376 14172
rect 12376 14116 12380 14172
rect 12316 14112 12380 14116
rect 12396 14172 12460 14176
rect 12396 14116 12400 14172
rect 12400 14116 12456 14172
rect 12456 14116 12460 14172
rect 12396 14112 12460 14116
rect 12476 14172 12540 14176
rect 12476 14116 12480 14172
rect 12480 14116 12536 14172
rect 12536 14116 12540 14172
rect 12476 14112 12540 14116
rect 19319 14172 19383 14176
rect 19319 14116 19323 14172
rect 19323 14116 19379 14172
rect 19379 14116 19383 14172
rect 19319 14112 19383 14116
rect 19399 14172 19463 14176
rect 19399 14116 19403 14172
rect 19403 14116 19459 14172
rect 19459 14116 19463 14172
rect 19399 14112 19463 14116
rect 19479 14172 19543 14176
rect 19479 14116 19483 14172
rect 19483 14116 19539 14172
rect 19539 14116 19543 14172
rect 19479 14112 19543 14116
rect 19559 14172 19623 14176
rect 19559 14116 19563 14172
rect 19563 14116 19619 14172
rect 19619 14116 19623 14172
rect 19559 14112 19623 14116
rect 26402 14172 26466 14176
rect 26402 14116 26406 14172
rect 26406 14116 26462 14172
rect 26462 14116 26466 14172
rect 26402 14112 26466 14116
rect 26482 14172 26546 14176
rect 26482 14116 26486 14172
rect 26486 14116 26542 14172
rect 26542 14116 26546 14172
rect 26482 14112 26546 14116
rect 26562 14172 26626 14176
rect 26562 14116 26566 14172
rect 26566 14116 26622 14172
rect 26622 14116 26626 14172
rect 26562 14112 26626 14116
rect 26642 14172 26706 14176
rect 26642 14116 26646 14172
rect 26646 14116 26702 14172
rect 26702 14116 26706 14172
rect 26642 14112 26706 14116
rect 10548 13832 10612 13836
rect 10548 13776 10562 13832
rect 10562 13776 10612 13832
rect 10548 13772 10612 13776
rect 4493 13628 4557 13632
rect 4493 13572 4497 13628
rect 4497 13572 4553 13628
rect 4553 13572 4557 13628
rect 4493 13568 4557 13572
rect 4573 13628 4637 13632
rect 4573 13572 4577 13628
rect 4577 13572 4633 13628
rect 4633 13572 4637 13628
rect 4573 13568 4637 13572
rect 4653 13628 4717 13632
rect 4653 13572 4657 13628
rect 4657 13572 4713 13628
rect 4713 13572 4717 13628
rect 4653 13568 4717 13572
rect 4733 13628 4797 13632
rect 4733 13572 4737 13628
rect 4737 13572 4793 13628
rect 4793 13572 4797 13628
rect 4733 13568 4797 13572
rect 11576 13628 11640 13632
rect 11576 13572 11580 13628
rect 11580 13572 11636 13628
rect 11636 13572 11640 13628
rect 11576 13568 11640 13572
rect 11656 13628 11720 13632
rect 11656 13572 11660 13628
rect 11660 13572 11716 13628
rect 11716 13572 11720 13628
rect 11656 13568 11720 13572
rect 11736 13628 11800 13632
rect 11736 13572 11740 13628
rect 11740 13572 11796 13628
rect 11796 13572 11800 13628
rect 11736 13568 11800 13572
rect 11816 13628 11880 13632
rect 11816 13572 11820 13628
rect 11820 13572 11876 13628
rect 11876 13572 11880 13628
rect 11816 13568 11880 13572
rect 18659 13628 18723 13632
rect 18659 13572 18663 13628
rect 18663 13572 18719 13628
rect 18719 13572 18723 13628
rect 18659 13568 18723 13572
rect 18739 13628 18803 13632
rect 18739 13572 18743 13628
rect 18743 13572 18799 13628
rect 18799 13572 18803 13628
rect 18739 13568 18803 13572
rect 18819 13628 18883 13632
rect 18819 13572 18823 13628
rect 18823 13572 18879 13628
rect 18879 13572 18883 13628
rect 18819 13568 18883 13572
rect 18899 13628 18963 13632
rect 18899 13572 18903 13628
rect 18903 13572 18959 13628
rect 18959 13572 18963 13628
rect 18899 13568 18963 13572
rect 25742 13628 25806 13632
rect 25742 13572 25746 13628
rect 25746 13572 25802 13628
rect 25802 13572 25806 13628
rect 25742 13568 25806 13572
rect 25822 13628 25886 13632
rect 25822 13572 25826 13628
rect 25826 13572 25882 13628
rect 25882 13572 25886 13628
rect 25822 13568 25886 13572
rect 25902 13628 25966 13632
rect 25902 13572 25906 13628
rect 25906 13572 25962 13628
rect 25962 13572 25966 13628
rect 25902 13568 25966 13572
rect 25982 13628 26046 13632
rect 25982 13572 25986 13628
rect 25986 13572 26042 13628
rect 26042 13572 26046 13628
rect 25982 13568 26046 13572
rect 10732 13228 10796 13292
rect 5153 13084 5217 13088
rect 5153 13028 5157 13084
rect 5157 13028 5213 13084
rect 5213 13028 5217 13084
rect 5153 13024 5217 13028
rect 5233 13084 5297 13088
rect 5233 13028 5237 13084
rect 5237 13028 5293 13084
rect 5293 13028 5297 13084
rect 5233 13024 5297 13028
rect 5313 13084 5377 13088
rect 5313 13028 5317 13084
rect 5317 13028 5373 13084
rect 5373 13028 5377 13084
rect 5313 13024 5377 13028
rect 5393 13084 5457 13088
rect 5393 13028 5397 13084
rect 5397 13028 5453 13084
rect 5453 13028 5457 13084
rect 5393 13024 5457 13028
rect 12236 13084 12300 13088
rect 12236 13028 12240 13084
rect 12240 13028 12296 13084
rect 12296 13028 12300 13084
rect 12236 13024 12300 13028
rect 12316 13084 12380 13088
rect 12316 13028 12320 13084
rect 12320 13028 12376 13084
rect 12376 13028 12380 13084
rect 12316 13024 12380 13028
rect 12396 13084 12460 13088
rect 12396 13028 12400 13084
rect 12400 13028 12456 13084
rect 12456 13028 12460 13084
rect 12396 13024 12460 13028
rect 12476 13084 12540 13088
rect 12476 13028 12480 13084
rect 12480 13028 12536 13084
rect 12536 13028 12540 13084
rect 12476 13024 12540 13028
rect 19319 13084 19383 13088
rect 19319 13028 19323 13084
rect 19323 13028 19379 13084
rect 19379 13028 19383 13084
rect 19319 13024 19383 13028
rect 19399 13084 19463 13088
rect 19399 13028 19403 13084
rect 19403 13028 19459 13084
rect 19459 13028 19463 13084
rect 19399 13024 19463 13028
rect 19479 13084 19543 13088
rect 19479 13028 19483 13084
rect 19483 13028 19539 13084
rect 19539 13028 19543 13084
rect 19479 13024 19543 13028
rect 19559 13084 19623 13088
rect 19559 13028 19563 13084
rect 19563 13028 19619 13084
rect 19619 13028 19623 13084
rect 19559 13024 19623 13028
rect 26402 13084 26466 13088
rect 26402 13028 26406 13084
rect 26406 13028 26462 13084
rect 26462 13028 26466 13084
rect 26402 13024 26466 13028
rect 26482 13084 26546 13088
rect 26482 13028 26486 13084
rect 26486 13028 26542 13084
rect 26542 13028 26546 13084
rect 26482 13024 26546 13028
rect 26562 13084 26626 13088
rect 26562 13028 26566 13084
rect 26566 13028 26622 13084
rect 26622 13028 26626 13084
rect 26562 13024 26626 13028
rect 26642 13084 26706 13088
rect 26642 13028 26646 13084
rect 26646 13028 26702 13084
rect 26702 13028 26706 13084
rect 26642 13024 26706 13028
rect 4493 12540 4557 12544
rect 4493 12484 4497 12540
rect 4497 12484 4553 12540
rect 4553 12484 4557 12540
rect 4493 12480 4557 12484
rect 4573 12540 4637 12544
rect 4573 12484 4577 12540
rect 4577 12484 4633 12540
rect 4633 12484 4637 12540
rect 4573 12480 4637 12484
rect 4653 12540 4717 12544
rect 4653 12484 4657 12540
rect 4657 12484 4713 12540
rect 4713 12484 4717 12540
rect 4653 12480 4717 12484
rect 4733 12540 4797 12544
rect 4733 12484 4737 12540
rect 4737 12484 4793 12540
rect 4793 12484 4797 12540
rect 4733 12480 4797 12484
rect 11576 12540 11640 12544
rect 11576 12484 11580 12540
rect 11580 12484 11636 12540
rect 11636 12484 11640 12540
rect 11576 12480 11640 12484
rect 11656 12540 11720 12544
rect 11656 12484 11660 12540
rect 11660 12484 11716 12540
rect 11716 12484 11720 12540
rect 11656 12480 11720 12484
rect 11736 12540 11800 12544
rect 11736 12484 11740 12540
rect 11740 12484 11796 12540
rect 11796 12484 11800 12540
rect 11736 12480 11800 12484
rect 11816 12540 11880 12544
rect 11816 12484 11820 12540
rect 11820 12484 11876 12540
rect 11876 12484 11880 12540
rect 11816 12480 11880 12484
rect 18659 12540 18723 12544
rect 18659 12484 18663 12540
rect 18663 12484 18719 12540
rect 18719 12484 18723 12540
rect 18659 12480 18723 12484
rect 18739 12540 18803 12544
rect 18739 12484 18743 12540
rect 18743 12484 18799 12540
rect 18799 12484 18803 12540
rect 18739 12480 18803 12484
rect 18819 12540 18883 12544
rect 18819 12484 18823 12540
rect 18823 12484 18879 12540
rect 18879 12484 18883 12540
rect 18819 12480 18883 12484
rect 18899 12540 18963 12544
rect 18899 12484 18903 12540
rect 18903 12484 18959 12540
rect 18959 12484 18963 12540
rect 18899 12480 18963 12484
rect 25742 12540 25806 12544
rect 25742 12484 25746 12540
rect 25746 12484 25802 12540
rect 25802 12484 25806 12540
rect 25742 12480 25806 12484
rect 25822 12540 25886 12544
rect 25822 12484 25826 12540
rect 25826 12484 25882 12540
rect 25882 12484 25886 12540
rect 25822 12480 25886 12484
rect 25902 12540 25966 12544
rect 25902 12484 25906 12540
rect 25906 12484 25962 12540
rect 25962 12484 25966 12540
rect 25902 12480 25966 12484
rect 25982 12540 26046 12544
rect 25982 12484 25986 12540
rect 25986 12484 26042 12540
rect 26042 12484 26046 12540
rect 25982 12480 26046 12484
rect 5153 11996 5217 12000
rect 5153 11940 5157 11996
rect 5157 11940 5213 11996
rect 5213 11940 5217 11996
rect 5153 11936 5217 11940
rect 5233 11996 5297 12000
rect 5233 11940 5237 11996
rect 5237 11940 5293 11996
rect 5293 11940 5297 11996
rect 5233 11936 5297 11940
rect 5313 11996 5377 12000
rect 5313 11940 5317 11996
rect 5317 11940 5373 11996
rect 5373 11940 5377 11996
rect 5313 11936 5377 11940
rect 5393 11996 5457 12000
rect 5393 11940 5397 11996
rect 5397 11940 5453 11996
rect 5453 11940 5457 11996
rect 5393 11936 5457 11940
rect 12236 11996 12300 12000
rect 12236 11940 12240 11996
rect 12240 11940 12296 11996
rect 12296 11940 12300 11996
rect 12236 11936 12300 11940
rect 12316 11996 12380 12000
rect 12316 11940 12320 11996
rect 12320 11940 12376 11996
rect 12376 11940 12380 11996
rect 12316 11936 12380 11940
rect 12396 11996 12460 12000
rect 12396 11940 12400 11996
rect 12400 11940 12456 11996
rect 12456 11940 12460 11996
rect 12396 11936 12460 11940
rect 12476 11996 12540 12000
rect 12476 11940 12480 11996
rect 12480 11940 12536 11996
rect 12536 11940 12540 11996
rect 12476 11936 12540 11940
rect 19319 11996 19383 12000
rect 19319 11940 19323 11996
rect 19323 11940 19379 11996
rect 19379 11940 19383 11996
rect 19319 11936 19383 11940
rect 19399 11996 19463 12000
rect 19399 11940 19403 11996
rect 19403 11940 19459 11996
rect 19459 11940 19463 11996
rect 19399 11936 19463 11940
rect 19479 11996 19543 12000
rect 19479 11940 19483 11996
rect 19483 11940 19539 11996
rect 19539 11940 19543 11996
rect 19479 11936 19543 11940
rect 19559 11996 19623 12000
rect 19559 11940 19563 11996
rect 19563 11940 19619 11996
rect 19619 11940 19623 11996
rect 19559 11936 19623 11940
rect 26402 11996 26466 12000
rect 26402 11940 26406 11996
rect 26406 11940 26462 11996
rect 26462 11940 26466 11996
rect 26402 11936 26466 11940
rect 26482 11996 26546 12000
rect 26482 11940 26486 11996
rect 26486 11940 26542 11996
rect 26542 11940 26546 11996
rect 26482 11936 26546 11940
rect 26562 11996 26626 12000
rect 26562 11940 26566 11996
rect 26566 11940 26622 11996
rect 26622 11940 26626 11996
rect 26562 11936 26626 11940
rect 26642 11996 26706 12000
rect 26642 11940 26646 11996
rect 26646 11940 26702 11996
rect 26702 11940 26706 11996
rect 26642 11936 26706 11940
rect 27660 11732 27724 11796
rect 4493 11452 4557 11456
rect 4493 11396 4497 11452
rect 4497 11396 4553 11452
rect 4553 11396 4557 11452
rect 4493 11392 4557 11396
rect 4573 11452 4637 11456
rect 4573 11396 4577 11452
rect 4577 11396 4633 11452
rect 4633 11396 4637 11452
rect 4573 11392 4637 11396
rect 4653 11452 4717 11456
rect 4653 11396 4657 11452
rect 4657 11396 4713 11452
rect 4713 11396 4717 11452
rect 4653 11392 4717 11396
rect 4733 11452 4797 11456
rect 4733 11396 4737 11452
rect 4737 11396 4793 11452
rect 4793 11396 4797 11452
rect 4733 11392 4797 11396
rect 11576 11452 11640 11456
rect 11576 11396 11580 11452
rect 11580 11396 11636 11452
rect 11636 11396 11640 11452
rect 11576 11392 11640 11396
rect 11656 11452 11720 11456
rect 11656 11396 11660 11452
rect 11660 11396 11716 11452
rect 11716 11396 11720 11452
rect 11656 11392 11720 11396
rect 11736 11452 11800 11456
rect 11736 11396 11740 11452
rect 11740 11396 11796 11452
rect 11796 11396 11800 11452
rect 11736 11392 11800 11396
rect 11816 11452 11880 11456
rect 11816 11396 11820 11452
rect 11820 11396 11876 11452
rect 11876 11396 11880 11452
rect 11816 11392 11880 11396
rect 18659 11452 18723 11456
rect 18659 11396 18663 11452
rect 18663 11396 18719 11452
rect 18719 11396 18723 11452
rect 18659 11392 18723 11396
rect 18739 11452 18803 11456
rect 18739 11396 18743 11452
rect 18743 11396 18799 11452
rect 18799 11396 18803 11452
rect 18739 11392 18803 11396
rect 18819 11452 18883 11456
rect 18819 11396 18823 11452
rect 18823 11396 18879 11452
rect 18879 11396 18883 11452
rect 18819 11392 18883 11396
rect 18899 11452 18963 11456
rect 18899 11396 18903 11452
rect 18903 11396 18959 11452
rect 18959 11396 18963 11452
rect 18899 11392 18963 11396
rect 25742 11452 25806 11456
rect 25742 11396 25746 11452
rect 25746 11396 25802 11452
rect 25802 11396 25806 11452
rect 25742 11392 25806 11396
rect 25822 11452 25886 11456
rect 25822 11396 25826 11452
rect 25826 11396 25882 11452
rect 25882 11396 25886 11452
rect 25822 11392 25886 11396
rect 25902 11452 25966 11456
rect 25902 11396 25906 11452
rect 25906 11396 25962 11452
rect 25962 11396 25966 11452
rect 25902 11392 25966 11396
rect 25982 11452 26046 11456
rect 25982 11396 25986 11452
rect 25986 11396 26042 11452
rect 26042 11396 26046 11452
rect 25982 11392 26046 11396
rect 5153 10908 5217 10912
rect 5153 10852 5157 10908
rect 5157 10852 5213 10908
rect 5213 10852 5217 10908
rect 5153 10848 5217 10852
rect 5233 10908 5297 10912
rect 5233 10852 5237 10908
rect 5237 10852 5293 10908
rect 5293 10852 5297 10908
rect 5233 10848 5297 10852
rect 5313 10908 5377 10912
rect 5313 10852 5317 10908
rect 5317 10852 5373 10908
rect 5373 10852 5377 10908
rect 5313 10848 5377 10852
rect 5393 10908 5457 10912
rect 5393 10852 5397 10908
rect 5397 10852 5453 10908
rect 5453 10852 5457 10908
rect 5393 10848 5457 10852
rect 12236 10908 12300 10912
rect 12236 10852 12240 10908
rect 12240 10852 12296 10908
rect 12296 10852 12300 10908
rect 12236 10848 12300 10852
rect 12316 10908 12380 10912
rect 12316 10852 12320 10908
rect 12320 10852 12376 10908
rect 12376 10852 12380 10908
rect 12316 10848 12380 10852
rect 12396 10908 12460 10912
rect 12396 10852 12400 10908
rect 12400 10852 12456 10908
rect 12456 10852 12460 10908
rect 12396 10848 12460 10852
rect 12476 10908 12540 10912
rect 12476 10852 12480 10908
rect 12480 10852 12536 10908
rect 12536 10852 12540 10908
rect 12476 10848 12540 10852
rect 19319 10908 19383 10912
rect 19319 10852 19323 10908
rect 19323 10852 19379 10908
rect 19379 10852 19383 10908
rect 19319 10848 19383 10852
rect 19399 10908 19463 10912
rect 19399 10852 19403 10908
rect 19403 10852 19459 10908
rect 19459 10852 19463 10908
rect 19399 10848 19463 10852
rect 19479 10908 19543 10912
rect 19479 10852 19483 10908
rect 19483 10852 19539 10908
rect 19539 10852 19543 10908
rect 19479 10848 19543 10852
rect 19559 10908 19623 10912
rect 19559 10852 19563 10908
rect 19563 10852 19619 10908
rect 19619 10852 19623 10908
rect 19559 10848 19623 10852
rect 26402 10908 26466 10912
rect 26402 10852 26406 10908
rect 26406 10852 26462 10908
rect 26462 10852 26466 10908
rect 26402 10848 26466 10852
rect 26482 10908 26546 10912
rect 26482 10852 26486 10908
rect 26486 10852 26542 10908
rect 26542 10852 26546 10908
rect 26482 10848 26546 10852
rect 26562 10908 26626 10912
rect 26562 10852 26566 10908
rect 26566 10852 26622 10908
rect 26622 10852 26626 10908
rect 26562 10848 26626 10852
rect 26642 10908 26706 10912
rect 26642 10852 26646 10908
rect 26646 10852 26702 10908
rect 26702 10852 26706 10908
rect 26642 10848 26706 10852
rect 4493 10364 4557 10368
rect 4493 10308 4497 10364
rect 4497 10308 4553 10364
rect 4553 10308 4557 10364
rect 4493 10304 4557 10308
rect 4573 10364 4637 10368
rect 4573 10308 4577 10364
rect 4577 10308 4633 10364
rect 4633 10308 4637 10364
rect 4573 10304 4637 10308
rect 4653 10364 4717 10368
rect 4653 10308 4657 10364
rect 4657 10308 4713 10364
rect 4713 10308 4717 10364
rect 4653 10304 4717 10308
rect 4733 10364 4797 10368
rect 4733 10308 4737 10364
rect 4737 10308 4793 10364
rect 4793 10308 4797 10364
rect 4733 10304 4797 10308
rect 11576 10364 11640 10368
rect 11576 10308 11580 10364
rect 11580 10308 11636 10364
rect 11636 10308 11640 10364
rect 11576 10304 11640 10308
rect 11656 10364 11720 10368
rect 11656 10308 11660 10364
rect 11660 10308 11716 10364
rect 11716 10308 11720 10364
rect 11656 10304 11720 10308
rect 11736 10364 11800 10368
rect 11736 10308 11740 10364
rect 11740 10308 11796 10364
rect 11796 10308 11800 10364
rect 11736 10304 11800 10308
rect 11816 10364 11880 10368
rect 11816 10308 11820 10364
rect 11820 10308 11876 10364
rect 11876 10308 11880 10364
rect 11816 10304 11880 10308
rect 18659 10364 18723 10368
rect 18659 10308 18663 10364
rect 18663 10308 18719 10364
rect 18719 10308 18723 10364
rect 18659 10304 18723 10308
rect 18739 10364 18803 10368
rect 18739 10308 18743 10364
rect 18743 10308 18799 10364
rect 18799 10308 18803 10364
rect 18739 10304 18803 10308
rect 18819 10364 18883 10368
rect 18819 10308 18823 10364
rect 18823 10308 18879 10364
rect 18879 10308 18883 10364
rect 18819 10304 18883 10308
rect 18899 10364 18963 10368
rect 18899 10308 18903 10364
rect 18903 10308 18959 10364
rect 18959 10308 18963 10364
rect 18899 10304 18963 10308
rect 25742 10364 25806 10368
rect 25742 10308 25746 10364
rect 25746 10308 25802 10364
rect 25802 10308 25806 10364
rect 25742 10304 25806 10308
rect 25822 10364 25886 10368
rect 25822 10308 25826 10364
rect 25826 10308 25882 10364
rect 25882 10308 25886 10364
rect 25822 10304 25886 10308
rect 25902 10364 25966 10368
rect 25902 10308 25906 10364
rect 25906 10308 25962 10364
rect 25962 10308 25966 10364
rect 25902 10304 25966 10308
rect 25982 10364 26046 10368
rect 25982 10308 25986 10364
rect 25986 10308 26042 10364
rect 26042 10308 26046 10364
rect 25982 10304 26046 10308
rect 5153 9820 5217 9824
rect 5153 9764 5157 9820
rect 5157 9764 5213 9820
rect 5213 9764 5217 9820
rect 5153 9760 5217 9764
rect 5233 9820 5297 9824
rect 5233 9764 5237 9820
rect 5237 9764 5293 9820
rect 5293 9764 5297 9820
rect 5233 9760 5297 9764
rect 5313 9820 5377 9824
rect 5313 9764 5317 9820
rect 5317 9764 5373 9820
rect 5373 9764 5377 9820
rect 5313 9760 5377 9764
rect 5393 9820 5457 9824
rect 5393 9764 5397 9820
rect 5397 9764 5453 9820
rect 5453 9764 5457 9820
rect 5393 9760 5457 9764
rect 12236 9820 12300 9824
rect 12236 9764 12240 9820
rect 12240 9764 12296 9820
rect 12296 9764 12300 9820
rect 12236 9760 12300 9764
rect 12316 9820 12380 9824
rect 12316 9764 12320 9820
rect 12320 9764 12376 9820
rect 12376 9764 12380 9820
rect 12316 9760 12380 9764
rect 12396 9820 12460 9824
rect 12396 9764 12400 9820
rect 12400 9764 12456 9820
rect 12456 9764 12460 9820
rect 12396 9760 12460 9764
rect 12476 9820 12540 9824
rect 12476 9764 12480 9820
rect 12480 9764 12536 9820
rect 12536 9764 12540 9820
rect 12476 9760 12540 9764
rect 19319 9820 19383 9824
rect 19319 9764 19323 9820
rect 19323 9764 19379 9820
rect 19379 9764 19383 9820
rect 19319 9760 19383 9764
rect 19399 9820 19463 9824
rect 19399 9764 19403 9820
rect 19403 9764 19459 9820
rect 19459 9764 19463 9820
rect 19399 9760 19463 9764
rect 19479 9820 19543 9824
rect 19479 9764 19483 9820
rect 19483 9764 19539 9820
rect 19539 9764 19543 9820
rect 19479 9760 19543 9764
rect 19559 9820 19623 9824
rect 19559 9764 19563 9820
rect 19563 9764 19619 9820
rect 19619 9764 19623 9820
rect 19559 9760 19623 9764
rect 26402 9820 26466 9824
rect 26402 9764 26406 9820
rect 26406 9764 26462 9820
rect 26462 9764 26466 9820
rect 26402 9760 26466 9764
rect 26482 9820 26546 9824
rect 26482 9764 26486 9820
rect 26486 9764 26542 9820
rect 26542 9764 26546 9820
rect 26482 9760 26546 9764
rect 26562 9820 26626 9824
rect 26562 9764 26566 9820
rect 26566 9764 26622 9820
rect 26622 9764 26626 9820
rect 26562 9760 26626 9764
rect 26642 9820 26706 9824
rect 26642 9764 26646 9820
rect 26646 9764 26702 9820
rect 26702 9764 26706 9820
rect 26642 9760 26706 9764
rect 4493 9276 4557 9280
rect 4493 9220 4497 9276
rect 4497 9220 4553 9276
rect 4553 9220 4557 9276
rect 4493 9216 4557 9220
rect 4573 9276 4637 9280
rect 4573 9220 4577 9276
rect 4577 9220 4633 9276
rect 4633 9220 4637 9276
rect 4573 9216 4637 9220
rect 4653 9276 4717 9280
rect 4653 9220 4657 9276
rect 4657 9220 4713 9276
rect 4713 9220 4717 9276
rect 4653 9216 4717 9220
rect 4733 9276 4797 9280
rect 4733 9220 4737 9276
rect 4737 9220 4793 9276
rect 4793 9220 4797 9276
rect 4733 9216 4797 9220
rect 11576 9276 11640 9280
rect 11576 9220 11580 9276
rect 11580 9220 11636 9276
rect 11636 9220 11640 9276
rect 11576 9216 11640 9220
rect 11656 9276 11720 9280
rect 11656 9220 11660 9276
rect 11660 9220 11716 9276
rect 11716 9220 11720 9276
rect 11656 9216 11720 9220
rect 11736 9276 11800 9280
rect 11736 9220 11740 9276
rect 11740 9220 11796 9276
rect 11796 9220 11800 9276
rect 11736 9216 11800 9220
rect 11816 9276 11880 9280
rect 11816 9220 11820 9276
rect 11820 9220 11876 9276
rect 11876 9220 11880 9276
rect 11816 9216 11880 9220
rect 18659 9276 18723 9280
rect 18659 9220 18663 9276
rect 18663 9220 18719 9276
rect 18719 9220 18723 9276
rect 18659 9216 18723 9220
rect 18739 9276 18803 9280
rect 18739 9220 18743 9276
rect 18743 9220 18799 9276
rect 18799 9220 18803 9276
rect 18739 9216 18803 9220
rect 18819 9276 18883 9280
rect 18819 9220 18823 9276
rect 18823 9220 18879 9276
rect 18879 9220 18883 9276
rect 18819 9216 18883 9220
rect 18899 9276 18963 9280
rect 18899 9220 18903 9276
rect 18903 9220 18959 9276
rect 18959 9220 18963 9276
rect 18899 9216 18963 9220
rect 25742 9276 25806 9280
rect 25742 9220 25746 9276
rect 25746 9220 25802 9276
rect 25802 9220 25806 9276
rect 25742 9216 25806 9220
rect 25822 9276 25886 9280
rect 25822 9220 25826 9276
rect 25826 9220 25882 9276
rect 25882 9220 25886 9276
rect 25822 9216 25886 9220
rect 25902 9276 25966 9280
rect 25902 9220 25906 9276
rect 25906 9220 25962 9276
rect 25962 9220 25966 9276
rect 25902 9216 25966 9220
rect 25982 9276 26046 9280
rect 25982 9220 25986 9276
rect 25986 9220 26042 9276
rect 26042 9220 26046 9276
rect 25982 9216 26046 9220
rect 5153 8732 5217 8736
rect 5153 8676 5157 8732
rect 5157 8676 5213 8732
rect 5213 8676 5217 8732
rect 5153 8672 5217 8676
rect 5233 8732 5297 8736
rect 5233 8676 5237 8732
rect 5237 8676 5293 8732
rect 5293 8676 5297 8732
rect 5233 8672 5297 8676
rect 5313 8732 5377 8736
rect 5313 8676 5317 8732
rect 5317 8676 5373 8732
rect 5373 8676 5377 8732
rect 5313 8672 5377 8676
rect 5393 8732 5457 8736
rect 5393 8676 5397 8732
rect 5397 8676 5453 8732
rect 5453 8676 5457 8732
rect 5393 8672 5457 8676
rect 12236 8732 12300 8736
rect 12236 8676 12240 8732
rect 12240 8676 12296 8732
rect 12296 8676 12300 8732
rect 12236 8672 12300 8676
rect 12316 8732 12380 8736
rect 12316 8676 12320 8732
rect 12320 8676 12376 8732
rect 12376 8676 12380 8732
rect 12316 8672 12380 8676
rect 12396 8732 12460 8736
rect 12396 8676 12400 8732
rect 12400 8676 12456 8732
rect 12456 8676 12460 8732
rect 12396 8672 12460 8676
rect 12476 8732 12540 8736
rect 12476 8676 12480 8732
rect 12480 8676 12536 8732
rect 12536 8676 12540 8732
rect 12476 8672 12540 8676
rect 19319 8732 19383 8736
rect 19319 8676 19323 8732
rect 19323 8676 19379 8732
rect 19379 8676 19383 8732
rect 19319 8672 19383 8676
rect 19399 8732 19463 8736
rect 19399 8676 19403 8732
rect 19403 8676 19459 8732
rect 19459 8676 19463 8732
rect 19399 8672 19463 8676
rect 19479 8732 19543 8736
rect 19479 8676 19483 8732
rect 19483 8676 19539 8732
rect 19539 8676 19543 8732
rect 19479 8672 19543 8676
rect 19559 8732 19623 8736
rect 19559 8676 19563 8732
rect 19563 8676 19619 8732
rect 19619 8676 19623 8732
rect 19559 8672 19623 8676
rect 26402 8732 26466 8736
rect 26402 8676 26406 8732
rect 26406 8676 26462 8732
rect 26462 8676 26466 8732
rect 26402 8672 26466 8676
rect 26482 8732 26546 8736
rect 26482 8676 26486 8732
rect 26486 8676 26542 8732
rect 26542 8676 26546 8732
rect 26482 8672 26546 8676
rect 26562 8732 26626 8736
rect 26562 8676 26566 8732
rect 26566 8676 26622 8732
rect 26622 8676 26626 8732
rect 26562 8672 26626 8676
rect 26642 8732 26706 8736
rect 26642 8676 26646 8732
rect 26646 8676 26702 8732
rect 26702 8676 26706 8732
rect 26642 8672 26706 8676
rect 10548 8196 10612 8260
rect 4493 8188 4557 8192
rect 4493 8132 4497 8188
rect 4497 8132 4553 8188
rect 4553 8132 4557 8188
rect 4493 8128 4557 8132
rect 4573 8188 4637 8192
rect 4573 8132 4577 8188
rect 4577 8132 4633 8188
rect 4633 8132 4637 8188
rect 4573 8128 4637 8132
rect 4653 8188 4717 8192
rect 4653 8132 4657 8188
rect 4657 8132 4713 8188
rect 4713 8132 4717 8188
rect 4653 8128 4717 8132
rect 4733 8188 4797 8192
rect 4733 8132 4737 8188
rect 4737 8132 4793 8188
rect 4793 8132 4797 8188
rect 4733 8128 4797 8132
rect 11576 8188 11640 8192
rect 11576 8132 11580 8188
rect 11580 8132 11636 8188
rect 11636 8132 11640 8188
rect 11576 8128 11640 8132
rect 11656 8188 11720 8192
rect 11656 8132 11660 8188
rect 11660 8132 11716 8188
rect 11716 8132 11720 8188
rect 11656 8128 11720 8132
rect 11736 8188 11800 8192
rect 11736 8132 11740 8188
rect 11740 8132 11796 8188
rect 11796 8132 11800 8188
rect 11736 8128 11800 8132
rect 11816 8188 11880 8192
rect 11816 8132 11820 8188
rect 11820 8132 11876 8188
rect 11876 8132 11880 8188
rect 11816 8128 11880 8132
rect 18659 8188 18723 8192
rect 18659 8132 18663 8188
rect 18663 8132 18719 8188
rect 18719 8132 18723 8188
rect 18659 8128 18723 8132
rect 18739 8188 18803 8192
rect 18739 8132 18743 8188
rect 18743 8132 18799 8188
rect 18799 8132 18803 8188
rect 18739 8128 18803 8132
rect 18819 8188 18883 8192
rect 18819 8132 18823 8188
rect 18823 8132 18879 8188
rect 18879 8132 18883 8188
rect 18819 8128 18883 8132
rect 18899 8188 18963 8192
rect 18899 8132 18903 8188
rect 18903 8132 18959 8188
rect 18959 8132 18963 8188
rect 18899 8128 18963 8132
rect 25742 8188 25806 8192
rect 25742 8132 25746 8188
rect 25746 8132 25802 8188
rect 25802 8132 25806 8188
rect 25742 8128 25806 8132
rect 25822 8188 25886 8192
rect 25822 8132 25826 8188
rect 25826 8132 25882 8188
rect 25882 8132 25886 8188
rect 25822 8128 25886 8132
rect 25902 8188 25966 8192
rect 25902 8132 25906 8188
rect 25906 8132 25962 8188
rect 25962 8132 25966 8188
rect 25902 8128 25966 8132
rect 25982 8188 26046 8192
rect 25982 8132 25986 8188
rect 25986 8132 26042 8188
rect 26042 8132 26046 8188
rect 25982 8128 26046 8132
rect 10732 8060 10796 8124
rect 5153 7644 5217 7648
rect 5153 7588 5157 7644
rect 5157 7588 5213 7644
rect 5213 7588 5217 7644
rect 5153 7584 5217 7588
rect 5233 7644 5297 7648
rect 5233 7588 5237 7644
rect 5237 7588 5293 7644
rect 5293 7588 5297 7644
rect 5233 7584 5297 7588
rect 5313 7644 5377 7648
rect 5313 7588 5317 7644
rect 5317 7588 5373 7644
rect 5373 7588 5377 7644
rect 5313 7584 5377 7588
rect 5393 7644 5457 7648
rect 5393 7588 5397 7644
rect 5397 7588 5453 7644
rect 5453 7588 5457 7644
rect 5393 7584 5457 7588
rect 12236 7644 12300 7648
rect 12236 7588 12240 7644
rect 12240 7588 12296 7644
rect 12296 7588 12300 7644
rect 12236 7584 12300 7588
rect 12316 7644 12380 7648
rect 12316 7588 12320 7644
rect 12320 7588 12376 7644
rect 12376 7588 12380 7644
rect 12316 7584 12380 7588
rect 12396 7644 12460 7648
rect 12396 7588 12400 7644
rect 12400 7588 12456 7644
rect 12456 7588 12460 7644
rect 12396 7584 12460 7588
rect 12476 7644 12540 7648
rect 12476 7588 12480 7644
rect 12480 7588 12536 7644
rect 12536 7588 12540 7644
rect 12476 7584 12540 7588
rect 19319 7644 19383 7648
rect 19319 7588 19323 7644
rect 19323 7588 19379 7644
rect 19379 7588 19383 7644
rect 19319 7584 19383 7588
rect 19399 7644 19463 7648
rect 19399 7588 19403 7644
rect 19403 7588 19459 7644
rect 19459 7588 19463 7644
rect 19399 7584 19463 7588
rect 19479 7644 19543 7648
rect 19479 7588 19483 7644
rect 19483 7588 19539 7644
rect 19539 7588 19543 7644
rect 19479 7584 19543 7588
rect 19559 7644 19623 7648
rect 19559 7588 19563 7644
rect 19563 7588 19619 7644
rect 19619 7588 19623 7644
rect 19559 7584 19623 7588
rect 26402 7644 26466 7648
rect 26402 7588 26406 7644
rect 26406 7588 26462 7644
rect 26462 7588 26466 7644
rect 26402 7584 26466 7588
rect 26482 7644 26546 7648
rect 26482 7588 26486 7644
rect 26486 7588 26542 7644
rect 26542 7588 26546 7644
rect 26482 7584 26546 7588
rect 26562 7644 26626 7648
rect 26562 7588 26566 7644
rect 26566 7588 26622 7644
rect 26622 7588 26626 7644
rect 26562 7584 26626 7588
rect 26642 7644 26706 7648
rect 26642 7588 26646 7644
rect 26646 7588 26702 7644
rect 26702 7588 26706 7644
rect 26642 7584 26706 7588
rect 4493 7100 4557 7104
rect 4493 7044 4497 7100
rect 4497 7044 4553 7100
rect 4553 7044 4557 7100
rect 4493 7040 4557 7044
rect 4573 7100 4637 7104
rect 4573 7044 4577 7100
rect 4577 7044 4633 7100
rect 4633 7044 4637 7100
rect 4573 7040 4637 7044
rect 4653 7100 4717 7104
rect 4653 7044 4657 7100
rect 4657 7044 4713 7100
rect 4713 7044 4717 7100
rect 4653 7040 4717 7044
rect 4733 7100 4797 7104
rect 4733 7044 4737 7100
rect 4737 7044 4793 7100
rect 4793 7044 4797 7100
rect 4733 7040 4797 7044
rect 11576 7100 11640 7104
rect 11576 7044 11580 7100
rect 11580 7044 11636 7100
rect 11636 7044 11640 7100
rect 11576 7040 11640 7044
rect 11656 7100 11720 7104
rect 11656 7044 11660 7100
rect 11660 7044 11716 7100
rect 11716 7044 11720 7100
rect 11656 7040 11720 7044
rect 11736 7100 11800 7104
rect 11736 7044 11740 7100
rect 11740 7044 11796 7100
rect 11796 7044 11800 7100
rect 11736 7040 11800 7044
rect 11816 7100 11880 7104
rect 11816 7044 11820 7100
rect 11820 7044 11876 7100
rect 11876 7044 11880 7100
rect 11816 7040 11880 7044
rect 18659 7100 18723 7104
rect 18659 7044 18663 7100
rect 18663 7044 18719 7100
rect 18719 7044 18723 7100
rect 18659 7040 18723 7044
rect 18739 7100 18803 7104
rect 18739 7044 18743 7100
rect 18743 7044 18799 7100
rect 18799 7044 18803 7100
rect 18739 7040 18803 7044
rect 18819 7100 18883 7104
rect 18819 7044 18823 7100
rect 18823 7044 18879 7100
rect 18879 7044 18883 7100
rect 18819 7040 18883 7044
rect 18899 7100 18963 7104
rect 18899 7044 18903 7100
rect 18903 7044 18959 7100
rect 18959 7044 18963 7100
rect 18899 7040 18963 7044
rect 25742 7100 25806 7104
rect 25742 7044 25746 7100
rect 25746 7044 25802 7100
rect 25802 7044 25806 7100
rect 25742 7040 25806 7044
rect 25822 7100 25886 7104
rect 25822 7044 25826 7100
rect 25826 7044 25882 7100
rect 25882 7044 25886 7100
rect 25822 7040 25886 7044
rect 25902 7100 25966 7104
rect 25902 7044 25906 7100
rect 25906 7044 25962 7100
rect 25962 7044 25966 7100
rect 25902 7040 25966 7044
rect 25982 7100 26046 7104
rect 25982 7044 25986 7100
rect 25986 7044 26042 7100
rect 26042 7044 26046 7100
rect 25982 7040 26046 7044
rect 28764 6700 28828 6764
rect 5153 6556 5217 6560
rect 5153 6500 5157 6556
rect 5157 6500 5213 6556
rect 5213 6500 5217 6556
rect 5153 6496 5217 6500
rect 5233 6556 5297 6560
rect 5233 6500 5237 6556
rect 5237 6500 5293 6556
rect 5293 6500 5297 6556
rect 5233 6496 5297 6500
rect 5313 6556 5377 6560
rect 5313 6500 5317 6556
rect 5317 6500 5373 6556
rect 5373 6500 5377 6556
rect 5313 6496 5377 6500
rect 5393 6556 5457 6560
rect 5393 6500 5397 6556
rect 5397 6500 5453 6556
rect 5453 6500 5457 6556
rect 5393 6496 5457 6500
rect 12236 6556 12300 6560
rect 12236 6500 12240 6556
rect 12240 6500 12296 6556
rect 12296 6500 12300 6556
rect 12236 6496 12300 6500
rect 12316 6556 12380 6560
rect 12316 6500 12320 6556
rect 12320 6500 12376 6556
rect 12376 6500 12380 6556
rect 12316 6496 12380 6500
rect 12396 6556 12460 6560
rect 12396 6500 12400 6556
rect 12400 6500 12456 6556
rect 12456 6500 12460 6556
rect 12396 6496 12460 6500
rect 12476 6556 12540 6560
rect 12476 6500 12480 6556
rect 12480 6500 12536 6556
rect 12536 6500 12540 6556
rect 12476 6496 12540 6500
rect 19319 6556 19383 6560
rect 19319 6500 19323 6556
rect 19323 6500 19379 6556
rect 19379 6500 19383 6556
rect 19319 6496 19383 6500
rect 19399 6556 19463 6560
rect 19399 6500 19403 6556
rect 19403 6500 19459 6556
rect 19459 6500 19463 6556
rect 19399 6496 19463 6500
rect 19479 6556 19543 6560
rect 19479 6500 19483 6556
rect 19483 6500 19539 6556
rect 19539 6500 19543 6556
rect 19479 6496 19543 6500
rect 19559 6556 19623 6560
rect 19559 6500 19563 6556
rect 19563 6500 19619 6556
rect 19619 6500 19623 6556
rect 19559 6496 19623 6500
rect 26402 6556 26466 6560
rect 26402 6500 26406 6556
rect 26406 6500 26462 6556
rect 26462 6500 26466 6556
rect 26402 6496 26466 6500
rect 26482 6556 26546 6560
rect 26482 6500 26486 6556
rect 26486 6500 26542 6556
rect 26542 6500 26546 6556
rect 26482 6496 26546 6500
rect 26562 6556 26626 6560
rect 26562 6500 26566 6556
rect 26566 6500 26622 6556
rect 26622 6500 26626 6556
rect 26562 6496 26626 6500
rect 26642 6556 26706 6560
rect 26642 6500 26646 6556
rect 26646 6500 26702 6556
rect 26702 6500 26706 6556
rect 26642 6496 26706 6500
rect 4493 6012 4557 6016
rect 4493 5956 4497 6012
rect 4497 5956 4553 6012
rect 4553 5956 4557 6012
rect 4493 5952 4557 5956
rect 4573 6012 4637 6016
rect 4573 5956 4577 6012
rect 4577 5956 4633 6012
rect 4633 5956 4637 6012
rect 4573 5952 4637 5956
rect 4653 6012 4717 6016
rect 4653 5956 4657 6012
rect 4657 5956 4713 6012
rect 4713 5956 4717 6012
rect 4653 5952 4717 5956
rect 4733 6012 4797 6016
rect 4733 5956 4737 6012
rect 4737 5956 4793 6012
rect 4793 5956 4797 6012
rect 4733 5952 4797 5956
rect 11576 6012 11640 6016
rect 11576 5956 11580 6012
rect 11580 5956 11636 6012
rect 11636 5956 11640 6012
rect 11576 5952 11640 5956
rect 11656 6012 11720 6016
rect 11656 5956 11660 6012
rect 11660 5956 11716 6012
rect 11716 5956 11720 6012
rect 11656 5952 11720 5956
rect 11736 6012 11800 6016
rect 11736 5956 11740 6012
rect 11740 5956 11796 6012
rect 11796 5956 11800 6012
rect 11736 5952 11800 5956
rect 11816 6012 11880 6016
rect 11816 5956 11820 6012
rect 11820 5956 11876 6012
rect 11876 5956 11880 6012
rect 11816 5952 11880 5956
rect 18659 6012 18723 6016
rect 18659 5956 18663 6012
rect 18663 5956 18719 6012
rect 18719 5956 18723 6012
rect 18659 5952 18723 5956
rect 18739 6012 18803 6016
rect 18739 5956 18743 6012
rect 18743 5956 18799 6012
rect 18799 5956 18803 6012
rect 18739 5952 18803 5956
rect 18819 6012 18883 6016
rect 18819 5956 18823 6012
rect 18823 5956 18879 6012
rect 18879 5956 18883 6012
rect 18819 5952 18883 5956
rect 18899 6012 18963 6016
rect 18899 5956 18903 6012
rect 18903 5956 18959 6012
rect 18959 5956 18963 6012
rect 18899 5952 18963 5956
rect 25742 6012 25806 6016
rect 25742 5956 25746 6012
rect 25746 5956 25802 6012
rect 25802 5956 25806 6012
rect 25742 5952 25806 5956
rect 25822 6012 25886 6016
rect 25822 5956 25826 6012
rect 25826 5956 25882 6012
rect 25882 5956 25886 6012
rect 25822 5952 25886 5956
rect 25902 6012 25966 6016
rect 25902 5956 25906 6012
rect 25906 5956 25962 6012
rect 25962 5956 25966 6012
rect 25902 5952 25966 5956
rect 25982 6012 26046 6016
rect 25982 5956 25986 6012
rect 25986 5956 26042 6012
rect 26042 5956 26046 6012
rect 25982 5952 26046 5956
rect 24348 5536 24412 5540
rect 24348 5480 24362 5536
rect 24362 5480 24412 5536
rect 24348 5476 24412 5480
rect 5153 5468 5217 5472
rect 5153 5412 5157 5468
rect 5157 5412 5213 5468
rect 5213 5412 5217 5468
rect 5153 5408 5217 5412
rect 5233 5468 5297 5472
rect 5233 5412 5237 5468
rect 5237 5412 5293 5468
rect 5293 5412 5297 5468
rect 5233 5408 5297 5412
rect 5313 5468 5377 5472
rect 5313 5412 5317 5468
rect 5317 5412 5373 5468
rect 5373 5412 5377 5468
rect 5313 5408 5377 5412
rect 5393 5468 5457 5472
rect 5393 5412 5397 5468
rect 5397 5412 5453 5468
rect 5453 5412 5457 5468
rect 5393 5408 5457 5412
rect 12236 5468 12300 5472
rect 12236 5412 12240 5468
rect 12240 5412 12296 5468
rect 12296 5412 12300 5468
rect 12236 5408 12300 5412
rect 12316 5468 12380 5472
rect 12316 5412 12320 5468
rect 12320 5412 12376 5468
rect 12376 5412 12380 5468
rect 12316 5408 12380 5412
rect 12396 5468 12460 5472
rect 12396 5412 12400 5468
rect 12400 5412 12456 5468
rect 12456 5412 12460 5468
rect 12396 5408 12460 5412
rect 12476 5468 12540 5472
rect 12476 5412 12480 5468
rect 12480 5412 12536 5468
rect 12536 5412 12540 5468
rect 12476 5408 12540 5412
rect 19319 5468 19383 5472
rect 19319 5412 19323 5468
rect 19323 5412 19379 5468
rect 19379 5412 19383 5468
rect 19319 5408 19383 5412
rect 19399 5468 19463 5472
rect 19399 5412 19403 5468
rect 19403 5412 19459 5468
rect 19459 5412 19463 5468
rect 19399 5408 19463 5412
rect 19479 5468 19543 5472
rect 19479 5412 19483 5468
rect 19483 5412 19539 5468
rect 19539 5412 19543 5468
rect 19479 5408 19543 5412
rect 19559 5468 19623 5472
rect 19559 5412 19563 5468
rect 19563 5412 19619 5468
rect 19619 5412 19623 5468
rect 19559 5408 19623 5412
rect 26402 5468 26466 5472
rect 26402 5412 26406 5468
rect 26406 5412 26462 5468
rect 26462 5412 26466 5468
rect 26402 5408 26466 5412
rect 26482 5468 26546 5472
rect 26482 5412 26486 5468
rect 26486 5412 26542 5468
rect 26542 5412 26546 5468
rect 26482 5408 26546 5412
rect 26562 5468 26626 5472
rect 26562 5412 26566 5468
rect 26566 5412 26622 5468
rect 26622 5412 26626 5468
rect 26562 5408 26626 5412
rect 26642 5468 26706 5472
rect 26642 5412 26646 5468
rect 26646 5412 26702 5468
rect 26702 5412 26706 5468
rect 26642 5408 26706 5412
rect 4493 4924 4557 4928
rect 4493 4868 4497 4924
rect 4497 4868 4553 4924
rect 4553 4868 4557 4924
rect 4493 4864 4557 4868
rect 4573 4924 4637 4928
rect 4573 4868 4577 4924
rect 4577 4868 4633 4924
rect 4633 4868 4637 4924
rect 4573 4864 4637 4868
rect 4653 4924 4717 4928
rect 4653 4868 4657 4924
rect 4657 4868 4713 4924
rect 4713 4868 4717 4924
rect 4653 4864 4717 4868
rect 4733 4924 4797 4928
rect 4733 4868 4737 4924
rect 4737 4868 4793 4924
rect 4793 4868 4797 4924
rect 4733 4864 4797 4868
rect 11576 4924 11640 4928
rect 11576 4868 11580 4924
rect 11580 4868 11636 4924
rect 11636 4868 11640 4924
rect 11576 4864 11640 4868
rect 11656 4924 11720 4928
rect 11656 4868 11660 4924
rect 11660 4868 11716 4924
rect 11716 4868 11720 4924
rect 11656 4864 11720 4868
rect 11736 4924 11800 4928
rect 11736 4868 11740 4924
rect 11740 4868 11796 4924
rect 11796 4868 11800 4924
rect 11736 4864 11800 4868
rect 11816 4924 11880 4928
rect 11816 4868 11820 4924
rect 11820 4868 11876 4924
rect 11876 4868 11880 4924
rect 11816 4864 11880 4868
rect 18659 4924 18723 4928
rect 18659 4868 18663 4924
rect 18663 4868 18719 4924
rect 18719 4868 18723 4924
rect 18659 4864 18723 4868
rect 18739 4924 18803 4928
rect 18739 4868 18743 4924
rect 18743 4868 18799 4924
rect 18799 4868 18803 4924
rect 18739 4864 18803 4868
rect 18819 4924 18883 4928
rect 18819 4868 18823 4924
rect 18823 4868 18879 4924
rect 18879 4868 18883 4924
rect 18819 4864 18883 4868
rect 18899 4924 18963 4928
rect 18899 4868 18903 4924
rect 18903 4868 18959 4924
rect 18959 4868 18963 4924
rect 18899 4864 18963 4868
rect 25742 4924 25806 4928
rect 25742 4868 25746 4924
rect 25746 4868 25802 4924
rect 25802 4868 25806 4924
rect 25742 4864 25806 4868
rect 25822 4924 25886 4928
rect 25822 4868 25826 4924
rect 25826 4868 25882 4924
rect 25882 4868 25886 4924
rect 25822 4864 25886 4868
rect 25902 4924 25966 4928
rect 25902 4868 25906 4924
rect 25906 4868 25962 4924
rect 25962 4868 25966 4924
rect 25902 4864 25966 4868
rect 25982 4924 26046 4928
rect 25982 4868 25986 4924
rect 25986 4868 26042 4924
rect 26042 4868 26046 4924
rect 25982 4864 26046 4868
rect 5153 4380 5217 4384
rect 5153 4324 5157 4380
rect 5157 4324 5213 4380
rect 5213 4324 5217 4380
rect 5153 4320 5217 4324
rect 5233 4380 5297 4384
rect 5233 4324 5237 4380
rect 5237 4324 5293 4380
rect 5293 4324 5297 4380
rect 5233 4320 5297 4324
rect 5313 4380 5377 4384
rect 5313 4324 5317 4380
rect 5317 4324 5373 4380
rect 5373 4324 5377 4380
rect 5313 4320 5377 4324
rect 5393 4380 5457 4384
rect 5393 4324 5397 4380
rect 5397 4324 5453 4380
rect 5453 4324 5457 4380
rect 5393 4320 5457 4324
rect 12236 4380 12300 4384
rect 12236 4324 12240 4380
rect 12240 4324 12296 4380
rect 12296 4324 12300 4380
rect 12236 4320 12300 4324
rect 12316 4380 12380 4384
rect 12316 4324 12320 4380
rect 12320 4324 12376 4380
rect 12376 4324 12380 4380
rect 12316 4320 12380 4324
rect 12396 4380 12460 4384
rect 12396 4324 12400 4380
rect 12400 4324 12456 4380
rect 12456 4324 12460 4380
rect 12396 4320 12460 4324
rect 12476 4380 12540 4384
rect 12476 4324 12480 4380
rect 12480 4324 12536 4380
rect 12536 4324 12540 4380
rect 12476 4320 12540 4324
rect 19319 4380 19383 4384
rect 19319 4324 19323 4380
rect 19323 4324 19379 4380
rect 19379 4324 19383 4380
rect 19319 4320 19383 4324
rect 19399 4380 19463 4384
rect 19399 4324 19403 4380
rect 19403 4324 19459 4380
rect 19459 4324 19463 4380
rect 19399 4320 19463 4324
rect 19479 4380 19543 4384
rect 19479 4324 19483 4380
rect 19483 4324 19539 4380
rect 19539 4324 19543 4380
rect 19479 4320 19543 4324
rect 19559 4380 19623 4384
rect 19559 4324 19563 4380
rect 19563 4324 19619 4380
rect 19619 4324 19623 4380
rect 19559 4320 19623 4324
rect 26402 4380 26466 4384
rect 26402 4324 26406 4380
rect 26406 4324 26462 4380
rect 26462 4324 26466 4380
rect 26402 4320 26466 4324
rect 26482 4380 26546 4384
rect 26482 4324 26486 4380
rect 26486 4324 26542 4380
rect 26542 4324 26546 4380
rect 26482 4320 26546 4324
rect 26562 4380 26626 4384
rect 26562 4324 26566 4380
rect 26566 4324 26622 4380
rect 26622 4324 26626 4380
rect 26562 4320 26626 4324
rect 26642 4380 26706 4384
rect 26642 4324 26646 4380
rect 26646 4324 26702 4380
rect 26702 4324 26706 4380
rect 26642 4320 26706 4324
rect 4493 3836 4557 3840
rect 4493 3780 4497 3836
rect 4497 3780 4553 3836
rect 4553 3780 4557 3836
rect 4493 3776 4557 3780
rect 4573 3836 4637 3840
rect 4573 3780 4577 3836
rect 4577 3780 4633 3836
rect 4633 3780 4637 3836
rect 4573 3776 4637 3780
rect 4653 3836 4717 3840
rect 4653 3780 4657 3836
rect 4657 3780 4713 3836
rect 4713 3780 4717 3836
rect 4653 3776 4717 3780
rect 4733 3836 4797 3840
rect 4733 3780 4737 3836
rect 4737 3780 4793 3836
rect 4793 3780 4797 3836
rect 4733 3776 4797 3780
rect 11576 3836 11640 3840
rect 11576 3780 11580 3836
rect 11580 3780 11636 3836
rect 11636 3780 11640 3836
rect 11576 3776 11640 3780
rect 11656 3836 11720 3840
rect 11656 3780 11660 3836
rect 11660 3780 11716 3836
rect 11716 3780 11720 3836
rect 11656 3776 11720 3780
rect 11736 3836 11800 3840
rect 11736 3780 11740 3836
rect 11740 3780 11796 3836
rect 11796 3780 11800 3836
rect 11736 3776 11800 3780
rect 11816 3836 11880 3840
rect 11816 3780 11820 3836
rect 11820 3780 11876 3836
rect 11876 3780 11880 3836
rect 11816 3776 11880 3780
rect 18659 3836 18723 3840
rect 18659 3780 18663 3836
rect 18663 3780 18719 3836
rect 18719 3780 18723 3836
rect 18659 3776 18723 3780
rect 18739 3836 18803 3840
rect 18739 3780 18743 3836
rect 18743 3780 18799 3836
rect 18799 3780 18803 3836
rect 18739 3776 18803 3780
rect 18819 3836 18883 3840
rect 18819 3780 18823 3836
rect 18823 3780 18879 3836
rect 18879 3780 18883 3836
rect 18819 3776 18883 3780
rect 18899 3836 18963 3840
rect 18899 3780 18903 3836
rect 18903 3780 18959 3836
rect 18959 3780 18963 3836
rect 18899 3776 18963 3780
rect 25742 3836 25806 3840
rect 25742 3780 25746 3836
rect 25746 3780 25802 3836
rect 25802 3780 25806 3836
rect 25742 3776 25806 3780
rect 25822 3836 25886 3840
rect 25822 3780 25826 3836
rect 25826 3780 25882 3836
rect 25882 3780 25886 3836
rect 25822 3776 25886 3780
rect 25902 3836 25966 3840
rect 25902 3780 25906 3836
rect 25906 3780 25962 3836
rect 25962 3780 25966 3836
rect 25902 3776 25966 3780
rect 25982 3836 26046 3840
rect 25982 3780 25986 3836
rect 25986 3780 26042 3836
rect 26042 3780 26046 3836
rect 25982 3776 26046 3780
rect 5153 3292 5217 3296
rect 5153 3236 5157 3292
rect 5157 3236 5213 3292
rect 5213 3236 5217 3292
rect 5153 3232 5217 3236
rect 5233 3292 5297 3296
rect 5233 3236 5237 3292
rect 5237 3236 5293 3292
rect 5293 3236 5297 3292
rect 5233 3232 5297 3236
rect 5313 3292 5377 3296
rect 5313 3236 5317 3292
rect 5317 3236 5373 3292
rect 5373 3236 5377 3292
rect 5313 3232 5377 3236
rect 5393 3292 5457 3296
rect 5393 3236 5397 3292
rect 5397 3236 5453 3292
rect 5453 3236 5457 3292
rect 5393 3232 5457 3236
rect 12236 3292 12300 3296
rect 12236 3236 12240 3292
rect 12240 3236 12296 3292
rect 12296 3236 12300 3292
rect 12236 3232 12300 3236
rect 12316 3292 12380 3296
rect 12316 3236 12320 3292
rect 12320 3236 12376 3292
rect 12376 3236 12380 3292
rect 12316 3232 12380 3236
rect 12396 3292 12460 3296
rect 12396 3236 12400 3292
rect 12400 3236 12456 3292
rect 12456 3236 12460 3292
rect 12396 3232 12460 3236
rect 12476 3292 12540 3296
rect 12476 3236 12480 3292
rect 12480 3236 12536 3292
rect 12536 3236 12540 3292
rect 12476 3232 12540 3236
rect 19319 3292 19383 3296
rect 19319 3236 19323 3292
rect 19323 3236 19379 3292
rect 19379 3236 19383 3292
rect 19319 3232 19383 3236
rect 19399 3292 19463 3296
rect 19399 3236 19403 3292
rect 19403 3236 19459 3292
rect 19459 3236 19463 3292
rect 19399 3232 19463 3236
rect 19479 3292 19543 3296
rect 19479 3236 19483 3292
rect 19483 3236 19539 3292
rect 19539 3236 19543 3292
rect 19479 3232 19543 3236
rect 19559 3292 19623 3296
rect 19559 3236 19563 3292
rect 19563 3236 19619 3292
rect 19619 3236 19623 3292
rect 19559 3232 19623 3236
rect 26402 3292 26466 3296
rect 26402 3236 26406 3292
rect 26406 3236 26462 3292
rect 26462 3236 26466 3292
rect 26402 3232 26466 3236
rect 26482 3292 26546 3296
rect 26482 3236 26486 3292
rect 26486 3236 26542 3292
rect 26542 3236 26546 3292
rect 26482 3232 26546 3236
rect 26562 3292 26626 3296
rect 26562 3236 26566 3292
rect 26566 3236 26622 3292
rect 26622 3236 26626 3292
rect 26562 3232 26626 3236
rect 26642 3292 26706 3296
rect 26642 3236 26646 3292
rect 26646 3236 26702 3292
rect 26702 3236 26706 3292
rect 26642 3232 26706 3236
rect 4493 2748 4557 2752
rect 4493 2692 4497 2748
rect 4497 2692 4553 2748
rect 4553 2692 4557 2748
rect 4493 2688 4557 2692
rect 4573 2748 4637 2752
rect 4573 2692 4577 2748
rect 4577 2692 4633 2748
rect 4633 2692 4637 2748
rect 4573 2688 4637 2692
rect 4653 2748 4717 2752
rect 4653 2692 4657 2748
rect 4657 2692 4713 2748
rect 4713 2692 4717 2748
rect 4653 2688 4717 2692
rect 4733 2748 4797 2752
rect 4733 2692 4737 2748
rect 4737 2692 4793 2748
rect 4793 2692 4797 2748
rect 4733 2688 4797 2692
rect 11576 2748 11640 2752
rect 11576 2692 11580 2748
rect 11580 2692 11636 2748
rect 11636 2692 11640 2748
rect 11576 2688 11640 2692
rect 11656 2748 11720 2752
rect 11656 2692 11660 2748
rect 11660 2692 11716 2748
rect 11716 2692 11720 2748
rect 11656 2688 11720 2692
rect 11736 2748 11800 2752
rect 11736 2692 11740 2748
rect 11740 2692 11796 2748
rect 11796 2692 11800 2748
rect 11736 2688 11800 2692
rect 11816 2748 11880 2752
rect 11816 2692 11820 2748
rect 11820 2692 11876 2748
rect 11876 2692 11880 2748
rect 11816 2688 11880 2692
rect 18659 2748 18723 2752
rect 18659 2692 18663 2748
rect 18663 2692 18719 2748
rect 18719 2692 18723 2748
rect 18659 2688 18723 2692
rect 18739 2748 18803 2752
rect 18739 2692 18743 2748
rect 18743 2692 18799 2748
rect 18799 2692 18803 2748
rect 18739 2688 18803 2692
rect 18819 2748 18883 2752
rect 18819 2692 18823 2748
rect 18823 2692 18879 2748
rect 18879 2692 18883 2748
rect 18819 2688 18883 2692
rect 18899 2748 18963 2752
rect 18899 2692 18903 2748
rect 18903 2692 18959 2748
rect 18959 2692 18963 2748
rect 18899 2688 18963 2692
rect 25742 2748 25806 2752
rect 25742 2692 25746 2748
rect 25746 2692 25802 2748
rect 25802 2692 25806 2748
rect 25742 2688 25806 2692
rect 25822 2748 25886 2752
rect 25822 2692 25826 2748
rect 25826 2692 25882 2748
rect 25882 2692 25886 2748
rect 25822 2688 25886 2692
rect 25902 2748 25966 2752
rect 25902 2692 25906 2748
rect 25906 2692 25962 2748
rect 25962 2692 25966 2748
rect 25902 2688 25966 2692
rect 25982 2748 26046 2752
rect 25982 2692 25986 2748
rect 25986 2692 26042 2748
rect 26042 2692 26046 2748
rect 25982 2688 26046 2692
rect 5153 2204 5217 2208
rect 5153 2148 5157 2204
rect 5157 2148 5213 2204
rect 5213 2148 5217 2204
rect 5153 2144 5217 2148
rect 5233 2204 5297 2208
rect 5233 2148 5237 2204
rect 5237 2148 5293 2204
rect 5293 2148 5297 2204
rect 5233 2144 5297 2148
rect 5313 2204 5377 2208
rect 5313 2148 5317 2204
rect 5317 2148 5373 2204
rect 5373 2148 5377 2204
rect 5313 2144 5377 2148
rect 5393 2204 5457 2208
rect 5393 2148 5397 2204
rect 5397 2148 5453 2204
rect 5453 2148 5457 2204
rect 5393 2144 5457 2148
rect 12236 2204 12300 2208
rect 12236 2148 12240 2204
rect 12240 2148 12296 2204
rect 12296 2148 12300 2204
rect 12236 2144 12300 2148
rect 12316 2204 12380 2208
rect 12316 2148 12320 2204
rect 12320 2148 12376 2204
rect 12376 2148 12380 2204
rect 12316 2144 12380 2148
rect 12396 2204 12460 2208
rect 12396 2148 12400 2204
rect 12400 2148 12456 2204
rect 12456 2148 12460 2204
rect 12396 2144 12460 2148
rect 12476 2204 12540 2208
rect 12476 2148 12480 2204
rect 12480 2148 12536 2204
rect 12536 2148 12540 2204
rect 12476 2144 12540 2148
rect 19319 2204 19383 2208
rect 19319 2148 19323 2204
rect 19323 2148 19379 2204
rect 19379 2148 19383 2204
rect 19319 2144 19383 2148
rect 19399 2204 19463 2208
rect 19399 2148 19403 2204
rect 19403 2148 19459 2204
rect 19459 2148 19463 2204
rect 19399 2144 19463 2148
rect 19479 2204 19543 2208
rect 19479 2148 19483 2204
rect 19483 2148 19539 2204
rect 19539 2148 19543 2204
rect 19479 2144 19543 2148
rect 19559 2204 19623 2208
rect 19559 2148 19563 2204
rect 19563 2148 19619 2204
rect 19619 2148 19623 2204
rect 19559 2144 19623 2148
rect 26402 2204 26466 2208
rect 26402 2148 26406 2204
rect 26406 2148 26462 2204
rect 26462 2148 26466 2204
rect 26402 2144 26466 2148
rect 26482 2204 26546 2208
rect 26482 2148 26486 2204
rect 26486 2148 26542 2204
rect 26542 2148 26546 2204
rect 26482 2144 26546 2148
rect 26562 2204 26626 2208
rect 26562 2148 26566 2204
rect 26566 2148 26622 2204
rect 26622 2148 26626 2204
rect 26562 2144 26626 2148
rect 26642 2204 26706 2208
rect 26642 2148 26646 2204
rect 26646 2148 26702 2204
rect 26702 2148 26706 2204
rect 26642 2144 26706 2148
<< metal4 >>
rect 4485 29952 4805 30512
rect 4485 29888 4493 29952
rect 4557 29888 4573 29952
rect 4637 29888 4653 29952
rect 4717 29888 4733 29952
rect 4797 29888 4805 29952
rect 4485 28864 4805 29888
rect 4485 28800 4493 28864
rect 4557 28800 4573 28864
rect 4637 28800 4653 28864
rect 4717 28800 4733 28864
rect 4797 28800 4805 28864
rect 4485 27776 4805 28800
rect 4485 27712 4493 27776
rect 4557 27712 4573 27776
rect 4637 27712 4653 27776
rect 4717 27712 4733 27776
rect 4797 27712 4805 27776
rect 4485 27046 4805 27712
rect 4485 26810 4527 27046
rect 4763 26810 4805 27046
rect 4485 26688 4805 26810
rect 4485 26624 4493 26688
rect 4557 26624 4573 26688
rect 4637 26624 4653 26688
rect 4717 26624 4733 26688
rect 4797 26624 4805 26688
rect 4485 25600 4805 26624
rect 4485 25536 4493 25600
rect 4557 25536 4573 25600
rect 4637 25536 4653 25600
rect 4717 25536 4733 25600
rect 4797 25536 4805 25600
rect 4485 24512 4805 25536
rect 4485 24448 4493 24512
rect 4557 24448 4573 24512
rect 4637 24448 4653 24512
rect 4717 24448 4733 24512
rect 4797 24448 4805 24512
rect 4485 23424 4805 24448
rect 4485 23360 4493 23424
rect 4557 23360 4573 23424
rect 4637 23360 4653 23424
rect 4717 23360 4733 23424
rect 4797 23360 4805 23424
rect 4485 22336 4805 23360
rect 4485 22272 4493 22336
rect 4557 22272 4573 22336
rect 4637 22272 4653 22336
rect 4717 22272 4733 22336
rect 4797 22272 4805 22336
rect 4485 21248 4805 22272
rect 4485 21184 4493 21248
rect 4557 21184 4573 21248
rect 4637 21184 4653 21248
rect 4717 21184 4733 21248
rect 4797 21184 4805 21248
rect 4485 20160 4805 21184
rect 4485 20096 4493 20160
rect 4557 20096 4573 20160
rect 4637 20096 4653 20160
rect 4717 20096 4733 20160
rect 4797 20096 4805 20160
rect 4485 19974 4805 20096
rect 4485 19738 4527 19974
rect 4763 19738 4805 19974
rect 4485 19072 4805 19738
rect 4485 19008 4493 19072
rect 4557 19008 4573 19072
rect 4637 19008 4653 19072
rect 4717 19008 4733 19072
rect 4797 19008 4805 19072
rect 4485 17984 4805 19008
rect 4485 17920 4493 17984
rect 4557 17920 4573 17984
rect 4637 17920 4653 17984
rect 4717 17920 4733 17984
rect 4797 17920 4805 17984
rect 4485 16896 4805 17920
rect 4485 16832 4493 16896
rect 4557 16832 4573 16896
rect 4637 16832 4653 16896
rect 4717 16832 4733 16896
rect 4797 16832 4805 16896
rect 4485 15808 4805 16832
rect 4485 15744 4493 15808
rect 4557 15744 4573 15808
rect 4637 15744 4653 15808
rect 4717 15744 4733 15808
rect 4797 15744 4805 15808
rect 4485 14720 4805 15744
rect 4485 14656 4493 14720
rect 4557 14656 4573 14720
rect 4637 14656 4653 14720
rect 4717 14656 4733 14720
rect 4797 14656 4805 14720
rect 4485 13632 4805 14656
rect 4485 13568 4493 13632
rect 4557 13568 4573 13632
rect 4637 13568 4653 13632
rect 4717 13568 4733 13632
rect 4797 13568 4805 13632
rect 4485 12902 4805 13568
rect 4485 12666 4527 12902
rect 4763 12666 4805 12902
rect 4485 12544 4805 12666
rect 4485 12480 4493 12544
rect 4557 12480 4573 12544
rect 4637 12480 4653 12544
rect 4717 12480 4733 12544
rect 4797 12480 4805 12544
rect 4485 11456 4805 12480
rect 4485 11392 4493 11456
rect 4557 11392 4573 11456
rect 4637 11392 4653 11456
rect 4717 11392 4733 11456
rect 4797 11392 4805 11456
rect 4485 10368 4805 11392
rect 4485 10304 4493 10368
rect 4557 10304 4573 10368
rect 4637 10304 4653 10368
rect 4717 10304 4733 10368
rect 4797 10304 4805 10368
rect 4485 9280 4805 10304
rect 4485 9216 4493 9280
rect 4557 9216 4573 9280
rect 4637 9216 4653 9280
rect 4717 9216 4733 9280
rect 4797 9216 4805 9280
rect 4485 8192 4805 9216
rect 4485 8128 4493 8192
rect 4557 8128 4573 8192
rect 4637 8128 4653 8192
rect 4717 8128 4733 8192
rect 4797 8128 4805 8192
rect 4485 7104 4805 8128
rect 4485 7040 4493 7104
rect 4557 7040 4573 7104
rect 4637 7040 4653 7104
rect 4717 7040 4733 7104
rect 4797 7040 4805 7104
rect 4485 6016 4805 7040
rect 4485 5952 4493 6016
rect 4557 5952 4573 6016
rect 4637 5952 4653 6016
rect 4717 5952 4733 6016
rect 4797 5952 4805 6016
rect 4485 5830 4805 5952
rect 4485 5594 4527 5830
rect 4763 5594 4805 5830
rect 4485 4928 4805 5594
rect 4485 4864 4493 4928
rect 4557 4864 4573 4928
rect 4637 4864 4653 4928
rect 4717 4864 4733 4928
rect 4797 4864 4805 4928
rect 4485 3840 4805 4864
rect 4485 3776 4493 3840
rect 4557 3776 4573 3840
rect 4637 3776 4653 3840
rect 4717 3776 4733 3840
rect 4797 3776 4805 3840
rect 4485 2752 4805 3776
rect 4485 2688 4493 2752
rect 4557 2688 4573 2752
rect 4637 2688 4653 2752
rect 4717 2688 4733 2752
rect 4797 2688 4805 2752
rect 4485 2128 4805 2688
rect 5145 30496 5465 30512
rect 5145 30432 5153 30496
rect 5217 30432 5233 30496
rect 5297 30432 5313 30496
rect 5377 30432 5393 30496
rect 5457 30432 5465 30496
rect 5145 29408 5465 30432
rect 5145 29344 5153 29408
rect 5217 29344 5233 29408
rect 5297 29344 5313 29408
rect 5377 29344 5393 29408
rect 5457 29344 5465 29408
rect 5145 28320 5465 29344
rect 5145 28256 5153 28320
rect 5217 28256 5233 28320
rect 5297 28256 5313 28320
rect 5377 28256 5393 28320
rect 5457 28256 5465 28320
rect 5145 27706 5465 28256
rect 5145 27470 5187 27706
rect 5423 27470 5465 27706
rect 5145 27232 5465 27470
rect 5145 27168 5153 27232
rect 5217 27168 5233 27232
rect 5297 27168 5313 27232
rect 5377 27168 5393 27232
rect 5457 27168 5465 27232
rect 5145 26144 5465 27168
rect 5145 26080 5153 26144
rect 5217 26080 5233 26144
rect 5297 26080 5313 26144
rect 5377 26080 5393 26144
rect 5457 26080 5465 26144
rect 5145 25056 5465 26080
rect 5145 24992 5153 25056
rect 5217 24992 5233 25056
rect 5297 24992 5313 25056
rect 5377 24992 5393 25056
rect 5457 24992 5465 25056
rect 5145 23968 5465 24992
rect 5145 23904 5153 23968
rect 5217 23904 5233 23968
rect 5297 23904 5313 23968
rect 5377 23904 5393 23968
rect 5457 23904 5465 23968
rect 5145 22880 5465 23904
rect 5145 22816 5153 22880
rect 5217 22816 5233 22880
rect 5297 22816 5313 22880
rect 5377 22816 5393 22880
rect 5457 22816 5465 22880
rect 5145 21792 5465 22816
rect 5145 21728 5153 21792
rect 5217 21728 5233 21792
rect 5297 21728 5313 21792
rect 5377 21728 5393 21792
rect 5457 21728 5465 21792
rect 5145 20704 5465 21728
rect 5145 20640 5153 20704
rect 5217 20640 5233 20704
rect 5297 20640 5313 20704
rect 5377 20640 5393 20704
rect 5457 20640 5465 20704
rect 5145 20634 5465 20640
rect 5145 20398 5187 20634
rect 5423 20398 5465 20634
rect 5145 19616 5465 20398
rect 5145 19552 5153 19616
rect 5217 19552 5233 19616
rect 5297 19552 5313 19616
rect 5377 19552 5393 19616
rect 5457 19552 5465 19616
rect 5145 18528 5465 19552
rect 5145 18464 5153 18528
rect 5217 18464 5233 18528
rect 5297 18464 5313 18528
rect 5377 18464 5393 18528
rect 5457 18464 5465 18528
rect 5145 17440 5465 18464
rect 5145 17376 5153 17440
rect 5217 17376 5233 17440
rect 5297 17376 5313 17440
rect 5377 17376 5393 17440
rect 5457 17376 5465 17440
rect 5145 16352 5465 17376
rect 5145 16288 5153 16352
rect 5217 16288 5233 16352
rect 5297 16288 5313 16352
rect 5377 16288 5393 16352
rect 5457 16288 5465 16352
rect 5145 15264 5465 16288
rect 5145 15200 5153 15264
rect 5217 15200 5233 15264
rect 5297 15200 5313 15264
rect 5377 15200 5393 15264
rect 5457 15200 5465 15264
rect 5145 14176 5465 15200
rect 5145 14112 5153 14176
rect 5217 14112 5233 14176
rect 5297 14112 5313 14176
rect 5377 14112 5393 14176
rect 5457 14112 5465 14176
rect 5145 13562 5465 14112
rect 11568 29952 11888 30512
rect 11568 29888 11576 29952
rect 11640 29888 11656 29952
rect 11720 29888 11736 29952
rect 11800 29888 11816 29952
rect 11880 29888 11888 29952
rect 11568 28864 11888 29888
rect 11568 28800 11576 28864
rect 11640 28800 11656 28864
rect 11720 28800 11736 28864
rect 11800 28800 11816 28864
rect 11880 28800 11888 28864
rect 11568 27776 11888 28800
rect 11568 27712 11576 27776
rect 11640 27712 11656 27776
rect 11720 27712 11736 27776
rect 11800 27712 11816 27776
rect 11880 27712 11888 27776
rect 11568 27046 11888 27712
rect 11568 26810 11610 27046
rect 11846 26810 11888 27046
rect 11568 26688 11888 26810
rect 11568 26624 11576 26688
rect 11640 26624 11656 26688
rect 11720 26624 11736 26688
rect 11800 26624 11816 26688
rect 11880 26624 11888 26688
rect 11568 25600 11888 26624
rect 11568 25536 11576 25600
rect 11640 25536 11656 25600
rect 11720 25536 11736 25600
rect 11800 25536 11816 25600
rect 11880 25536 11888 25600
rect 11568 24512 11888 25536
rect 11568 24448 11576 24512
rect 11640 24448 11656 24512
rect 11720 24448 11736 24512
rect 11800 24448 11816 24512
rect 11880 24448 11888 24512
rect 11568 23424 11888 24448
rect 11568 23360 11576 23424
rect 11640 23360 11656 23424
rect 11720 23360 11736 23424
rect 11800 23360 11816 23424
rect 11880 23360 11888 23424
rect 11568 22336 11888 23360
rect 11568 22272 11576 22336
rect 11640 22272 11656 22336
rect 11720 22272 11736 22336
rect 11800 22272 11816 22336
rect 11880 22272 11888 22336
rect 11568 21248 11888 22272
rect 11568 21184 11576 21248
rect 11640 21184 11656 21248
rect 11720 21184 11736 21248
rect 11800 21184 11816 21248
rect 11880 21184 11888 21248
rect 11568 20160 11888 21184
rect 11568 20096 11576 20160
rect 11640 20096 11656 20160
rect 11720 20096 11736 20160
rect 11800 20096 11816 20160
rect 11880 20096 11888 20160
rect 11568 19974 11888 20096
rect 11568 19738 11610 19974
rect 11846 19738 11888 19974
rect 11568 19072 11888 19738
rect 11568 19008 11576 19072
rect 11640 19008 11656 19072
rect 11720 19008 11736 19072
rect 11800 19008 11816 19072
rect 11880 19008 11888 19072
rect 11568 17984 11888 19008
rect 11568 17920 11576 17984
rect 11640 17920 11656 17984
rect 11720 17920 11736 17984
rect 11800 17920 11816 17984
rect 11880 17920 11888 17984
rect 11568 16896 11888 17920
rect 11568 16832 11576 16896
rect 11640 16832 11656 16896
rect 11720 16832 11736 16896
rect 11800 16832 11816 16896
rect 11880 16832 11888 16896
rect 11568 15808 11888 16832
rect 11568 15744 11576 15808
rect 11640 15744 11656 15808
rect 11720 15744 11736 15808
rect 11800 15744 11816 15808
rect 11880 15744 11888 15808
rect 11568 14720 11888 15744
rect 11568 14656 11576 14720
rect 11640 14656 11656 14720
rect 11720 14656 11736 14720
rect 11800 14656 11816 14720
rect 11880 14656 11888 14720
rect 10547 13836 10613 13837
rect 10547 13772 10548 13836
rect 10612 13772 10613 13836
rect 10547 13771 10613 13772
rect 5145 13326 5187 13562
rect 5423 13326 5465 13562
rect 5145 13088 5465 13326
rect 5145 13024 5153 13088
rect 5217 13024 5233 13088
rect 5297 13024 5313 13088
rect 5377 13024 5393 13088
rect 5457 13024 5465 13088
rect 5145 12000 5465 13024
rect 5145 11936 5153 12000
rect 5217 11936 5233 12000
rect 5297 11936 5313 12000
rect 5377 11936 5393 12000
rect 5457 11936 5465 12000
rect 5145 10912 5465 11936
rect 5145 10848 5153 10912
rect 5217 10848 5233 10912
rect 5297 10848 5313 10912
rect 5377 10848 5393 10912
rect 5457 10848 5465 10912
rect 5145 9824 5465 10848
rect 5145 9760 5153 9824
rect 5217 9760 5233 9824
rect 5297 9760 5313 9824
rect 5377 9760 5393 9824
rect 5457 9760 5465 9824
rect 5145 8736 5465 9760
rect 5145 8672 5153 8736
rect 5217 8672 5233 8736
rect 5297 8672 5313 8736
rect 5377 8672 5393 8736
rect 5457 8672 5465 8736
rect 5145 7648 5465 8672
rect 10550 8261 10610 13771
rect 11568 13632 11888 14656
rect 11568 13568 11576 13632
rect 11640 13568 11656 13632
rect 11720 13568 11736 13632
rect 11800 13568 11816 13632
rect 11880 13568 11888 13632
rect 10731 13292 10797 13293
rect 10731 13228 10732 13292
rect 10796 13228 10797 13292
rect 10731 13227 10797 13228
rect 10547 8260 10613 8261
rect 10547 8196 10548 8260
rect 10612 8196 10613 8260
rect 10547 8195 10613 8196
rect 10734 8125 10794 13227
rect 11568 12902 11888 13568
rect 11568 12666 11610 12902
rect 11846 12666 11888 12902
rect 11568 12544 11888 12666
rect 11568 12480 11576 12544
rect 11640 12480 11656 12544
rect 11720 12480 11736 12544
rect 11800 12480 11816 12544
rect 11880 12480 11888 12544
rect 11568 11456 11888 12480
rect 11568 11392 11576 11456
rect 11640 11392 11656 11456
rect 11720 11392 11736 11456
rect 11800 11392 11816 11456
rect 11880 11392 11888 11456
rect 11568 10368 11888 11392
rect 11568 10304 11576 10368
rect 11640 10304 11656 10368
rect 11720 10304 11736 10368
rect 11800 10304 11816 10368
rect 11880 10304 11888 10368
rect 11568 9280 11888 10304
rect 11568 9216 11576 9280
rect 11640 9216 11656 9280
rect 11720 9216 11736 9280
rect 11800 9216 11816 9280
rect 11880 9216 11888 9280
rect 11568 8192 11888 9216
rect 11568 8128 11576 8192
rect 11640 8128 11656 8192
rect 11720 8128 11736 8192
rect 11800 8128 11816 8192
rect 11880 8128 11888 8192
rect 10731 8124 10797 8125
rect 10731 8060 10732 8124
rect 10796 8060 10797 8124
rect 10731 8059 10797 8060
rect 5145 7584 5153 7648
rect 5217 7584 5233 7648
rect 5297 7584 5313 7648
rect 5377 7584 5393 7648
rect 5457 7584 5465 7648
rect 5145 6560 5465 7584
rect 5145 6496 5153 6560
rect 5217 6496 5233 6560
rect 5297 6496 5313 6560
rect 5377 6496 5393 6560
rect 5457 6496 5465 6560
rect 5145 6490 5465 6496
rect 5145 6254 5187 6490
rect 5423 6254 5465 6490
rect 5145 5472 5465 6254
rect 5145 5408 5153 5472
rect 5217 5408 5233 5472
rect 5297 5408 5313 5472
rect 5377 5408 5393 5472
rect 5457 5408 5465 5472
rect 5145 4384 5465 5408
rect 5145 4320 5153 4384
rect 5217 4320 5233 4384
rect 5297 4320 5313 4384
rect 5377 4320 5393 4384
rect 5457 4320 5465 4384
rect 5145 3296 5465 4320
rect 5145 3232 5153 3296
rect 5217 3232 5233 3296
rect 5297 3232 5313 3296
rect 5377 3232 5393 3296
rect 5457 3232 5465 3296
rect 5145 2208 5465 3232
rect 5145 2144 5153 2208
rect 5217 2144 5233 2208
rect 5297 2144 5313 2208
rect 5377 2144 5393 2208
rect 5457 2144 5465 2208
rect 5145 2128 5465 2144
rect 11568 7104 11888 8128
rect 11568 7040 11576 7104
rect 11640 7040 11656 7104
rect 11720 7040 11736 7104
rect 11800 7040 11816 7104
rect 11880 7040 11888 7104
rect 11568 6016 11888 7040
rect 11568 5952 11576 6016
rect 11640 5952 11656 6016
rect 11720 5952 11736 6016
rect 11800 5952 11816 6016
rect 11880 5952 11888 6016
rect 11568 5830 11888 5952
rect 11568 5594 11610 5830
rect 11846 5594 11888 5830
rect 11568 4928 11888 5594
rect 11568 4864 11576 4928
rect 11640 4864 11656 4928
rect 11720 4864 11736 4928
rect 11800 4864 11816 4928
rect 11880 4864 11888 4928
rect 11568 3840 11888 4864
rect 11568 3776 11576 3840
rect 11640 3776 11656 3840
rect 11720 3776 11736 3840
rect 11800 3776 11816 3840
rect 11880 3776 11888 3840
rect 11568 2752 11888 3776
rect 11568 2688 11576 2752
rect 11640 2688 11656 2752
rect 11720 2688 11736 2752
rect 11800 2688 11816 2752
rect 11880 2688 11888 2752
rect 11568 2128 11888 2688
rect 12228 30496 12548 30512
rect 12228 30432 12236 30496
rect 12300 30432 12316 30496
rect 12380 30432 12396 30496
rect 12460 30432 12476 30496
rect 12540 30432 12548 30496
rect 12228 29408 12548 30432
rect 12228 29344 12236 29408
rect 12300 29344 12316 29408
rect 12380 29344 12396 29408
rect 12460 29344 12476 29408
rect 12540 29344 12548 29408
rect 12228 28320 12548 29344
rect 12228 28256 12236 28320
rect 12300 28256 12316 28320
rect 12380 28256 12396 28320
rect 12460 28256 12476 28320
rect 12540 28256 12548 28320
rect 12228 27706 12548 28256
rect 12228 27470 12270 27706
rect 12506 27470 12548 27706
rect 12228 27232 12548 27470
rect 12228 27168 12236 27232
rect 12300 27168 12316 27232
rect 12380 27168 12396 27232
rect 12460 27168 12476 27232
rect 12540 27168 12548 27232
rect 12228 26144 12548 27168
rect 12228 26080 12236 26144
rect 12300 26080 12316 26144
rect 12380 26080 12396 26144
rect 12460 26080 12476 26144
rect 12540 26080 12548 26144
rect 12228 25056 12548 26080
rect 12228 24992 12236 25056
rect 12300 24992 12316 25056
rect 12380 24992 12396 25056
rect 12460 24992 12476 25056
rect 12540 24992 12548 25056
rect 12228 23968 12548 24992
rect 12228 23904 12236 23968
rect 12300 23904 12316 23968
rect 12380 23904 12396 23968
rect 12460 23904 12476 23968
rect 12540 23904 12548 23968
rect 12228 22880 12548 23904
rect 12228 22816 12236 22880
rect 12300 22816 12316 22880
rect 12380 22816 12396 22880
rect 12460 22816 12476 22880
rect 12540 22816 12548 22880
rect 12228 21792 12548 22816
rect 12228 21728 12236 21792
rect 12300 21728 12316 21792
rect 12380 21728 12396 21792
rect 12460 21728 12476 21792
rect 12540 21728 12548 21792
rect 12228 20704 12548 21728
rect 12228 20640 12236 20704
rect 12300 20640 12316 20704
rect 12380 20640 12396 20704
rect 12460 20640 12476 20704
rect 12540 20640 12548 20704
rect 12228 20634 12548 20640
rect 12228 20398 12270 20634
rect 12506 20398 12548 20634
rect 12228 19616 12548 20398
rect 12228 19552 12236 19616
rect 12300 19552 12316 19616
rect 12380 19552 12396 19616
rect 12460 19552 12476 19616
rect 12540 19552 12548 19616
rect 12228 18528 12548 19552
rect 12228 18464 12236 18528
rect 12300 18464 12316 18528
rect 12380 18464 12396 18528
rect 12460 18464 12476 18528
rect 12540 18464 12548 18528
rect 12228 17440 12548 18464
rect 12228 17376 12236 17440
rect 12300 17376 12316 17440
rect 12380 17376 12396 17440
rect 12460 17376 12476 17440
rect 12540 17376 12548 17440
rect 12228 16352 12548 17376
rect 12228 16288 12236 16352
rect 12300 16288 12316 16352
rect 12380 16288 12396 16352
rect 12460 16288 12476 16352
rect 12540 16288 12548 16352
rect 12228 15264 12548 16288
rect 12228 15200 12236 15264
rect 12300 15200 12316 15264
rect 12380 15200 12396 15264
rect 12460 15200 12476 15264
rect 12540 15200 12548 15264
rect 12228 14176 12548 15200
rect 12228 14112 12236 14176
rect 12300 14112 12316 14176
rect 12380 14112 12396 14176
rect 12460 14112 12476 14176
rect 12540 14112 12548 14176
rect 12228 13562 12548 14112
rect 12228 13326 12270 13562
rect 12506 13326 12548 13562
rect 12228 13088 12548 13326
rect 12228 13024 12236 13088
rect 12300 13024 12316 13088
rect 12380 13024 12396 13088
rect 12460 13024 12476 13088
rect 12540 13024 12548 13088
rect 12228 12000 12548 13024
rect 12228 11936 12236 12000
rect 12300 11936 12316 12000
rect 12380 11936 12396 12000
rect 12460 11936 12476 12000
rect 12540 11936 12548 12000
rect 12228 10912 12548 11936
rect 12228 10848 12236 10912
rect 12300 10848 12316 10912
rect 12380 10848 12396 10912
rect 12460 10848 12476 10912
rect 12540 10848 12548 10912
rect 12228 9824 12548 10848
rect 12228 9760 12236 9824
rect 12300 9760 12316 9824
rect 12380 9760 12396 9824
rect 12460 9760 12476 9824
rect 12540 9760 12548 9824
rect 12228 8736 12548 9760
rect 12228 8672 12236 8736
rect 12300 8672 12316 8736
rect 12380 8672 12396 8736
rect 12460 8672 12476 8736
rect 12540 8672 12548 8736
rect 12228 7648 12548 8672
rect 12228 7584 12236 7648
rect 12300 7584 12316 7648
rect 12380 7584 12396 7648
rect 12460 7584 12476 7648
rect 12540 7584 12548 7648
rect 12228 6560 12548 7584
rect 12228 6496 12236 6560
rect 12300 6496 12316 6560
rect 12380 6496 12396 6560
rect 12460 6496 12476 6560
rect 12540 6496 12548 6560
rect 12228 6490 12548 6496
rect 12228 6254 12270 6490
rect 12506 6254 12548 6490
rect 12228 5472 12548 6254
rect 12228 5408 12236 5472
rect 12300 5408 12316 5472
rect 12380 5408 12396 5472
rect 12460 5408 12476 5472
rect 12540 5408 12548 5472
rect 12228 4384 12548 5408
rect 12228 4320 12236 4384
rect 12300 4320 12316 4384
rect 12380 4320 12396 4384
rect 12460 4320 12476 4384
rect 12540 4320 12548 4384
rect 12228 3296 12548 4320
rect 12228 3232 12236 3296
rect 12300 3232 12316 3296
rect 12380 3232 12396 3296
rect 12460 3232 12476 3296
rect 12540 3232 12548 3296
rect 12228 2208 12548 3232
rect 12228 2144 12236 2208
rect 12300 2144 12316 2208
rect 12380 2144 12396 2208
rect 12460 2144 12476 2208
rect 12540 2144 12548 2208
rect 12228 2128 12548 2144
rect 18651 29952 18971 30512
rect 18651 29888 18659 29952
rect 18723 29888 18739 29952
rect 18803 29888 18819 29952
rect 18883 29888 18899 29952
rect 18963 29888 18971 29952
rect 18651 28864 18971 29888
rect 18651 28800 18659 28864
rect 18723 28800 18739 28864
rect 18803 28800 18819 28864
rect 18883 28800 18899 28864
rect 18963 28800 18971 28864
rect 18651 27776 18971 28800
rect 18651 27712 18659 27776
rect 18723 27712 18739 27776
rect 18803 27712 18819 27776
rect 18883 27712 18899 27776
rect 18963 27712 18971 27776
rect 18651 27046 18971 27712
rect 18651 26810 18693 27046
rect 18929 26810 18971 27046
rect 18651 26688 18971 26810
rect 18651 26624 18659 26688
rect 18723 26624 18739 26688
rect 18803 26624 18819 26688
rect 18883 26624 18899 26688
rect 18963 26624 18971 26688
rect 18651 25600 18971 26624
rect 18651 25536 18659 25600
rect 18723 25536 18739 25600
rect 18803 25536 18819 25600
rect 18883 25536 18899 25600
rect 18963 25536 18971 25600
rect 18651 24512 18971 25536
rect 18651 24448 18659 24512
rect 18723 24448 18739 24512
rect 18803 24448 18819 24512
rect 18883 24448 18899 24512
rect 18963 24448 18971 24512
rect 18651 23424 18971 24448
rect 18651 23360 18659 23424
rect 18723 23360 18739 23424
rect 18803 23360 18819 23424
rect 18883 23360 18899 23424
rect 18963 23360 18971 23424
rect 18651 22336 18971 23360
rect 18651 22272 18659 22336
rect 18723 22272 18739 22336
rect 18803 22272 18819 22336
rect 18883 22272 18899 22336
rect 18963 22272 18971 22336
rect 18651 21248 18971 22272
rect 18651 21184 18659 21248
rect 18723 21184 18739 21248
rect 18803 21184 18819 21248
rect 18883 21184 18899 21248
rect 18963 21184 18971 21248
rect 18651 20160 18971 21184
rect 18651 20096 18659 20160
rect 18723 20096 18739 20160
rect 18803 20096 18819 20160
rect 18883 20096 18899 20160
rect 18963 20096 18971 20160
rect 18651 19974 18971 20096
rect 18651 19738 18693 19974
rect 18929 19738 18971 19974
rect 18651 19072 18971 19738
rect 18651 19008 18659 19072
rect 18723 19008 18739 19072
rect 18803 19008 18819 19072
rect 18883 19008 18899 19072
rect 18963 19008 18971 19072
rect 18651 17984 18971 19008
rect 18651 17920 18659 17984
rect 18723 17920 18739 17984
rect 18803 17920 18819 17984
rect 18883 17920 18899 17984
rect 18963 17920 18971 17984
rect 18651 16896 18971 17920
rect 18651 16832 18659 16896
rect 18723 16832 18739 16896
rect 18803 16832 18819 16896
rect 18883 16832 18899 16896
rect 18963 16832 18971 16896
rect 18651 15808 18971 16832
rect 18651 15744 18659 15808
rect 18723 15744 18739 15808
rect 18803 15744 18819 15808
rect 18883 15744 18899 15808
rect 18963 15744 18971 15808
rect 18651 14720 18971 15744
rect 18651 14656 18659 14720
rect 18723 14656 18739 14720
rect 18803 14656 18819 14720
rect 18883 14656 18899 14720
rect 18963 14656 18971 14720
rect 18651 13632 18971 14656
rect 18651 13568 18659 13632
rect 18723 13568 18739 13632
rect 18803 13568 18819 13632
rect 18883 13568 18899 13632
rect 18963 13568 18971 13632
rect 18651 12902 18971 13568
rect 18651 12666 18693 12902
rect 18929 12666 18971 12902
rect 18651 12544 18971 12666
rect 18651 12480 18659 12544
rect 18723 12480 18739 12544
rect 18803 12480 18819 12544
rect 18883 12480 18899 12544
rect 18963 12480 18971 12544
rect 18651 11456 18971 12480
rect 18651 11392 18659 11456
rect 18723 11392 18739 11456
rect 18803 11392 18819 11456
rect 18883 11392 18899 11456
rect 18963 11392 18971 11456
rect 18651 10368 18971 11392
rect 18651 10304 18659 10368
rect 18723 10304 18739 10368
rect 18803 10304 18819 10368
rect 18883 10304 18899 10368
rect 18963 10304 18971 10368
rect 18651 9280 18971 10304
rect 18651 9216 18659 9280
rect 18723 9216 18739 9280
rect 18803 9216 18819 9280
rect 18883 9216 18899 9280
rect 18963 9216 18971 9280
rect 18651 8192 18971 9216
rect 18651 8128 18659 8192
rect 18723 8128 18739 8192
rect 18803 8128 18819 8192
rect 18883 8128 18899 8192
rect 18963 8128 18971 8192
rect 18651 7104 18971 8128
rect 18651 7040 18659 7104
rect 18723 7040 18739 7104
rect 18803 7040 18819 7104
rect 18883 7040 18899 7104
rect 18963 7040 18971 7104
rect 18651 6016 18971 7040
rect 18651 5952 18659 6016
rect 18723 5952 18739 6016
rect 18803 5952 18819 6016
rect 18883 5952 18899 6016
rect 18963 5952 18971 6016
rect 18651 5830 18971 5952
rect 18651 5594 18693 5830
rect 18929 5594 18971 5830
rect 18651 4928 18971 5594
rect 18651 4864 18659 4928
rect 18723 4864 18739 4928
rect 18803 4864 18819 4928
rect 18883 4864 18899 4928
rect 18963 4864 18971 4928
rect 18651 3840 18971 4864
rect 18651 3776 18659 3840
rect 18723 3776 18739 3840
rect 18803 3776 18819 3840
rect 18883 3776 18899 3840
rect 18963 3776 18971 3840
rect 18651 2752 18971 3776
rect 18651 2688 18659 2752
rect 18723 2688 18739 2752
rect 18803 2688 18819 2752
rect 18883 2688 18899 2752
rect 18963 2688 18971 2752
rect 18651 2128 18971 2688
rect 19311 30496 19631 30512
rect 19311 30432 19319 30496
rect 19383 30432 19399 30496
rect 19463 30432 19479 30496
rect 19543 30432 19559 30496
rect 19623 30432 19631 30496
rect 19311 29408 19631 30432
rect 19311 29344 19319 29408
rect 19383 29344 19399 29408
rect 19463 29344 19479 29408
rect 19543 29344 19559 29408
rect 19623 29344 19631 29408
rect 19311 28320 19631 29344
rect 19311 28256 19319 28320
rect 19383 28256 19399 28320
rect 19463 28256 19479 28320
rect 19543 28256 19559 28320
rect 19623 28256 19631 28320
rect 19311 27706 19631 28256
rect 19311 27470 19353 27706
rect 19589 27470 19631 27706
rect 19311 27232 19631 27470
rect 19311 27168 19319 27232
rect 19383 27168 19399 27232
rect 19463 27168 19479 27232
rect 19543 27168 19559 27232
rect 19623 27168 19631 27232
rect 19311 26144 19631 27168
rect 19311 26080 19319 26144
rect 19383 26080 19399 26144
rect 19463 26080 19479 26144
rect 19543 26080 19559 26144
rect 19623 26080 19631 26144
rect 19311 25056 19631 26080
rect 19311 24992 19319 25056
rect 19383 24992 19399 25056
rect 19463 24992 19479 25056
rect 19543 24992 19559 25056
rect 19623 24992 19631 25056
rect 19311 23968 19631 24992
rect 19311 23904 19319 23968
rect 19383 23904 19399 23968
rect 19463 23904 19479 23968
rect 19543 23904 19559 23968
rect 19623 23904 19631 23968
rect 19311 22880 19631 23904
rect 19311 22816 19319 22880
rect 19383 22816 19399 22880
rect 19463 22816 19479 22880
rect 19543 22816 19559 22880
rect 19623 22816 19631 22880
rect 19311 21792 19631 22816
rect 25734 29952 26054 30512
rect 25734 29888 25742 29952
rect 25806 29888 25822 29952
rect 25886 29888 25902 29952
rect 25966 29888 25982 29952
rect 26046 29888 26054 29952
rect 25734 28864 26054 29888
rect 25734 28800 25742 28864
rect 25806 28800 25822 28864
rect 25886 28800 25902 28864
rect 25966 28800 25982 28864
rect 26046 28800 26054 28864
rect 25734 27776 26054 28800
rect 25734 27712 25742 27776
rect 25806 27712 25822 27776
rect 25886 27712 25902 27776
rect 25966 27712 25982 27776
rect 26046 27712 26054 27776
rect 25734 27046 26054 27712
rect 25734 26810 25776 27046
rect 26012 26810 26054 27046
rect 25734 26688 26054 26810
rect 25734 26624 25742 26688
rect 25806 26624 25822 26688
rect 25886 26624 25902 26688
rect 25966 26624 25982 26688
rect 26046 26624 26054 26688
rect 25734 25600 26054 26624
rect 25734 25536 25742 25600
rect 25806 25536 25822 25600
rect 25886 25536 25902 25600
rect 25966 25536 25982 25600
rect 26046 25536 26054 25600
rect 25734 24512 26054 25536
rect 25734 24448 25742 24512
rect 25806 24448 25822 24512
rect 25886 24448 25902 24512
rect 25966 24448 25982 24512
rect 26046 24448 26054 24512
rect 25734 23424 26054 24448
rect 25734 23360 25742 23424
rect 25806 23360 25822 23424
rect 25886 23360 25902 23424
rect 25966 23360 25982 23424
rect 26046 23360 26054 23424
rect 24347 22540 24413 22541
rect 24347 22476 24348 22540
rect 24412 22476 24413 22540
rect 24347 22475 24413 22476
rect 19311 21728 19319 21792
rect 19383 21728 19399 21792
rect 19463 21728 19479 21792
rect 19543 21728 19559 21792
rect 19623 21728 19631 21792
rect 19311 20704 19631 21728
rect 19311 20640 19319 20704
rect 19383 20640 19399 20704
rect 19463 20640 19479 20704
rect 19543 20640 19559 20704
rect 19623 20640 19631 20704
rect 19311 20634 19631 20640
rect 19311 20398 19353 20634
rect 19589 20398 19631 20634
rect 19311 19616 19631 20398
rect 19311 19552 19319 19616
rect 19383 19552 19399 19616
rect 19463 19552 19479 19616
rect 19543 19552 19559 19616
rect 19623 19552 19631 19616
rect 19311 18528 19631 19552
rect 19311 18464 19319 18528
rect 19383 18464 19399 18528
rect 19463 18464 19479 18528
rect 19543 18464 19559 18528
rect 19623 18464 19631 18528
rect 19311 17440 19631 18464
rect 19311 17376 19319 17440
rect 19383 17376 19399 17440
rect 19463 17376 19479 17440
rect 19543 17376 19559 17440
rect 19623 17376 19631 17440
rect 19311 16352 19631 17376
rect 19311 16288 19319 16352
rect 19383 16288 19399 16352
rect 19463 16288 19479 16352
rect 19543 16288 19559 16352
rect 19623 16288 19631 16352
rect 19311 15264 19631 16288
rect 19311 15200 19319 15264
rect 19383 15200 19399 15264
rect 19463 15200 19479 15264
rect 19543 15200 19559 15264
rect 19623 15200 19631 15264
rect 19311 14176 19631 15200
rect 19311 14112 19319 14176
rect 19383 14112 19399 14176
rect 19463 14112 19479 14176
rect 19543 14112 19559 14176
rect 19623 14112 19631 14176
rect 19311 13562 19631 14112
rect 19311 13326 19353 13562
rect 19589 13326 19631 13562
rect 19311 13088 19631 13326
rect 19311 13024 19319 13088
rect 19383 13024 19399 13088
rect 19463 13024 19479 13088
rect 19543 13024 19559 13088
rect 19623 13024 19631 13088
rect 19311 12000 19631 13024
rect 19311 11936 19319 12000
rect 19383 11936 19399 12000
rect 19463 11936 19479 12000
rect 19543 11936 19559 12000
rect 19623 11936 19631 12000
rect 19311 10912 19631 11936
rect 19311 10848 19319 10912
rect 19383 10848 19399 10912
rect 19463 10848 19479 10912
rect 19543 10848 19559 10912
rect 19623 10848 19631 10912
rect 19311 9824 19631 10848
rect 19311 9760 19319 9824
rect 19383 9760 19399 9824
rect 19463 9760 19479 9824
rect 19543 9760 19559 9824
rect 19623 9760 19631 9824
rect 19311 8736 19631 9760
rect 19311 8672 19319 8736
rect 19383 8672 19399 8736
rect 19463 8672 19479 8736
rect 19543 8672 19559 8736
rect 19623 8672 19631 8736
rect 19311 7648 19631 8672
rect 19311 7584 19319 7648
rect 19383 7584 19399 7648
rect 19463 7584 19479 7648
rect 19543 7584 19559 7648
rect 19623 7584 19631 7648
rect 19311 6560 19631 7584
rect 19311 6496 19319 6560
rect 19383 6496 19399 6560
rect 19463 6496 19479 6560
rect 19543 6496 19559 6560
rect 19623 6496 19631 6560
rect 19311 6490 19631 6496
rect 19311 6254 19353 6490
rect 19589 6254 19631 6490
rect 19311 5472 19631 6254
rect 24350 5541 24410 22475
rect 25734 22336 26054 23360
rect 25734 22272 25742 22336
rect 25806 22272 25822 22336
rect 25886 22272 25902 22336
rect 25966 22272 25982 22336
rect 26046 22272 26054 22336
rect 25734 21248 26054 22272
rect 25734 21184 25742 21248
rect 25806 21184 25822 21248
rect 25886 21184 25902 21248
rect 25966 21184 25982 21248
rect 26046 21184 26054 21248
rect 25734 20160 26054 21184
rect 25734 20096 25742 20160
rect 25806 20096 25822 20160
rect 25886 20096 25902 20160
rect 25966 20096 25982 20160
rect 26046 20096 26054 20160
rect 25734 19974 26054 20096
rect 25734 19738 25776 19974
rect 26012 19738 26054 19974
rect 25734 19072 26054 19738
rect 25734 19008 25742 19072
rect 25806 19008 25822 19072
rect 25886 19008 25902 19072
rect 25966 19008 25982 19072
rect 26046 19008 26054 19072
rect 25734 17984 26054 19008
rect 25734 17920 25742 17984
rect 25806 17920 25822 17984
rect 25886 17920 25902 17984
rect 25966 17920 25982 17984
rect 26046 17920 26054 17984
rect 25734 16896 26054 17920
rect 25734 16832 25742 16896
rect 25806 16832 25822 16896
rect 25886 16832 25902 16896
rect 25966 16832 25982 16896
rect 26046 16832 26054 16896
rect 25734 15808 26054 16832
rect 25734 15744 25742 15808
rect 25806 15744 25822 15808
rect 25886 15744 25902 15808
rect 25966 15744 25982 15808
rect 26046 15744 26054 15808
rect 25734 14720 26054 15744
rect 25734 14656 25742 14720
rect 25806 14656 25822 14720
rect 25886 14656 25902 14720
rect 25966 14656 25982 14720
rect 26046 14656 26054 14720
rect 25734 13632 26054 14656
rect 25734 13568 25742 13632
rect 25806 13568 25822 13632
rect 25886 13568 25902 13632
rect 25966 13568 25982 13632
rect 26046 13568 26054 13632
rect 25734 12902 26054 13568
rect 25734 12666 25776 12902
rect 26012 12666 26054 12902
rect 25734 12544 26054 12666
rect 25734 12480 25742 12544
rect 25806 12480 25822 12544
rect 25886 12480 25902 12544
rect 25966 12480 25982 12544
rect 26046 12480 26054 12544
rect 25734 11456 26054 12480
rect 25734 11392 25742 11456
rect 25806 11392 25822 11456
rect 25886 11392 25902 11456
rect 25966 11392 25982 11456
rect 26046 11392 26054 11456
rect 25734 10368 26054 11392
rect 25734 10304 25742 10368
rect 25806 10304 25822 10368
rect 25886 10304 25902 10368
rect 25966 10304 25982 10368
rect 26046 10304 26054 10368
rect 25734 9280 26054 10304
rect 25734 9216 25742 9280
rect 25806 9216 25822 9280
rect 25886 9216 25902 9280
rect 25966 9216 25982 9280
rect 26046 9216 26054 9280
rect 25734 8192 26054 9216
rect 25734 8128 25742 8192
rect 25806 8128 25822 8192
rect 25886 8128 25902 8192
rect 25966 8128 25982 8192
rect 26046 8128 26054 8192
rect 25734 7104 26054 8128
rect 25734 7040 25742 7104
rect 25806 7040 25822 7104
rect 25886 7040 25902 7104
rect 25966 7040 25982 7104
rect 26046 7040 26054 7104
rect 25734 6016 26054 7040
rect 25734 5952 25742 6016
rect 25806 5952 25822 6016
rect 25886 5952 25902 6016
rect 25966 5952 25982 6016
rect 26046 5952 26054 6016
rect 25734 5830 26054 5952
rect 25734 5594 25776 5830
rect 26012 5594 26054 5830
rect 24347 5540 24413 5541
rect 24347 5476 24348 5540
rect 24412 5476 24413 5540
rect 24347 5475 24413 5476
rect 19311 5408 19319 5472
rect 19383 5408 19399 5472
rect 19463 5408 19479 5472
rect 19543 5408 19559 5472
rect 19623 5408 19631 5472
rect 19311 4384 19631 5408
rect 19311 4320 19319 4384
rect 19383 4320 19399 4384
rect 19463 4320 19479 4384
rect 19543 4320 19559 4384
rect 19623 4320 19631 4384
rect 19311 3296 19631 4320
rect 19311 3232 19319 3296
rect 19383 3232 19399 3296
rect 19463 3232 19479 3296
rect 19543 3232 19559 3296
rect 19623 3232 19631 3296
rect 19311 2208 19631 3232
rect 19311 2144 19319 2208
rect 19383 2144 19399 2208
rect 19463 2144 19479 2208
rect 19543 2144 19559 2208
rect 19623 2144 19631 2208
rect 19311 2128 19631 2144
rect 25734 4928 26054 5594
rect 25734 4864 25742 4928
rect 25806 4864 25822 4928
rect 25886 4864 25902 4928
rect 25966 4864 25982 4928
rect 26046 4864 26054 4928
rect 25734 3840 26054 4864
rect 25734 3776 25742 3840
rect 25806 3776 25822 3840
rect 25886 3776 25902 3840
rect 25966 3776 25982 3840
rect 26046 3776 26054 3840
rect 25734 2752 26054 3776
rect 25734 2688 25742 2752
rect 25806 2688 25822 2752
rect 25886 2688 25902 2752
rect 25966 2688 25982 2752
rect 26046 2688 26054 2752
rect 25734 2128 26054 2688
rect 26394 30496 26714 30512
rect 26394 30432 26402 30496
rect 26466 30432 26482 30496
rect 26546 30432 26562 30496
rect 26626 30432 26642 30496
rect 26706 30432 26714 30496
rect 26394 29408 26714 30432
rect 26394 29344 26402 29408
rect 26466 29344 26482 29408
rect 26546 29344 26562 29408
rect 26626 29344 26642 29408
rect 26706 29344 26714 29408
rect 26394 28320 26714 29344
rect 28763 29068 28829 29069
rect 28763 29004 28764 29068
rect 28828 29004 28829 29068
rect 28763 29003 28829 29004
rect 26394 28256 26402 28320
rect 26466 28256 26482 28320
rect 26546 28256 26562 28320
rect 26626 28256 26642 28320
rect 26706 28256 26714 28320
rect 26394 27706 26714 28256
rect 26394 27470 26436 27706
rect 26672 27470 26714 27706
rect 26394 27232 26714 27470
rect 26394 27168 26402 27232
rect 26466 27168 26482 27232
rect 26546 27168 26562 27232
rect 26626 27168 26642 27232
rect 26706 27168 26714 27232
rect 26394 26144 26714 27168
rect 26394 26080 26402 26144
rect 26466 26080 26482 26144
rect 26546 26080 26562 26144
rect 26626 26080 26642 26144
rect 26706 26080 26714 26144
rect 26394 25056 26714 26080
rect 26394 24992 26402 25056
rect 26466 24992 26482 25056
rect 26546 24992 26562 25056
rect 26626 24992 26642 25056
rect 26706 24992 26714 25056
rect 26394 23968 26714 24992
rect 26394 23904 26402 23968
rect 26466 23904 26482 23968
rect 26546 23904 26562 23968
rect 26626 23904 26642 23968
rect 26706 23904 26714 23968
rect 26394 22880 26714 23904
rect 26394 22816 26402 22880
rect 26466 22816 26482 22880
rect 26546 22816 26562 22880
rect 26626 22816 26642 22880
rect 26706 22816 26714 22880
rect 26394 21792 26714 22816
rect 26394 21728 26402 21792
rect 26466 21728 26482 21792
rect 26546 21728 26562 21792
rect 26626 21728 26642 21792
rect 26706 21728 26714 21792
rect 26394 20704 26714 21728
rect 26394 20640 26402 20704
rect 26466 20640 26482 20704
rect 26546 20640 26562 20704
rect 26626 20640 26642 20704
rect 26706 20640 26714 20704
rect 26394 20634 26714 20640
rect 26394 20398 26436 20634
rect 26672 20398 26714 20634
rect 26394 19616 26714 20398
rect 26394 19552 26402 19616
rect 26466 19552 26482 19616
rect 26546 19552 26562 19616
rect 26626 19552 26642 19616
rect 26706 19552 26714 19616
rect 26394 18528 26714 19552
rect 26394 18464 26402 18528
rect 26466 18464 26482 18528
rect 26546 18464 26562 18528
rect 26626 18464 26642 18528
rect 26706 18464 26714 18528
rect 26394 17440 26714 18464
rect 27659 18052 27725 18053
rect 27659 17988 27660 18052
rect 27724 17988 27725 18052
rect 27659 17987 27725 17988
rect 26394 17376 26402 17440
rect 26466 17376 26482 17440
rect 26546 17376 26562 17440
rect 26626 17376 26642 17440
rect 26706 17376 26714 17440
rect 26394 16352 26714 17376
rect 26394 16288 26402 16352
rect 26466 16288 26482 16352
rect 26546 16288 26562 16352
rect 26626 16288 26642 16352
rect 26706 16288 26714 16352
rect 26394 15264 26714 16288
rect 26394 15200 26402 15264
rect 26466 15200 26482 15264
rect 26546 15200 26562 15264
rect 26626 15200 26642 15264
rect 26706 15200 26714 15264
rect 26394 14176 26714 15200
rect 26394 14112 26402 14176
rect 26466 14112 26482 14176
rect 26546 14112 26562 14176
rect 26626 14112 26642 14176
rect 26706 14112 26714 14176
rect 26394 13562 26714 14112
rect 26394 13326 26436 13562
rect 26672 13326 26714 13562
rect 26394 13088 26714 13326
rect 26394 13024 26402 13088
rect 26466 13024 26482 13088
rect 26546 13024 26562 13088
rect 26626 13024 26642 13088
rect 26706 13024 26714 13088
rect 26394 12000 26714 13024
rect 26394 11936 26402 12000
rect 26466 11936 26482 12000
rect 26546 11936 26562 12000
rect 26626 11936 26642 12000
rect 26706 11936 26714 12000
rect 26394 10912 26714 11936
rect 27662 11797 27722 17987
rect 27659 11796 27725 11797
rect 27659 11732 27660 11796
rect 27724 11732 27725 11796
rect 27659 11731 27725 11732
rect 26394 10848 26402 10912
rect 26466 10848 26482 10912
rect 26546 10848 26562 10912
rect 26626 10848 26642 10912
rect 26706 10848 26714 10912
rect 26394 9824 26714 10848
rect 26394 9760 26402 9824
rect 26466 9760 26482 9824
rect 26546 9760 26562 9824
rect 26626 9760 26642 9824
rect 26706 9760 26714 9824
rect 26394 8736 26714 9760
rect 26394 8672 26402 8736
rect 26466 8672 26482 8736
rect 26546 8672 26562 8736
rect 26626 8672 26642 8736
rect 26706 8672 26714 8736
rect 26394 7648 26714 8672
rect 26394 7584 26402 7648
rect 26466 7584 26482 7648
rect 26546 7584 26562 7648
rect 26626 7584 26642 7648
rect 26706 7584 26714 7648
rect 26394 6560 26714 7584
rect 28766 6765 28826 29003
rect 28763 6764 28829 6765
rect 28763 6700 28764 6764
rect 28828 6700 28829 6764
rect 28763 6699 28829 6700
rect 26394 6496 26402 6560
rect 26466 6496 26482 6560
rect 26546 6496 26562 6560
rect 26626 6496 26642 6560
rect 26706 6496 26714 6560
rect 26394 6490 26714 6496
rect 26394 6254 26436 6490
rect 26672 6254 26714 6490
rect 26394 5472 26714 6254
rect 26394 5408 26402 5472
rect 26466 5408 26482 5472
rect 26546 5408 26562 5472
rect 26626 5408 26642 5472
rect 26706 5408 26714 5472
rect 26394 4384 26714 5408
rect 26394 4320 26402 4384
rect 26466 4320 26482 4384
rect 26546 4320 26562 4384
rect 26626 4320 26642 4384
rect 26706 4320 26714 4384
rect 26394 3296 26714 4320
rect 26394 3232 26402 3296
rect 26466 3232 26482 3296
rect 26546 3232 26562 3296
rect 26626 3232 26642 3296
rect 26706 3232 26714 3296
rect 26394 2208 26714 3232
rect 26394 2144 26402 2208
rect 26466 2144 26482 2208
rect 26546 2144 26562 2208
rect 26626 2144 26642 2208
rect 26706 2144 26714 2208
rect 26394 2128 26714 2144
<< via4 >>
rect 4527 26810 4763 27046
rect 4527 19738 4763 19974
rect 4527 12666 4763 12902
rect 4527 5594 4763 5830
rect 5187 27470 5423 27706
rect 5187 20398 5423 20634
rect 11610 26810 11846 27046
rect 11610 19738 11846 19974
rect 5187 13326 5423 13562
rect 11610 12666 11846 12902
rect 5187 6254 5423 6490
rect 11610 5594 11846 5830
rect 12270 27470 12506 27706
rect 12270 20398 12506 20634
rect 12270 13326 12506 13562
rect 12270 6254 12506 6490
rect 18693 26810 18929 27046
rect 18693 19738 18929 19974
rect 18693 12666 18929 12902
rect 18693 5594 18929 5830
rect 19353 27470 19589 27706
rect 25776 26810 26012 27046
rect 19353 20398 19589 20634
rect 19353 13326 19589 13562
rect 19353 6254 19589 6490
rect 25776 19738 26012 19974
rect 25776 12666 26012 12902
rect 25776 5594 26012 5830
rect 26436 27470 26672 27706
rect 26436 20398 26672 20634
rect 26436 13326 26672 13562
rect 26436 6254 26672 6490
<< metal5 >>
rect 1056 27706 29488 27748
rect 1056 27470 5187 27706
rect 5423 27470 12270 27706
rect 12506 27470 19353 27706
rect 19589 27470 26436 27706
rect 26672 27470 29488 27706
rect 1056 27428 29488 27470
rect 1056 27046 29488 27088
rect 1056 26810 4527 27046
rect 4763 26810 11610 27046
rect 11846 26810 18693 27046
rect 18929 26810 25776 27046
rect 26012 26810 29488 27046
rect 1056 26768 29488 26810
rect 1056 20634 29488 20676
rect 1056 20398 5187 20634
rect 5423 20398 12270 20634
rect 12506 20398 19353 20634
rect 19589 20398 26436 20634
rect 26672 20398 29488 20634
rect 1056 20356 29488 20398
rect 1056 19974 29488 20016
rect 1056 19738 4527 19974
rect 4763 19738 11610 19974
rect 11846 19738 18693 19974
rect 18929 19738 25776 19974
rect 26012 19738 29488 19974
rect 1056 19696 29488 19738
rect 1056 13562 29488 13604
rect 1056 13326 5187 13562
rect 5423 13326 12270 13562
rect 12506 13326 19353 13562
rect 19589 13326 26436 13562
rect 26672 13326 29488 13562
rect 1056 13284 29488 13326
rect 1056 12902 29488 12944
rect 1056 12666 4527 12902
rect 4763 12666 11610 12902
rect 11846 12666 18693 12902
rect 18929 12666 25776 12902
rect 26012 12666 29488 12902
rect 1056 12624 29488 12666
rect 1056 6490 29488 6532
rect 1056 6254 5187 6490
rect 5423 6254 12270 6490
rect 12506 6254 19353 6490
rect 19589 6254 26436 6490
rect 26672 6254 29488 6490
rect 1056 6212 29488 6254
rect 1056 5830 29488 5872
rect 1056 5594 4527 5830
rect 4763 5594 11610 5830
rect 11846 5594 18693 5830
rect 18929 5594 25776 5830
rect 26012 5594 29488 5830
rect 1056 5552 29488 5594
use sky130_fd_sc_hd__or4b_1  _0462_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0463_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0464_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0465_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0466_
timestamp 1688980957
transform 1 0 10212 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0467_
timestamp 1688980957
transform 1 0 21252 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0468_
timestamp 1688980957
transform 1 0 17296 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0469_
timestamp 1688980957
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0470_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0471_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0472_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22080 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_4  _0473_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__or4bb_4  _0474_
timestamp 1688980957
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_8  _0475_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  _0476_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _0477_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9936 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0478_
timestamp 1688980957
transform 1 0 10580 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _0479_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _0480_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0481_
timestamp 1688980957
transform 1 0 7544 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0482_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0483_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_4  _0484_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__nor3b_2  _0485_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0486_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0487_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13892 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand4b_4  _0488_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__or4b_1  _0489_
timestamp 1688980957
transform 1 0 22080 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0490_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23276 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_8  _0491_
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__nor3b_4  _0492_
timestamp 1688980957
transform 1 0 20148 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _0493_
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0494_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _0495_
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0496_
timestamp 1688980957
transform 1 0 14076 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0497_
timestamp 1688980957
transform 1 0 16928 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _0498_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_2  _0499_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0500_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _0501_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0502_
timestamp 1688980957
transform 1 0 5244 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0503_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0504_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0505_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0506_
timestamp 1688980957
transform 1 0 16376 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _0507_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0508_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0509_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0510_
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _0511_
timestamp 1688980957
transform 1 0 5520 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0512_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0513_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0514_
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0515_
timestamp 1688980957
transform 1 0 17572 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0516_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _0517_
timestamp 1688980957
transform 1 0 17112 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0518_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _0519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0520_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0521_
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _0522_
timestamp 1688980957
transform 1 0 6992 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0523_
timestamp 1688980957
transform 1 0 5336 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0524_
timestamp 1688980957
transform 1 0 4232 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0525_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0526_
timestamp 1688980957
transform 1 0 17664 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0527_
timestamp 1688980957
transform 1 0 16100 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _0528_
timestamp 1688980957
transform 1 0 16836 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0529_
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0530_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0531_
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0532_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0533_
timestamp 1688980957
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0534_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0535_
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0536_
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _0537_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__o21ai_1  _0538_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _0539_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0540_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0542_
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1688980957
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0544_
timestamp 1688980957
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0545_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0546_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0547_
timestamp 1688980957
transform 1 0 20056 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0548_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0549_
timestamp 1688980957
transform 1 0 8188 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0550_
timestamp 1688980957
transform 1 0 4416 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0551_
timestamp 1688980957
transform 1 0 4968 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0552_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0553_
timestamp 1688980957
transform 1 0 7084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0554_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6532 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0555_
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0556_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0557_
timestamp 1688980957
transform 1 0 5704 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0558_
timestamp 1688980957
transform 1 0 4968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0559_
timestamp 1688980957
transform 1 0 4692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0560_
timestamp 1688980957
transform 1 0 3864 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0561_
timestamp 1688980957
transform 1 0 4232 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1688980957
transform 1 0 3404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0563_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0564_
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0565_
timestamp 1688980957
transform 1 0 5244 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0566_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0568_
timestamp 1688980957
transform 1 0 7360 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0569_
timestamp 1688980957
transform 1 0 7084 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0570_
timestamp 1688980957
transform 1 0 7176 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1688980957
transform 1 0 6624 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0572_
timestamp 1688980957
transform 1 0 7636 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0573_
timestamp 1688980957
transform 1 0 8740 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0574_
timestamp 1688980957
transform 1 0 6900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0575_
timestamp 1688980957
transform 1 0 9476 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0576_
timestamp 1688980957
transform 1 0 10304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0577_
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0578_
timestamp 1688980957
transform 1 0 9936 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0579_
timestamp 1688980957
transform 1 0 11040 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0580_
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1688980957
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0582_
timestamp 1688980957
transform 1 0 10488 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0583_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0584_
timestamp 1688980957
transform 1 0 11960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0585_
timestamp 1688980957
transform 1 0 11316 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0586_
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0587_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0588_
timestamp 1688980957
transform 1 0 12972 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0589_
timestamp 1688980957
transform 1 0 14352 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0590_
timestamp 1688980957
transform 1 0 16008 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0591_
timestamp 1688980957
transform 1 0 15456 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0592_
timestamp 1688980957
transform 1 0 13156 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0593_
timestamp 1688980957
transform 1 0 14904 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0594_
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0595_
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0596_
timestamp 1688980957
transform 1 0 16100 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1688980957
transform 1 0 17296 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0598_
timestamp 1688980957
transform 1 0 16652 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0599_
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0600_
timestamp 1688980957
transform 1 0 18032 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0601_
timestamp 1688980957
transform 1 0 17112 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1688980957
transform 1 0 16192 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0603_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0604_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0605_
timestamp 1688980957
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0606_
timestamp 1688980957
transform 1 0 20792 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0607_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0608_
timestamp 1688980957
transform 1 0 22172 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0609_
timestamp 1688980957
transform 1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0610_
timestamp 1688980957
transform 1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0611_
timestamp 1688980957
transform 1 0 22448 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0612_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0613_
timestamp 1688980957
transform 1 0 20608 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0614_
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1688980957
transform 1 0 20608 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0616_
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0617_
timestamp 1688980957
transform 1 0 6992 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0618_
timestamp 1688980957
transform 1 0 15732 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0619_
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _0620_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1688980957
transform 1 0 6164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0622_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0623_
timestamp 1688980957
transform 1 0 5612 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0624_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0625_
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0626_
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0627_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0628_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0629_
timestamp 1688980957
transform 1 0 11408 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0630_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0631_
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0632_
timestamp 1688980957
transform 1 0 19320 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _0633_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_1  _0634_
timestamp 1688980957
transform 1 0 10396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0635_
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0636_
timestamp 1688980957
transform 1 0 17940 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0637_
timestamp 1688980957
transform 1 0 20240 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0638_
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0639_
timestamp 1688980957
transform 1 0 18584 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0640_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0641_
timestamp 1688980957
transform 1 0 7268 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0642_
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0643_
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0644_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _0645_
timestamp 1688980957
transform 1 0 18676 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _0646_
timestamp 1688980957
transform 1 0 21896 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1688980957
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0648_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0649_
timestamp 1688980957
transform 1 0 18492 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0650_
timestamp 1688980957
transform 1 0 20884 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0651_
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0652_
timestamp 1688980957
transform 1 0 25024 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0653_
timestamp 1688980957
transform 1 0 23092 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 1688980957
transform 1 0 22724 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _0655_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23276 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0656_
timestamp 1688980957
transform 1 0 23460 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0657_
timestamp 1688980957
transform 1 0 24932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0658_
timestamp 1688980957
transform 1 0 21252 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0659_
timestamp 1688980957
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0660_
timestamp 1688980957
transform 1 0 24564 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0661_
timestamp 1688980957
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0662_
timestamp 1688980957
transform 1 0 21712 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0663_
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0664_
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0665_
timestamp 1688980957
transform 1 0 23460 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0667_
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 1688980957
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0669_
timestamp 1688980957
transform 1 0 24840 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0671_
timestamp 1688980957
transform 1 0 24380 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1688980957
transform 1 0 21068 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0673_
timestamp 1688980957
transform 1 0 20792 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_4  _0675_
timestamp 1688980957
transform 1 0 19780 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__nand2b_4  _0676_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11684 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_8  _0677_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _0678_
timestamp 1688980957
transform 1 0 22080 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0679_
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  _0680_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23184 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _0681_
timestamp 1688980957
transform 1 0 16008 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0682_
timestamp 1688980957
transform 1 0 14996 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0683_
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0684_
timestamp 1688980957
transform 1 0 17296 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0685_
timestamp 1688980957
transform 1 0 18216 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0686_
timestamp 1688980957
transform 1 0 14904 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0687_
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0688_
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0689_
timestamp 1688980957
transform 1 0 15640 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0690_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0691_
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0692_
timestamp 1688980957
transform 1 0 17940 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0693_
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0694_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _0695_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _0696_
timestamp 1688980957
transform 1 0 10304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _0698_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0699_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0700_
timestamp 1688980957
transform 1 0 10212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0701_
timestamp 1688980957
transform 1 0 9384 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0702_
timestamp 1688980957
transform 1 0 8648 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0703_
timestamp 1688980957
transform 1 0 9016 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0704_
timestamp 1688980957
transform 1 0 4600 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0705_
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0706_
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0707_
timestamp 1688980957
transform 1 0 5244 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0708_
timestamp 1688980957
transform 1 0 5612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0709_
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0710_
timestamp 1688980957
transform 1 0 11500 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0711_
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0712_
timestamp 1688980957
transform 1 0 9844 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0713_
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0714_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0715_
timestamp 1688980957
transform 1 0 6716 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0716_
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0717_
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0718_
timestamp 1688980957
transform 1 0 12052 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0719_
timestamp 1688980957
transform 1 0 6164 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0720_
timestamp 1688980957
transform 1 0 6348 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0721_
timestamp 1688980957
transform 1 0 7268 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0722_
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0723_
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0724_
timestamp 1688980957
transform 1 0 6808 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0725_
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0726_
timestamp 1688980957
transform 1 0 7452 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0727_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0728_
timestamp 1688980957
transform 1 0 10856 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0729_
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0730_
timestamp 1688980957
transform 1 0 3956 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0731_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0732_
timestamp 1688980957
transform 1 0 12788 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0733_
timestamp 1688980957
transform 1 0 14352 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0734_
timestamp 1688980957
transform 1 0 4968 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0735_
timestamp 1688980957
transform 1 0 3312 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0736_
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0737_
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0738_
timestamp 1688980957
transform 1 0 4600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0739_
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0740_
timestamp 1688980957
transform 1 0 14812 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0741_
timestamp 1688980957
transform 1 0 5060 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1688980957
transform 1 0 11868 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0744_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0745_
timestamp 1688980957
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0746_
timestamp 1688980957
transform 1 0 3956 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0747_
timestamp 1688980957
transform 1 0 10028 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0748_
timestamp 1688980957
transform 1 0 12236 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0749_
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0750_
timestamp 1688980957
transform 1 0 3956 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0751_
timestamp 1688980957
transform 1 0 3128 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0752_
timestamp 1688980957
transform 1 0 6716 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0753_
timestamp 1688980957
transform 1 0 3312 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0754_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0755_
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0756_
timestamp 1688980957
transform 1 0 9844 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0757_
timestamp 1688980957
transform 1 0 3956 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0758_
timestamp 1688980957
transform 1 0 9844 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0759_
timestamp 1688980957
transform 1 0 11408 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0760_
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0761_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0762_
timestamp 1688980957
transform 1 0 20332 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1688980957
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0764_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24656 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0765_
timestamp 1688980957
transform 1 0 27232 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0766_
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0767_
timestamp 1688980957
transform 1 0 23460 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0768_
timestamp 1688980957
transform 1 0 20516 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0769_
timestamp 1688980957
transform 1 0 20056 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0770_
timestamp 1688980957
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0771_
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0772_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0773_
timestamp 1688980957
transform 1 0 21068 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0774_
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0775_
timestamp 1688980957
transform 1 0 23460 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0776_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _0777_
timestamp 1688980957
transform 1 0 24104 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0778_
timestamp 1688980957
transform 1 0 27508 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0779_
timestamp 1688980957
transform 1 0 27048 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0780_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 1688980957
transform 1 0 22724 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0782_
timestamp 1688980957
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0783_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0784_
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0786_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0787_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0788_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0789_
timestamp 1688980957
transform 1 0 25300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0790_
timestamp 1688980957
transform 1 0 27048 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0791_
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0792_
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0793_
timestamp 1688980957
transform 1 0 27600 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0794_
timestamp 1688980957
transform 1 0 27416 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0795_
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0796_
timestamp 1688980957
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0797_
timestamp 1688980957
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0798_
timestamp 1688980957
transform 1 0 28244 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0799_
timestamp 1688980957
transform 1 0 28336 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0800_
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0801_
timestamp 1688980957
transform 1 0 15548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0803_
timestamp 1688980957
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0804_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1688980957
transform 1 0 17480 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1688980957
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0807_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0808_
timestamp 1688980957
transform 1 0 16376 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _0809_
timestamp 1688980957
transform 1 0 18492 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0810_
timestamp 1688980957
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0811_
timestamp 1688980957
transform 1 0 16560 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0812_
timestamp 1688980957
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0813_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1688980957
transform 1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 1688980957
transform 1 0 16744 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0816_
timestamp 1688980957
transform 1 0 17848 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0817_
timestamp 1688980957
transform 1 0 16928 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0818_
timestamp 1688980957
transform 1 0 17204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0819_
timestamp 1688980957
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0820_
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0821_
timestamp 1688980957
transform 1 0 8372 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0822_
timestamp 1688980957
transform 1 0 14812 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0823_
timestamp 1688980957
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1688980957
transform 1 0 14352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0825_
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0826_
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0827_
timestamp 1688980957
transform 1 0 12880 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0828_
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0829_
timestamp 1688980957
transform 1 0 14812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0830_
timestamp 1688980957
transform 1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0831_
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 1688980957
transform 1 0 2208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1688980957
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0834_
timestamp 1688980957
transform 1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0835_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0836_
timestamp 1688980957
transform 1 0 13156 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _0838_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_2  _0839_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0840_
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0842_
timestamp 1688980957
transform 1 0 19688 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0843_
timestamp 1688980957
transform 1 0 19228 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0844_
timestamp 1688980957
transform 1 0 23552 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0845_
timestamp 1688980957
transform 1 0 22448 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_2  _0846_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0847_
timestamp 1688980957
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0848_
timestamp 1688980957
transform 1 0 17664 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _0849_
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0850_
timestamp 1688980957
transform 1 0 21620 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0851_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0852_
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0853_
timestamp 1688980957
transform 1 0 20700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _0854_
timestamp 1688980957
transform 1 0 15732 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1688980957
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0856_
timestamp 1688980957
transform 1 0 18768 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0857_
timestamp 1688980957
transform 1 0 18308 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0858_
timestamp 1688980957
transform 1 0 19044 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0859_
timestamp 1688980957
transform 1 0 18400 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0860_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0861_
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0862_
timestamp 1688980957
transform 1 0 19964 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0863_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0864_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0865_
timestamp 1688980957
transform 1 0 19780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0866_
timestamp 1688980957
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0867_
timestamp 1688980957
transform 1 0 23000 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0868_
timestamp 1688980957
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0870_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1688980957
transform 1 0 24932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0872_
timestamp 1688980957
transform 1 0 25392 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1688980957
transform 1 0 27416 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1688980957
transform 1 0 28244 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0875_
timestamp 1688980957
transform 1 0 23184 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0876_
timestamp 1688980957
transform 1 0 23092 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0877_
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0878_
timestamp 1688980957
transform 1 0 22816 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0879_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0880_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0881_
timestamp 1688980957
transform 1 0 23552 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0882_
timestamp 1688980957
transform 1 0 23276 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0883_
timestamp 1688980957
transform 1 0 23460 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0884_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0885_
timestamp 1688980957
transform 1 0 21712 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1688980957
transform 1 0 22816 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0890_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0891_
timestamp 1688980957
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0892_
timestamp 1688980957
transform 1 0 22356 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0893_
timestamp 1688980957
transform 1 0 23920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0895_
timestamp 1688980957
transform 1 0 23368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0896_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23368 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0897_
timestamp 1688980957
transform 1 0 24472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0898_
timestamp 1688980957
transform 1 0 23828 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0899_
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1688980957
transform 1 0 25852 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0901_
timestamp 1688980957
transform 1 0 24840 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0902_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0903_
timestamp 1688980957
transform 1 0 27232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0904_
timestamp 1688980957
transform 1 0 25576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0905_
timestamp 1688980957
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0906_
timestamp 1688980957
transform 1 0 28152 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0907_
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _0908_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0909_
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0910_
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0911_
timestamp 1688980957
transform 1 0 25484 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0912_
timestamp 1688980957
transform 1 0 25852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0913_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0914_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25392 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0915_
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0916_
timestamp 1688980957
transform 1 0 14168 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0917_
timestamp 1688980957
transform 1 0 15640 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0918_
timestamp 1688980957
transform 1 0 17572 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0919_
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0920_
timestamp 1688980957
transform 1 0 16376 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 1688980957
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0922_
timestamp 1688980957
transform 1 0 2576 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0923_
timestamp 1688980957
transform 1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1688980957
transform 1 0 3864 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0925_
timestamp 1688980957
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0926_
timestamp 1688980957
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0927_
timestamp 1688980957
transform 1 0 13892 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0928_
timestamp 1688980957
transform 1 0 13524 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0929_
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1688980957
transform 1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0931_
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0932_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0933_
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0934_
timestamp 1688980957
transform 1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0935_
timestamp 1688980957
transform 1 0 12972 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0936_
timestamp 1688980957
transform 1 0 13524 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0937_
timestamp 1688980957
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0938_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0939_
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0940_
timestamp 1688980957
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0941_
timestamp 1688980957
transform 1 0 26128 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1688980957
transform 1 0 22264 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0943_
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0944_
timestamp 1688980957
transform 1 0 22724 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0945_
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0946_
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0947_
timestamp 1688980957
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0948_
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1688980957
transform 1 0 26128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0950_
timestamp 1688980957
transform 1 0 25668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1688980957
transform 1 0 26680 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0952_
timestamp 1688980957
transform 1 0 26036 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0953_
timestamp 1688980957
transform 1 0 26496 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0954_
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0955_
timestamp 1688980957
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0956_
timestamp 1688980957
transform 1 0 26864 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0957_
timestamp 1688980957
transform 1 0 28152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0958_
timestamp 1688980957
transform 1 0 27232 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0959_
timestamp 1688980957
transform 1 0 27232 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0960_
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0961_
timestamp 1688980957
transform 1 0 26404 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1688980957
transform 1 0 27876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0963_
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 1688980957
transform 1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0965_
timestamp 1688980957
transform 1 0 27784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0966_
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0967_
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0968_
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0969_
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0970_
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0971_
timestamp 1688980957
transform 1 0 23644 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0972_
timestamp 1688980957
transform 1 0 18584 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 1688980957
transform 1 0 9016 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _0974_
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 1688980957
transform 1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0976_
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _0977_
timestamp 1688980957
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0978_
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0979_
timestamp 1688980957
transform 1 0 10304 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0980_
timestamp 1688980957
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1688980957
transform 1 0 10672 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0982_
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0983_
timestamp 1688980957
transform 1 0 8464 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0984_
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0985_
timestamp 1688980957
transform 1 0 21988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0986_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1688980957
transform 1 0 20792 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0988_
timestamp 1688980957
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0990_
timestamp 1688980957
transform 1 0 9200 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0991_
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0992_
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0993_
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0994_
timestamp 1688980957
transform 1 0 11224 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0995_
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0996_
timestamp 1688980957
transform 1 0 19320 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0997_
timestamp 1688980957
transform 1 0 17664 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0998_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0999_
timestamp 1688980957
transform 1 0 19780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1000_
timestamp 1688980957
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1001_
timestamp 1688980957
transform 1 0 17572 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1002_
timestamp 1688980957
transform 1 0 16928 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1688980957
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1004_
timestamp 1688980957
transform 1 0 15640 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1005_
timestamp 1688980957
transform 1 0 15640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1688980957
transform 1 0 15640 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1688980957
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1008_
timestamp 1688980957
transform 1 0 14904 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1009_
timestamp 1688980957
transform 1 0 15272 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1010_
timestamp 1688980957
transform 1 0 15088 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1688980957
transform 1 0 14720 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1012_
timestamp 1688980957
transform 1 0 14076 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1688980957
transform 1 0 12972 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1688980957
transform 1 0 11868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1016_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1017_
timestamp 1688980957
transform 1 0 16468 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1018_
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1019_
timestamp 1688980957
transform 1 0 1840 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1020_
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1021_
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1022_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1023_
timestamp 1688980957
transform 1 0 6992 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1024_
timestamp 1688980957
transform 1 0 3128 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1025_
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1026_
timestamp 1688980957
transform 1 0 4692 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1027_
timestamp 1688980957
transform 1 0 3220 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1028_
timestamp 1688980957
transform 1 0 3680 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1029_
timestamp 1688980957
transform 1 0 4324 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1030_
timestamp 1688980957
transform 1 0 6900 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1031_
timestamp 1688980957
transform 1 0 7636 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1032_
timestamp 1688980957
transform 1 0 7912 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1033_
timestamp 1688980957
transform 1 0 10396 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1034_
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1035_
timestamp 1688980957
transform 1 0 10764 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1036_
timestamp 1688980957
transform 1 0 12512 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1037_
timestamp 1688980957
transform 1 0 13432 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1038_
timestamp 1688980957
transform 1 0 13432 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1039_
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1040_
timestamp 1688980957
transform 1 0 16744 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1041_
timestamp 1688980957
transform 1 0 16468 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1042_
timestamp 1688980957
transform 1 0 18952 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1043_
timestamp 1688980957
transform 1 0 19872 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1044_
timestamp 1688980957
transform 1 0 22448 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1045_
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1046_
timestamp 1688980957
transform 1 0 19872 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1047_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1048_
timestamp 1688980957
transform 1 0 20516 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1049_
timestamp 1688980957
transform 1 0 22448 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1050_
timestamp 1688980957
transform 1 0 24932 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1051_
timestamp 1688980957
transform 1 0 26220 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1052_
timestamp 1688980957
transform 1 0 24932 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1053_
timestamp 1688980957
transform 1 0 14444 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1054_
timestamp 1688980957
transform 1 0 1564 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1055_
timestamp 1688980957
transform 1 0 1748 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1056_
timestamp 1688980957
transform 1 0 13248 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1057_
timestamp 1688980957
transform 1 0 13524 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1058_
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1059_
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1060_
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1061_
timestamp 1688980957
transform 1 0 24472 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1062_
timestamp 1688980957
transform 1 0 26772 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1063_
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1064_
timestamp 1688980957
transform 1 0 23460 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1065_
timestamp 1688980957
transform 1 0 24472 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1066_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1067_
timestamp 1688980957
transform 1 0 8648 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1068_
timestamp 1688980957
transform 1 0 6164 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1069_
timestamp 1688980957
transform 1 0 20056 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1070_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1071_
timestamp 1688980957
transform 1 0 8464 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1072_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1073_
timestamp 1688980957
transform 1 0 18768 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1074_
timestamp 1688980957
transform 1 0 18400 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1075_
timestamp 1688980957
transform 1 0 16376 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1076_
timestamp 1688980957
transform 1 0 14996 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1077_
timestamp 1688980957
transform 1 0 11592 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1078_
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1079_
timestamp 1688980957
transform 1 0 9568 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1080_
timestamp 1688980957
transform 1 0 9200 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1081_
timestamp 1688980957
transform 1 0 9016 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1082_
timestamp 1688980957
transform 1 0 1840 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1083_
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1084_
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1085_
timestamp 1688980957
transform 1 0 1840 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1086_
timestamp 1688980957
transform 1 0 2300 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1087_
timestamp 1688980957
transform 1 0 1656 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1088_
timestamp 1688980957
transform 1 0 9200 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1089_
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1090_
timestamp 1688980957
transform 1 0 9200 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1091_
timestamp 1688980957
transform 1 0 12144 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1092_
timestamp 1688980957
transform 1 0 12880 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1093_
timestamp 1688980957
transform 1 0 12144 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1094_
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 1688980957
transform 1 0 1840 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1096_
timestamp 1688980957
transform 1 0 7912 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 1688980957
transform 1 0 6624 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1098_
timestamp 1688980957
transform 1 0 1840 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1099_
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 1688980957
transform 1 0 12144 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 1688980957
transform 1 0 1840 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1688980957
transform 1 0 12144 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 1688980957
transform 1 0 12144 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1688980957
transform 1 0 10120 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1688980957
transform 1 0 11776 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1688980957
transform 1 0 5244 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 1688980957
transform 1 0 6992 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1688980957
transform 1 0 6532 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1688980957
transform 1 0 5428 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1688980957
transform 1 0 6256 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1688980957
transform 1 0 12052 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 1688980957
transform 1 0 11592 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1115_
timestamp 1688980957
transform 1 0 9568 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1116_
timestamp 1688980957
transform 1 0 9016 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1117_
timestamp 1688980957
transform 1 0 9292 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1688980957
transform 1 0 3680 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1688980957
transform 1 0 3772 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 1688980957
transform 1 0 4232 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 1688980957
transform 1 0 5152 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1124_
timestamp 1688980957
transform 1 0 9200 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1688980957
transform 1 0 9200 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1688980957
transform 1 0 14720 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1688980957
transform 1 0 16560 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1688980957
transform 1 0 17296 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1131_
timestamp 1688980957
transform 1 0 14168 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1132_
timestamp 1688980957
transform 1 0 17020 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1133_
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1688980957
transform 1 0 14720 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1688980957
transform 1 0 14444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1139_
timestamp 1688980957
transform 1 0 19872 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1140_
timestamp 1688980957
transform 1 0 18032 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1141_
timestamp 1688980957
transform 1 0 19964 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1142_
timestamp 1688980957
transform 1 0 22816 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform 1 0 9936 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 11040 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 10396 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform 1 0 10856 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 18216 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform 1 0 21988 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 22632 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 15364 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform 1 0 14536 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 19596 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout35
timestamp 1688980957
transform 1 0 7820 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout36
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout37
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp 1688980957
transform 1 0 14628 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout39
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout40
timestamp 1688980957
transform 1 0 27968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout41
timestamp 1688980957
transform 1 0 24288 0 -1 29376
box -38 -48 866 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_35
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_47 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_72
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_119
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_131
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_156
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_203
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_225 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_233
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_245
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_265 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_275
timestamp 1688980957
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_147
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_159
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_187
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_199
timestamp 1688980957
transform 1 0 19412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_211
timestamp 1688980957
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_9
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_135
timestamp 1688980957
transform 1 0 13524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_158
timestamp 1688980957
transform 1 0 15640 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_174
timestamp 1688980957
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_261
timestamp 1688980957
transform 1 0 25116 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_11
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_147
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_155
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1688980957
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_184
timestamp 1688980957
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_188
timestamp 1688980957
transform 1 0 18400 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_209
timestamp 1688980957
transform 1 0 20332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_221
timestamp 1688980957
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_254
timestamp 1688980957
transform 1 0 24472 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_260
timestamp 1688980957
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_272
timestamp 1688980957
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_113
timestamp 1688980957
transform 1 0 11500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_125
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_134
timestamp 1688980957
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_187
timestamp 1688980957
transform 1 0 18308 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_214
timestamp 1688980957
transform 1 0 20792 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_226
timestamp 1688980957
transform 1 0 21896 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_238
timestamp 1688980957
transform 1 0 23000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_77
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1688980957
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_134
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_146
timestamp 1688980957
transform 1 0 14536 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_158
timestamp 1688980957
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 1688980957
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_197
timestamp 1688980957
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_211
timestamp 1688980957
transform 1 0 20516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_296
timestamp 1688980957
transform 1 0 28336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_304
timestamp 1688980957
transform 1 0 29072 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_51
timestamp 1688980957
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_55
timestamp 1688980957
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 1688980957
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_117
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_50
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_84
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_119
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_131
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_157
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_176
timestamp 1688980957
transform 1 0 17296 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_188
timestamp 1688980957
transform 1 0 18400 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_200
timestamp 1688980957
transform 1 0 19504 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_218
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_44
timestamp 1688980957
transform 1 0 5152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_60
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_76
timestamp 1688980957
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_122
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_134
timestamp 1688980957
transform 1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_147
timestamp 1688980957
transform 1 0 14628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_159
timestamp 1688980957
transform 1 0 15732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_185
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_231
timestamp 1688980957
transform 1 0 22356 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_256
timestamp 1688980957
transform 1 0 24656 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_268
timestamp 1688980957
transform 1 0 25760 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_280
timestamp 1688980957
transform 1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_292
timestamp 1688980957
transform 1 0 27968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_304
timestamp 1688980957
transform 1 0 29072 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_47
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_99
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_122
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_128
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_158
timestamp 1688980957
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_189
timestamp 1688980957
transform 1 0 18492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_201
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_213
timestamp 1688980957
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_257
timestamp 1688980957
transform 1 0 24748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_290
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_298
timestamp 1688980957
transform 1 0 28520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1688980957
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_45
timestamp 1688980957
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_70
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_149
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_161
timestamp 1688980957
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_190
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_205
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_263
timestamp 1688980957
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_274
timestamp 1688980957
transform 1 0 26312 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_291
timestamp 1688980957
transform 1 0 27876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_303
timestamp 1688980957
transform 1 0 28980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_38
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_64
timestamp 1688980957
transform 1 0 6992 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_75
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_99
timestamp 1688980957
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_129
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_165
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_183
timestamp 1688980957
transform 1 0 17940 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_191
timestamp 1688980957
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_213
timestamp 1688980957
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_218
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_233
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_241
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_251
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_263
timestamp 1688980957
transform 1 0 25300 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_291
timestamp 1688980957
transform 1 0 27876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_303
timestamp 1688980957
transform 1 0 28980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_42
timestamp 1688980957
transform 1 0 4968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1688980957
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_120
timestamp 1688980957
transform 1 0 12144 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_128
timestamp 1688980957
transform 1 0 12880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_132
timestamp 1688980957
transform 1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_145
timestamp 1688980957
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_154
timestamp 1688980957
transform 1 0 15272 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_166
timestamp 1688980957
transform 1 0 16376 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_178
timestamp 1688980957
transform 1 0 17480 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_182
timestamp 1688980957
transform 1 0 17848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_190
timestamp 1688980957
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_205
timestamp 1688980957
transform 1 0 19964 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_217
timestamp 1688980957
transform 1 0 21068 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_223
timestamp 1688980957
transform 1 0 21620 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_239
timestamp 1688980957
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_299
timestamp 1688980957
transform 1 0 28612 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_67
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_79
timestamp 1688980957
transform 1 0 8372 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_155
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_176
timestamp 1688980957
transform 1 0 17296 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_195
timestamp 1688980957
transform 1 0 19044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_207
timestamp 1688980957
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_219
timestamp 1688980957
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 1688980957
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_296
timestamp 1688980957
transform 1 0 28336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_304
timestamp 1688980957
transform 1 0 29072 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_40
timestamp 1688980957
transform 1 0 4784 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_52
timestamp 1688980957
transform 1 0 5888 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_64
timestamp 1688980957
transform 1 0 6992 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_76
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_113
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_144
timestamp 1688980957
transform 1 0 14352 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_152
timestamp 1688980957
transform 1 0 15088 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_163
timestamp 1688980957
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_167
timestamp 1688980957
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_215
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_227
timestamp 1688980957
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_242
timestamp 1688980957
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1688980957
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_273
timestamp 1688980957
transform 1 0 26220 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_285
timestamp 1688980957
transform 1 0 27324 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_297
timestamp 1688980957
transform 1 0 28428 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_36
timestamp 1688980957
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_45
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_63
timestamp 1688980957
transform 1 0 6900 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_75
timestamp 1688980957
transform 1 0 8004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_87
timestamp 1688980957
transform 1 0 9108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_133
timestamp 1688980957
transform 1 0 13340 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_188
timestamp 1688980957
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 1688980957
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_259
timestamp 1688980957
transform 1 0 24932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_263
timestamp 1688980957
transform 1 0 25300 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_7
timestamp 1688980957
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_44
timestamp 1688980957
transform 1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_74
timestamp 1688980957
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_107
timestamp 1688980957
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_119
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 1688980957
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_157
timestamp 1688980957
transform 1 0 15548 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_185
timestamp 1688980957
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_288
timestamp 1688980957
transform 1 0 27600 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_296
timestamp 1688980957
transform 1 0 28336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1688980957
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_67
timestamp 1688980957
transform 1 0 7268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_78
timestamp 1688980957
transform 1 0 8280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_144
timestamp 1688980957
transform 1 0 14352 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_156
timestamp 1688980957
transform 1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_160
timestamp 1688980957
transform 1 0 15824 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_180
timestamp 1688980957
transform 1 0 17664 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_186
timestamp 1688980957
transform 1 0 18216 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_218
timestamp 1688980957
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_255
timestamp 1688980957
transform 1 0 24564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_263
timestamp 1688980957
transform 1 0 25300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_272
timestamp 1688980957
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_33
timestamp 1688980957
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_75
timestamp 1688980957
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_119
timestamp 1688980957
transform 1 0 12052 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_156
timestamp 1688980957
transform 1 0 15456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_160
timestamp 1688980957
transform 1 0 15824 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_174
timestamp 1688980957
transform 1 0 17112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_186
timestamp 1688980957
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_206
timestamp 1688980957
transform 1 0 20056 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_218
timestamp 1688980957
transform 1 0 21160 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_230
timestamp 1688980957
transform 1 0 22264 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_35
timestamp 1688980957
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_76
timestamp 1688980957
transform 1 0 8096 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_108
timestamp 1688980957
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_132
timestamp 1688980957
transform 1 0 13248 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_176
timestamp 1688980957
transform 1 0 17296 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_207
timestamp 1688980957
transform 1 0 20148 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_215
timestamp 1688980957
transform 1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_243
timestamp 1688980957
transform 1 0 23460 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_255
timestamp 1688980957
transform 1 0 24564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_267
timestamp 1688980957
transform 1 0 25668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_11
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_66
timestamp 1688980957
transform 1 0 7176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_100
timestamp 1688980957
transform 1 0 10304 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_120
timestamp 1688980957
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_203
timestamp 1688980957
transform 1 0 19780 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_215
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_223
timestamp 1688980957
transform 1 0 21620 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_227
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_247
timestamp 1688980957
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_269
timestamp 1688980957
transform 1 0 25852 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_281
timestamp 1688980957
transform 1 0 26956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_293
timestamp 1688980957
transform 1 0 28060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_28
timestamp 1688980957
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_40
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_52
timestamp 1688980957
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_64
timestamp 1688980957
transform 1 0 6992 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_76
timestamp 1688980957
transform 1 0 8096 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_88
timestamp 1688980957
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_94
timestamp 1688980957
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_102
timestamp 1688980957
transform 1 0 10488 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_146
timestamp 1688980957
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_157
timestamp 1688980957
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1688980957
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_187
timestamp 1688980957
transform 1 0 18308 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_212
timestamp 1688980957
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_216
timestamp 1688980957
transform 1 0 20976 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_233
timestamp 1688980957
transform 1 0 22540 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_253
timestamp 1688980957
transform 1 0 24380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_274
timestamp 1688980957
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_289
timestamp 1688980957
transform 1 0 27692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_304
timestamp 1688980957
transform 1 0 29072 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_113
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_150
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_171
timestamp 1688980957
transform 1 0 16836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_183
timestamp 1688980957
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_216
timestamp 1688980957
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_240
timestamp 1688980957
transform 1 0 23184 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_302
timestamp 1688980957
transform 1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_31
timestamp 1688980957
transform 1 0 3956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 1688980957
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_87
timestamp 1688980957
transform 1 0 9108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 1688980957
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_140
timestamp 1688980957
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_144
timestamp 1688980957
transform 1 0 14352 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_203
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_234
timestamp 1688980957
transform 1 0 22632 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_250
timestamp 1688980957
transform 1 0 24104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_262
timestamp 1688980957
transform 1 0 25208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_7
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_33
timestamp 1688980957
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_54
timestamp 1688980957
transform 1 0 6072 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_80
timestamp 1688980957
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_108
timestamp 1688980957
transform 1 0 11040 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_116
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_164
timestamp 1688980957
transform 1 0 16192 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_208
timestamp 1688980957
transform 1 0 20240 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_220
timestamp 1688980957
transform 1 0 21344 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_232
timestamp 1688980957
transform 1 0 22448 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_238
timestamp 1688980957
transform 1 0 23000 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_287
timestamp 1688980957
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_299
timestamp 1688980957
transform 1 0 28612 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_6
timestamp 1688980957
transform 1 0 1656 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_14
timestamp 1688980957
transform 1 0 2392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_43
timestamp 1688980957
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_47
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_72
timestamp 1688980957
transform 1 0 7728 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_90
timestamp 1688980957
transform 1 0 9384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_94
timestamp 1688980957
transform 1 0 9752 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1688980957
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_121
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_136
timestamp 1688980957
transform 1 0 13616 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_148
timestamp 1688980957
transform 1 0 14720 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1688980957
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_246
timestamp 1688980957
transform 1 0 23736 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_258
timestamp 1688980957
transform 1 0 24840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_266
timestamp 1688980957
transform 1 0 25576 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_270
timestamp 1688980957
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_278
timestamp 1688980957
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_23
timestamp 1688980957
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_37
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_57
timestamp 1688980957
transform 1 0 6348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_69
timestamp 1688980957
transform 1 0 7452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_102
timestamp 1688980957
transform 1 0 10488 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_111
timestamp 1688980957
transform 1 0 11316 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_123
timestamp 1688980957
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_135
timestamp 1688980957
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_148
timestamp 1688980957
transform 1 0 14720 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_157
timestamp 1688980957
transform 1 0 15548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_169
timestamp 1688980957
transform 1 0 16652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_181
timestamp 1688980957
transform 1 0 17756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_248
timestamp 1688980957
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_262
timestamp 1688980957
transform 1 0 25208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_268
timestamp 1688980957
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_283
timestamp 1688980957
transform 1 0 27140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_297
timestamp 1688980957
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_23
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1688980957
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_89
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 1688980957
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_148
timestamp 1688980957
transform 1 0 14720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_158
timestamp 1688980957
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_177
timestamp 1688980957
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_198
timestamp 1688980957
transform 1 0 19320 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_210
timestamp 1688980957
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_234
timestamp 1688980957
transform 1 0 22632 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_300
timestamp 1688980957
transform 1 0 28704 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_304
timestamp 1688980957
transform 1 0 29072 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_43
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_72
timestamp 1688980957
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_91
timestamp 1688980957
transform 1 0 9476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_170
timestamp 1688980957
transform 1 0 16744 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_204
timestamp 1688980957
transform 1 0 19872 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_227
timestamp 1688980957
transform 1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_239
timestamp 1688980957
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1688980957
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_284
timestamp 1688980957
transform 1 0 27232 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_297
timestamp 1688980957
transform 1 0 28428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_7
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_48
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_78
timestamp 1688980957
transform 1 0 8280 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_121
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_141
timestamp 1688980957
transform 1 0 14076 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_147
timestamp 1688980957
transform 1 0 14628 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_218
timestamp 1688980957
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_268
timestamp 1688980957
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_304
timestamp 1688980957
transform 1 0 29072 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_40
timestamp 1688980957
transform 1 0 4784 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_52
timestamp 1688980957
transform 1 0 5888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_62
timestamp 1688980957
transform 1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_118
timestamp 1688980957
transform 1 0 11960 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_128
timestamp 1688980957
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_184
timestamp 1688980957
transform 1 0 18032 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_9
timestamp 1688980957
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_21
timestamp 1688980957
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_33
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_45
timestamp 1688980957
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_94
timestamp 1688980957
transform 1 0 9752 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_106
timestamp 1688980957
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_121
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_134
timestamp 1688980957
transform 1 0 13432 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_146
timestamp 1688980957
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_157
timestamp 1688980957
transform 1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_176
timestamp 1688980957
transform 1 0 17296 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_188
timestamp 1688980957
transform 1 0 18400 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_212
timestamp 1688980957
transform 1 0 20608 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_285
timestamp 1688980957
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_291
timestamp 1688980957
transform 1 0 27876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_303
timestamp 1688980957
transform 1 0 28980 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_37
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_49
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_72
timestamp 1688980957
transform 1 0 7728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_93
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_110
timestamp 1688980957
transform 1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_118
timestamp 1688980957
transform 1 0 11960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_126
timestamp 1688980957
transform 1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1688980957
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_164
timestamp 1688980957
transform 1 0 16192 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_176
timestamp 1688980957
transform 1 0 17296 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_188
timestamp 1688980957
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_281
timestamp 1688980957
transform 1 0 26956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_297
timestamp 1688980957
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_23
timestamp 1688980957
transform 1 0 3220 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_40
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_52
timestamp 1688980957
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_85
timestamp 1688980957
transform 1 0 8924 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_151
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp 1688980957
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_189
timestamp 1688980957
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_203
timestamp 1688980957
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_215
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_230
timestamp 1688980957
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_234
timestamp 1688980957
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_240
timestamp 1688980957
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1688980957
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1688980957
transform 1 0 25484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_303
timestamp 1688980957
transform 1 0 28980 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_49
timestamp 1688980957
transform 1 0 5612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_61
timestamp 1688980957
transform 1 0 6716 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_75
timestamp 1688980957
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_99
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_157
timestamp 1688980957
transform 1 0 15548 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_224
timestamp 1688980957
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_273
timestamp 1688980957
transform 1 0 26220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_300
timestamp 1688980957
transform 1 0 28704 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_304
timestamp 1688980957
transform 1 0 29072 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_21
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_84
timestamp 1688980957
transform 1 0 8832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1688980957
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_127
timestamp 1688980957
transform 1 0 12788 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_148
timestamp 1688980957
transform 1 0 14720 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_160
timestamp 1688980957
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_201
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_266
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1688980957
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_284
timestamp 1688980957
transform 1 0 27232 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_290
timestamp 1688980957
transform 1 0 27784 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_302
timestamp 1688980957
transform 1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_40
timestamp 1688980957
transform 1 0 4784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_44
timestamp 1688980957
transform 1 0 5152 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_173
timestamp 1688980957
transform 1 0 17020 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_183
timestamp 1688980957
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_205
timestamp 1688980957
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_215
timestamp 1688980957
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_271
timestamp 1688980957
transform 1 0 26036 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_283
timestamp 1688980957
transform 1 0 27140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_295
timestamp 1688980957
transform 1 0 28244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_303
timestamp 1688980957
transform 1 0 28980 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_35
timestamp 1688980957
transform 1 0 4324 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_44
timestamp 1688980957
transform 1 0 5152 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_68
timestamp 1688980957
transform 1 0 7360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_78
timestamp 1688980957
transform 1 0 8280 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1688980957
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_128
timestamp 1688980957
transform 1 0 12880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_140
timestamp 1688980957
transform 1 0 13984 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_148
timestamp 1688980957
transform 1 0 14720 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1688980957
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_177
timestamp 1688980957
transform 1 0 17388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_189
timestamp 1688980957
transform 1 0 18492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_201
timestamp 1688980957
transform 1 0 19596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_209
timestamp 1688980957
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_216
timestamp 1688980957
transform 1 0 20976 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_228
timestamp 1688980957
transform 1 0 22080 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_234
timestamp 1688980957
transform 1 0 22632 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_238
timestamp 1688980957
transform 1 0 23000 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_242
timestamp 1688980957
transform 1 0 23368 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_265
timestamp 1688980957
transform 1 0 25484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_35
timestamp 1688980957
transform 1 0 4324 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_44
timestamp 1688980957
transform 1 0 5152 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_52
timestamp 1688980957
transform 1 0 5888 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_64
timestamp 1688980957
transform 1 0 6992 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_76
timestamp 1688980957
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_117
timestamp 1688980957
transform 1 0 11868 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_129
timestamp 1688980957
transform 1 0 12972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1688980957
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_163
timestamp 1688980957
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_175
timestamp 1688980957
transform 1 0 17204 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_182
timestamp 1688980957
transform 1 0 17848 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_220
timestamp 1688980957
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_232
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1688980957
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_263
timestamp 1688980957
transform 1 0 25300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_275
timestamp 1688980957
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_287
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_299
timestamp 1688980957
transform 1 0 28612 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_9
timestamp 1688980957
transform 1 0 1932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_21
timestamp 1688980957
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_33
timestamp 1688980957
transform 1 0 4140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_45
timestamp 1688980957
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_53
timestamp 1688980957
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_87
timestamp 1688980957
transform 1 0 9108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_108
timestamp 1688980957
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_121
timestamp 1688980957
transform 1 0 12236 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_138
timestamp 1688980957
transform 1 0 13800 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_164
timestamp 1688980957
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_186
timestamp 1688980957
transform 1 0 18216 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_198
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_210
timestamp 1688980957
transform 1 0 20424 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1688980957
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_35
timestamp 1688980957
transform 1 0 4324 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_43
timestamp 1688980957
transform 1 0 5060 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_68
timestamp 1688980957
transform 1 0 7360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_80
timestamp 1688980957
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_104
timestamp 1688980957
transform 1 0 10672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_112
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_145
timestamp 1688980957
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_157
timestamp 1688980957
transform 1 0 15548 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_207
timestamp 1688980957
transform 1 0 20148 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_219
timestamp 1688980957
transform 1 0 21252 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_231
timestamp 1688980957
transform 1 0 22356 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_243
timestamp 1688980957
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_21
timestamp 1688980957
transform 1 0 3036 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_47
timestamp 1688980957
transform 1 0 5428 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_72
timestamp 1688980957
transform 1 0 7728 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_100
timestamp 1688980957
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_136
timestamp 1688980957
transform 1 0 13616 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_148
timestamp 1688980957
transform 1 0 14720 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_166
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_174
timestamp 1688980957
transform 1 0 17112 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_220
timestamp 1688980957
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_7
timestamp 1688980957
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_35
timestamp 1688980957
transform 1 0 4324 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_120
timestamp 1688980957
transform 1 0 12144 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_132
timestamp 1688980957
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_149
timestamp 1688980957
transform 1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_235
timestamp 1688980957
transform 1 0 22724 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_247
timestamp 1688980957
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_80
timestamp 1688980957
transform 1 0 8464 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_92
timestamp 1688980957
transform 1 0 9568 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_104
timestamp 1688980957
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_189
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_212
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_11
timestamp 1688980957
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_49
timestamp 1688980957
transform 1 0 5612 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_63
timestamp 1688980957
transform 1 0 6900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_75
timestamp 1688980957
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_125
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_137
timestamp 1688980957
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_202
timestamp 1688980957
transform 1 0 19688 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_214
timestamp 1688980957
transform 1 0 20792 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_226
timestamp 1688980957
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_238
timestamp 1688980957
transform 1 0 23000 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_250
timestamp 1688980957
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_73
timestamp 1688980957
transform 1 0 7820 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_94
timestamp 1688980957
transform 1 0 9752 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_106
timestamp 1688980957
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_119
timestamp 1688980957
transform 1 0 12052 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_123
timestamp 1688980957
transform 1 0 12420 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_148
timestamp 1688980957
transform 1 0 14720 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_160
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_173
timestamp 1688980957
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_180
timestamp 1688980957
transform 1 0 17664 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_192
timestamp 1688980957
transform 1 0 18768 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_204
timestamp 1688980957
transform 1 0 19872 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_212
timestamp 1688980957
transform 1 0 20608 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_219
timestamp 1688980957
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_9
timestamp 1688980957
transform 1 0 1932 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_25
timestamp 1688980957
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_33
timestamp 1688980957
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_42
timestamp 1688980957
transform 1 0 4968 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_54
timestamp 1688980957
transform 1 0 6072 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_66
timestamp 1688980957
transform 1 0 7176 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_91
timestamp 1688980957
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_103
timestamp 1688980957
transform 1 0 10580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_130
timestamp 1688980957
transform 1 0 13064 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_150
timestamp 1688980957
transform 1 0 14904 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_162
timestamp 1688980957
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_187
timestamp 1688980957
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_201
timestamp 1688980957
transform 1 0 19596 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_228
timestamp 1688980957
transform 1 0 22080 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1688980957
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_301
timestamp 1688980957
transform 1 0 28796 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_23
timestamp 1688980957
transform 1 0 3220 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_54
timestamp 1688980957
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_68
timestamp 1688980957
transform 1 0 7360 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_96
timestamp 1688980957
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_120
timestamp 1688980957
transform 1 0 12144 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_128
timestamp 1688980957
transform 1 0 12880 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_165
timestamp 1688980957
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_191
timestamp 1688980957
transform 1 0 18676 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_257
timestamp 1688980957
transform 1 0 24748 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_269
timestamp 1688980957
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_277
timestamp 1688980957
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_62
timestamp 1688980957
transform 1 0 6808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_95
timestamp 1688980957
transform 1 0 9844 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_126
timestamp 1688980957
transform 1 0 12696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_130
timestamp 1688980957
transform 1 0 13064 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_149
timestamp 1688980957
transform 1 0 14812 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_161
timestamp 1688980957
transform 1 0 15916 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_190
timestamp 1688980957
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_201
timestamp 1688980957
transform 1 0 19596 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_270
timestamp 1688980957
transform 1 0 25944 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_282
timestamp 1688980957
transform 1 0 27048 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_294
timestamp 1688980957
transform 1 0 28152 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_302
timestamp 1688980957
transform 1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_87
timestamp 1688980957
transform 1 0 9108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_99
timestamp 1688980957
transform 1 0 10212 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_133
timestamp 1688980957
transform 1 0 13340 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_162
timestamp 1688980957
transform 1 0 16008 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_197
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_203
timestamp 1688980957
transform 1 0 19780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_231
timestamp 1688980957
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_250
timestamp 1688980957
transform 1 0 24104 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_44
timestamp 1688980957
transform 1 0 5152 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_52
timestamp 1688980957
transform 1 0 5888 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_64
timestamp 1688980957
transform 1 0 6992 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_73
timestamp 1688980957
transform 1 0 7820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 1688980957
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_94
timestamp 1688980957
transform 1 0 9752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_106
timestamp 1688980957
transform 1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_117
timestamp 1688980957
transform 1 0 11868 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_129
timestamp 1688980957
transform 1 0 12972 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_137
timestamp 1688980957
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_156
timestamp 1688980957
transform 1 0 15456 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_168
timestamp 1688980957
transform 1 0 16560 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_179
timestamp 1688980957
transform 1 0 17572 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_191
timestamp 1688980957
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_215
timestamp 1688980957
transform 1 0 20884 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_227
timestamp 1688980957
transform 1 0 21988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_239
timestamp 1688980957
transform 1 0 23092 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_248
timestamp 1688980957
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_6
timestamp 1688980957
transform 1 0 1656 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_14
timestamp 1688980957
transform 1 0 2392 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_23
timestamp 1688980957
transform 1 0 3220 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_29
timestamp 1688980957
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_41
timestamp 1688980957
transform 1 0 4876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_53
timestamp 1688980957
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_77
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_83
timestamp 1688980957
transform 1 0 8740 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_85
timestamp 1688980957
transform 1 0 8924 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_100
timestamp 1688980957
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_147
timestamp 1688980957
transform 1 0 14628 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_159
timestamp 1688980957
transform 1 0 15732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_177
timestamp 1688980957
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_184
timestamp 1688980957
transform 1 0 18032 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_197
timestamp 1688980957
transform 1 0 19228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_209
timestamp 1688980957
transform 1 0 20332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_221
timestamp 1688980957
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_231
timestamp 1688980957
transform 1 0 22356 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_243
timestamp 1688980957
transform 1 0 23460 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_251
timestamp 1688980957
transform 1 0 24196 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_253
timestamp 1688980957
transform 1 0 24380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_268
timestamp 1688980957
transform 1 0 25760 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 2668 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 16192 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 16928 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 7544 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 14996 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 8188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 4048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 13340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 8648 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 7544 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 13616 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 7544 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 14996 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 4416 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 8096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 12880 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 9476 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 17204 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 4232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 4416 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 4324 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 5612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 9936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 4048 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 4416 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 15272 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 15272 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 3864 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 9568 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 18492 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 25116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform 1 0 9108 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 8096 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 6164 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 5060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 23368 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 25208 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 26496 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 14536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 25392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 26864 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform 1 0 23092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 25024 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 28336 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap33
timestamp 1688980957
transform 1 0 8280 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap34
timestamp 1688980957
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1688980957
transform 1 0 9752 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1688980957
transform -1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1688980957
transform 1 0 28612 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1688980957
transform 1 0 17480 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1688980957
transform 1 0 28796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1688980957
transform 1 0 25208 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 6532 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1688980957
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform 1 0 2668 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform 1 0 28612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1688980957
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform 1 0 28612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 14076 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 29440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 29440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 29440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 29440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 29440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 29440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 29440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 29440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 29440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 29440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 29440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 29440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 29440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 29440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 29440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 29440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 29440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 29440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 29440 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 29440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 29440 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 29440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 29440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 29440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 29440 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 29440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 29440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 29440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 29440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 29440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 29440 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 29440 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 29440 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 29440 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 29440 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 29440 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 29440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 29440 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 29440 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 29440 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 29440 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 29440 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 29440 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 29440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 29440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 3680 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
<< labels >>
flabel metal4 s 5145 2128 5465 30512 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12228 2128 12548 30512 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19311 2128 19631 30512 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 26394 2128 26714 30512 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6212 29488 6532 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13284 29488 13604 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 20356 29488 20676 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 27428 29488 27748 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4485 2128 4805 30512 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11568 2128 11888 30512 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 18651 2128 18971 30512 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 25734 2128 26054 30512 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5552 29488 5872 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12624 29488 12944 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 19696 29488 20016 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 26768 29488 27088 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 28998 31925 29054 32725 0 FreeSans 224 90 0 0 nrst
port 3 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 out_0[0]
port 4 nsew signal tristate
flabel metal2 s 9678 31925 9734 32725 0 FreeSans 224 90 0 0 out_0[1]
port 5 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 out_0[2]
port 6 nsew signal tristate
flabel metal3 s 29781 10888 30581 11008 0 FreeSans 480 0 0 0 out_0[3]
port 7 nsew signal tristate
flabel metal2 s 17406 31925 17462 32725 0 FreeSans 224 90 0 0 out_0[4]
port 8 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 out_0[5]
port 9 nsew signal tristate
flabel metal3 s 29781 18368 30581 18488 0 FreeSans 480 0 0 0 out_0[6]
port 10 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 out_1[0]
port 11 nsew signal tristate
flabel metal3 s 29781 22448 30581 22568 0 FreeSans 480 0 0 0 out_1[1]
port 12 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 out_1[2]
port 13 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 out_1[3]
port 14 nsew signal tristate
flabel metal2 s 21270 31925 21326 32725 0 FreeSans 224 90 0 0 out_1[4]
port 15 nsew signal tristate
flabel metal2 s 25134 31925 25190 32725 0 FreeSans 224 90 0 0 out_1[5]
port 16 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 out_1[6]
port 17 nsew signal tristate
flabel metal2 s 6458 31925 6514 32725 0 FreeSans 224 90 0 0 out_2[0]
port 18 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 out_2[1]
port 19 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 out_2[2]
port 20 nsew signal tristate
flabel metal3 s 29781 2728 30581 2848 0 FreeSans 480 0 0 0 out_2[3]
port 21 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 out_2[4]
port 22 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 out_2[5]
port 23 nsew signal tristate
flabel metal2 s 2594 31925 2650 32725 0 FreeSans 224 90 0 0 out_2[6]
port 24 nsew signal tristate
flabel metal3 s 29781 6808 30581 6928 0 FreeSans 480 0 0 0 out_3[0]
port 25 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 out_3[1]
port 26 nsew signal tristate
flabel metal3 s 29781 26528 30581 26648 0 FreeSans 480 0 0 0 out_3[2]
port 27 nsew signal tristate
flabel metal3 s 29781 30608 30581 30728 0 FreeSans 480 0 0 0 out_3[3]
port 28 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 out_3[4]
port 29 nsew signal tristate
flabel metal2 s 13542 31925 13598 32725 0 FreeSans 224 90 0 0 out_3[5]
port 30 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 out_3[6]
port 31 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 pb_0
port 32 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 pb_1
port 33 nsew signal input
flabel metal3 s 29781 14288 30581 14408 0 FreeSans 480 0 0 0 time_done
port 34 nsew signal tristate
rlabel metal1 15272 30464 15272 30464 0 VGND
rlabel metal1 15272 29920 15272 29920 0 VPWR
rlabel metal1 7590 25738 7590 25738 0 CLKDIV.count\[0\]
rlabel metal2 11730 28254 11730 28254 0 CLKDIV.count\[10\]
rlabel metal2 13294 29444 13294 29444 0 CLKDIV.count\[11\]
rlabel metal1 12052 27506 12052 27506 0 CLKDIV.count\[12\]
rlabel metal1 13202 27506 13202 27506 0 CLKDIV.count\[13\]
rlabel metal1 14398 27846 14398 27846 0 CLKDIV.count\[14\]
rlabel metal2 15502 28016 15502 28016 0 CLKDIV.count\[15\]
rlabel metal2 18354 28458 18354 28458 0 CLKDIV.count\[16\]
rlabel metal1 18492 29070 18492 29070 0 CLKDIV.count\[17\]
rlabel metal1 17296 27982 17296 27982 0 CLKDIV.count\[18\]
rlabel metal1 20792 28050 20792 28050 0 CLKDIV.count\[19\]
rlabel metal1 7176 24854 7176 24854 0 CLKDIV.count\[1\]
rlabel metal1 21344 27302 21344 27302 0 CLKDIV.count\[20\]
rlabel viali 21850 28527 21850 28527 0 CLKDIV.count\[21\]
rlabel metal1 22908 29002 22908 29002 0 CLKDIV.count\[22\]
rlabel metal1 21666 28968 21666 28968 0 CLKDIV.count\[23\]
rlabel metal1 5658 24718 5658 24718 0 CLKDIV.count\[2\]
rlabel metal2 6486 25024 6486 25024 0 CLKDIV.count\[3\]
rlabel metal2 6394 28118 6394 28118 0 CLKDIV.count\[4\]
rlabel metal1 6532 28458 6532 28458 0 CLKDIV.count\[5\]
rlabel metal1 5934 28730 5934 28730 0 CLKDIV.count\[6\]
rlabel metal1 7268 28050 7268 28050 0 CLKDIV.count\[7\]
rlabel metal1 9154 28628 9154 28628 0 CLKDIV.count\[8\]
rlabel metal1 9660 27982 9660 27982 0 CLKDIV.count\[9\]
rlabel metal1 19826 24208 19826 24208 0 CLKDIV.secpulse
rlabel metal1 16376 21862 16376 21862 0 CTR.minutes
rlabel metal1 20792 24786 20792 24786 0 CTR.time_out\[0\]
rlabel metal1 8004 6698 8004 6698 0 CTR.time_out\[10\]
rlabel metal1 15594 8534 15594 8534 0 CTR.time_out\[11\]
rlabel metal1 20286 24786 20286 24786 0 CTR.time_out\[1\]
rlabel via1 19366 19363 19366 19363 0 CTR.time_out\[2\]
rlabel metal1 16882 25194 16882 25194 0 CTR.time_out\[3\]
rlabel metal1 5658 21488 5658 21488 0 CTR.time_out\[4\]
rlabel metal1 17618 18734 17618 18734 0 CTR.time_out\[5\]
rlabel metal2 7406 16150 7406 16150 0 CTR.time_out\[6\]
rlabel metal1 7590 11016 7590 11016 0 CTR.time_out\[7\]
rlabel metal1 7130 6800 7130 6800 0 CTR.time_out\[8\]
rlabel via1 14122 8058 14122 8058 0 CTR.time_out\[9\]
rlabel metal1 20470 14586 20470 14586 0 FSM.next_state\[0\]
rlabel metal1 18354 12920 18354 12920 0 FSM.next_state\[1\]
rlabel metal1 20046 11322 20046 11322 0 FSM.next_state\[2\]
rlabel metal1 23138 10744 23138 10744 0 FSM.next_state\[3\]
rlabel metal1 22126 14960 22126 14960 0 FSM.state\[0\]
rlabel metal1 24288 11050 24288 11050 0 FSM.state\[1\]
rlabel metal1 23736 11730 23736 11730 0 FSM.state\[2\]
rlabel metal1 19734 10540 19734 10540 0 FSM.state\[3\]
rlabel metal1 10672 8942 10672 8942 0 MEM.addr\[0\]
rlabel metal1 10856 9010 10856 9010 0 MEM.addr\[1\]
rlabel metal2 12604 5134 12604 5134 0 MEM.addr\[2\]
rlabel metal2 16146 17442 16146 17442 0 MEM.mem1\[0\]
rlabel metal1 20010 8942 20010 8942 0 MEM.mem1\[10\]
rlabel metal1 15686 14450 15686 14450 0 MEM.mem1\[11\]
rlabel metal2 18446 21828 18446 21828 0 MEM.mem1\[1\]
rlabel metal1 18860 20978 18860 20978 0 MEM.mem1\[2\]
rlabel metal1 18906 17272 18906 17272 0 MEM.mem1\[3\]
rlabel metal2 15870 19108 15870 19108 0 MEM.mem1\[4\]
rlabel metal1 18860 18734 18860 18734 0 MEM.mem1\[5\]
rlabel metal1 15640 16014 15640 16014 0 MEM.mem1\[6\]
rlabel metal2 18078 11492 18078 11492 0 MEM.mem1\[7\]
rlabel metal2 18354 9724 18354 9724 0 MEM.mem1\[8\]
rlabel metal1 16652 13294 16652 13294 0 MEM.mem1\[9\]
rlabel viali 11546 17646 11546 17646 0 MEM.mem2\[0\]
rlabel metal1 6072 6222 6072 6222 0 MEM.mem2\[10\]
rlabel metal2 10994 15878 10994 15878 0 MEM.mem2\[11\]
rlabel via1 10534 21998 10534 21998 0 MEM.mem2\[1\]
rlabel metal2 11500 21114 11500 21114 0 MEM.mem2\[2\]
rlabel metal1 5336 18054 5336 18054 0 MEM.mem2\[3\]
rlabel metal2 5566 21828 5566 21828 0 MEM.mem2\[4\]
rlabel metal1 7774 21318 7774 21318 0 MEM.mem2\[5\]
rlabel metal1 5888 15674 5888 15674 0 MEM.mem2\[6\]
rlabel metal2 6946 12852 6946 12852 0 MEM.mem2\[7\]
rlabel metal1 5658 6834 5658 6834 0 MEM.mem2\[8\]
rlabel via1 10534 13294 10534 13294 0 MEM.mem2\[9\]
rlabel metal1 13662 18190 13662 18190 0 MEM.mem3\[0\]
rlabel metal2 8234 7344 8234 7344 0 MEM.mem3\[10\]
rlabel metal1 12650 15436 12650 15436 0 MEM.mem3\[11\]
rlabel metal1 11914 19278 11914 19278 0 MEM.mem3\[1\]
rlabel metal1 13984 20434 13984 20434 0 MEM.mem3\[2\]
rlabel metal1 7406 17680 7406 17680 0 MEM.mem3\[3\]
rlabel metal1 7682 20230 7682 20230 0 MEM.mem3\[4\]
rlabel metal1 8878 18938 8878 18938 0 MEM.mem3\[5\]
rlabel metal1 8234 14790 8234 14790 0 MEM.mem3\[6\]
rlabel metal1 7268 11730 7268 11730 0 MEM.mem3\[7\]
rlabel metal1 7314 6290 7314 6290 0 MEM.mem3\[8\]
rlabel metal1 13800 12818 13800 12818 0 MEM.mem3\[9\]
rlabel metal2 13938 18088 13938 18088 0 MEM.mem4\[0\]
rlabel metal1 4738 9010 4738 9010 0 MEM.mem4\[10\]
rlabel metal1 13662 15470 13662 15470 0 MEM.mem4\[11\]
rlabel metal1 12650 21590 12650 21590 0 MEM.mem4\[1\]
rlabel metal1 14490 20808 14490 20808 0 MEM.mem4\[2\]
rlabel metal1 5750 15130 5750 15130 0 MEM.mem4\[3\]
rlabel metal1 3910 19754 3910 19754 0 MEM.mem4\[4\]
rlabel metal1 9292 19278 9292 19278 0 MEM.mem4\[5\]
rlabel metal1 8556 15674 8556 15674 0 MEM.mem4\[6\]
rlabel metal1 4554 11084 4554 11084 0 MEM.mem4\[7\]
rlabel metal2 4094 9826 4094 9826 0 MEM.mem4\[8\]
rlabel metal1 14306 12206 14306 12206 0 MEM.mem4\[9\]
rlabel metal2 11362 17986 11362 17986 0 MEM.mem5\[0\]
rlabel metal1 4186 8330 4186 8330 0 MEM.mem5\[10\]
rlabel metal1 10948 15674 10948 15674 0 MEM.mem5\[11\]
rlabel metal1 10948 21658 10948 21658 0 MEM.mem5\[1\]
rlabel metal2 10810 21148 10810 21148 0 MEM.mem5\[2\]
rlabel metal1 4830 18734 4830 18734 0 MEM.mem5\[3\]
rlabel metal1 5658 21114 5658 21114 0 MEM.mem5\[4\]
rlabel metal1 7728 22202 7728 22202 0 MEM.mem5\[5\]
rlabel metal1 4462 15980 4462 15980 0 MEM.mem5\[6\]
rlabel metal1 4370 11730 4370 11730 0 MEM.mem5\[7\]
rlabel metal1 4232 7854 4232 7854 0 MEM.mem5\[8\]
rlabel metal2 10810 13566 10810 13566 0 MEM.mem5\[9\]
rlabel metal1 15548 17034 15548 17034 0 MEM.next_mem1\[0\]
rlabel metal1 18860 8398 18860 8398 0 MEM.next_mem1\[10\]
rlabel metal2 15502 14348 15502 14348 0 MEM.next_mem1\[11\]
rlabel metal1 16744 21114 16744 21114 0 MEM.next_mem1\[1\]
rlabel metal2 17894 20094 17894 20094 0 MEM.next_mem1\[2\]
rlabel metal1 18216 17306 18216 17306 0 MEM.next_mem1\[3\]
rlabel metal1 14996 18802 14996 18802 0 MEM.next_mem1\[4\]
rlabel metal1 17342 18360 17342 18360 0 MEM.next_mem1\[5\]
rlabel metal1 15502 15538 15502 15538 0 MEM.next_mem1\[6\]
rlabel metal1 16422 11050 16422 11050 0 MEM.next_mem1\[7\]
rlabel metal1 17066 9690 17066 9690 0 MEM.next_mem1\[8\]
rlabel metal1 16146 12750 16146 12750 0 MEM.next_mem1\[9\]
rlabel metal2 9890 17578 9890 17578 0 MEM.next_mem2\[0\]
rlabel metal1 5421 5882 5421 5882 0 MEM.next_mem2\[10\]
rlabel metal1 9522 15096 9522 15096 0 MEM.next_mem2\[11\]
rlabel metal1 9292 22746 9292 22746 0 MEM.next_mem2\[1\]
rlabel metal1 9614 21930 9614 21930 0 MEM.next_mem2\[2\]
rlabel metal1 5152 17306 5152 17306 0 MEM.next_mem2\[3\]
rlabel metal1 5382 23086 5382 23086 0 MEM.next_mem2\[4\]
rlabel metal1 7452 21454 7452 21454 0 MEM.next_mem2\[5\]
rlabel metal1 5198 15538 5198 15538 0 MEM.next_mem2\[6\]
rlabel metal1 5842 12274 5842 12274 0 MEM.next_mem2\[7\]
rlabel metal1 4186 6392 4186 6392 0 MEM.next_mem2\[8\]
rlabel metal1 10948 13430 10948 13430 0 MEM.next_mem2\[9\]
rlabel metal1 12466 17272 12466 17272 0 MEM.next_mem3\[0\]
rlabel metal1 7360 5134 7360 5134 0 MEM.next_mem3\[10\]
rlabel metal1 11999 14586 11999 14586 0 MEM.next_mem3\[11\]
rlabel metal1 10810 18802 10810 18802 0 MEM.next_mem3\[1\]
rlabel metal2 12098 20196 12098 20196 0 MEM.next_mem3\[2\]
rlabel metal1 5704 17578 5704 17578 0 MEM.next_mem3\[3\]
rlabel metal1 6808 20026 6808 20026 0 MEM.next_mem3\[4\]
rlabel metal1 7590 18802 7590 18802 0 MEM.next_mem3\[5\]
rlabel metal1 7268 14586 7268 14586 0 MEM.next_mem3\[6\]
rlabel metal1 6801 11322 6801 11322 0 MEM.next_mem3\[7\]
rlabel metal1 6946 5746 6946 5746 0 MEM.next_mem3\[8\]
rlabel metal2 12834 12517 12834 12517 0 MEM.next_mem3\[9\]
rlabel metal2 14674 17136 14674 17136 0 MEM.next_mem4\[0\]
rlabel metal2 5658 9248 5658 9248 0 MEM.next_mem4\[10\]
rlabel metal1 12466 15096 12466 15096 0 MEM.next_mem4\[11\]
rlabel metal1 13340 19482 13340 19482 0 MEM.next_mem4\[1\]
rlabel metal1 14444 20570 14444 20570 0 MEM.next_mem4\[2\]
rlabel metal1 4370 15096 4370 15096 0 MEM.next_mem4\[3\]
rlabel metal1 3910 19958 3910 19958 0 MEM.next_mem4\[4\]
rlabel metal1 8372 19414 8372 19414 0 MEM.next_mem4\[5\]
rlabel metal1 7314 15538 7314 15538 0 MEM.next_mem4\[6\]
rlabel metal1 5244 10778 5244 10778 0 MEM.next_mem4\[7\]
rlabel metal2 4186 9962 4186 9962 0 MEM.next_mem4\[8\]
rlabel metal1 14582 12342 14582 12342 0 MEM.next_mem4\[9\]
rlabel metal1 10028 17578 10028 17578 0 MEM.next_mem5\[0\]
rlabel metal1 4554 8364 4554 8364 0 MEM.next_mem5\[10\]
rlabel metal1 9745 15674 9745 15674 0 MEM.next_mem5\[11\]
rlabel metal2 12834 23222 12834 23222 0 MEM.next_mem5\[1\]
rlabel metal1 10488 20570 10488 20570 0 MEM.next_mem5\[2\]
rlabel metal2 4554 17442 4554 17442 0 MEM.next_mem5\[3\]
rlabel metal1 3900 21114 3900 21114 0 MEM.next_mem5\[4\]
rlabel metal1 6801 22202 6801 22202 0 MEM.next_mem5\[5\]
rlabel metal2 3358 16252 3358 16252 0 MEM.next_mem5\[6\]
rlabel metal2 4370 11492 4370 11492 0 MEM.next_mem5\[7\]
rlabel metal1 4002 7990 4002 7990 0 MEM.next_mem5\[8\]
rlabel metal1 9522 12920 9522 12920 0 MEM.next_mem5\[9\]
rlabel metal1 9246 8568 9246 8568 0 MEM.raddr\[0\]
rlabel metal1 10557 11730 10557 11730 0 MEM.raddr\[1\]
rlabel metal1 6394 9622 6394 9622 0 MEM.raddr\[2\]
rlabel metal1 21298 17714 21298 17714 0 TIM.cnt\[0\]
rlabel metal1 18722 7786 18722 7786 0 TIM.cnt\[10\]
rlabel metal1 16238 12104 16238 12104 0 TIM.cnt\[11\]
rlabel metal1 21482 19414 21482 19414 0 TIM.cnt\[1\]
rlabel metal1 19918 19720 19918 19720 0 TIM.cnt\[2\]
rlabel metal1 25944 17510 25944 17510 0 TIM.cnt\[3\]
rlabel metal2 20010 19584 20010 19584 0 TIM.cnt\[4\]
rlabel metal2 23322 17714 23322 17714 0 TIM.cnt\[5\]
rlabel metal1 18262 9928 18262 9928 0 TIM.cnt\[6\]
rlabel metal1 23000 8466 23000 8466 0 TIM.cnt\[7\]
rlabel metal2 17526 8806 17526 8806 0 TIM.cnt\[8\]
rlabel metal2 17434 7905 17434 7905 0 TIM.cnt\[9\]
rlabel metal1 7537 25466 7537 25466 0 _0000_
rlabel metal1 10948 28594 10948 28594 0 _0001_
rlabel metal1 11270 29002 11270 29002 0 _0002_
rlabel metal1 11171 26554 11171 26554 0 _0003_
rlabel metal1 13018 27438 13018 27438 0 _0004_
rlabel metal1 14352 27982 14352 27982 0 _0005_
rlabel metal1 14352 28730 14352 28730 0 _0006_
rlabel metal1 16974 29240 16974 29240 0 _0007_
rlabel metal1 17112 28594 17112 28594 0 _0008_
rlabel metal1 16790 27336 16790 27336 0 _0009_
rlabel metal1 19320 27982 19320 27982 0 _0010_
rlabel metal1 3772 24378 3772 24378 0 _0011_
rlabel metal2 22586 27744 22586 27744 0 _0012_
rlabel metal1 22954 28594 22954 28594 0 _0013_
rlabel metal1 23138 28118 23138 28118 0 _0014_
rlabel metal1 20332 29206 20332 29206 0 _0015_
rlabel metal1 7038 24106 7038 24106 0 _0016_
rlabel metal2 5014 25500 5014 25500 0 _0017_
rlabel metal1 3496 28186 3496 28186 0 _0018_
rlabel metal1 4002 28152 4002 28152 0 _0019_
rlabel metal1 4784 28458 4784 28458 0 _0020_
rlabel metal1 7222 29240 7222 29240 0 _0021_
rlabel metal1 7498 27982 7498 27982 0 _0022_
rlabel metal1 8234 27064 8234 27064 0 _0023_
rlabel metal2 21942 26656 21942 26656 0 _0024_
rlabel metal1 20654 7922 20654 7922 0 _0025_
rlabel metal2 22402 7344 22402 7344 0 _0026_
rlabel metal1 23591 6970 23591 6970 0 _0027_
rlabel metal1 25438 7446 25438 7446 0 _0028_
rlabel metal1 26542 8840 26542 8840 0 _0029_
rlabel metal1 25346 10778 25346 10778 0 _0030_
rlabel metal1 14805 22202 14805 22202 0 _0031_
rlabel metal1 2070 13498 2070 13498 0 _0032_
rlabel metal1 2392 12410 2392 12410 0 _0033_
rlabel metal1 13708 9622 13708 9622 0 _0034_
rlabel metal1 13432 7446 13432 7446 0 _0035_
rlabel metal1 13754 6392 13754 6392 0 _0036_
rlabel via1 13665 8806 13665 8806 0 _0037_
rlabel metal1 23276 17850 23276 17850 0 _0038_
rlabel metal1 24646 14586 24646 14586 0 _0039_
rlabel metal2 27094 14620 27094 14620 0 _0040_
rlabel metal1 27232 17850 27232 17850 0 _0041_
rlabel metal1 23782 17272 23782 17272 0 _0042_
rlabel metal1 24564 13838 24564 13838 0 _0043_
rlabel metal1 9246 9010 9246 9010 0 _0044_
rlabel metal1 9752 10778 9752 10778 0 _0045_
rlabel metal2 6578 9180 6578 9180 0 _0046_
rlabel metal1 20608 17306 20608 17306 0 _0047_
rlabel metal2 9338 5100 9338 5100 0 _0048_
rlabel metal1 9338 5134 9338 5134 0 _0049_
rlabel metal1 11868 5202 11868 5202 0 _0050_
rlabel metal1 17986 24650 17986 24650 0 _0051_
rlabel metal1 18584 24854 18584 24854 0 _0052_
rlabel metal1 16274 24378 16274 24378 0 _0053_
rlabel metal2 14950 25058 14950 25058 0 _0054_
rlabel metal1 13294 23800 13294 23800 0 _0055_
rlabel metal1 11868 24854 11868 24854 0 _0056_
rlabel metal1 6164 25806 6164 25806 0 _0057_
rlabel metal2 5658 25228 5658 25228 0 _0058_
rlabel metal1 7084 26010 7084 26010 0 _0059_
rlabel metal1 14444 27574 14444 27574 0 _0060_
rlabel metal2 12926 28458 12926 28458 0 _0061_
rlabel via2 13662 28611 13662 28611 0 _0062_
rlabel metal2 17986 28033 17986 28033 0 _0063_
rlabel metal2 13662 27047 13662 27047 0 _0064_
rlabel metal1 19688 28594 19688 28594 0 _0065_
rlabel metal1 20378 10132 20378 10132 0 _0066_
rlabel metal1 18998 13260 18998 13260 0 _0067_
rlabel metal1 18952 10778 18952 10778 0 _0068_
rlabel metal1 15364 16558 15364 16558 0 _0069_
rlabel metal2 10258 20366 10258 20366 0 _0070_
rlabel metal1 15548 19822 15548 19822 0 _0071_
rlabel metal1 9430 13226 9430 13226 0 _0072_
rlabel metal1 5244 9078 5244 9078 0 _0073_
rlabel metal1 7774 12410 7774 12410 0 _0074_
rlabel viali 7776 20910 7776 20910 0 _0075_
rlabel metal2 10718 13770 10718 13770 0 _0076_
rlabel metal1 11086 13974 11086 13974 0 _0077_
rlabel metal1 14490 13294 14490 13294 0 _0078_
rlabel metal2 7314 18700 7314 18700 0 _0079_
rlabel metal1 14214 13940 14214 13940 0 _0080_
rlabel metal2 16790 12750 16790 12750 0 _0081_
rlabel metal1 22011 13294 22011 13294 0 _0082_
rlabel metal1 22908 10778 22908 10778 0 _0083_
rlabel metal1 23736 12070 23736 12070 0 _0084_
rlabel metal1 21988 13430 21988 13430 0 _0085_
rlabel metal1 15916 14382 15916 14382 0 _0086_
rlabel metal1 16330 11866 16330 11866 0 _0087_
rlabel metal1 16744 12342 16744 12342 0 _0088_
rlabel metal1 16146 13192 16146 13192 0 _0089_
rlabel metal1 15226 12954 15226 12954 0 _0090_
rlabel metal1 15594 13328 15594 13328 0 _0091_
rlabel metal1 16744 13430 16744 13430 0 _0092_
rlabel metal1 17296 6766 17296 6766 0 _0093_
rlabel metal1 5382 8466 5382 8466 0 _0094_
rlabel metal1 5382 7514 5382 7514 0 _0095_
rlabel metal2 5106 8602 5106 8602 0 _0096_
rlabel metal1 5336 8534 5336 8534 0 _0097_
rlabel metal1 5520 8602 5520 8602 0 _0098_
rlabel via1 17968 7854 17968 7854 0 _0099_
rlabel metal1 17158 7412 17158 7412 0 _0100_
rlabel metal2 17434 6970 17434 6970 0 _0101_
rlabel metal1 17342 4998 17342 4998 0 _0102_
rlabel metal1 18722 5168 18722 5168 0 _0103_
rlabel metal1 6946 7854 6946 7854 0 _0104_
rlabel metal1 5842 8058 5842 8058 0 _0105_
rlabel metal1 6762 7922 6762 7922 0 _0106_
rlabel metal1 6164 7786 6164 7786 0 _0107_
rlabel metal1 14398 6936 14398 6936 0 _0108_
rlabel metal1 17324 8466 17324 8466 0 _0109_
rlabel metal1 17112 8466 17112 8466 0 _0110_
rlabel metal2 18538 4352 18538 4352 0 _0111_
rlabel metal1 18216 5542 18216 5542 0 _0112_
rlabel metal1 17434 6358 17434 6358 0 _0113_
rlabel metal1 6946 10642 6946 10642 0 _0114_
rlabel metal1 6578 10506 6578 10506 0 _0115_
rlabel metal1 6348 10574 6348 10574 0 _0116_
rlabel metal1 5980 10710 5980 10710 0 _0117_
rlabel metal1 9614 10608 9614 10608 0 _0118_
rlabel metal1 17048 10642 17048 10642 0 _0119_
rlabel metal1 16698 10642 16698 10642 0 _0120_
rlabel metal1 17480 10438 17480 10438 0 _0121_
rlabel metal2 16974 5338 16974 5338 0 _0122_
rlabel metal1 17526 4726 17526 4726 0 _0123_
rlabel metal1 16238 4794 16238 4794 0 _0124_
rlabel metal2 18630 4641 18630 4641 0 _0125_
rlabel metal1 19182 4590 19182 4590 0 _0126_
rlabel metal1 18078 2992 18078 2992 0 _0127_
rlabel metal1 19780 4590 19780 4590 0 _0128_
rlabel metal1 17480 6426 17480 6426 0 _0129_
rlabel metal1 20516 4590 20516 4590 0 _0130_
rlabel metal1 19642 5134 19642 5134 0 _0131_
rlabel metal1 20194 5202 20194 5202 0 _0132_
rlabel metal2 20194 3740 20194 3740 0 _0133_
rlabel metal1 19274 4556 19274 4556 0 _0134_
rlabel metal2 28106 4998 28106 4998 0 _0135_
rlabel metal1 5198 24820 5198 24820 0 _0136_
rlabel metal1 4278 24242 4278 24242 0 _0137_
rlabel metal1 6486 25772 6486 25772 0 _0138_
rlabel metal1 6992 25466 6992 25466 0 _0139_
rlabel metal1 5152 25874 5152 25874 0 _0140_
rlabel metal1 5014 25908 5014 25908 0 _0141_
rlabel metal2 4278 28050 4278 28050 0 _0142_
rlabel metal1 4416 27438 4416 27438 0 _0143_
rlabel metal1 4646 27608 4646 27608 0 _0144_
rlabel metal1 7406 29512 7406 29512 0 _0145_
rlabel metal2 5842 28696 5842 28696 0 _0146_
rlabel metal2 6026 28866 6026 28866 0 _0147_
rlabel metal1 7590 28730 7590 28730 0 _0148_
rlabel metal1 7452 28186 7452 28186 0 _0149_
rlabel metal1 7360 28662 7360 28662 0 _0150_
rlabel metal1 7590 28390 7590 28390 0 _0151_
rlabel metal1 8510 28594 8510 28594 0 _0152_
rlabel metal1 9936 28186 9936 28186 0 _0153_
rlabel metal1 9154 27404 9154 27404 0 _0154_
rlabel metal1 11408 28730 11408 28730 0 _0155_
rlabel metal1 11040 29070 11040 29070 0 _0156_
rlabel metal2 12650 29002 12650 29002 0 _0157_
rlabel metal1 11960 27438 11960 27438 0 _0158_
rlabel metal2 12742 27183 12742 27183 0 _0159_
rlabel metal2 11914 27132 11914 27132 0 _0160_
rlabel metal1 15318 28458 15318 28458 0 _0161_
rlabel metal1 14858 26826 14858 26826 0 _0162_
rlabel metal1 14536 28662 14536 28662 0 _0163_
rlabel metal1 15134 28492 15134 28492 0 _0164_
rlabel metal2 16238 29410 16238 29410 0 _0165_
rlabel metal2 16698 28968 16698 28968 0 _0166_
rlabel metal2 16514 29410 16514 29410 0 _0167_
rlabel metal1 17204 27846 17204 27846 0 _0168_
rlabel metal1 17802 26826 17802 26826 0 _0169_
rlabel metal1 17020 27098 17020 27098 0 _0170_
rlabel metal1 19504 27370 19504 27370 0 _0171_
rlabel metal2 22678 27744 22678 27744 0 _0172_
rlabel metal1 21068 27098 21068 27098 0 _0173_
rlabel metal1 22172 28458 22172 28458 0 _0174_
rlabel metal1 22770 27540 22770 27540 0 _0175_
rlabel metal1 20378 28696 20378 28696 0 _0176_
rlabel metal1 20532 28458 20532 28458 0 _0177_
rlabel metal1 20700 28730 20700 28730 0 _0178_
rlabel metal1 6992 19822 6992 19822 0 _0179_
rlabel metal1 7682 19720 7682 19720 0 _0180_
rlabel metal1 16514 20026 16514 20026 0 _0181_
rlabel metal2 17250 19958 17250 19958 0 _0182_
rlabel metal2 21114 20774 21114 20774 0 _0183_
rlabel metal1 6486 13498 6486 13498 0 _0184_
rlabel metal2 6394 15776 6394 15776 0 _0185_
rlabel metal2 7682 17850 7682 17850 0 _0186_
rlabel metal2 19458 17935 19458 17935 0 _0187_
rlabel metal2 19274 17748 19274 17748 0 _0188_
rlabel metal2 14260 20332 14260 20332 0 _0189_
rlabel metal2 19826 18054 19826 18054 0 _0190_
rlabel metal1 20608 18122 20608 18122 0 _0191_
rlabel metal1 13754 20842 13754 20842 0 _0192_
rlabel metal1 19826 20876 19826 20876 0 _0193_
rlabel metal1 19458 20944 19458 20944 0 _0194_
rlabel metal2 20378 21216 20378 21216 0 _0195_
rlabel metal2 23874 20604 23874 20604 0 _0196_
rlabel metal1 11592 21862 11592 21862 0 _0197_
rlabel metal1 19136 20434 19136 20434 0 _0198_
rlabel metal1 18722 20502 18722 20502 0 _0199_
rlabel metal2 8694 22406 8694 22406 0 _0200_
rlabel metal2 20562 19924 20562 19924 0 _0201_
rlabel metal2 19182 20536 19182 20536 0 _0202_
rlabel metal2 22218 20961 22218 20961 0 _0203_
rlabel metal1 8786 18734 8786 18734 0 _0204_
rlabel metal1 18492 19482 18492 19482 0 _0205_
rlabel metal2 20286 19091 20286 19091 0 _0206_
rlabel metal1 19642 18938 19642 18938 0 _0207_
rlabel metal1 18722 19176 18722 19176 0 _0208_
rlabel metal2 22862 21522 22862 21522 0 _0209_
rlabel metal1 20378 21998 20378 21998 0 _0210_
rlabel metal2 20838 21828 20838 21828 0 _0211_
rlabel metal1 21022 21454 21022 21454 0 _0212_
rlabel metal1 21206 21386 21206 21386 0 _0213_
rlabel via2 20378 21845 20378 21845 0 _0214_
rlabel metal1 24288 4182 24288 4182 0 _0215_
rlabel metal1 23368 21998 23368 21998 0 _0216_
rlabel viali 24610 21995 24610 21995 0 _0217_
rlabel metal1 23736 21522 23736 21522 0 _0218_
rlabel metal1 25208 21862 25208 21862 0 _0219_
rlabel metal1 21574 22644 21574 22644 0 _0220_
rlabel metal1 24564 4114 24564 4114 0 _0221_
rlabel metal1 25208 3502 25208 3502 0 _0222_
rlabel metal1 24886 21930 24886 21930 0 _0223_
rlabel metal1 25622 21998 25622 21998 0 _0224_
rlabel metal1 25438 20978 25438 20978 0 _0225_
rlabel metal2 2438 4063 2438 4063 0 _0226_
rlabel metal1 2599 3502 2599 3502 0 _0227_
rlabel metal2 25254 26452 25254 26452 0 _0228_
rlabel metal2 19780 21556 19780 21556 0 _0229_
rlabel metal1 11546 9622 11546 9622 0 _0230_
rlabel metal1 9430 10098 9430 10098 0 _0231_
rlabel metal1 11546 7174 11546 7174 0 _0232_
rlabel metal3 14628 9588 14628 9588 0 _0233_
rlabel metal1 21942 14280 21942 14280 0 _0234_
rlabel metal1 24150 11118 24150 11118 0 _0235_
rlabel metal1 19274 13974 19274 13974 0 _0236_
rlabel metal2 16882 9214 16882 9214 0 _0237_
rlabel metal1 19918 15436 19918 15436 0 _0238_
rlabel metal1 10350 7412 10350 7412 0 _0239_
rlabel metal1 11776 13294 11776 13294 0 _0240_
rlabel metal1 10580 6358 10580 6358 0 _0241_
rlabel metal1 12466 9894 12466 9894 0 _0242_
rlabel metal1 10580 6426 10580 6426 0 _0243_
rlabel metal1 10074 16456 10074 16456 0 _0244_
rlabel metal1 11868 6290 11868 6290 0 _0245_
rlabel metal1 7682 14382 7682 14382 0 _0246_
rlabel metal1 7222 6698 7222 6698 0 _0247_
rlabel metal1 11592 8942 11592 8942 0 _0248_
rlabel metal2 13202 19584 13202 19584 0 _0249_
rlabel metal1 13938 19346 13938 19346 0 _0250_
rlabel metal2 11086 6324 11086 6324 0 _0251_
rlabel metal2 11362 7140 11362 7140 0 _0252_
rlabel metal2 12650 22406 12650 22406 0 _0253_
rlabel metal1 12466 22712 12466 22712 0 _0254_
rlabel metal2 12650 18054 12650 18054 0 _0255_
rlabel metal1 17342 17238 17342 17238 0 _0256_
rlabel metal1 17526 17102 17526 17102 0 _0257_
rlabel metal1 25622 20842 25622 20842 0 _0258_
rlabel metal1 27370 20876 27370 20876 0 _0259_
rlabel metal1 25944 20774 25944 20774 0 _0260_
rlabel metal1 28290 20978 28290 20978 0 _0261_
rlabel metal2 23690 20876 23690 20876 0 _0262_
rlabel metal1 24104 20570 24104 20570 0 _0263_
rlabel metal1 20838 22746 20838 22746 0 _0264_
rlabel metal1 20700 21930 20700 21930 0 _0265_
rlabel metal1 21298 22032 21298 22032 0 _0266_
rlabel metal1 23046 21658 23046 21658 0 _0267_
rlabel metal2 21114 22202 21114 22202 0 _0268_
rlabel metal2 21666 22338 21666 22338 0 _0269_
rlabel via1 23899 22610 23899 22610 0 _0270_
rlabel metal2 24978 21420 24978 21420 0 _0271_
rlabel metal1 24380 21522 24380 21522 0 _0272_
rlabel metal1 26220 20910 26220 20910 0 _0273_
rlabel metal1 27554 19686 27554 19686 0 _0274_
rlabel metal2 27554 20026 27554 20026 0 _0275_
rlabel metal1 22264 21998 22264 21998 0 _0276_
rlabel metal1 22862 21930 22862 21930 0 _0277_
rlabel metal1 22678 22032 22678 22032 0 _0278_
rlabel metal2 22494 21692 22494 21692 0 _0279_
rlabel metal1 21804 20230 21804 20230 0 _0280_
rlabel metal1 21720 20570 21720 20570 0 _0281_
rlabel metal1 22402 20570 22402 20570 0 _0282_
rlabel metal1 21850 21488 21850 21488 0 _0283_
rlabel metal2 21850 21471 21850 21471 0 _0284_
rlabel metal2 27278 20570 27278 20570 0 _0285_
rlabel metal1 27048 21114 27048 21114 0 _0286_
rlabel metal1 27876 20026 27876 20026 0 _0287_
rlabel metal1 28290 19822 28290 19822 0 _0288_
rlabel viali 28567 20456 28567 20456 0 _0289_
rlabel metal1 16790 3570 16790 3570 0 _0290_
rlabel metal1 18078 5678 18078 5678 0 _0291_
rlabel metal1 18400 3162 18400 3162 0 _0292_
rlabel metal1 18170 3366 18170 3366 0 _0293_
rlabel metal1 17388 3026 17388 3026 0 _0294_
rlabel metal1 17204 2958 17204 2958 0 _0295_
rlabel metal1 16882 3468 16882 3468 0 _0296_
rlabel metal1 16008 3502 16008 3502 0 _0297_
rlabel metal1 14628 4114 14628 4114 0 _0298_
rlabel metal1 13079 4114 13079 4114 0 _0299_
rlabel metal1 16330 4148 16330 4148 0 _0300_
rlabel metal1 17079 5338 17079 5338 0 _0301_
rlabel metal1 17618 4658 17618 4658 0 _0302_
rlabel metal1 16790 7344 16790 7344 0 _0303_
rlabel metal1 17848 6766 17848 6766 0 _0304_
rlabel metal1 17618 6290 17618 6290 0 _0305_
rlabel metal2 17618 5440 17618 5440 0 _0306_
rlabel metal1 16744 4046 16744 4046 0 _0307_
rlabel metal1 13708 2414 13708 2414 0 _0308_
rlabel metal1 8372 14994 8372 14994 0 _0309_
rlabel via1 12558 15045 12558 15045 0 _0310_
rlabel metal2 15180 16422 15180 16422 0 _0311_
rlabel metal1 15640 9894 15640 9894 0 _0312_
rlabel metal2 14858 3876 14858 3876 0 _0313_
rlabel metal1 13386 2618 13386 2618 0 _0314_
rlabel metal2 14030 3774 14030 3774 0 _0315_
rlabel metal1 14858 3162 14858 3162 0 _0316_
rlabel metal2 15318 3230 15318 3230 0 _0317_
rlabel metal2 2438 5575 2438 5575 0 _0318_
rlabel metal1 14076 3366 14076 3366 0 _0319_
rlabel metal2 12650 3978 12650 3978 0 _0320_
rlabel metal1 20792 13770 20792 13770 0 _0321_
rlabel metal1 20516 14382 20516 14382 0 _0322_
rlabel metal1 19688 15470 19688 15470 0 _0323_
rlabel metal1 19458 14960 19458 14960 0 _0324_
rlabel metal2 19274 14688 19274 14688 0 _0325_
rlabel metal1 21390 12716 21390 12716 0 _0326_
rlabel metal1 22862 8432 22862 8432 0 _0327_
rlabel metal1 19090 14484 19090 14484 0 _0328_
rlabel viali 21758 14382 21758 14382 0 _0329_
rlabel metal1 18492 14586 18492 14586 0 _0330_
rlabel metal1 21436 12954 21436 12954 0 _0331_
rlabel metal1 20286 14484 20286 14484 0 _0332_
rlabel metal1 20286 14042 20286 14042 0 _0333_
rlabel viali 20930 14381 20930 14381 0 _0334_
rlabel metal1 16284 14994 16284 14994 0 _0335_
rlabel metal1 17572 14382 17572 14382 0 _0336_
rlabel metal1 18676 13498 18676 13498 0 _0337_
rlabel metal1 18906 13940 18906 13940 0 _0338_
rlabel metal1 19044 13906 19044 13906 0 _0339_
rlabel metal1 19780 13294 19780 13294 0 _0340_
rlabel metal1 19964 13770 19964 13770 0 _0341_
rlabel metal1 19458 14416 19458 14416 0 _0342_
rlabel metal2 19274 13770 19274 13770 0 _0343_
rlabel metal1 19780 13158 19780 13158 0 _0344_
rlabel metal2 21850 12988 21850 12988 0 _0345_
rlabel metal1 23460 12614 23460 12614 0 _0346_
rlabel metal1 22264 8942 22264 8942 0 _0347_
rlabel metal1 26358 16626 26358 16626 0 _0348_
rlabel metal1 24886 16524 24886 16524 0 _0349_
rlabel metal2 26542 16796 26542 16796 0 _0350_
rlabel metal1 27738 17510 27738 17510 0 _0351_
rlabel metal1 28336 16422 28336 16422 0 _0352_
rlabel metal1 23230 16456 23230 16456 0 _0353_
rlabel metal1 23276 14994 23276 14994 0 _0354_
rlabel metal1 22954 9146 22954 9146 0 _0355_
rlabel metal1 23046 14042 23046 14042 0 _0356_
rlabel metal1 23276 14586 23276 14586 0 _0357_
rlabel metal1 25829 17646 25829 17646 0 _0358_
rlabel metal2 23598 16320 23598 16320 0 _0359_
rlabel metal1 27370 17170 27370 17170 0 _0360_
rlabel metal2 24012 11628 24012 11628 0 _0361_
rlabel metal1 26358 10710 26358 10710 0 _0362_
rlabel metal1 21436 8466 21436 8466 0 _0363_
rlabel metal2 25898 8577 25898 8577 0 _0364_
rlabel metal2 22954 7888 22954 7888 0 _0365_
rlabel metal1 23046 7310 23046 7310 0 _0366_
rlabel metal2 22540 7514 22540 7514 0 _0367_
rlabel via1 22586 7852 22586 7852 0 _0368_
rlabel metal1 23828 8330 23828 8330 0 _0369_
rlabel metal2 23782 8126 23782 8126 0 _0370_
rlabel metal1 24702 7446 24702 7446 0 _0371_
rlabel metal1 24794 7854 24794 7854 0 _0372_
rlabel metal1 23874 7344 23874 7344 0 _0373_
rlabel metal1 27554 7956 27554 7956 0 _0374_
rlabel metal1 27968 8466 27968 8466 0 _0375_
rlabel metal2 26634 8194 26634 8194 0 _0376_
rlabel metal1 26542 7514 26542 7514 0 _0377_
rlabel metal1 25806 7786 25806 7786 0 _0378_
rlabel metal1 27554 8432 27554 8432 0 _0379_
rlabel metal1 28520 8874 28520 8874 0 _0380_
rlabel metal1 26772 9486 26772 9486 0 _0381_
rlabel metal2 25806 8704 25806 8704 0 _0382_
rlabel metal1 25668 8942 25668 8942 0 _0383_
rlabel metal1 26266 10642 26266 10642 0 _0384_
rlabel metal2 25622 10404 25622 10404 0 _0385_
rlabel metal1 25668 10642 25668 10642 0 _0386_
rlabel metal1 14628 23290 14628 23290 0 _0387_
rlabel metal1 15686 23800 15686 23800 0 _0388_
rlabel metal1 18216 24854 18216 24854 0 _0389_
rlabel metal1 15916 23562 15916 23562 0 _0390_
rlabel metal2 16744 14246 16744 14246 0 _0391_
rlabel metal1 3312 13158 3312 13158 0 _0392_
rlabel metal1 2530 13294 2530 13294 0 _0393_
rlabel metal1 2990 12274 2990 12274 0 _0394_
rlabel metal1 2898 12308 2898 12308 0 _0395_
rlabel metal2 14582 11152 14582 11152 0 _0396_
rlabel via1 13581 10234 13581 10234 0 _0397_
rlabel metal1 14306 7888 14306 7888 0 _0398_
rlabel metal2 13110 9520 13110 9520 0 _0399_
rlabel metal1 14030 10030 14030 10030 0 _0400_
rlabel metal2 14490 7344 14490 7344 0 _0401_
rlabel metal1 13064 7378 13064 7378 0 _0402_
rlabel metal2 13938 7310 13938 7310 0 _0403_
rlabel metal1 14306 6800 14306 6800 0 _0404_
rlabel metal1 13340 8602 13340 8602 0 _0405_
rlabel metal1 25530 17578 25530 17578 0 _0406_
rlabel metal1 22678 17782 22678 17782 0 _0407_
rlabel metal2 23138 17238 23138 17238 0 _0408_
rlabel metal1 23000 16762 23000 16762 0 _0409_
rlabel metal1 23506 17306 23506 17306 0 _0410_
rlabel metal1 23828 16762 23828 16762 0 _0411_
rlabel metal1 26634 16524 26634 16524 0 _0412_
rlabel metal2 26818 15708 26818 15708 0 _0413_
rlabel metal1 26220 15674 26220 15674 0 _0414_
rlabel metal1 27140 16422 27140 16422 0 _0415_
rlabel metal1 26542 15368 26542 15368 0 _0416_
rlabel viali 24702 15016 24702 15016 0 _0417_
rlabel metal2 27738 15198 27738 15198 0 _0418_
rlabel metal1 27140 15062 27140 15062 0 _0419_
rlabel metal1 27876 16558 27876 16558 0 _0420_
rlabel metal2 27278 15946 27278 15946 0 _0421_
rlabel metal1 27186 14960 27186 14960 0 _0422_
rlabel metal2 27922 17476 27922 17476 0 _0423_
rlabel metal2 27278 17170 27278 17170 0 _0424_
rlabel metal1 27370 17068 27370 17068 0 _0425_
rlabel metal2 28106 17034 28106 17034 0 _0426_
rlabel metal1 27738 17170 27738 17170 0 _0427_
rlabel metal1 26818 18054 26818 18054 0 _0428_
rlabel metal1 25668 17306 25668 17306 0 _0429_
rlabel metal1 24886 16762 24886 16762 0 _0430_
rlabel metal1 10948 10030 10948 10030 0 _0431_
rlabel metal1 9200 9554 9200 9554 0 _0432_
rlabel metal1 10442 10098 10442 10098 0 _0433_
rlabel metal1 10396 10234 10396 10234 0 _0434_
rlabel metal1 10258 10574 10258 10574 0 _0435_
rlabel metal1 10166 9656 10166 9656 0 _0436_
rlabel metal1 11040 9418 11040 9418 0 _0437_
rlabel metal1 10557 9622 10557 9622 0 _0438_
rlabel metal1 8970 9452 8970 9452 0 _0439_
rlabel metal1 22356 16762 22356 16762 0 _0440_
rlabel metal2 22218 16966 22218 16966 0 _0441_
rlabel metal1 21022 17204 21022 17204 0 _0442_
rlabel metal1 10626 5746 10626 5746 0 _0443_
rlabel metal1 9430 5780 9430 5780 0 _0444_
rlabel metal1 10350 5678 10350 5678 0 _0445_
rlabel metal1 11408 4794 11408 4794 0 _0446_
rlabel metal2 17986 25568 17986 25568 0 _0447_
rlabel metal1 17894 24820 17894 24820 0 _0448_
rlabel metal2 19274 24854 19274 24854 0 _0449_
rlabel metal1 19734 25364 19734 25364 0 _0450_
rlabel metal1 17204 23834 17204 23834 0 _0451_
rlabel metal2 15686 24582 15686 24582 0 _0452_
rlabel metal1 15824 24174 15824 24174 0 _0453_
rlabel metal1 15364 23698 15364 23698 0 _0454_
rlabel metal1 15226 24752 15226 24752 0 _0455_
rlabel metal1 15134 24718 15134 24718 0 _0456_
rlabel metal2 15594 23460 15594 23460 0 _0457_
rlabel metal1 14030 23698 14030 23698 0 _0458_
rlabel metal2 15226 23392 15226 23392 0 _0459_
rlabel metal1 13386 23630 13386 23630 0 _0460_
rlabel metal2 13018 24548 13018 24548 0 _0461_
rlabel metal2 14214 12784 14214 12784 0 clk
rlabel metal1 15824 17850 15824 17850 0 clknet_0_clk
rlabel metal1 2714 5712 2714 5712 0 clknet_4_0_0_clk
rlabel metal1 19642 11186 19642 11186 0 clknet_4_10_0_clk
rlabel metal1 26864 14450 26864 14450 0 clknet_4_11_0_clk
rlabel metal1 14766 18326 14766 18326 0 clknet_4_12_0_clk
rlabel metal2 15042 24786 15042 24786 0 clknet_4_13_0_clk
rlabel metal1 17388 25262 17388 25262 0 clknet_4_14_0_clk
rlabel metal1 19918 29036 19918 29036 0 clknet_4_15_0_clk
rlabel metal1 1656 15538 1656 15538 0 clknet_4_1_0_clk
rlabel metal1 13064 6222 13064 6222 0 clknet_4_2_0_clk
rlabel metal2 9246 13838 9246 13838 0 clknet_4_3_0_clk
rlabel metal2 1886 20366 1886 20366 0 clknet_4_4_0_clk
rlabel metal1 5934 24242 5934 24242 0 clknet_4_5_0_clk
rlabel metal1 9062 21590 9062 21590 0 clknet_4_6_0_clk
rlabel metal1 11546 26418 11546 26418 0 clknet_4_7_0_clk
rlabel metal2 17434 15300 17434 15300 0 clknet_4_8_0_clk
rlabel metal1 14766 17714 14766 17714 0 clknet_4_9_0_clk
rlabel metal1 18216 15334 18216 15334 0 e1.edge_d
rlabel metal1 3496 16626 3496 16626 0 e1.intermediate
rlabel via1 17986 15538 17986 15538 0 e1.sync
rlabel metal1 9706 24582 9706 24582 0 e2.edge_d
rlabel metal2 3174 28254 3174 28254 0 e2.intermediate
rlabel metal2 6394 25126 6394 25126 0 e2.sync
rlabel metal1 26496 29138 26496 29138 0 net1
rlabel metal1 28290 18734 28290 18734 0 net10
rlabel metal2 10166 21964 10166 21964 0 net100
rlabel metal1 10258 22066 10258 22066 0 net101
rlabel metal1 19872 27302 19872 27302 0 net102
rlabel metal1 12236 22610 12236 22610 0 net103
rlabel metal1 5014 16490 5014 16490 0 net104
rlabel metal1 14582 27030 14582 27030 0 net105
rlabel metal1 16008 28050 16008 28050 0 net106
rlabel metal1 3358 20400 3358 20400 0 net107
rlabel metal1 12006 12954 12006 12954 0 net108
rlabel metal1 15686 28594 15686 28594 0 net109
rlabel metal1 25622 2414 25622 2414 0 net11
rlabel metal1 4600 7854 4600 7854 0 net110
rlabel metal1 12650 27506 12650 27506 0 net111
rlabel metal1 3404 17170 3404 17170 0 net112
rlabel metal1 9844 27506 9844 27506 0 net113
rlabel metal1 7774 25874 7774 25874 0 net114
rlabel metal2 19182 29478 19182 29478 0 net115
rlabel metal1 10994 29138 10994 29138 0 net116
rlabel metal1 25392 13498 25392 13498 0 net117
rlabel metal1 16330 22610 16330 22610 0 net118
rlabel metal2 9798 28900 9798 28900 0 net119
rlabel metal1 28842 21964 28842 21964 0 net12
rlabel metal1 6992 28526 6992 28526 0 net120
rlabel metal1 5934 26384 5934 26384 0 net121
rlabel metal1 3266 28628 3266 28628 0 net122
rlabel metal1 22678 29172 22678 29172 0 net123
rlabel metal1 23644 27438 23644 27438 0 net124
rlabel metal1 6578 24650 6578 24650 0 net125
rlabel metal2 7314 24922 7314 24922 0 net126
rlabel metal1 26726 7922 26726 7922 0 net127
rlabel metal2 26174 9180 26174 9180 0 net128
rlabel metal1 25806 17782 25806 17782 0 net129
rlabel metal1 1886 3502 1886 3502 0 net13
rlabel metal1 14490 8806 14490 8806 0 net130
rlabel metal2 22494 27608 22494 27608 0 net131
rlabel metal1 25622 14994 25622 14994 0 net132
rlabel metal1 26358 10574 26358 10574 0 net133
rlabel metal1 22770 7446 22770 7446 0 net134
rlabel metal1 10396 5066 10396 5066 0 net135
rlabel metal1 23966 7446 23966 7446 0 net136
rlabel metal1 24426 17714 24426 17714 0 net137
rlabel metal1 1886 2414 1886 2414 0 net14
rlabel metal2 21942 30022 21942 30022 0 net15
rlabel metal1 24886 22746 24886 22746 0 net16
rlabel metal2 1518 23375 1518 23375 0 net17
rlabel metal2 6210 17204 6210 17204 0 net18
rlabel metal2 22126 2890 22126 2890 0 net19
rlabel metal1 1564 16218 1564 16218 0 net2
rlabel metal1 1886 26554 1886 26554 0 net20
rlabel metal1 22080 2958 22080 2958 0 net21
rlabel metal1 5405 2414 5405 2414 0 net22
rlabel metal1 7314 2414 7314 2414 0 net23
rlabel metal1 8280 3978 8280 3978 0 net24
rlabel metal2 28750 6902 28750 6902 0 net25
rlabel metal1 19826 4080 19826 4080 0 net26
rlabel metal1 28566 26962 28566 26962 0 net27
rlabel metal2 20102 6579 20102 6579 0 net28
rlabel metal2 1518 12835 1518 12835 0 net29
rlabel metal1 1656 29206 1656 29206 0 net3
rlabel metal1 18814 4454 18814 4454 0 net30
rlabel metal2 20102 3230 20102 3230 0 net31
rlabel metal1 25116 13362 25116 13362 0 net32
rlabel metal2 13294 13226 13294 13226 0 net33
rlabel metal1 16882 19414 16882 19414 0 net34
rlabel metal2 7130 7242 7130 7242 0 net35
rlabel metal1 13347 14314 13347 14314 0 net36
rlabel metal1 3411 19754 3411 19754 0 net37
rlabel metal1 13570 17129 13570 17129 0 net38
rlabel metal1 20141 25874 20141 25874 0 net39
rlabel metal1 22218 2380 22218 2380 0 net4
rlabel metal1 19550 8568 19550 8568 0 net40
rlabel metal2 14352 18836 14352 18836 0 net41
rlabel metal1 2806 16184 2806 16184 0 net42
rlabel metal1 2162 25160 2162 25160 0 net43
rlabel metal1 8050 24718 8050 24718 0 net44
rlabel metal1 13478 15912 13478 15912 0 net45
rlabel metal1 17434 18768 17434 18768 0 net46
rlabel metal1 18216 17170 18216 17170 0 net47
rlabel metal1 14950 19278 14950 19278 0 net48
rlabel metal1 16698 9588 16698 9588 0 net49
rlabel metal3 9959 21964 9959 21964 0 net5
rlabel metal1 17388 20434 17388 20434 0 net50
rlabel metal1 16652 12818 16652 12818 0 net51
rlabel metal1 15824 11118 15824 11118 0 net52
rlabel via1 11914 15453 11914 15453 0 net53
rlabel metal1 7360 11118 7360 11118 0 net54
rlabel metal1 15732 16082 15732 16082 0 net55
rlabel metal1 6854 6698 6854 6698 0 net56
rlabel metal1 15042 17238 15042 17238 0 net57
rlabel metal1 5934 12920 5934 12920 0 net58
rlabel metal1 7314 19414 7314 19414 0 net59
rlabel via2 2254 11747 2254 11747 0 net6
rlabel metal1 10074 18292 10074 18292 0 net60
rlabel metal1 9890 13940 9890 13940 0 net61
rlabel metal1 7130 14314 7130 14314 0 net62
rlabel metal1 14444 20434 14444 20434 0 net63
rlabel metal1 18032 8942 18032 8942 0 net64
rlabel metal1 6394 19856 6394 19856 0 net65
rlabel metal2 11546 15062 11546 15062 0 net66
rlabel metal1 3818 10540 3818 10540 0 net67
rlabel metal1 12282 12852 12282 12852 0 net68
rlabel metal1 14812 12206 14812 12206 0 net69
rlabel metal1 28336 19686 28336 19686 0 net7
rlabel metal1 9246 20026 9246 20026 0 net70
rlabel metal1 9890 16048 9890 16048 0 net71
rlabel metal2 14122 16762 14122 16762 0 net72
rlabel metal1 5382 6698 5382 6698 0 net73
rlabel metal1 7130 16116 7130 16116 0 net74
rlabel metal1 6762 22644 6762 22644 0 net75
rlabel metal1 14306 19958 14306 19958 0 net76
rlabel metal1 6210 18700 6210 18700 0 net77
rlabel metal1 14950 13974 14950 13974 0 net78
rlabel metal1 4646 10710 4646 10710 0 net79
rlabel metal2 17664 26180 17664 26180 0 net8
rlabel metal1 13386 18394 13386 18394 0 net80
rlabel metal1 5060 9554 5060 9554 0 net81
rlabel metal1 3772 11118 3772 11118 0 net82
rlabel metal1 6670 6426 6670 6426 0 net83
rlabel metal2 7498 6596 7498 6596 0 net84
rlabel metal1 12880 19346 12880 19346 0 net85
rlabel metal1 10258 20434 10258 20434 0 net86
rlabel metal1 15962 20944 15962 20944 0 net87
rlabel metal1 4002 8500 4002 8500 0 net88
rlabel metal1 3174 21590 3174 21590 0 net89
rlabel metal1 28658 2414 28658 2414 0 net9
rlabel metal1 4876 17170 4876 17170 0 net90
rlabel metal1 5934 16762 5934 16762 0 net91
rlabel metal1 10626 19754 10626 19754 0 net92
rlabel metal1 9338 22678 9338 22678 0 net93
rlabel metal2 8510 21726 8510 21726 0 net94
rlabel metal2 4002 17884 4002 17884 0 net95
rlabel metal1 5934 21590 5934 21590 0 net96
rlabel metal1 4600 21454 4600 21454 0 net97
rlabel metal1 10718 16490 10718 16490 0 net98
rlabel metal1 9706 18224 9706 18224 0 net99
rlabel metal1 28382 30260 28382 30260 0 nrst
rlabel metal2 14858 959 14858 959 0 out_0[0]
rlabel metal1 9982 30294 9982 30294 0 out_0[1]
rlabel metal3 820 11628 820 11628 0 out_0[2]
rlabel metal1 28980 11186 28980 11186 0 out_0[3]
rlabel metal1 17618 30090 17618 30090 0 out_0[4]
rlabel metal2 29670 1554 29670 1554 0 out_0[5]
rlabel metal2 29026 18513 29026 18513 0 out_0[6]
rlabel metal2 25806 823 25806 823 0 out_1[0]
rlabel via2 29026 22491 29026 22491 0 out_1[1]
rlabel metal3 820 3468 820 3468 0 out_1[2]
rlabel metal2 46 1520 46 1520 0 out_1[3]
rlabel metal2 21298 31154 21298 31154 0 out_1[4]
rlabel metal1 25576 30294 25576 30294 0 out_1[5]
rlabel metal3 751 23188 751 23188 0 out_1[6]
rlabel metal2 6762 31195 6762 31195 0 out_2[0]
rlabel metal2 21942 1571 21942 1571 0 out_2[1]
rlabel metal3 820 27268 820 27268 0 out_2[2]
rlabel via2 29026 2805 29026 2805 0 out_2[3]
rlabel metal2 3266 1520 3266 1520 0 out_2[4]
rlabel metal2 7130 1520 7130 1520 0 out_2[5]
rlabel metal2 2714 31144 2714 31144 0 out_2[6]
rlabel metal1 28980 7174 28980 7174 0 out_3[0]
rlabel metal2 10994 1095 10994 1095 0 out_3[1]
rlabel metal2 29026 26673 29026 26673 0 out_3[2]
rlabel metal1 28980 30158 28980 30158 0 out_3[3]
rlabel metal3 751 19788 751 19788 0 out_3[4]
rlabel metal1 14122 30090 14122 30090 0 out_3[5]
rlabel metal2 18722 959 18722 959 0 out_3[6]
rlabel metal3 820 15708 820 15708 0 pb_0
rlabel metal3 751 31348 751 31348 0 pb_1
rlabel metal1 28980 13498 28980 13498 0 time_done
<< properties >>
string FIXED_BBOX 0 0 30581 32725
<< end >>
